module s1196(G1,G12,G550,VDD,G542,G532,G0,G7,G2,G547,G539,G548,G552,G13,G4,G6,VSS,G3,G5,G9,G11,G549,G546,G530,G535,G537,CLOCK,G8,G10,G551,G45);
input G1,G4,G6,VSS,VDD,G3,G5,G9,G0,G7,G11,G2,CLOCK,G12,G8,G10,G13;
output G550,G549,G542,G546,G532,G530,G535,G537,G547,G539,G551,G548,G552,G45;

  wire G273,G521,G196,G339,G435,G472,G419,G518,G36,G528,I374,G470,G61,G59,G350,I662,G403,G288,G53,G81,G139,G35,I330,G359,G188,G33,G68,G490,G512,G272,G498,G74,G317,G217,G79,G392,G355,G484,G255,G211,G212,G164,G439,G161,G93,G46,G357,G70,G516,G242,I280,G325,G209,I276,G459,G75,G534,G230,G136,G257,G321,G433,G369,G292,G375,G502,G483,G343,G464,G153,G443,G334,G383,G38,G203,G360,G144,G201,G554,G51,G300,G531,G235,G446,G30,G135,G227,G251,G290,G346,G143,G387,G441,G452,G128,G49,G244,G52,G269,I631,G428,G178,G326,G494,G386,G208,I156,G123,G394,G241,G57,G333,G458,G510,G154,G460,G90,G39,G214,G191,G545,G294,G373,G491,G440,G306,G195,G486,G482,G377,G331,G425,G259,G171,G92,G220,G83,G236,G505,G89,G129,G388,G457,G519,G268,G311,G40,G462,G199,G32,G529,G310,G165,I493,G329,G137,G378,G302,G270,G473,G180,G499,G474,G485,G181,G100,G297,G356,G189,G522,G351,G145,G338,G500,G157,G332,G316,G309,G322,G151,G192,G335,G232,G286,G216,G418,G399,G506,G318,G215,G152,G487,I576,G308,G376,G400,G86,G285,G501,G281,G219,G225,G345,G543,G73,G102,G461,G43,G96,G34,G237,G454,G252,G97,G374,I536,G194,G233,G525,G489,G156,G71,G80,G234,G540,G385,G398,G226,G434,G438,G160,G469,G368,G303,G337,G132,G475,G456,G246,G238,G396,G64,G221,G240,G94,G223,G478,G204,I249,G414,G495,G361,G341,G41,G130,G250,G106,G218,I573,G72,G275,G342,G397,G116,I316,G389,G371,G450,G29,G60,G520,G85,G210,G37,G283,G312,I386,G515,G436,I272,G497,G393,G173,G182,G426,G176,G508,G54,G88,G362,G111,G126,G406,G249,G107,G276,G62,G553,G271,G158,G390,G131,G42,G253,G193,G496,G168,G305,G455,G149,G48,G364,G202,G507,G536,G323,G247,G314,G365,G379,G183,G231,G422,G284,I692,G134,G417,G122,G492,G488,G476,G544,G504,G63,G256,G174,G517,G55,G289,G291,G121,G261,G118,G104,G146,G444,G77,G190,G363,G409,G293,I287,G348,G437,G447,G523,G327,G430,I624,G105,G155,G99,G480,G367,G243,G84,G463,G56,G101,G296,G91,G429,G280,G527,G533,G31,I529,G479,G315,G254,G405,G114,G119,G112,G298,G87,G526,G213,G328,G172,G224,G222,G103,G349,G395,G465,G313,G167,G207,G513,G200,G82,G248,G142,G69,G299,G503,G427,G266,G380,G415,G471,G262,G493,G170,G477,G423,G370,G169,G468,G179,G353,G115,G133,G206,G120,G245,G432,G267,G150,G344,G524,G514,G198,G239,G184,G141,G277,G47,G295,G78,G411,G410,G175,G304,G445,G420,G264,G347,G449,G109,G66,G324,I295,G453,G148,G147,G187,G162,G229,G58,G401,G108,G442,G408,G205,G541,G320,G509,G307,G354,G197,G424,G260,G358,I218,G413,G416,G159,G407,G278,G274,G330,G287,G319,G228,G127,G301,I371,G138,I327,G166,G352,G366,G185,G448,G113,G431,G67,G50,G279,G265,G372,G76,G382,G340,G95,G412,G511,G451,G384,G163,G186,G124,G282,G44,G140,G381,G110,I502,G538,I352,G263,G177,G125,G98,G391,G404,G117,G258,G402,G421,G336;
//# 14 inputs
//# 14 outputs
//# 18 D-type flipflops
//# 141 inverters
//# 388 gates (118 ANDs + 119 NANDs + 101 ORs + 50 NORs)
//
//
//
  MSFF DFF_0(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G29),.DATA(G502));
  MSFF DFF_1(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G30),.DATA(G503));
  MSFF DFF_2(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G31),.DATA(G504));
  MSFF DFF_3(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G32),.DATA(G505));
  MSFF DFF_4(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G33),.DATA(G506));
  MSFF DFF_5(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G34),.DATA(G507));
  MSFF DFF_6(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G35),.DATA(G508));
  MSFF DFF_7(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G36),.DATA(G509));
  MSFF DFF_8(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G37),.DATA(G510));
  MSFF DFF_9(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G38),.DATA(G511));
  MSFF DFF_10(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G39),.DATA(G512));
  MSFF DFF_11(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G40),.DATA(G513));
  MSFF DFF_12(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G41),.DATA(G514));
  MSFF DFF_13(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G42),.DATA(G515));
  MSFF DFF_14(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G43),.DATA(G516));
  MSFF DFF_15(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G44),.DATA(G517));
  MSFF DFF_16(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G45),.DATA(G518));
  MSFF DFF_17(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G46),.DATA(G519));
//
  NOT NOT1_0(.VSS(VSS),.VDD(VDD),.Y(G520),.A(G0));
  NOT NOT1_1(.VSS(VSS),.VDD(VDD),.Y(G521),.A(G1));
  NOT NOT1_2(.VSS(VSS),.VDD(VDD),.Y(G522),.A(G2));
  NOT NOT1_3(.VSS(VSS),.VDD(VDD),.Y(G524),.A(G3));
  NOT NOT1_4(.VSS(VSS),.VDD(VDD),.Y(I156),.A(G4));
  NOT NOT1_5(.VSS(VSS),.VDD(VDD),.Y(G334),.A(I156));
  NOT NOT1_6(.VSS(VSS),.VDD(VDD),.Y(G527),.A(G4));
  NOT NOT1_7(.VSS(VSS),.VDD(VDD),.Y(G528),.A(G5));
  NOT NOT1_8(.VSS(VSS),.VDD(VDD),.Y(G529),.A(G6));
  NOT NOT1_9(.VSS(VSS),.VDD(VDD),.Y(G531),.A(G7));
  NOT NOT1_10(.VSS(VSS),.VDD(VDD),.Y(G533),.A(G8));
  NOT NOT1_11(.VSS(VSS),.VDD(VDD),.Y(G536),.A(G9));
  NOT NOT1_12(.VSS(VSS),.VDD(VDD),.Y(G538),.A(G10));
  NOT NOT1_13(.VSS(VSS),.VDD(VDD),.Y(G540),.A(G11));
  NOT NOT1_14(.VSS(VSS),.VDD(VDD),.Y(G541),.A(G12));
  NOT NOT1_15(.VSS(VSS),.VDD(VDD),.Y(G543),.A(G13));
  NOT NOT1_16(.VSS(VSS),.VDD(VDD),.Y(G476),.A(G30));
  NOT NOT1_17(.VSS(VSS),.VDD(VDD),.Y(G484),.A(G30));
  NOT NOT1_18(.VSS(VSS),.VDD(VDD),.Y(G125),.A(G40));
  NOT NOT1_19(.VSS(VSS),.VDD(VDD),.Y(G140),.A(G33));
  NOT NOT1_20(.VSS(VSS),.VDD(VDD),.Y(G546),.A(G41));
  NOT NOT1_21(.VSS(VSS),.VDD(VDD),.Y(G132),.A(G42));
  NOT NOT1_22(.VSS(VSS),.VDD(VDD),.Y(G70),.A(G43));
  NOT NOT1_23(.VSS(VSS),.VDD(VDD),.Y(G67),.A(G44));
  NOT NOT1_24(.VSS(VSS),.VDD(VDD),.Y(G99),.A(G29));
  NOT NOT1_25(.VSS(VSS),.VDD(VDD),.Y(G475),.A(G57));
  NOT NOT1_26(.VSS(VSS),.VDD(VDD),.Y(G59),.A(G58));
  NOT NOT1_27(.VSS(VSS),.VDD(VDD),.Y(G228),.A(G524));
  NOT NOT1_28(.VSS(VSS),.VDD(VDD),.Y(G272),.A(G271));
  NOT NOT1_29(.VSS(VSS),.VDD(VDD),.Y(G98),.A(G97));
  NOT NOT1_30(.VSS(VSS),.VDD(VDD),.Y(G135),.A(G134));
  NOT NOT1_31(.VSS(VSS),.VDD(VDD),.Y(I218),.A(G528));
  NOT NOT1_32(.VSS(VSS),.VDD(VDD),.Y(G333),.A(I218));
  NOT NOT1_33(.VSS(VSS),.VDD(VDD),.Y(G55),.A(G54));
  NOT NOT1_34(.VSS(VSS),.VDD(VDD),.Y(G165),.A(G529));
  NOT NOT1_35(.VSS(VSS),.VDD(VDD),.Y(G72),.A(G71));
  NOT NOT1_36(.VSS(VSS),.VDD(VDD),.Y(G236),.A(G274));
  NOT NOT1_37(.VSS(VSS),.VDD(VDD),.Y(G275),.A(G274));
  NOT NOT1_38(.VSS(VSS),.VDD(VDD),.Y(I249),.A(G538));
  NOT NOT1_39(.VSS(VSS),.VDD(VDD),.Y(G370),.A(I249));
  NOT NOT1_40(.VSS(VSS),.VDD(VDD),.Y(G75),.A(G74));
  NOT NOT1_41(.VSS(VSS),.VDD(VDD),.Y(G490),.A(G190));
  NOT NOT1_42(.VSS(VSS),.VDD(VDD),.Y(G482),.A(G241));
  NOT NOT1_43(.VSS(VSS),.VDD(VDD),.Y(G153),.A(G522));
  NOT NOT1_44(.VSS(VSS),.VDD(VDD),.Y(G192),.A(G193));
  NOT NOT1_45(.VSS(VSS),.VDD(VDD),.Y(G123),.A(G122));
  NOT NOT1_46(.VSS(VSS),.VDD(VDD),.Y(I272),.A(G209));
  NOT NOT1_47(.VSS(VSS),.VDD(VDD),.Y(G458),.A(I272));
  NOT NOT1_48(.VSS(VSS),.VDD(VDD),.Y(I276),.A(G238));
  NOT NOT1_49(.VSS(VSS),.VDD(VDD),.Y(G332),.A(I276));
  NOT NOT1_50(.VSS(VSS),.VDD(VDD),.Y(I280),.A(G272));
  NOT NOT1_51(.VSS(VSS),.VDD(VDD),.Y(G309),.A(I280));
  NOT NOT1_52(.VSS(VSS),.VDD(VDD),.Y(I287),.A(G135));
  NOT NOT1_53(.VSS(VSS),.VDD(VDD),.Y(G347),.A(I287));
  NOT NOT1_54(.VSS(VSS),.VDD(VDD),.Y(G498),.A(G195));
  NOT NOT1_55(.VSS(VSS),.VDD(VDD),.Y(G78),.A(G77));
  NOT NOT1_56(.VSS(VSS),.VDD(VDD),.Y(I295),.A(G198));
  NOT NOT1_57(.VSS(VSS),.VDD(VDD),.Y(G459),.A(I295));
  NOT NOT1_58(.VSS(VSS),.VDD(VDD),.Y(G199),.A(G200));
  NOT NOT1_59(.VSS(VSS),.VDD(VDD),.Y(G90),.A(G89));
  NOT NOT1_60(.VSS(VSS),.VDD(VDD),.Y(G221),.A(G222));
  NOT NOT1_61(.VSS(VSS),.VDD(VDD),.Y(G223),.A(G224));
  NOT NOT1_62(.VSS(VSS),.VDD(VDD),.Y(I316),.A(G239));
  NOT NOT1_63(.VSS(VSS),.VDD(VDD),.Y(G369),.A(I316));
  NOT NOT1_64(.VSS(VSS),.VDD(VDD),.Y(G234),.A(G235));
  NOT NOT1_65(.VSS(VSS),.VDD(VDD),.Y(I327),.A(G135));
  NOT NOT1_66(.VSS(VSS),.VDD(VDD),.Y(G435),.A(I327));
  NOT NOT1_67(.VSS(VSS),.VDD(VDD),.Y(I330),.A(G236));
  NOT NOT1_68(.VSS(VSS),.VDD(VDD),.Y(G441),.A(I330));
  NOT NOT1_69(.VSS(VSS),.VDD(VDD),.Y(G50),.A(G49));
  NOT NOT1_70(.VSS(VSS),.VDD(VDD),.Y(G130),.A(G9));
  NOT NOT1_71(.VSS(VSS),.VDD(VDD),.Y(G501),.A(G156));
  NOT NOT1_72(.VSS(VSS),.VDD(VDD),.Y(G477),.A(G276));
  NOT NOT1_73(.VSS(VSS),.VDD(VDD),.Y(G485),.A(G276));
  NOT NOT1_74(.VSS(VSS),.VDD(VDD),.Y(I352),.A(G77));
  NOT NOT1_75(.VSS(VSS),.VDD(VDD),.Y(G299),.A(I352));
  NOT NOT1_76(.VSS(VSS),.VDD(VDD),.Y(G497),.A(G205));
  NOT NOT1_77(.VSS(VSS),.VDD(VDD),.Y(I371),.A(G1));
  NOT NOT1_78(.VSS(VSS),.VDD(VDD),.Y(G335),.A(I371));
  NOT NOT1_79(.VSS(VSS),.VDD(VDD),.Y(I374),.A(G520));
  NOT NOT1_80(.VSS(VSS),.VDD(VDD),.Y(G456),.A(I374));
  NOT NOT1_81(.VSS(VSS),.VDD(VDD),.Y(G87),.A(G86));
  NOT NOT1_82(.VSS(VSS),.VDD(VDD),.Y(I386),.A(G199));
  NOT NOT1_83(.VSS(VSS),.VDD(VDD),.Y(G414),.A(I386));
  NOT NOT1_84(.VSS(VSS),.VDD(VDD),.Y(G486),.A(G68));
  NOT NOT1_85(.VSS(VSS),.VDD(VDD),.Y(G231),.A(G232));
  NOT NOT1_86(.VSS(VSS),.VDD(VDD),.Y(G160),.A(G161));
  NOT NOT1_87(.VSS(VSS),.VDD(VDD),.Y(G265),.A(G50));
  NOT NOT1_88(.VSS(VSS),.VDD(VDD),.Y(G64),.A(G63));
  NOT NOT1_89(.VSS(VSS),.VDD(VDD),.Y(G180),.A(G181));
  NOT NOT1_90(.VSS(VSS),.VDD(VDD),.Y(G107),.A(G456));
  NOT NOT1_91(.VSS(VSS),.VDD(VDD),.Y(G207),.A(G208));
  NOT NOT1_92(.VSS(VSS),.VDD(VDD),.Y(G167),.A(G168));
  NOT NOT1_93(.VSS(VSS),.VDD(VDD),.Y(G124),.A(G206));
  NOT NOT1_94(.VSS(VSS),.VDD(VDD),.Y(G203),.A(G204));
  NOT NOT1_95(.VSS(VSS),.VDD(VDD),.Y(G489),.A(G273));
  NOT NOT1_96(.VSS(VSS),.VDD(VDD),.Y(G495),.A(G273));
  NOT NOT1_97(.VSS(VSS),.VDD(VDD),.Y(G177),.A(G357));
  NOT NOT1_98(.VSS(VSS),.VDD(VDD),.Y(G212),.A(G213));
  NOT NOT1_99(.VSS(VSS),.VDD(VDD),.Y(I493),.A(G218));
  NOT NOT1_100(.VSS(VSS),.VDD(VDD),.Y(G404),.A(I493));
  NOT NOT1_101(.VSS(VSS),.VDD(VDD),.Y(I502),.A(G124));
  NOT NOT1_102(.VSS(VSS),.VDD(VDD),.Y(G468),.A(I502));
  NOT NOT1_103(.VSS(VSS),.VDD(VDD),.Y(G173),.A(G495));
  NOT NOT1_104(.VSS(VSS),.VDD(VDD),.Y(G487),.A(G534));
  NOT NOT1_105(.VSS(VSS),.VDD(VDD),.Y(I529),.A(G468));
  NOT NOT1_106(.VSS(VSS),.VDD(VDD),.Y(G149),.A(I529));
  NOT NOT1_107(.VSS(VSS),.VDD(VDD),.Y(I536),.A(G79));
  NOT NOT1_108(.VSS(VSS),.VDD(VDD),.Y(G446),.A(I536));
  NOT NOT1_109(.VSS(VSS),.VDD(VDD),.Y(G494),.A(G173));
  NOT NOT1_110(.VSS(VSS),.VDD(VDD),.Y(G500),.A(G173));
  NOT NOT1_111(.VSS(VSS),.VDD(VDD),.Y(G214),.A(G215));
  NOT NOT1_112(.VSS(VSS),.VDD(VDD),.Y(G492),.A(G62));
  NOT NOT1_113(.VSS(VSS),.VDD(VDD),.Y(G483),.A(G182));
  NOT NOT1_114(.VSS(VSS),.VDD(VDD),.Y(G282),.A(G281));
  NOT NOT1_115(.VSS(VSS),.VDD(VDD),.Y(I573),.A(G176));
  NOT NOT1_116(.VSS(VSS),.VDD(VDD),.Y(G403),.A(I573));
  NOT NOT1_117(.VSS(VSS),.VDD(VDD),.Y(I576),.A(G175));
  NOT NOT1_118(.VSS(VSS),.VDD(VDD),.Y(G447),.A(I576));
  NOT NOT1_119(.VSS(VSS),.VDD(VDD),.Y(G479),.A(G194));
  NOT NOT1_120(.VSS(VSS),.VDD(VDD),.Y(G491),.A(G194));
  NOT NOT1_121(.VSS(VSS),.VDD(VDD),.Y(G554),.A(G553));
  NOT NOT1_122(.VSS(VSS),.VDD(VDD),.Y(G170),.A(G171));
  NOT NOT1_123(.VSS(VSS),.VDD(VDD),.Y(G172),.A(G171));
  NOT NOT1_124(.VSS(VSS),.VDD(VDD),.Y(G525),.A(G526));
  NOT NOT1_125(.VSS(VSS),.VDD(VDD),.Y(G493),.A(G544));
  NOT NOT1_126(.VSS(VSS),.VDD(VDD),.Y(G545),.A(G544));
  NOT NOT1_127(.VSS(VSS),.VDD(VDD),.Y(G488),.A(G172));
  NOT NOT1_128(.VSS(VSS),.VDD(VDD),.Y(G499),.A(G280));
  NOT NOT1_129(.VSS(VSS),.VDD(VDD),.Y(I624),.A(G120));
  NOT NOT1_130(.VSS(VSS),.VDD(VDD),.Y(G303),.A(I624));
  NOT NOT1_131(.VSS(VSS),.VDD(VDD),.Y(G480),.A(G179));
  NOT NOT1_132(.VSS(VSS),.VDD(VDD),.Y(I631),.A(G188));
  NOT NOT1_133(.VSS(VSS),.VDD(VDD),.Y(G336),.A(I631));
  NOT NOT1_134(.VSS(VSS),.VDD(VDD),.Y(G496),.A(G188));
  NOT NOT1_135(.VSS(VSS),.VDD(VDD),.Y(G174),.A(G496));
  NOT NOT1_136(.VSS(VSS),.VDD(VDD),.Y(I662),.A(G174));
  NOT NOT1_137(.VSS(VSS),.VDD(VDD),.Y(G405),.A(I662));
  NOT NOT1_138(.VSS(VSS),.VDD(VDD),.Y(G478),.A(G279));
  NOT NOT1_139(.VSS(VSS),.VDD(VDD),.Y(I692),.A(G145));
  NOT NOT1_140(.VSS(VSS),.VDD(VDD),.Y(G432),.A(I692));
//
  AND2 AND2_0(.VSS(VSS),.VDD(VDD),.Y(G359),.A(G6),.B(G31));
  AND2 AND2_1(.VSS(VSS),.VDD(VDD),.Y(G469),.A(G163),.B(G3));
  AND2 AND2_2(.VSS(VSS),.VDD(VDD),.Y(G461),.A(G529),.B(G531));
  AND2 AND2_3(.VSS(VSS),.VDD(VDD),.Y(G431),.A(G524),.B(G67));
  AND2 AND2_4(.VSS(VSS),.VDD(VDD),.Y(G362),.A(G129),.B(G77));
  AND2 AND2_5(.VSS(VSS),.VDD(VDD),.Y(G81),.A(G288),.B(G240));
  AND2 AND2_6(.VSS(VSS),.VDD(VDD),.Y(G348),.A(G97),.B(G55));
  AND4 AND4_0(.VSS(VSS),.VDD(VDD),.Y(G352),.A(G8),.B(G135),.C(G37),.D(G164));
  AND2 AND2_7(.VSS(VSS),.VDD(VDD),.Y(G511),.A(G163),.B(G164));
  AND2 AND2_8(.VSS(VSS),.VDD(VDD),.Y(G379),.A(G9),.B(G211));
  AND3 AND3_0(.VSS(VSS),.VDD(VDD),.Y(G385),.A(G529),.B(G7),.C(G49));
  AND2 AND2_9(.VSS(VSS),.VDD(VDD),.Y(G376),.A(G533),.B(G75));
  AND3 AND3_1(.VSS(VSS),.VDD(VDD),.Y(G387),.A(G6),.B(G274),.C(G75));
  AND2 AND2_10(.VSS(VSS),.VDD(VDD),.Y(G462),.A(G192),.B(G538));
  AND2 AND2_11(.VSS(VSS),.VDD(VDD),.Y(G436),.A(G123),.B(G77));
  AND2 AND2_12(.VSS(VSS),.VDD(VDD),.Y(G363),.A(G77),.B(G205));
  AND2 AND2_13(.VSS(VSS),.VDD(VDD),.Y(G410),.A(G1),.B(G205));
  AND2 AND2_14(.VSS(VSS),.VDD(VDD),.Y(G399),.A(G520),.B(G1));
  AND2 AND2_15(.VSS(VSS),.VDD(VDD),.Y(G437),.A(G66),.B(G229));
  AND2 AND2_16(.VSS(VSS),.VDD(VDD),.Y(G307),.A(G6),.B(G104));
  AND2 AND2_17(.VSS(VSS),.VDD(VDD),.Y(G306),.A(G524),.B(G78));
  AND2 AND2_18(.VSS(VSS),.VDD(VDD),.Y(G283),.A(G122),.B(G219));
  AND3 AND3_2(.VSS(VSS),.VDD(VDD),.Y(G339),.A(G533),.B(G199),.C(G209));
  AND3 AND3_3(.VSS(VSS),.VDD(VDD),.Y(G472),.A(G136),.B(G9),.C(G190));
  AND4 AND4_1(.VSS(VSS),.VDD(VDD),.Y(G351),.A(G524),.B(G169),.C(G221),.D(G234));
  AND2 AND2_19(.VSS(VSS),.VDD(VDD),.Y(G440),.A(G38),.B(G234));
  AND3 AND3_4(.VSS(VSS),.VDD(VDD),.Y(G382),.A(G9),.B(G100),.C(G34));
  AND2 AND2_20(.VSS(VSS),.VDD(VDD),.Y(G386),.A(G536),.B(G85));
  AND2 AND2_21(.VSS(VSS),.VDD(VDD),.Y(G321),.A(G90),.B(G50));
  AND2 AND2_22(.VSS(VSS),.VDD(VDD),.Y(G378),.A(G89),.B(G50));
  AND3 AND3_5(.VSS(VSS),.VDD(VDD),.Y(G471),.A(G191),.B(G103),.C(G112));
  AND2 AND2_23(.VSS(VSS),.VDD(VDD),.Y(G377),.A(G90),.B(G56));
  AND2 AND2_24(.VSS(VSS),.VDD(VDD),.Y(G358),.A(G7),.B(G83));
  AND2 AND2_25(.VSS(VSS),.VDD(VDD),.Y(G400),.A(G0),.B(G277));
  AND2 AND2_26(.VSS(VSS),.VDD(VDD),.Y(G308),.A(G5),.B(G151));
  AND2 AND2_27(.VSS(VSS),.VDD(VDD),.Y(G411),.A(G48),.B(G59));
  AND2 AND2_28(.VSS(VSS),.VDD(VDD),.Y(G413),.A(G197),.B(G201));
  AND2 AND2_29(.VSS(VSS),.VDD(VDD),.Y(G434),.A(G165),.B(G231));
  AND2 AND2_30(.VSS(VSS),.VDD(VDD),.Y(G373),.A(G34),.B(G160));
  AND2 AND2_31(.VSS(VSS),.VDD(VDD),.Y(G357),.A(G265),.B(G232));
  AND3 AND3_6(.VSS(VSS),.VDD(VDD),.Y(G444),.A(G64),.B(G78),.C(G211));
  AND2 AND2_32(.VSS(VSS),.VDD(VDD),.Y(G361),.A(G6),.B(G202));
  AND2 AND2_33(.VSS(VSS),.VDD(VDD),.Y(G346),.A(G2),.B(G82));
  AND2 AND2_34(.VSS(VSS),.VDD(VDD),.Y(G457),.A(G4),.B(G107));
  AND2 AND2_35(.VSS(VSS),.VDD(VDD),.Y(G364),.A(G2),.B(G109));
  AND2 AND2_36(.VSS(VSS),.VDD(VDD),.Y(G445),.A(G53),.B(G225));
  AND2 AND2_37(.VSS(VSS),.VDD(VDD),.Y(G412),.A(G3),.B(G207));
  AND3 AND3_7(.VSS(VSS),.VDD(VDD),.Y(G371),.A(G161),.B(G168),.C(G267));
  AND3 AND3_8(.VSS(VSS),.VDD(VDD),.Y(G353),.A(G11),.B(G92),.C(G163));
  AND2 AND2_38(.VSS(VSS),.VDD(VDD),.Y(G388),.A(G11),.B(G114));
  AND2 AND2_39(.VSS(VSS),.VDD(VDD),.Y(G473),.A(G11),.B(G143));
  AND2 AND2_40(.VSS(VSS),.VDD(VDD),.Y(G331),.A(G213),.B(G257));
  AND2 AND2_41(.VSS(VSS),.VDD(VDD),.Y(G429),.A(G51),.B(G225));
  AND2 AND2_42(.VSS(VSS),.VDD(VDD),.Y(G380),.A(G6),.B(G93));
  AND2 AND2_43(.VSS(VSS),.VDD(VDD),.Y(G360),.A(G8),.B(G106));
  AND2 AND2_44(.VSS(VSS),.VDD(VDD),.Y(G338),.A(G202),.B(G203));
  AND2 AND2_45(.VSS(VSS),.VDD(VDD),.Y(G337),.A(G270),.B(G167));
  AND2 AND2_46(.VSS(VSS),.VDD(VDD),.Y(G340),.A(G8),.B(G270));
  AND3 AND3_9(.VSS(VSS),.VDD(VDD),.Y(G322),.A(G522),.B(G105),.C(G196));
  AND2 AND2_47(.VSS(VSS),.VDD(VDD),.Y(G330),.A(G248),.B(G249));
  AND2 AND2_48(.VSS(VSS),.VDD(VDD),.Y(G430),.A(G177),.B(G196));
  AND3 AND3_10(.VSS(VSS),.VDD(VDD),.Y(G344),.A(G111),.B(G189),.C(G195));
  AND2 AND2_49(.VSS(VSS),.VDD(VDD),.Y(G428),.A(G212),.B(G227));
  AND2 AND2_50(.VSS(VSS),.VDD(VDD),.Y(G349),.A(G6),.B(G108));
  AND3 AND3_11(.VSS(VSS),.VDD(VDD),.Y(G460),.A(G2),.B(G81),.C(G115));
  AND2 AND2_51(.VSS(VSS),.VDD(VDD),.Y(G463),.A(G521),.B(G148));
  AND2 AND2_52(.VSS(VSS),.VDD(VDD),.Y(G393),.A(G127),.B(G34));
  AND2 AND2_53(.VSS(VSS),.VDD(VDD),.Y(G470),.A(G528),.B(G149));
  AND2 AND2_54(.VSS(VSS),.VDD(VDD),.Y(G341),.A(G531),.B(G118));
  AND2 AND2_55(.VSS(VSS),.VDD(VDD),.Y(G342),.A(G73),.B(G197));
  AND2 AND2_56(.VSS(VSS),.VDD(VDD),.Y(G324),.A(G522),.B(G183));
  AND2 AND2_57(.VSS(VSS),.VDD(VDD),.Y(G323),.A(G2),.B(G144));
  AND2 AND2_58(.VSS(VSS),.VDD(VDD),.Y(G354),.A(G0),.B(G214));
  AND2 AND2_59(.VSS(VSS),.VDD(VDD),.Y(G312),.A(G180),.B(G182));
  AND2 AND2_60(.VSS(VSS),.VDD(VDD),.Y(G315),.A(G250),.B(G251));
  AND2 AND2_61(.VSS(VSS),.VDD(VDD),.Y(G474),.A(G242),.B(G77));
  AND3 AND3_12(.VSS(VSS),.VDD(VDD),.Y(G343),.A(G2),.B(G528),.C(G147));
  AND2 AND2_62(.VSS(VSS),.VDD(VDD),.Y(G304),.A(G52),.B(G158));
  AND3 AND3_13(.VSS(VSS),.VDD(VDD),.Y(G398),.A(G94),.B(G156),.C(G158));
  AND3 AND3_14(.VSS(VSS),.VDD(VDD),.Y(G365),.A(G282),.B(G137),.C(G156));
  AND3 AND3_15(.VSS(VSS),.VDD(VDD),.Y(G417),.A(G13),.B(G282),.C(G70));
  AND3 AND3_16(.VSS(VSS),.VDD(VDD),.Y(G290),.A(G117),.B(G135),.C(G157));
  AND3 AND3_17(.VSS(VSS),.VDD(VDD),.Y(G327),.A(G4),.B(G39),.C(G157));
  AND2 AND2_63(.VSS(VSS),.VDD(VDD),.Y(G367),.A(G126),.B(G157));
  AND3 AND3_18(.VSS(VSS),.VDD(VDD),.Y(G397),.A(G101),.B(G98),.C(G157));
  AND3 AND3_19(.VSS(VSS),.VDD(VDD),.Y(G451),.A(G541),.B(G554),.C(G187));
  AND2 AND2_64(.VSS(VSS),.VDD(VDD),.Y(G406),.A(G87),.B(G172));
  AND3 AND3_20(.VSS(VSS),.VDD(VDD),.Y(G418),.A(G524),.B(G60),.C(G172));
  AND2 AND2_65(.VSS(VSS),.VDD(VDD),.Y(G453),.A(G545),.B(G186));
  AND3 AND3_21(.VSS(VSS),.VDD(VDD),.Y(G289),.A(G2),.B(G119),.C(G156));
  AND3 AND3_22(.VSS(VSS),.VDD(VDD),.Y(G311),.A(G0),.B(G178),.C(G179));
  AND2 AND2_66(.VSS(VSS),.VDD(VDD),.Y(G402),.A(G154),.B(G183));
  AND2 AND2_67(.VSS(VSS),.VDD(VDD),.Y(G433),.A(G91),.B(G154));
  AND2 AND2_68(.VSS(VSS),.VDD(VDD),.Y(G449),.A(G88),.B(G154));
  AND2 AND2_69(.VSS(VSS),.VDD(VDD),.Y(G452),.A(G526),.B(G184));
  AND2 AND2_70(.VSS(VSS),.VDD(VDD),.Y(G329),.A(G150),.B(G156));
  AND2 AND2_71(.VSS(VSS),.VDD(VDD),.Y(G291),.A(G138),.B(G155));
  AND3 AND3_23(.VSS(VSS),.VDD(VDD),.Y(G328),.A(G5),.B(G102),.C(G155));
  AND2 AND2_72(.VSS(VSS),.VDD(VDD),.Y(G366),.A(G125),.B(G155));
  AND3 AND3_24(.VSS(VSS),.VDD(VDD),.Y(G372),.A(G116),.B(G275),.C(G155));
  AND2 AND2_73(.VSS(VSS),.VDD(VDD),.Y(G383),.A(G131),.B(G155));
  AND2 AND2_74(.VSS(VSS),.VDD(VDD),.Y(G392),.A(G132),.B(G155));
  AND3 AND3_25(.VSS(VSS),.VDD(VDD),.Y(G396),.A(G76),.B(G272),.C(G155));
  AND3 AND3_26(.VSS(VSS),.VDD(VDD),.Y(G401),.A(G2),.B(G110),.C(G155));
  AND3 AND3_27(.VSS(VSS),.VDD(VDD),.Y(G422),.A(G0),.B(G80),.C(G155));
  AND3 AND3_28(.VSS(VSS),.VDD(VDD),.Y(G415),.A(G146),.B(G142),.C(G165));
  AND2 AND2_75(.VSS(VSS),.VDD(VDD),.Y(G425),.A(G146),.B(G176));
  AND3 AND3_29(.VSS(VSS),.VDD(VDD),.Y(G438),.A(G8),.B(G146),.C(G133));
  AND3 AND3_30(.VSS(VSS),.VDD(VDD),.Y(G424),.A(G78),.B(G174),.C(G177));
  AND2 AND2_76(.VSS(VSS),.VDD(VDD),.Y(G439),.A(G174),.B(G175));
  AND2 AND2_77(.VSS(VSS),.VDD(VDD),.Y(G317),.A(G159),.B(G245));
  AND3 AND3_31(.VSS(VSS),.VDD(VDD),.Y(G426),.A(G37),.B(G162),.C(G38));
  AND2 AND2_78(.VSS(VSS),.VDD(VDD),.Y(G443),.A(G47),.B(G162));
  AND2 AND2_79(.VSS(VSS),.VDD(VDD),.Y(G416),.A(G61),.B(G167));
  AND3 AND3_32(.VSS(VSS),.VDD(VDD),.Y(G427),.A(G541),.B(G95),.C(G165));
  AND2 AND2_80(.VSS(VSS),.VDD(VDD),.Y(G442),.A(G541),.B(G121));
  AND2 AND2_81(.VSS(VSS),.VDD(VDD),.Y(G423),.A(G541),.B(G128));
  AND2 AND2_82(.VSS(VSS),.VDD(VDD),.Y(G448),.A(G139),.B(G153));
//
  OR2 OR2_0(.VSS(VSS),.VDD(VDD),.Y(G419),.A(G3),.B(G5));
  OR2 OR2_1(.VSS(VSS),.VDD(VDD),.Y(G193),.A(G6),.B(G30));
  OR2 OR2_2(.VSS(VSS),.VDD(VDD),.Y(G394),.A(G5),.B(G58));
  OR2 OR2_3(.VSS(VSS),.VDD(VDD),.Y(G407),.A(G6),.B(G117));
  OR2 OR2_4(.VSS(VSS),.VDD(VDD),.Y(G314),.A(G527),.B(G57));
  OR2 OR2_5(.VSS(VSS),.VDD(VDD),.Y(G395),.A(G4),.B(G134));
  OR2 OR2_6(.VSS(VSS),.VDD(VDD),.Y(G288),.A(G1),.B(G528));
  OR2 OR2_7(.VSS(VSS),.VDD(VDD),.Y(G302),.A(G4),.B(G529));
  OR2 OR2_8(.VSS(VSS),.VDD(VDD),.Y(G224),.A(G533),.B(G31));
  OR2 OR2_9(.VSS(VSS),.VDD(VDD),.Y(G355),.A(G11),.B(G116));
  OR2 OR2_10(.VSS(VSS),.VDD(VDD),.Y(G316),.A(G531),.B(G536));
  OR2 OR2_11(.VSS(VSS),.VDD(VDD),.Y(G350),.A(G6),.B(G536));
  OR2 OR2_12(.VSS(VSS),.VDD(VDD),.Y(G368),.A(G533),.B(G536));
  OR2 OR2_13(.VSS(VSS),.VDD(VDD),.Y(G381),.A(G7),.B(G71));
  OR2 OR2_14(.VSS(VSS),.VDD(VDD),.Y(G384),.A(G529),.B(G71));
  OR2 OR2_15(.VSS(VSS),.VDD(VDD),.Y(G389),.A(G9),.B(G274));
  OR2 OR2_16(.VSS(VSS),.VDD(VDD),.Y(G374),.A(G536),.B(G538));
  OR2 OR2_17(.VSS(VSS),.VDD(VDD),.Y(G286),.A(G9),.B(G540));
  OR2 OR2_18(.VSS(VSS),.VDD(VDD),.Y(G293),.A(G7),.B(G540));
  OR2 OR2_19(.VSS(VSS),.VDD(VDD),.Y(G375),.A(G10),.B(G540));
  OR2 OR2_20(.VSS(VSS),.VDD(VDD),.Y(G356),.A(G6),.B(G476));
  OR2 OR2_21(.VSS(VSS),.VDD(VDD),.Y(G313),.A(G521),.B(G475));
  OR2 OR2_22(.VSS(VSS),.VDD(VDD),.Y(G420),.A(G522),.B(G59));
  OR3 OR3_0(.VSS(VSS),.VDD(VDD),.Y(G421),.A(G521),.B(G2),.C(G228));
  OR2 OR2_23(.VSS(VSS),.VDD(VDD),.Y(G320),.A(G76),.B(G272));
  OR2 OR2_24(.VSS(VSS),.VDD(VDD),.Y(G310),.A(G522),.B(G135));
  OR2 OR2_25(.VSS(VSS),.VDD(VDD),.Y(G408),.A(G529),.B(G77));
  OR2 OR2_26(.VSS(VSS),.VDD(VDD),.Y(G305),.A(G524),.B(G55));
  OR2 OR2_27(.VSS(VSS),.VDD(VDD),.Y(G409),.A(G528),.B(G55));
  OR2 OR2_28(.VSS(VSS),.VDD(VDD),.Y(G296),.A(G89),.B(G484));
  OR3 OR3_1(.VSS(VSS),.VDD(VDD),.Y(G325),.A(G7),.B(G536),.C(G222));
  OR2 OR2_29(.VSS(VSS),.VDD(VDD),.Y(G464),.A(G72),.B(G536));
  OR2 OR2_30(.VSS(VSS),.VDD(VDD),.Y(G391),.A(G74),.B(G220));
  OR2 OR2_31(.VSS(VSS),.VDD(VDD),.Y(G292),.A(G538),.B(G75));
  OR2 OR2_32(.VSS(VSS),.VDD(VDD),.Y(G345),.A(G529),.B(G226));
  OR2 OR2_33(.VSS(VSS),.VDD(VDD),.Y(G465),.A(G524),.B(G210));
  OR2 OR2_34(.VSS(VSS),.VDD(VDD),.Y(G454),.A(G122),.B(G77));
  OR2 OR2_35(.VSS(VSS),.VDD(VDD),.Y(G269),.A(G362),.B(G529));
  OR2 OR2_36(.VSS(VSS),.VDD(VDD),.Y(G287),.A(G522),.B(G81));
  OR3 OR3_2(.VSS(VSS),.VDD(VDD),.Y(G318),.A(G6),.B(G8),.C(G232));
  OR2 OR2_37(.VSS(VSS),.VDD(VDD),.Y(G326),.A(G533),.B(G232));
  OR2 OR2_38(.VSS(VSS),.VDD(VDD),.Y(G390),.A(G89),.B(G50));
  OR2 OR2_39(.VSS(VSS),.VDD(VDD),.Y(G298),.A(G5),.B(G497));
  OR2 OR2_40(.VSS(VSS),.VDD(VDD),.Y(G300),.A(G87),.B(G97));
  OR2 OR2_41(.VSS(VSS),.VDD(VDD),.Y(G261),.A(G283),.B(G528));
  OR2 OR2_42(.VSS(VSS),.VDD(VDD),.Y(G301),.A(G122),.B(G486));
  OR2 OR2_43(.VSS(VSS),.VDD(VDD),.Y(G92),.A(G351),.B(G352));
  OR2 OR2_44(.VSS(VSS),.VDD(VDD),.Y(G47),.A(G440),.B(G441));
  OR2 OR2_45(.VSS(VSS),.VDD(VDD),.Y(G114),.A(G385),.B(G386));
  OR2 OR2_46(.VSS(VSS),.VDD(VDD),.Y(G297),.A(G64),.B(G274));
  OR3 OR3_3(.VSS(VSS),.VDD(VDD),.Y(G93),.A(G376),.B(G377),.C(G378));
  OR2 OR2_47(.VSS(VSS),.VDD(VDD),.Y(G106),.A(G358),.B(G359));
  OR2 OR2_48(.VSS(VSS),.VDD(VDD),.Y(G110),.A(G399),.B(G400));
  OR2 OR2_49(.VSS(VSS),.VDD(VDD),.Y(G455),.A(G78),.B(G206));
  OR3 OR3_4(.VSS(VSS),.VDD(VDD),.Y(G152),.A(G306),.B(G307),.C(G308));
  OR2 OR2_50(.VSS(VSS),.VDD(VDD),.Y(G60),.A(G413),.B(G414));
  OR2 OR2_51(.VSS(VSS),.VDD(VDD),.Y(G133),.A(G434),.B(G435));
  OR2 OR2_52(.VSS(VSS),.VDD(VDD),.Y(G105),.A(G321),.B(G273));
  OR2 OR2_53(.VSS(VSS),.VDD(VDD),.Y(G108),.A(G346),.B(G347));
  OR3 OR3_5(.VSS(VSS),.VDD(VDD),.Y(G115),.A(G457),.B(G458),.C(G459));
  OR2 OR2_54(.VSS(VSS),.VDD(VDD),.Y(G126),.A(G363),.B(G364));
  OR2 OR2_55(.VSS(VSS),.VDD(VDD),.Y(G79),.A(G444),.B(G445));
  OR2 OR2_56(.VSS(VSS),.VDD(VDD),.Y(G319),.A(G529),.B(G489));
  OR2 OR2_57(.VSS(VSS),.VDD(VDD),.Y(G131),.A(G379),.B(G380));
  OR2 OR2_58(.VSS(VSS),.VDD(VDD),.Y(G118),.A(G337),.B(G338));
  OR2 OR2_59(.VSS(VSS),.VDD(VDD),.Y(G73),.A(G339),.B(G340));
  OR2 OR2_60(.VSS(VSS),.VDD(VDD),.Y(G91),.A(G430),.B(G431));
  OR2 OR2_61(.VSS(VSS),.VDD(VDD),.Y(G137),.A(G348),.B(G349));
  OR2 OR2_62(.VSS(VSS),.VDD(VDD),.Y(G242),.A(G469),.B(G470));
  OR2 OR2_63(.VSS(VSS),.VDD(VDD),.Y(G147),.A(G341),.B(G342));
  OR3 OR3_6(.VSS(VSS),.VDD(VDD),.Y(G284),.A(G528),.B(G272),.C(G281));
  OR3 OR3_7(.VSS(VSS),.VDD(VDD),.Y(G294),.A(G1),.B(G117),.C(G281));
  OR3 OR3_8(.VSS(VSS),.VDD(VDD),.Y(G553),.A(G322),.B(G323),.C(G324));
  OR2 OR2_64(.VSS(VSS),.VDD(VDD),.Y(G141),.A(G353),.B(G354));
  OR2 OR2_65(.VSS(VSS),.VDD(VDD),.Y(G142),.A(G403),.B(G404));
  OR2 OR2_66(.VSS(VSS),.VDD(VDD),.Y(G88),.A(G446),.B(G447));
  OR2 OR2_67(.VSS(VSS),.VDD(VDD),.Y(G544),.A(G343),.B(G344));
  OR2 OR2_68(.VSS(VSS),.VDD(VDD),.Y(G285),.A(G5),.B(G479));
  OR2 OR2_69(.VSS(VSS),.VDD(VDD),.Y(G295),.A(G122),.B(G491));
  OR2 OR2_70(.VSS(VSS),.VDD(VDD),.Y(G450),.A(G12),.B(G171));
  OR2 OR2_71(.VSS(VSS),.VDD(VDD),.Y(G150),.A(G303),.B(G304));
  OR2 OR2_72(.VSS(VSS),.VDD(VDD),.Y(G146),.A(G336),.B(G170));
  OR3 OR3_9(.VSS(VSS),.VDD(VDD),.Y(G539),.A(G451),.B(G452),.C(G453));
  OR2 OR2_73(.VSS(VSS),.VDD(VDD),.Y(G244),.A(G371),.B(G159));
  OR4 OR4_0(.VSS(VSS),.VDD(VDD),.Y(G550),.A(G289),.B(G290),.C(G291),.D(G485));
  OR3 OR3_10(.VSS(VSS),.VDD(VDD),.Y(G551),.A(G327),.B(G328),.C(G329));
  OR3 OR3_11(.VSS(VSS),.VDD(VDD),.Y(G552),.A(G365),.B(G366),.C(G367));
  OR2 OR2_74(.VSS(VSS),.VDD(VDD),.Y(G547),.A(G382),.B(G383));
  OR2 OR2_75(.VSS(VSS),.VDD(VDD),.Y(G548),.A(G392),.B(G393));
  OR4 OR4_1(.VSS(VSS),.VDD(VDD),.Y(G549),.A(G396),.B(G397),.C(G398),.D(G477));
  OR2 OR2_76(.VSS(VSS),.VDD(VDD),.Y(G530),.A(G401),.B(G402));
  OR2 OR2_77(.VSS(VSS),.VDD(VDD),.Y(G61),.A(G405),.B(G406));
  OR2 OR2_78(.VSS(VSS),.VDD(VDD),.Y(G95),.A(G424),.B(G425));
  OR2 OR2_79(.VSS(VSS),.VDD(VDD),.Y(G121),.A(G438),.B(G439));
  OR2 OR2_80(.VSS(VSS),.VDD(VDD),.Y(G279),.A(G317),.B(G166));
  OR4 OR4_2(.VSS(VSS),.VDD(VDD),.Y(G128),.A(G415),.B(G416),.C(G417),.D(G418));
  OR2 OR2_81(.VSS(VSS),.VDD(VDD),.Y(G145),.A(G426),.B(G427));
  OR2 OR2_82(.VSS(VSS),.VDD(VDD),.Y(G139),.A(G442),.B(G443));
  OR2 OR2_83(.VSS(VSS),.VDD(VDD),.Y(G532),.A(G422),.B(G423));
  OR2 OR2_84(.VSS(VSS),.VDD(VDD),.Y(G535),.A(G432),.B(G433));
  OR2 OR2_85(.VSS(VSS),.VDD(VDD),.Y(G537),.A(G448),.B(G449));
//
  NAND2 NAND2_0(.VSS(VSS),.VDD(VDD),.Y(G57),.A(G0),.B(G2));
  NAND2 NAND2_1(.VSS(VSS),.VDD(VDD),.Y(G58),.A(G1),.B(G3));
  NAND2 NAND2_2(.VSS(VSS),.VDD(VDD),.Y(G76),.A(G0),.B(G3));
  NAND2 NAND2_3(.VSS(VSS),.VDD(VDD),.Y(G101),.A(G3),.B(G4));
  NAND2 NAND2_4(.VSS(VSS),.VDD(VDD),.Y(G117),.A(G2),.B(G4));
  NAND2 NAND2_5(.VSS(VSS),.VDD(VDD),.Y(G271),.A(G1),.B(G4));
  NAND2 NAND2_6(.VSS(VSS),.VDD(VDD),.Y(G97),.A(G2),.B(G5));
  NAND2 NAND2_7(.VSS(VSS),.VDD(VDD),.Y(G134),.A(G3),.B(G5));
  NAND2 NAND2_8(.VSS(VSS),.VDD(VDD),.Y(G54),.A(G4),.B(G6));
  NAND2 NAND2_9(.VSS(VSS),.VDD(VDD),.Y(G116),.A(G6),.B(G9));
  NAND2 NAND2_10(.VSS(VSS),.VDD(VDD),.Y(G71),.A(G8),.B(G10));
  NAND2 NAND2_11(.VSS(VSS),.VDD(VDD),.Y(G274),.A(G7),.B(G10));
  NAND2 NAND2_12(.VSS(VSS),.VDD(VDD),.Y(G74),.A(G9),.B(G11));
  NAND2 NAND2_13(.VSS(VSS),.VDD(VDD),.Y(G112),.A(G8),.B(G31));
  NAND2 NAND2_14(.VSS(VSS),.VDD(VDD),.Y(G245),.A(G8),.B(G34));
  NAND2 NAND2_15(.VSS(VSS),.VDD(VDD),.Y(G122),.A(G522),.B(G3));
  NAND2 NAND2_16(.VSS(VSS),.VDD(VDD),.Y(G238),.A(G2),.B(G524));
  NAND2 NAND2_17(.VSS(VSS),.VDD(VDD),.Y(G129),.A(G527),.B(G5));
  NAND2 NAND2_18(.VSS(VSS),.VDD(VDD),.Y(G240),.A(G4),.B(G134));
  NAND4 NAND4_0(.VSS(VSS),.VDD(VDD),.Y(G252),.A(G3),.B(G11),.C(G35),.D(G216));
  NAND2 NAND2_19(.VSS(VSS),.VDD(VDD),.Y(G77),.A(G4),.B(G528));
  NAND3 NAND3_0(.VSS(VSS),.VDD(VDD),.Y(G103),.A(G529),.B(G7),.C(G30));
  NAND2 NAND2_20(.VSS(VSS),.VDD(VDD),.Y(G200),.A(G527),.B(G529));
  NAND2 NAND2_21(.VSS(VSS),.VDD(VDD),.Y(G248),.A(G529),.B(G36));
  NAND2 NAND2_22(.VSS(VSS),.VDD(VDD),.Y(G89),.A(G531),.B(G8));
  NAND2 NAND2_23(.VSS(VSS),.VDD(VDD),.Y(G222),.A(G533),.B(G10));
  NAND2 NAND2_24(.VSS(VSS),.VDD(VDD),.Y(G239),.A(G7),.B(G533));
  NAND2 NAND2_25(.VSS(VSS),.VDD(VDD),.Y(G235),.A(G6),.B(G536));
  NAND2 NAND2_26(.VSS(VSS),.VDD(VDD),.Y(G220),.A(G7),.B(G71));
  NAND2 NAND2_27(.VSS(VSS),.VDD(VDD),.Y(G49),.A(G9),.B(G538));
  NAND2 NAND2_28(.VSS(VSS),.VDD(VDD),.Y(G251),.A(G543),.B(G32));
  NAND3 NAND3_1(.VSS(VSS),.VDD(VDD),.Y(G276),.A(G3),.B(G543),.C(G140));
  NAND2 NAND2_29(.VSS(VSS),.VDD(VDD),.Y(G263),.A(G0),.B(G99));
  NAND2 NAND2_30(.VSS(VSS),.VDD(VDD),.Y(G226),.A(G527),.B(G59));
  NAND2 NAND2_31(.VSS(VSS),.VDD(VDD),.Y(G210),.A(G520),.B(G272));
  NAND2 NAND2_32(.VSS(VSS),.VDD(VDD),.Y(G66),.A(G129),.B(G101));
  NAND2 NAND2_33(.VSS(VSS),.VDD(VDD),.Y(G233),.A(G522),.B(G135));
  NAND3 NAND3_2(.VSS(VSS),.VDD(VDD),.Y(G104),.A(G122),.B(G238),.C(G240));
  NAND2 NAND2_34(.VSS(VSS),.VDD(VDD),.Y(G86),.A(G55),.B(G3));
  NAND2 NAND2_35(.VSS(VSS),.VDD(VDD),.Y(G219),.A(G524),.B(G55));
  NAND2 NAND2_36(.VSS(VSS),.VDD(VDD),.Y(G68),.A(G302),.B(G528));
  NAND2 NAND2_37(.VSS(VSS),.VDD(VDD),.Y(G232),.A(G536),.B(G164));
  NAND2 NAND2_38(.VSS(VSS),.VDD(VDD),.Y(G136),.A(G222),.B(G224));
  NAND2 NAND2_39(.VSS(VSS),.VDD(VDD),.Y(G510),.A(G350),.B(G235));
  NAND2 NAND2_40(.VSS(VSS),.VDD(VDD),.Y(G161),.A(G316),.B(G72));
  NAND2 NAND2_41(.VSS(VSS),.VDD(VDD),.Y(G100),.A(G381),.B(G220));
  NAND2 NAND2_42(.VSS(VSS),.VDD(VDD),.Y(G85),.A(G384),.B(G239));
  NAND3 NAND3_3(.VSS(VSS),.VDD(VDD),.Y(G243),.A(G368),.B(G275),.C(G34));
  NAND2 NAND2_43(.VSS(VSS),.VDD(VDD),.Y(G63),.A(G75),.B(G8));
  NAND3 NAND3_4(.VSS(VSS),.VDD(VDD),.Y(G237),.A(G10),.B(G75),.C(G201));
  NAND2 NAND2_44(.VSS(VSS),.VDD(VDD),.Y(G503),.A(G286),.B(G538));
  NAND2 NAND2_45(.VSS(VSS),.VDD(VDD),.Y(G56),.A(G374),.B(G375));
  NAND2 NAND2_46(.VSS(VSS),.VDD(VDD),.Y(G83),.A(G355),.B(G356));
  NAND2 NAND2_47(.VSS(VSS),.VDD(VDD),.Y(G96),.A(G313),.B(G314));
  NAND2 NAND2_48(.VSS(VSS),.VDD(VDD),.Y(G278),.A(G332),.B(G333));
  NAND3 NAND3_5(.VSS(VSS),.VDD(VDD),.Y(G255),.A(G309),.B(G2),.C(G529));
  NAND3 NAND3_6(.VSS(VSS),.VDD(VDD),.Y(G69),.A(G419),.B(G420),.C(G233));
  NAND2 NAND2_49(.VSS(VSS),.VDD(VDD),.Y(G512),.A(G310),.B(G233));
  NAND2 NAND2_50(.VSS(VSS),.VDD(VDD),.Y(G181),.A(G2),.B(G78));
  NAND3 NAND3_7(.VSS(VSS),.VDD(VDD),.Y(G277),.A(G394),.B(G395),.C(G81));
  NAND2 NAND2_51(.VSS(VSS),.VDD(VDD),.Y(G151),.A(G305),.B(G200));
  NAND3 NAND3_8(.VSS(VSS),.VDD(VDD),.Y(G48),.A(G407),.B(G408),.C(G409));
  NAND2 NAND2_52(.VSS(VSS),.VDD(VDD),.Y(G264),.A(G227),.B(G241));
  NAND2 NAND2_53(.VSS(VSS),.VDD(VDD),.Y(G208),.A(G68),.B(G229));
  NAND2 NAND2_54(.VSS(VSS),.VDD(VDD),.Y(G168),.A(G75),.B(G221));
  NAND2 NAND2_55(.VSS(VSS),.VDD(VDD),.Y(G84),.A(G369),.B(G370));
  NAND3 NAND3_9(.VSS(VSS),.VDD(VDD),.Y(G258),.A(G464),.B(G103),.C(G223));
  NAND2 NAND2_56(.VSS(VSS),.VDD(VDD),.Y(G166),.A(G7),.B(G50));
  NAND2 NAND2_57(.VSS(VSS),.VDD(VDD),.Y(G259),.A(G130),.B(G225));
  NAND2 NAND2_58(.VSS(VSS),.VDD(VDD),.Y(G504),.A(G292),.B(G293));
  NAND2 NAND2_59(.VSS(VSS),.VDD(VDD),.Y(G217),.A(G50),.B(G230));
  NAND2 NAND2_60(.VSS(VSS),.VDD(VDD),.Y(G257),.A(G538),.B(G230));
  NAND3 NAND3_10(.VSS(VSS),.VDD(VDD),.Y(G260),.A(G528),.B(G529),.C(G191));
  NAND2 NAND2_61(.VSS(VSS),.VDD(VDD),.Y(G266),.A(G524),.B(G96));
  NAND2 NAND2_62(.VSS(VSS),.VDD(VDD),.Y(G262),.A(G527),.B(G278));
  NAND2 NAND2_63(.VSS(VSS),.VDD(VDD),.Y(G138),.A(G465),.B(G263));
  NAND2 NAND2_64(.VSS(VSS),.VDD(VDD),.Y(G256),.A(G4),.B(G69));
  NAND2 NAND2_65(.VSS(VSS),.VDD(VDD),.Y(G82),.A(G334),.B(G335));
  NAND2 NAND2_66(.VSS(VSS),.VDD(VDD),.Y(G109),.A(G269),.B(G219));
  NAND2 NAND2_67(.VSS(VSS),.VDD(VDD),.Y(G206),.A(G287),.B(G524));
  NAND2 NAND2_68(.VSS(VSS),.VDD(VDD),.Y(G204),.A(G521),.B(G87));
  NAND2 NAND2_69(.VSS(VSS),.VDD(VDD),.Y(G53),.A(G264),.B(G237));
  NAND2 NAND2_70(.VSS(VSS),.VDD(VDD),.Y(G273),.A(G325),.B(G326));
  NAND2 NAND2_71(.VSS(VSS),.VDD(VDD),.Y(G267),.A(G536),.B(G84));
  NAND2 NAND2_72(.VSS(VSS),.VDD(VDD),.Y(G113),.A(G389),.B(G390));
  NAND3 NAND3_11(.VSS(VSS),.VDD(VDD),.Y(G143),.A(G258),.B(G193),.C(G259));
  NAND2 NAND2_73(.VSS(VSS),.VDD(VDD),.Y(G213),.A(G64),.B(G275));
  NAND2 NAND2_74(.VSS(VSS),.VDD(VDD),.Y(G51),.A(G260),.B(G237));
  NAND3 NAND3_12(.VSS(VSS),.VDD(VDD),.Y(G102),.A(G320),.B(G266),.C(G210));
  NAND3 NAND3_13(.VSS(VSS),.VDD(VDD),.Y(G52),.A(G298),.B(G299),.C(G219));
  NAND3 NAND3_14(.VSS(VSS),.VDD(VDD),.Y(G80),.A(G421),.B(G226),.C(G256));
  NAND2 NAND2_75(.VSS(VSS),.VDD(VDD),.Y(G270),.A(G345),.B(G204));
  NAND3 NAND3_15(.VSS(VSS),.VDD(VDD),.Y(G94),.A(G261),.B(G181),.C(G262));
  NAND3 NAND3_16(.VSS(VSS),.VDD(VDD),.Y(G505),.A(G300),.B(G301),.C(G181));
  NAND3 NAND3_17(.VSS(VSS),.VDD(VDD),.Y(G249),.A(G11),.B(G273),.C(G201));
  NAND2 NAND2_76(.VSS(VSS),.VDD(VDD),.Y(G268),.A(G11),.B(G113));
  NAND2 NAND2_77(.VSS(VSS),.VDD(VDD),.Y(G111),.A(G213),.B(G217));
  NAND3 NAND3_18(.VSS(VSS),.VDD(VDD),.Y(G534),.A(G296),.B(G297),.C(G166));
  NAND2 NAND2_78(.VSS(VSS),.VDD(VDD),.Y(G253),.A(G87),.B(G218));
  NAND3 NAND3_19(.VSS(VSS),.VDD(VDD),.Y(G148),.A(G454),.B(G455),.C(G0));
  NAND2 NAND2_79(.VSS(VSS),.VDD(VDD),.Y(G254),.A(G1),.B(G152));
  NAND2 NAND2_80(.VSS(VSS),.VDD(VDD),.Y(G127),.A(G391),.B(G268));
  NAND3 NAND3_20(.VSS(VSS),.VDD(VDD),.Y(G215),.A(G135),.B(G55),.C(G212));
  NAND2 NAND2_81(.VSS(VSS),.VDD(VDD),.Y(G62),.A(G534),.B(G32));
  NAND3 NAND3_21(.VSS(VSS),.VDD(VDD),.Y(G523),.A(G254),.B(G255),.C(G208));
  NAND2 NAND2_82(.VSS(VSS),.VDD(VDD),.Y(G508),.A(G318),.B(G319));
  NAND3 NAND3_22(.VSS(VSS),.VDD(VDD),.Y(G144),.A(G215),.B(G252),.C(G253));
  NAND2 NAND2_83(.VSS(VSS),.VDD(VDD),.Y(G250),.A(G13),.B(G523));
  NAND2 NAND2_84(.VSS(VSS),.VDD(VDD),.Y(G281),.A(G523),.B(G534));
  NAND2 NAND2_85(.VSS(VSS),.VDD(VDD),.Y(G171),.A(G553),.B(G187));
  NAND3 NAND3_23(.VSS(VSS),.VDD(VDD),.Y(G526),.A(G1),.B(G2),.C(G141));
  NAND2 NAND2_86(.VSS(VSS),.VDD(VDD),.Y(G280),.A(G46),.B(G247));
  NAND2 NAND2_87(.VSS(VSS),.VDD(VDD),.Y(G246),.A(G544),.B(G186));
  NAND2 NAND2_88(.VSS(VSS),.VDD(VDD),.Y(G119),.A(G284),.B(G285));
  NAND2 NAND2_89(.VSS(VSS),.VDD(VDD),.Y(G120),.A(G294),.B(G295));
  NAND2 NAND2_90(.VSS(VSS),.VDD(VDD),.Y(G185),.A(G525),.B(G184));
  NAND2 NAND2_91(.VSS(VSS),.VDD(VDD),.Y(G159),.A(G6),.B(G155));
  NAND3 NAND3_24(.VSS(VSS),.VDD(VDD),.Y(G518),.A(G450),.B(G185),.C(G246));
  NAND3 NAND3_25(.VSS(VSS),.VDD(VDD),.Y(G542),.A(G243),.B(G244),.C(G279));
//
  NOR2 NOR2_0(.VSS(VSS),.VDD(VDD),.Y(G163),.A(G0),.B(G4));
  NOR2 NOR2_1(.VSS(VSS),.VDD(VDD),.Y(G216),.A(G4),.B(G5));
  NOR2 NOR2_2(.VSS(VSS),.VDD(VDD),.Y(G169),.A(G5),.B(G7));
  NOR2 NOR2_3(.VSS(VSS),.VDD(VDD),.Y(G225),.A(G7),.B(G8));
  NOR2 NOR2_4(.VSS(VSS),.VDD(VDD),.Y(G190),.A(G7),.B(G11));
  NOR2 NOR2_5(.VSS(VSS),.VDD(VDD),.Y(G241),.A(G10),.B(G11));
  NOR2 NOR2_6(.VSS(VSS),.VDD(VDD),.Y(G198),.A(G520),.B(G3));
  NOR2 NOR2_7(.VSS(VSS),.VDD(VDD),.Y(G178),.A(G521),.B(G4));
  NOR2 NOR2_8(.VSS(VSS),.VDD(VDD),.Y(G229),.A(G1),.B(G522));
  NOR2 NOR2_9(.VSS(VSS),.VDD(VDD),.Y(G209),.A(G1),.B(G524));
  NOR2 NOR2_10(.VSS(VSS),.VDD(VDD),.Y(G195),.A(G521),.B(G134));
  NOR2 NOR2_11(.VSS(VSS),.VDD(VDD),.Y(G189),.A(G522),.B(G54));
  NOR2 NOR2_12(.VSS(VSS),.VDD(VDD),.Y(G201),.A(G528),.B(G54));
  NOR2 NOR2_13(.VSS(VSS),.VDD(VDD),.Y(G164),.A(G531),.B(G10));
  NOR2 NOR2_14(.VSS(VSS),.VDD(VDD),.Y(G211),.A(G6),.B(G274));
  NOR2 NOR2_15(.VSS(VSS),.VDD(VDD),.Y(G156),.A(G12),.B(G543));
  NOR2 NOR2_16(.VSS(VSS),.VDD(VDD),.Y(G205),.A(G529),.B(G122));
  NOR2 NOR2_17(.VSS(VSS),.VDD(VDD),.Y(G227),.A(G5),.B(G200));
  NOR2 NOR2_18(.VSS(VSS),.VDD(VDD),.Y(G230),.A(G8),.B(G490));
  NOR2 NOR2_19(.VSS(VSS),.VDD(VDD),.Y(G191),.A(G9),.B(G482));
  NOR3 NOR3_0(.VSS(VSS),.VDD(VDD),.Y(G196),.A(G5),.B(G540),.C(G86));
  NOR2 NOR2_20(.VSS(VSS),.VDD(VDD),.Y(G197),.A(G540),.B(G232));
  NOR2 NOR2_21(.VSS(VSS),.VDD(VDD),.Y(G202),.A(G10),.B(G63));
  NOR2 NOR2_22(.VSS(VSS),.VDD(VDD),.Y(G502),.A(G436),.B(G437));
  NOR2 NOR2_23(.VSS(VSS),.VDD(VDD),.Y(G218),.A(G528),.B(G217));
  NOR3 NOR3_1(.VSS(VSS),.VDD(VDD),.Y(G516),.A(G410),.B(G411),.C(G412));
  NOR2 NOR2_24(.VSS(VSS),.VDD(VDD),.Y(G515),.A(G387),.B(G388));
  NOR2 NOR2_25(.VSS(VSS),.VDD(VDD),.Y(G509),.A(G331),.B(G5));
  NOR2 NOR2_26(.VSS(VSS),.VDD(VDD),.Y(G513),.A(G360),.B(G361));
  NOR2 NOR2_27(.VSS(VSS),.VDD(VDD),.Y(G183),.A(G330),.B(G3));
  NOR2 NOR2_28(.VSS(VSS),.VDD(VDD),.Y(G517),.A(G428),.B(G429));
  NOR2 NOR2_29(.VSS(VSS),.VDD(VDD),.Y(G182),.A(G12),.B(G62));
  NOR4 NOR4_0(.VSS(VSS),.VDD(VDD),.Y(G519),.A(G460),.B(G461),.C(G462),.D(G463));
  NOR2 NOR2_30(.VSS(VSS),.VDD(VDD),.Y(G176),.A(G4),.B(G494));
  NOR2 NOR2_31(.VSS(VSS),.VDD(VDD),.Y(G175),.A(G86),.B(G500));
  NOR2 NOR2_32(.VSS(VSS),.VDD(VDD),.Y(G187),.A(G13),.B(G492));
  NOR2 NOR2_33(.VSS(VSS),.VDD(VDD),.Y(G158),.A(G521),.B(G281));
  NOR2 NOR2_34(.VSS(VSS),.VDD(VDD),.Y(G194),.A(G281),.B(G271));
  NOR2 NOR2_35(.VSS(VSS),.VDD(VDD),.Y(G157),.A(G13),.B(G483));
  NOR3 NOR3_2(.VSS(VSS),.VDD(VDD),.Y(G507),.A(G315),.B(G12),.C(G487));
  NOR2 NOR2_36(.VSS(VSS),.VDD(VDD),.Y(G186),.A(G282),.B(G501));
  NOR4 NOR4_1(.VSS(VSS),.VDD(VDD),.Y(G247),.A(G471),.B(G472),.C(G473),.D(G474));
  NOR2 NOR2_37(.VSS(VSS),.VDD(VDD),.Y(G179),.A(G541),.B(G280));
  NOR2 NOR2_38(.VSS(VSS),.VDD(VDD),.Y(G188),.A(G543),.B(G493));
  NOR2 NOR2_39(.VSS(VSS),.VDD(VDD),.Y(G154),.A(G12),.B(G488));
  NOR3 NOR3_3(.VSS(VSS),.VDD(VDD),.Y(G184),.A(G541),.B(G13),.C(G499));
  NOR2 NOR2_40(.VSS(VSS),.VDD(VDD),.Y(G506),.A(G311),.B(G312));
  NOR2 NOR2_41(.VSS(VSS),.VDD(VDD),.Y(G155),.A(G13),.B(G480));
  NOR2 NOR2_42(.VSS(VSS),.VDD(VDD),.Y(G162),.A(G185),.B(G498));
  NOR3 NOR3_4(.VSS(VSS),.VDD(VDD),.Y(G514),.A(G372),.B(G373),.C(G478));

endmodule