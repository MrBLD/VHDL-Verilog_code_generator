module s526w(G2,G148,G147,VDD,G0,G198,G213,CLOCK,G214,G199,G1,VSS);
input G2,VDD,G0,CLOCK,G1,VSS;
output G148,G147,G198,G213,G214,G199;

  wire G125,G146,G144,G195,G23,G113,G67,G31,G111,G183,G201,G39,G36,G17,G208,G171,G72,G155,G121,G211,G73,G139,G33,G70,G212,G128,G127,G196,G22,G37,G48,I288,G194,G180,G76,G40,G74,G119,G207,G130,G53,G82,G43,G182,G30,G138,G169,G206,G12,G20,G96,I359,G178,I285,G59,G116,G19,G97,G174,G65,G42,G88,G205,G164,G188,G54,G159,G145,G133,G38,G63,G149,G18,G102,G34,G115,G176,G80,G172,G78,G11,G179,G143,G24,G175,G204,G105,G190,G58,G47,G120,G151,G85,G136,G135,G92,G185,G71,G87,G93,G55,G165,G14,G142,G131,G161,G50,G177,G103,G61,G21,G25,G62,G173,G160,G122,G90,G106,G189,G32,G15,G163,G81,G27,G132,G191,G86,G79,G129,G35,G52,G210,G83,G193,G68,G60,G91,G154,G57,G158,G181,G101,G150,G16,G41,G202,G94,G134,I362,G186,G187,G166,G56,G29,G51,G140,G200,G66,G46,G89,G184,I343,G98,G13,G95,G137,I368,G104,G110,G100,G49,G26,G114,G45,G162,G167,I351,G209,G69,G99,G64,G203,G156,G28,G118,G157,G44,G10,G168,G141,G152,G126,G117,G124,G109,G84,G197,G112,G192,G123,G108,I365,I340,G153,G75,G107,G77,G170;
//# 3 inputs
//# 6 outputs
//# 21 D-type flipflops
//# 52 inverters
//# 141 gates (56 ANDs + 22 NANDs + 28 ORs + 35 NORs)
//
//
//
  MSFF DFF_0(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G10),.DATA(G60));
  MSFF DFF_1(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G11),.DATA(G61));
  MSFF DFF_2(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G12),.DATA(G62));
  MSFF DFF_3(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G13),.DATA(G69));
  MSFF DFF_4(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G14),.DATA(G79));
  MSFF DFF_5(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G15),.DATA(G84));
  MSFF DFF_6(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G16),.DATA(G89));
  MSFF DFF_7(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G17),.DATA(G96));
  MSFF DFF_8(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G18),.DATA(G101));
  MSFF DFF_9(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G19),.DATA(G106));
  MSFF DFF_10(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G20),.DATA(G115));
  MSFF DFF_11(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G21),.DATA(G127));
  MSFF DFF_12(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G22),.DATA(G137));
  MSFF DFF_13(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G23),.DATA(G167));
  MSFF DFF_14(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G24),.DATA(G173));
  MSFF DFF_15(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G25),.DATA(G179));
  MSFF DFF_16(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G26),.DATA(G183));
  MSFF DFF_17(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G27),.DATA(G188));
  MSFF DFF_18(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G28),.DATA(G194));
  MSFF DFF_19(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G29),.DATA(G200));
  MSFF DFF_20(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G30),.DATA(G206));
//
  NOT NOT1_0(.VSS(VSS),.VDD(VDD),.Y(G59),.A(G211));
  NOT NOT1_1(.VSS(VSS),.VDD(VDD),.Y(G65),.A(G12));
  NOT NOT1_2(.VSS(VSS),.VDD(VDD),.Y(G72),.A(G13));
  NOT NOT1_3(.VSS(VSS),.VDD(VDD),.Y(G83),.A(G10));
  NOT NOT1_4(.VSS(VSS),.VDD(VDD),.Y(G85),.A(G15));
  NOT NOT1_5(.VSS(VSS),.VDD(VDD),.Y(G90),.A(G14));
  NOT NOT1_6(.VSS(VSS),.VDD(VDD),.Y(G94),.A(G16));
  NOT NOT1_7(.VSS(VSS),.VDD(VDD),.Y(G104),.A(G18));
  NOT NOT1_8(.VSS(VSS),.VDD(VDD),.Y(G107),.A(G11));
  NOT NOT1_9(.VSS(VSS),.VDD(VDD),.Y(G112),.A(G19));
  NOT NOT1_10(.VSS(VSS),.VDD(VDD),.Y(G116),.A(G17));
  NOT NOT1_11(.VSS(VSS),.VDD(VDD),.Y(G122),.A(G30));
  NOT NOT1_12(.VSS(VSS),.VDD(VDD),.Y(G124),.A(G20));
  NOT NOT1_13(.VSS(VSS),.VDD(VDD),.Y(G126),.A(G59));
  NOT NOT1_14(.VSS(VSS),.VDD(VDD),.Y(G131),.A(G21));
  NOT NOT1_15(.VSS(VSS),.VDD(VDD),.Y(G135),.A(G20));
  NOT NOT1_16(.VSS(VSS),.VDD(VDD),.Y(G136),.A(G12));
  NOT NOT1_17(.VSS(VSS),.VDD(VDD),.Y(G140),.A(G21));
  NOT NOT1_18(.VSS(VSS),.VDD(VDD),.Y(G141),.A(G29));
  NOT NOT1_19(.VSS(VSS),.VDD(VDD),.Y(G145),.A(G22));
  NOT NOT1_20(.VSS(VSS),.VDD(VDD),.Y(I285),.A(G23));
  NOT NOT1_21(.VSS(VSS),.VDD(VDD),.Y(G147),.A(I285));
  NOT NOT1_22(.VSS(VSS),.VDD(VDD),.Y(I288),.A(G24));
  NOT NOT1_23(.VSS(VSS),.VDD(VDD),.Y(G148),.A(I288));
  NOT NOT1_24(.VSS(VSS),.VDD(VDD),.Y(G157),.A(G18));
  NOT NOT1_25(.VSS(VSS),.VDD(VDD),.Y(G163),.A(G20));
  NOT NOT1_26(.VSS(VSS),.VDD(VDD),.Y(G168),.A(G23));
  NOT NOT1_27(.VSS(VSS),.VDD(VDD),.Y(G172),.A(G21));
  NOT NOT1_28(.VSS(VSS),.VDD(VDD),.Y(G174),.A(G24));
  NOT NOT1_29(.VSS(VSS),.VDD(VDD),.Y(G177),.A(G13));
  NOT NOT1_30(.VSS(VSS),.VDD(VDD),.Y(G180),.A(G25));
  NOT NOT1_31(.VSS(VSS),.VDD(VDD),.Y(G184),.A(G12));
  NOT NOT1_32(.VSS(VSS),.VDD(VDD),.Y(G189),.A(G193));
  NOT NOT1_33(.VSS(VSS),.VDD(VDD),.Y(G195),.A(G28));
  NOT NOT1_34(.VSS(VSS),.VDD(VDD),.Y(I340),.A(G25));
  NOT NOT1_35(.VSS(VSS),.VDD(VDD),.Y(G198),.A(I340));
  NOT NOT1_36(.VSS(VSS),.VDD(VDD),.Y(I343),.A(G26));
  NOT NOT1_37(.VSS(VSS),.VDD(VDD),.Y(G199),.A(I343));
  NOT NOT1_38(.VSS(VSS),.VDD(VDD),.Y(G201),.A(G205));
  NOT NOT1_39(.VSS(VSS),.VDD(VDD),.Y(G202),.A(G29));
  NOT NOT1_40(.VSS(VSS),.VDD(VDD),.Y(I351),.A(G2));
  NOT NOT1_41(.VSS(VSS),.VDD(VDD),.Y(G205),.A(I351));
  NOT NOT1_42(.VSS(VSS),.VDD(VDD),.Y(G207),.A(G212));
  NOT NOT1_43(.VSS(VSS),.VDD(VDD),.Y(G208),.A(G30));
  NOT NOT1_44(.VSS(VSS),.VDD(VDD),.Y(I359),.A(G0));
  NOT NOT1_45(.VSS(VSS),.VDD(VDD),.Y(G211),.A(I359));
  NOT NOT1_46(.VSS(VSS),.VDD(VDD),.Y(I362),.A(G1));
  NOT NOT1_47(.VSS(VSS),.VDD(VDD),.Y(G212),.A(I362));
  NOT NOT1_48(.VSS(VSS),.VDD(VDD),.Y(I365),.A(G27));
  NOT NOT1_49(.VSS(VSS),.VDD(VDD),.Y(G213),.A(I365));
  NOT NOT1_50(.VSS(VSS),.VDD(VDD),.Y(I368),.A(G28));
  NOT NOT1_51(.VSS(VSS),.VDD(VDD),.Y(G214),.A(I368));
//
  AND2 AND2_0(.VSS(VSS),.VDD(VDD),.Y(G34),.A(G122),.B(G123));
  AND4 AND4_0(.VSS(VSS),.VDD(VDD),.Y(G35),.A(G10),.B(G107),.C(G90),.D(G15));
  AND2 AND2_1(.VSS(VSS),.VDD(VDD),.Y(G36),.A(G122),.B(G123));
  AND2 AND2_2(.VSS(VSS),.VDD(VDD),.Y(G38),.A(G122),.B(G123));
  AND2 AND2_3(.VSS(VSS),.VDD(VDD),.Y(G39),.A(G65),.B(G21));
  AND2 AND2_4(.VSS(VSS),.VDD(VDD),.Y(G40),.A(G12),.B(G131));
  AND2 AND2_5(.VSS(VSS),.VDD(VDD),.Y(G44),.A(G59),.B(G94));
  AND2 AND2_6(.VSS(VSS),.VDD(VDD),.Y(G45),.A(G122),.B(G59));
  AND2 AND2_7(.VSS(VSS),.VDD(VDD),.Y(G46),.A(G116),.B(G112));
  AND2 AND2_8(.VSS(VSS),.VDD(VDD),.Y(G47),.A(G116),.B(G18));
  AND3 AND3_0(.VSS(VSS),.VDD(VDD),.Y(G51),.A(G59),.B(G16),.C(G17));
  AND2 AND2_9(.VSS(VSS),.VDD(VDD),.Y(G52),.A(G59),.B(G18));
  AND2 AND2_10(.VSS(VSS),.VDD(VDD),.Y(G54),.A(G17),.B(G104));
  AND2 AND2_11(.VSS(VSS),.VDD(VDD),.Y(G55),.A(G116),.B(G18));
  AND2 AND2_12(.VSS(VSS),.VDD(VDD),.Y(G56),.A(G17),.B(G112));
  AND4 AND4_1(.VSS(VSS),.VDD(VDD),.Y(G57),.A(G59),.B(G16),.C(G17),.D(G18));
  AND2 AND2_13(.VSS(VSS),.VDD(VDD),.Y(G58),.A(G59),.B(G19));
  AND3 AND3_1(.VSS(VSS),.VDD(VDD),.Y(G76),.A(G10),.B(G90),.C(G15));
  AND2 AND2_14(.VSS(VSS),.VDD(VDD),.Y(G77),.A(G10),.B(G11));
  AND2 AND2_15(.VSS(VSS),.VDD(VDD),.Y(G78),.A(G83),.B(G107));
  AND3 AND3_2(.VSS(VSS),.VDD(VDD),.Y(G80),.A(G10),.B(G11),.C(G14));
  AND2 AND2_16(.VSS(VSS),.VDD(VDD),.Y(G81),.A(G83),.B(G90));
  AND2 AND2_17(.VSS(VSS),.VDD(VDD),.Y(G82),.A(G107),.B(G90));
  AND2 AND2_18(.VSS(VSS),.VDD(VDD),.Y(G87),.A(G85),.B(G86));
  AND4 AND4_2(.VSS(VSS),.VDD(VDD),.Y(G92),.A(G90),.B(G107),.C(G10),.D(G91));
  AND3 AND3_3(.VSS(VSS),.VDD(VDD),.Y(G93),.A(G94),.B(G122),.C(G123));
  AND4 AND4_3(.VSS(VSS),.VDD(VDD),.Y(G98),.A(G107),.B(G10),.C(G108),.D(G97));
  AND3 AND3_4(.VSS(VSS),.VDD(VDD),.Y(G99),.A(G116),.B(G122),.C(G123));
  AND4 AND4_4(.VSS(VSS),.VDD(VDD),.Y(G102),.A(G18),.B(G17),.C(G16),.D(G118));
  AND3 AND3_5(.VSS(VSS),.VDD(VDD),.Y(G103),.A(G104),.B(G122),.C(G123));
  AND4 AND4_5(.VSS(VSS),.VDD(VDD),.Y(G109),.A(G107),.B(G10),.C(G108),.D(G113));
  AND3 AND3_6(.VSS(VSS),.VDD(VDD),.Y(G110),.A(G112),.B(G122),.C(G123));
  AND3 AND3_7(.VSS(VSS),.VDD(VDD),.Y(G111),.A(G16),.B(G30),.C(G113));
  AND4 AND4_6(.VSS(VSS),.VDD(VDD),.Y(G119),.A(G116),.B(G16),.C(G117),.D(G118));
  AND3 AND3_8(.VSS(VSS),.VDD(VDD),.Y(G120),.A(G124),.B(G122),.C(G123));
  AND2 AND2_19(.VSS(VSS),.VDD(VDD),.Y(G121),.A(G124),.B(G125));
  AND4 AND4_7(.VSS(VSS),.VDD(VDD),.Y(G138),.A(G140),.B(G20),.C(G141),.D(G142));
  AND2 AND2_20(.VSS(VSS),.VDD(VDD),.Y(G139),.A(G145),.B(G146));
  AND4 AND4_8(.VSS(VSS),.VDD(VDD),.Y(G143),.A(G140),.B(G20),.C(G141),.D(G142));
  AND2 AND2_21(.VSS(VSS),.VDD(VDD),.Y(G144),.A(G145),.B(G146));
  AND3 AND3_9(.VSS(VSS),.VDD(VDD),.Y(G155),.A(G21),.B(G13),.C(G26));
  AND3 AND3_10(.VSS(VSS),.VDD(VDD),.Y(G156),.A(G163),.B(G172),.C(G13));
  AND2 AND2_22(.VSS(VSS),.VDD(VDD),.Y(G169),.A(G13),.B(G168));
  AND2 AND2_23(.VSS(VSS),.VDD(VDD),.Y(G170),.A(G184),.B(G177));
  AND2 AND2_24(.VSS(VSS),.VDD(VDD),.Y(G171),.A(G172),.B(G184));
  AND2 AND2_25(.VSS(VSS),.VDD(VDD),.Y(G175),.A(G174),.B(G12));
  AND2 AND2_26(.VSS(VSS),.VDD(VDD),.Y(G176),.A(G177),.B(G12));
  AND3 AND3_11(.VSS(VSS),.VDD(VDD),.Y(G181),.A(G180),.B(G13),.C(G21));
  AND3 AND3_12(.VSS(VSS),.VDD(VDD),.Y(G186),.A(G184),.B(G189),.C(G185));
  AND2 AND2_27(.VSS(VSS),.VDD(VDD),.Y(G191),.A(G189),.B(G190));
  AND2 AND2_28(.VSS(VSS),.VDD(VDD),.Y(G192),.A(G18),.B(G193));
  AND2 AND2_29(.VSS(VSS),.VDD(VDD),.Y(G196),.A(G195),.B(G13));
  AND2 AND2_30(.VSS(VSS),.VDD(VDD),.Y(G203),.A(G201),.B(G202));
  AND2 AND2_31(.VSS(VSS),.VDD(VDD),.Y(G204),.A(G205),.B(G29));
  AND2 AND2_32(.VSS(VSS),.VDD(VDD),.Y(G209),.A(G207),.B(G208));
  AND2 AND2_33(.VSS(VSS),.VDD(VDD),.Y(G210),.A(G212),.B(G30));
//
  OR2 OR2_0(.VSS(VSS),.VDD(VDD),.Y(G32),.A(G30),.B(G31));
  OR2 OR2_1(.VSS(VSS),.VDD(VDD),.Y(G33),.A(G72),.B(G12));
  OR4 OR4_0(.VSS(VSS),.VDD(VDD),.Y(G42),.A(G83),.B(G107),.C(G90),.D(G85));
  OR3 OR3_0(.VSS(VSS),.VDD(VDD),.Y(G43),.A(G83),.B(G11),.C(G14));
  OR4 OR4_1(.VSS(VSS),.VDD(VDD),.Y(G48),.A(G122),.B(G94),.C(G18),.D(G112));
  OR3 OR3_1(.VSS(VSS),.VDD(VDD),.Y(G49),.A(G122),.B(G94),.C(G116));
  OR2 OR2_2(.VSS(VSS),.VDD(VDD),.Y(G50),.A(G16),.B(G17));
  OR4 OR4_2(.VSS(VSS),.VDD(VDD),.Y(G53),.A(G83),.B(G11),.C(G14),.D(G85));
  OR4 OR4_3(.VSS(VSS),.VDD(VDD),.Y(G67),.A(G211),.B(G63),.C(G64),.D(G71));
  OR3 OR3_2(.VSS(VSS),.VDD(VDD),.Y(G68),.A(G65),.B(G211),.C(G66));
  OR4 OR4_4(.VSS(VSS),.VDD(VDD),.Y(G74),.A(G211),.B(G125),.C(G70),.D(G71));
  OR3 OR3_3(.VSS(VSS),.VDD(VDD),.Y(G75),.A(G72),.B(G211),.C(G73));
  OR4 OR4_5(.VSS(VSS),.VDD(VDD),.Y(G133),.A(G211),.B(G128),.C(G129),.D(G130));
  OR3 OR3_4(.VSS(VSS),.VDD(VDD),.Y(G134),.A(G131),.B(G211),.C(G132));
  OR4 OR4_6(.VSS(VSS),.VDD(VDD),.Y(G149),.A(G20),.B(G21),.C(G12),.D(G177));
  OR2 OR2_3(.VSS(VSS),.VDD(VDD),.Y(G150),.A(G184),.B(G25));
  OR2 OR2_4(.VSS(VSS),.VDD(VDD),.Y(G151),.A(G184),.B(G13));
  OR3 OR3_5(.VSS(VSS),.VDD(VDD),.Y(G152),.A(G163),.B(G21),.C(G12));
  OR2 OR2_5(.VSS(VSS),.VDD(VDD),.Y(G153),.A(G172),.B(G27));
  OR2 OR2_6(.VSS(VSS),.VDD(VDD),.Y(G154),.A(G184),.B(G27));
  OR4 OR4_7(.VSS(VSS),.VDD(VDD),.Y(G158),.A(G193),.B(G184),.C(G177),.D(G26));
  OR2 OR2_7(.VSS(VSS),.VDD(VDD),.Y(G159),.A(G189),.B(G157));
  OR2 OR2_8(.VSS(VSS),.VDD(VDD),.Y(G160),.A(G184),.B(G13));
  OR2 OR2_9(.VSS(VSS),.VDD(VDD),.Y(G161),.A(G20),.B(G13));
  OR2 OR2_10(.VSS(VSS),.VDD(VDD),.Y(G162),.A(G21),.B(G12));
  OR4 OR4_8(.VSS(VSS),.VDD(VDD),.Y(G164),.A(G20),.B(G21),.C(G12),.D(G177));
  OR3 OR3_6(.VSS(VSS),.VDD(VDD),.Y(G165),.A(G163),.B(G172),.C(G13));
  OR3 OR3_7(.VSS(VSS),.VDD(VDD),.Y(G166),.A(G172),.B(G177),.C(G24));
//
  NAND4 NAND4_0(.VSS(VSS),.VDD(VDD),.Y(G41),.A(G104),.B(G116),.C(G16),.D(G37));
  NAND2 NAND2_0(.VSS(VSS),.VDD(VDD),.Y(G62),.A(G67),.B(G68));
  NAND3 NAND3_0(.VSS(VSS),.VDD(VDD),.Y(G63),.A(G104),.B(G116),.C(G16));
  NAND4 NAND4_1(.VSS(VSS),.VDD(VDD),.Y(G64),.A(G65),.B(G21),.C(G20),.D(G19));
  NAND2 NAND2_1(.VSS(VSS),.VDD(VDD),.Y(G69),.A(G74),.B(G75));
  NAND4 NAND4_2(.VSS(VSS),.VDD(VDD),.Y(G70),.A(G72),.B(G12),.C(G21),.D(G20));
  NAND3 NAND3_1(.VSS(VSS),.VDD(VDD),.Y(G86),.A(G14),.B(G11),.C(G10));
  NAND3 NAND3_2(.VSS(VSS),.VDD(VDD),.Y(G88),.A(G42),.B(G43),.C(G59));
  NAND4 NAND4_3(.VSS(VSS),.VDD(VDD),.Y(G100),.A(G48),.B(G49),.C(G50),.D(G59));
  NAND2 NAND2_2(.VSS(VSS),.VDD(VDD),.Y(G118),.A(G53),.B(G122));
  NAND4 NAND4_4(.VSS(VSS),.VDD(VDD),.Y(G123),.A(G15),.B(G90),.C(G107),.D(G10));
  NAND4 NAND4_5(.VSS(VSS),.VDD(VDD),.Y(G125),.A(G19),.B(G104),.C(G116),.D(G16));
  NAND2 NAND2_3(.VSS(VSS),.VDD(VDD),.Y(G127),.A(G133),.B(G134));
  NAND2 NAND2_4(.VSS(VSS),.VDD(VDD),.Y(G128),.A(G116),.B(G16));
  NAND4 NAND4_6(.VSS(VSS),.VDD(VDD),.Y(G129),.A(G131),.B(G20),.C(G19),.D(G104));
  NAND2 NAND2_5(.VSS(VSS),.VDD(VDD),.Y(G130),.A(G32),.B(G33));
  NAND4 NAND4_7(.VSS(VSS),.VDD(VDD),.Y(G146),.A(G140),.B(G135),.C(G29),.D(G142));
  NAND4 NAND4_8(.VSS(VSS),.VDD(VDD),.Y(G178),.A(G164),.B(G165),.C(G166),.D(G189));
  NAND4 NAND4_9(.VSS(VSS),.VDD(VDD),.Y(G182),.A(G149),.B(G150),.C(G151),.D(G189));
  NAND2 NAND2_6(.VSS(VSS),.VDD(VDD),.Y(G187),.A(G158),.B(G159));
  NAND4 NAND4_10(.VSS(VSS),.VDD(VDD),.Y(G190),.A(G152),.B(G153),.C(G154),.D(G13));
  NAND4 NAND4_11(.VSS(VSS),.VDD(VDD),.Y(G197),.A(G160),.B(G161),.C(G162),.D(G189));
//
  NOR4 NOR4_0(.VSS(VSS),.VDD(VDD),.Y(G31),.A(G85),.B(G14),.C(G11),.D(G83));
  NOR2 NOR2_0(.VSS(VSS),.VDD(VDD),.Y(G37),.A(G124),.B(G112));
  NOR2 NOR2_1(.VSS(VSS),.VDD(VDD),.Y(G60),.A(G10),.B(G211));
  NOR4 NOR4_1(.VSS(VSS),.VDD(VDD),.Y(G61),.A(G76),.B(G77),.C(G78),.D(G211));
  NOR4 NOR4_2(.VSS(VSS),.VDD(VDD),.Y(G66),.A(G36),.B(G131),.C(G124),.D(G125));
  NOR2 NOR2_2(.VSS(VSS),.VDD(VDD),.Y(G71),.A(G35),.B(G30));
  NOR4 NOR4_3(.VSS(VSS),.VDD(VDD),.Y(G73),.A(G38),.B(G39),.C(G40),.D(G41));
  NOR4 NOR4_4(.VSS(VSS),.VDD(VDD),.Y(G79),.A(G80),.B(G81),.C(G82),.D(G211));
  NOR2 NOR2_3(.VSS(VSS),.VDD(VDD),.Y(G84),.A(G87),.B(G88));
  NOR3 NOR3_0(.VSS(VSS),.VDD(VDD),.Y(G89),.A(G92),.B(G93),.C(G95));
  NOR2 NOR2_4(.VSS(VSS),.VDD(VDD),.Y(G91),.A(G94),.B(G85));
  NOR2 NOR2_5(.VSS(VSS),.VDD(VDD),.Y(G95),.A(G44),.B(G45));
  NOR3 NOR3_1(.VSS(VSS),.VDD(VDD),.Y(G96),.A(G98),.B(G99),.C(G100));
  NOR2 NOR2_6(.VSS(VSS),.VDD(VDD),.Y(G97),.A(G46),.B(G47));
  NOR3 NOR3_2(.VSS(VSS),.VDD(VDD),.Y(G101),.A(G102),.B(G103),.C(G105));
  NOR2 NOR2_7(.VSS(VSS),.VDD(VDD),.Y(G105),.A(G51),.B(G52));
  NOR4 NOR4_5(.VSS(VSS),.VDD(VDD),.Y(G106),.A(G109),.B(G110),.C(G111),.D(G114));
  NOR3 NOR3_3(.VSS(VSS),.VDD(VDD),.Y(G108),.A(G94),.B(G85),.C(G14));
  NOR3 NOR3_4(.VSS(VSS),.VDD(VDD),.Y(G113),.A(G54),.B(G55),.C(G56));
  NOR2 NOR2_8(.VSS(VSS),.VDD(VDD),.Y(G114),.A(G57),.B(G58));
  NOR4 NOR4_6(.VSS(VSS),.VDD(VDD),.Y(G115),.A(G119),.B(G120),.C(G121),.D(G126));
  NOR3 NOR3_5(.VSS(VSS),.VDD(VDD),.Y(G117),.A(G124),.B(G112),.C(G18));
  NOR3 NOR3_6(.VSS(VSS),.VDD(VDD),.Y(G132),.A(G34),.B(G124),.C(G125));
  NOR3 NOR3_7(.VSS(VSS),.VDD(VDD),.Y(G137),.A(G138),.B(G139),.C(G211));
  NOR2 NOR2_9(.VSS(VSS),.VDD(VDD),.Y(G142),.A(G13),.B(G136));
  NOR4 NOR4_7(.VSS(VSS),.VDD(VDD),.Y(G167),.A(G169),.B(G170),.C(G171),.D(G193));
  NOR3 NOR3_8(.VSS(VSS),.VDD(VDD),.Y(G173),.A(G175),.B(G176),.C(G178));
  NOR2 NOR2_10(.VSS(VSS),.VDD(VDD),.Y(G179),.A(G181),.B(G182));
  NOR2 NOR2_11(.VSS(VSS),.VDD(VDD),.Y(G183),.A(G186),.B(G187));
  NOR2 NOR2_12(.VSS(VSS),.VDD(VDD),.Y(G185),.A(G155),.B(G156));
  NOR2 NOR2_13(.VSS(VSS),.VDD(VDD),.Y(G188),.A(G191),.B(G192));
  NOR2 NOR2_14(.VSS(VSS),.VDD(VDD),.Y(G193),.A(G143),.B(G144));
  NOR2 NOR2_15(.VSS(VSS),.VDD(VDD),.Y(G194),.A(G196),.B(G197));
  NOR3 NOR3_9(.VSS(VSS),.VDD(VDD),.Y(G200),.A(G203),.B(G204),.C(G211));
  NOR3 NOR3_10(.VSS(VSS),.VDD(VDD),.Y(G206),.A(G209),.B(G210),.C(G211));
//

endmodule