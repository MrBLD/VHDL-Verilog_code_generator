module s5378(n3065gat,n3110gat,n3074gat,n3121gat,n3079gat,n3148gat,n3127gat,n3105gat,n3141gat,n3146gat,n3094gat,n3137gat,n3104gat,n3067gat,n3069gat,n3089gat,n3108gat,n3143gat,n3132gat,n3147gat,n3129gat,n3091gat,n3124gat,n3134gat,VDD,n3070gat,n3117gat,n3068gat,n3093gat,n3099gat,n3098gat,n3100gat,n3151gat,n3073gat,n3138gat,n3144gat,n3097gat,n3084gat,n3066gat,n3109gat,n3088gat,n3083gat,n3072gat,n3082gat,n3115gat,n3120gat,n3118gat,n3114gat,n3113gat,n3106gat,n3142gat,n3145gat,n3077gat,n3090gat,n3107gat,n3123gat,n3150gat,n3111gat,n3130gat,n3081gat,n3126gat,n3131gat,n3135gat,n3087gat,n3119gat,n3086gat,n3152gat,n3133gat,n3080gat,n3095gat,n3116gat,n3122gat,n3085gat,n3112gat,n3125gat,n3128gat,VSS,n3139gat,n3140gat,n3136gat,n3078gat,CLOCK,n3076gat,n3075gat,n3149gat,n3092gat,n3071gat);
input n3065gat,n3074gat,n3088gat,n3083gat,n3072gat,n3082gat,n3079gat,n3077gat,n3090gat,n3094gat,n3067gat,n3069gat,n3089gat,n3081gat,n3087gat,n3086gat,n3091gat,n3080gat,VDD,n3070gat,n3095gat,n3068gat,n3093gat,n3099gat,n3098gat,n3100gat,n3073gat,n3085gat,VSS,n3078gat,n3097gat,CLOCK,n3076gat,n3084gat,n3066gat,n3075gat,n3092gat,n3071gat;
output n3110gat,n3115gat,n3120gat,n3118gat,n3114gat,n3148gat,n3113gat,n3106gat,n3105gat,n3127gat,n3141gat,n3142gat,n3145gat,n3107gat,n3123gat,n3146gat,n3137gat,n3150gat,n3111gat,n3104gat,n3130gat,n3108gat,n3126gat,n3131gat,n3132gat,n3135gat,n3143gat,n3119gat,n3147gat,n3129gat,n3152gat,n3124gat,n3133gat,n3134gat,n3117gat,n3116gat,n3151gat,n3122gat,n3112gat,n3138gat,n3125gat,n3128gat,n3139gat,n3140gat,n3144gat,n3136gat,n3149gat,n3121gat,n3109gat;

  wire n2756gat,n2729gat,n3020gat,n296gat,n2622gat,n2867gat,n1150gat,n1304gat,n2602gat,I2238,n334gat,n2637gat,I62,I658,I3191,n583gat,n1298gat,I44,n2726gat,n2782gat,n1269gat,n2979gat,n2827gat,n734gat,n811gat,I3000,n2237gat,n1503gat,n1259gat,n511gat,I2989,I2934,n595gat,n228gat,I729,n2143gat,n3032gat,n1686gat,I1981,n1055gat,n1717gat,n2123gat,n1230gat,n2669gat,n2364gat,n834gat,n733gat,n662gat,I4750,n1816gat,n1439gat,n2852gat,n390gat,n2470gat,n567gat,n2903gat,n1481gat,I3713,I4475,n1712gat,I2130,n2780gat,n1146gat,n1644gat,n1175gat,n1389gat,n2843gat,n2595gat,n2218gat,I2890,n1458gat,n858gat,n2419gat,n807gat,n3053gat,n1606gat,n1387gat,n983gat,n661gat,n2574gat,I334,n2363gat,n2358gat,n782gat,n1157gat,n1280gat,n2701gat,n1846gat,n1962gat,I3287,n1460gat,I206,I1769,n368gat,n2350gat,n297gat,n242gat,n2886gat,n652gat,n2760gat,n769gat,n1559gat,n2487gat,n229gat,n837gat,n2751gat,n2281gat,n1030gat,n2891gat,n2325gat,n1880gat,n899gat,n164gat,n2706gat,I317,I1302,n1470gat,I796,n1791gat,n2789gat,n1082gat,I4720,n2764gat,n195gat,n2410gat,n2731gat,n520gat,n1115gat,n3064gat,I1278,n3003gat,I4690,n2150gat,I746,n2282gat,n3037gat,n2707gat,n1043gat,n2401gat,n2854gat,n2044gat,n758gat,n1329gat,I4573,n169gat,n784gat,I1371,n1351gat,n2243gat,n1281gat,n38gat,n1869gat,n3034gat,n1217gat,n795gat,n337gat,n1467gat,I1860,n148gat,n749gat,n2895gat,n77gat,n483gat,n2839gat,n1419gat,n1765gat,I453,I4774,n844gat,n751gat,n374gat,n2879gat,n2508gat,n561gat,n1279gat,n2681gat,n620gat,n2433gat,n1334gat,n1260gat,n470gat,n3016gat,n664gat,n1208gat,n132gat,n912gat,n1698gat,n759gat,n2672gat,I256,n176gat,n1192gat,n339gat,n1548gat,n634gat,n2201gat,n366gat,I3491,n2207gat,I1667,n2900gat,I579,n1215gat,n532gat,n1349gat,n1632gat,n2474gat,I793,n2746gat,n1410gat,n1842gat,n2270gat,I977,I2169,n2004gat,n1286gat,n2601gat,I1255,n2338gat,n1604gat,n768gat,I753,n2884gat,n1239gat,n1926gat,n1414gat,I4753,n2440gat,n2000gat,n881gat,n1971gat,I4672,n874gat,n233gat,n1551gat,n2422gat,n2648gat,n1836gat,n2658gat,n1568gat,n1957gat,n2941gat,n1461gat,I1500,I512,n1305gat,n2853gat,I259,n1284gat,I1248,I1734,I2847,n1702gat,n655gat,n908gat,n1620gat,n1838gat,n1740gat,n1003gat,I921,I100,n724gat,I661,n743gat,n2524gat,n1479gat,n1671gat,n1495gat,n69gat,I4708,n259gat,I715,n1179gat,n659gat,n1967gat,n1747gat,I4759,n1119gat,I203,n2359gat,n261gat,n2781gat,n2695gat,I4626,n1466gat,n2093gat,I14,I1488,n2625gat,n219gat,n1552gat,n2396gat,n988gat,n2355gat,I2162,n476gat,n126gat,n1237gat,n313gat,n1258gat,n788gat,n1486gat,n1308gat,n89gat,n2168gat,n572gat,I4660,n1600gat,n716gat,n2561gat,n144gat,n1670gat,n1888gat,n2629gat,n199gat,n2806gat,n1076gat,I3290,I2235,n336gat,n913gat,n1892gat,n1978gat,n2824gat,n2656gat,n2838gat,I1388,n2533gat,n410gat,n2146gat,n333gat,n2986gat,n1871gat,n1314gat,I846,I1899,n2947gat,n2138gat,n2943gat,n1555gat,n2630gat,I4506,I1584,I4738,n391gat,n1515gat,I4524,n2682gat,I2831,n2709gat,n54gat,n1358gat,n1197gat,n2506gat,n2031gat,n2697gat,I223,n1123gat,n1316gat,n2749gat,n650gat,n1099gat,n2293gat,n1771gat,n401gat,I1996,n2570gat,n2766gat,n903gat,n2551gat,I1894,n3045gat,n375gat,I1795,n521gat,I863,I675,I1216,n2025gat,I65,n1801gat,n989gat,n2097gat,n2209gat,n2878gat,n648gat,I936,n1575gat,n2931gat,n855gat,I1118,n964gat,n2449gat,n1285gat,n1080gat,n2090gat,n2951gat,n197gat,n1665gat,n1599gat,n2812gat,n756gat,n1229gat,n1074gat,n2223gat,n2926gat,n1525gat,n930gat,n1054gat,I1999,n331gat,n992gat,n1988gat,n1769gat,n1622gat,n910gat,n416gat,n2823gat,n1490gat,n1118gat,n757gat,n442gat,n1724gat,I1002,n3017gat,n1161gat,n1659gat,n1582gat,n1827gat,n1441gat,n959gat,n1462gat,n498gat,n168gat,n2399gat,n510gat,n1011gat,I620,n3018gat,n2967gat,n2699gat,n2054gat,n345gat,n741gat,I4105,n1218gat,I2109,I395,n225gat,n1058gat,n2841gat,I248,I3143,n3061gat,I2394,I692,n1327gat,n1104gat,n840gat,n3030gat,n1401gat,n2571gat,n522gat,n484gat,n1918gat,I1515,n1927gat,n1159gat,I4678,n1761gat,n1270gat,n1196gat,n1639gat,n1886gat,n2952gat,n1645gat,I1439,I2935,n1634gat,n2197gat,n925gat,I4798,n93gat,n810gat,I2837,I3635,n1963gat,n364gat,I468,I980,n1834gat,I4312,n935gat,n2999gat,n1176gat,n3052gat,n2617gat,n2807gat,I1877,n2418gat,n127gat,n1685gat,I4309,n2797gat,n2389gat,n791gat,n696gat,n2438gat,n2995gat,n686gat,n965gat,n761gat,n2864gat,n1268gat,n2741gat,n2135gat,n808gat,n2162gat,I3703,n1375gat,n820gat,n822gat,I4558,n314gat,I815,n1646gat,n1309gat,n1829gat,n2317gat,I3336,I3742,n1455gat,n996gat,n372gat,n861gat,n629gat,n656gat,n2115gat,n2971gat,n325gat,n1112gat,n1057gat,n2255gat,n2119gat,I1655,n1550gat,n2125gat,I2014,n1691gat,I4792,n2924gat,n617gat,n2633gat,n1415gat,n125gat,I1152,I1115,n2258gat,n2611gat,I3867,n409gat,n2753gat,n902gat,n848gat,n2021gat,I1082,n2705gat,n1453gat,n698gat,n2846gat,n159gat,I4780,n2565gat,n1819gat,I3530,n40gat,n905gat,n2536gat,n2252gat,n760gat,I3293,n354gat,n1338gat,n657gat,n2494gat,n2820gat,n1012gat,n2997gat,n1532gat,n957gat,I3315,n349gat,n1079gat,I812,I2251,I3954,n796gat,n1790gat,n898gat,n2961gat,n2950gat,n1895gat,n1009gat,n1096gat,n2139gat,n2329gat,n2430gat,n946gat,n2844gat,n1570gat,n977gat,n3001gat,I3390,n2765gat,n360gat,n2804gat,n852gat,I1703,n2516gat,n1422gat,n460gat,n414gat,n13gat,n1696gat,n907gat,n2557gat,n155gat,I1183,n1785gat,I282,n568gat,n2052gat,n962gat,n1915gat,n960gat,n1271gat,n1859gat,n2257gat,n343gat,n2330gat,n2450gat,n1026gat,n2203gat,n1133gat,n1417gat,n2662gat,I1496,n1718gat,n2176gat,n1034gat,n677gat,n1850gat,n1478gat,n392gat,n1394gat,n1024gat,n2916gat,n2194gat,I1791,n2929gat,n1233gat,I3935,n1381gat,I4777,n871gat,n2499gat,n174gat,n2628gat,n701gat,n423gat,n680gat,n1091gat,n2579gat,I178,I300,n2205gat,n2253gat,n2974gat,n2215gat,n979gat,n2946gat,n2634gat,n1986gat,n801gat,n591gat,I4744,n1778gat,n2269gat,n2417gat,n859gat,I3149,n279gat,n85gat,I2735,n417gat,n2720gat,I340,n1100gat,I4726,I1121,I2873,n1651gat,n1521gat,n2761gat,n1318gat,n1821gat,n457gat,n65gat,n2860gat,n1716gat,n2689gat,I4108,n273gat,n1658gat,n1640gat,n555gat,n991gat,n2152gat,n3011gat,I1630,I3610,I4729,n945gat,n1307gat,I4485,n2414gat,I955,I4222,n445gat,n22gat,n967gat,n2014gat,n779gat,n1576gat,n2996gat,I2812,I2084,n667gat,n2492gat,n2249gat,n2640gat,I4702,n1336gat,n509gat,n137gat,n1204gat,I985,n1315gat,n1655gat,I440,n2124gat,n2035gat,n793gat,n880gat,n1340gat,n188gat,n2351gat,n2745gat,I2439,n2942gat,n2890gat,I1344,n16gat,n3050gat,n250gat,n1523gat,I3429,n2017gat,n1060gat,n121gat,n997gat,n170gat,n1887gat,n361gat,n1248gat,n987gat,n833gat,n1823gat,n204gat,n1733gat,n1253gat,n641gat,n867gat,n922gat,n984gat,n2596gat,n1408gat,n2169gat,I1422,n350gat,n2288gat,n2456gat,n1224gat,n2050gat,n1013gat,n1653gat,n2290gat,n574gat,n1891gat,n2163gat,n1719gat,n2060gat,n865gat,n1392gat,n1332gat,n1683gat,n2514gat,I240,n2646gat,n2994gat,n1999gat,n2624gat,n683gat,n2885gat,n948gat,I2254,n365gat,I1169,n1424gat,n3023gat,I4236,n1714gat,n2918gat,n1017gat,I623,n856gat,n711gat,n864gat,n2559gat,n37gat,n2468gat,I4409,n1383gat,n1748gat,n1556gat,n2650gat,n1114gat,I5,I3509,n295gat,n2842gat,n854gat,n1662gat,I3817,I3841,n1435gat,I1079,I47,I331,n985gat,I3962,I1,n1581gat,I2088,n255gat,n2606gat,n2416gat,n777gat,n2292gat,I1927,n2552gat,n179gat,I4554,I3342,n2845gat,n587gat,I76,I2056,n566gat,I1243,n1958gat,n263gat,I476,n1173gat,n34gat,n2694gat,n62gat,n151gat,n1407gat,n573gat,n2018gat,n2758gat,n2822gat,I3273,n2588gat,n1090gat,I726,n462gat,n2538gat,n702gat,n2202gat,I278,n1045gat,n1739gat,n3040gat,n2913gat,n972gat,I4693,n1379gat,n1593gat,n2732gat,n17gat,I930,n2486gat,n1730gat,n2985gat,n2614gat,I381,n1400gat,n2917gat,n2887gat,n2110gat,I2696,n2575gat,I456,I1476,n1845gat,I409,I2420,n2921gat,n3049gat,n49gat,n1010gat,n1077gat,n1643gat,n2808gat,I1411,n2934gat,n815gat,n1565gat,n1707gat,n136gat,I1857,I3303,n671gat,n450gat,n413gat,n785gat,n3057gat,n519gat,n1584gat,n2027gat,I842,n330gat,n2250gat,n719gat,I480,I2324,n1557gat,I4518,n2920gat,n1369gat,n451gat,I2925,I3999,n1219gat,n2577gat,n2677gat,n1870gat,I3472,n653gat,I443,n1202gat,n2737gat,n2402gat,n883gat,I4135,n485gat,n2964gat,n1817gat,n1623gat,I1493,n496gat,n2531gat,n2919gat,I790,n1257gat,I4212,n222gat,n978gat,n2905gat,n505gat,n1372gat,n2541gat,n398gat,n2767gat,n823gat,I734,n1106gat,n980gat,n2638gat,n2403gat,I1011,n2306gat,n2684gat,n2965gat,n2214gat,n775gat,n891gat,n73gat,n804gat,n982gat,n2837gat,n684gat,n726gat,n2794gat,n1737gat,n501gat,n396gat,n1533gat,n1420gat,n327gat,n2703gat,n134gat,n2944gat,n240gat,n1631gat,n3056gat,I1227,n2245gat,I4512,I576,I899,I4705,n970gat,n2084gat,n1605gat,n1642gat,n358gat,I3056,n177gat,n1885gat,n335gat,n873gat,n2117gat,I3539,n2992gat,I1399,n1633gat,I426,n2597gat,n441gat,n2819gat,n2700gat,I111,n1147gat,n495gat,n776gat,n1430gat,n934gat,n2131gat,n1068gat,n1443gat,n243gat,n968gat,n2738gat,I1067,n1174gat,n2636gat,n1553gat,n165gat,n1201gat,n1195gat,n513gat,n1216gat,I449,n2346gat,I2049,n690gat,n915gat,n84gat,n2882gat,n2059gat,n2504gat,n963gat,n713gat,I3621,n1367gat,n766gat,n1194gat,n1828gat,n377gat,n2095gat,n2564gat,I297,n2573gat,n882gat,n2642gat,I437,n2639gat,n406gat,I2915,n1002gat,I4372,n1200gat,n1275gat,n66gat,n1615gat,n1694gat,n1498gat,I4081,n1669gat,n929gat,n1203gat,n1767gat,n2265gat,n2925gat,n703gat,I4765,I4117,n2101gat,I4771,n341gat,n2158gat,n1641gat,n819gat,I4723,n1916gat,n1236gat,n1228gat,I2044,n1832gat,n1507gat,n878gat,n2883gat,n1711gat,n1960gat,I4194,n1773gat,n1021gat,n2073gat,n1654gat,n931gat,I858,n224gat,I1837,I401,n1879gat,n805gat,n2482gat,n1690gat,n2547gat,I4129,n194gat,n2877gat,I606,n2159gat,n2480gat,n2534gat,n1373gat,I718,n294gat,I3765,n1544gat,n1775gat,n755gat,n2409gat,I4217,n737gat,n2518gat,I1724,I3660,n961gat,n2955gat,I741,I3646,n637gat,n851gat,n2151gat,n3002gat,n2522gat,n857gat,n1207gat,n2384gat,n1961gat,n941gat,n1974gat,n682gat,n2129gat,n2619gat,n2686gat,n2341gat,n2266gat,n2553gat,n763gat,n1413gat,n1894gat,I1190,n1849gat,n299gat,I721,n317gat,n1396gat,n636gat,I2721,n2680gat,n2928gat,n1085gat,n2998gat,n3008gat,n504gat,n2413gat,I2157,n2615gat,n1756gat,n531gat,n2128gat,I958,n1807gat,n2783gat,n927gat,n2815gat,n628gat,n387gat,n480gat,I651,n900gat,n1841gat,n2910gat,n1089gat,n1447gat,n1468gat,n1878gat,n1162gat,n830gat,n2710gat,I1028,I4227,I270,n738gat,n1135gat,n1163gat,n577gat,n670gat,n2821gat,I4786,n966gat,n1053gat,n110gat,n1431gat,n1735gat,n2616gat,n1487gat,n1734gat,n672gat,n52gat,I1023,n1182gat,n1274gat,n2938gat,n12gat,n1483gat,n2436gat,n732gat,n58gat,n1044gat,n802gat,n292gat,n2716gat,n2219gat,n1595gat,I1091,I2433,I1209,n2353gat,n2592gat,n2127gat,n725gat,n1543gat,I4233,I1178,I171,n1745gat,n2973gat,I311,n2356gat,n3042gat,n3005gat,n2647gat,I749,n2560gat,I1585,I1749,I4014,I4768,I594,n1244gat,n754gat,I3339,n853gat,I3677,n1072gat,n394gat,n1231gat,I818,n378gat,n1172gat,I243,n1678gat,I851,n1882gat,I2112,n2796gat,n753gat,n171gat,I2885,I1550,I1920,n2082gat,n2566gat,n936gat,n2691gat,n2002gat,n2757gat,I4714,n322gat,n1220gat,n2612gat,I4623,n2476gat,n1225gat,n1459gat,n824gat,n1618gat,n422gat,n1366gat,I1908,n645gat,n2426gat,n3063gat,n1502gat,n909gat,n278gat,n163gat,n2847gat,n1416gat,n818gat,n1656gat,n2949gat,n76gat,n2079gat,I4747,n1252gat,n1603gat,n2167gat,n386gat,n1831gat,n649gat,n842gat,n316gat,n1784gat,I192,n2978gat,n863gat,n2407gat,n1370gat,n408gat,n589gat,n2569gat,n926gat,I1277,n2825gat,I2344,n2805gat,n1451gat,n1371gat,n1352gat,n2862gat,n1494gat,n288gat,I768,n491gat,n1477gat,n1667gat,n2609gat,n1728gat,n933gat,n1294gat,I3513,n1223gat,n2936gat,n1428gat,n1528gat,n1406gat,n901gat,n2490gat,n59gat,n1291gat,I3549,I3309,n2537gat,n2309gat,n707gat,n2954gat,n2029gat,n2289gat,n1374gat,n1625gat,n499gat,n1798gat,n1554gat,n2190gat,n986gat,n586gat,n1577gat,n924gat,n173gat,I398,n2793gat,n718gat,n2261gat,I2177,n1704gat,n841gat,n2196gat,n15gat,n1348gat,n1266gat,I642,n571gat,n2056gat,n814gat,n2586gat,n750gat,I50,I3387,n2590gat,n2448gat,n180gat,n357gat,n1699gat,n689gat,n2387gat,n373gat,n2005gat,n2784gat,n3029gat,n2762gat,n1324gat,I230,n2498gat,n3014gat,n2826gat,n621gat,n1117gat,n167gat,I1007,n21gat,n1193gat,n890gat,n172gat,n1403gat,n1263gat,n189gat,I210,n588gat,n2532gat,n2715gat,n2187gat,n1531gat,n2264gat,n2246gat,n1035gat,n1994gat,n917gat,I913,n489gat,n2935gat,n1945gat,n2460gat,I2181,n954gat,I678,n1580gat,n1619gat,n2053gat,n482gat,n1695gat,n1360gat,n3026gat,n829gat,n1014gat,n1598gat,n493gat,n2755gat,I1708,n673gat,n1325gat,n974gat,n200gat,n448gat,n2055gat,n1925gat,I877,n1652gat,n748gat,n836gat,n1613gat,I4789,n2328gat,n797gat,n643gat,n1889gat,n584gat,n593gat,n479gat,I834,n530gat,I1723,n551gat,I1138,n631gat,n1970gat,n35gat,I687,I3318,n897gat,n2959gat,n1732gat,n2058gat,n518gat,I2385,n2493gat,n2698gat,n237gat,I1683,n1023gat,n2892gat,n503gat,I2417,n2256gat,n226gat,I4144,n765gat,n2217gat,n1276gat,I591,n687gat,I3882,n1660gat,I2953,n2134gat,n2652gat,n129gat,n553gat,I3461,n320gat,n2906gat,n2786gat,n158gat,I4530,I2672,n3051gat,n2427gat,n916gat,n1703gat,n2932gat,n565gat,n1616gat,n1454gat,n1339gat,n1626gat,I2785,n2049gat,n281gat,n2966gat,n885gat,n370gat,I2271,n1095gat,n1742gat,n2200gat,I3494,n2443gat,n2608gat,n380gat,I3945,n2776gat,n39gat,n3007gat,n1425gat,n1205gat,n2660gat,n1028gat,n2181gat,n1847gat,n1418gat,n3025gat,n2802gat,I1166,n1191gat,n1006gat,n415gat,n207gat,n2894gat,n781gat,n2081gat,n1649gat,n1347gat,n580gat,n1001gat,I275,n2983gat,I1103,n79gat,n502gat,n447gat,I2978,n1380gat,I2257,n1361gat,n624gat,n944gat,n1446gat,n111gat,I237,n2520gat,n3059gat,n1614gat,I217,n481gat,n2858gat,I1353,n1862gat,n2343gat,I1807,n1774gat,n2785gat,n3022gat,I3394,n1763gat,n1213gat,n2620gat,n45gat,n1675gat,n876gat,n2958gat,n1608gat,I3179,n1956gat,n2037gat,n256gat,n2702gat,n120gat,n1226gat,n2184gat,n904gat,n1518gat,I314,n2500gat,n3038gat,n1016gat,n646gat,n1154gat,I3777,n2863gat,n2724gat,n2721gat,n2896gat,n2610gat,n508gat,n355gat,n3010gat,I1085,n618gat,n1485gat,n1519gat,n894gat,n2193gat,n262gat,n2182gat,n918gat,n2963gat,n407gat,n2690gat,n1760gat,n141gat,n2859gat,n1602gat,n1350gat,n1444gat,n2881gat,n2599gat,n1189gat,n590gat,n2868gat,n3048gat,n2719gat,n2723gat,I2228,n458gat,I637,n635gat,n2478gat,n1376gat,I149,n1601gat,n1520gat,I1031,n1594gat,n735gat,n1241gat,n1032gat,n1701gat,I1903,n2284gat,n622gat,n130gat,n2133gat,n1668gat,n2437gat,n1731gat,n1105gat,n351gat,n1848gat,n247gat,n2613gat,n658gat,n614gat,n666gat,n348gat,n1178gat,I2771,n745gat,n2555gat,n1427gat,n2632gat,n1673gat,n1924gat,n2816gat,n1705gat,n2211gat,n632gat,I4783,n238gat,I4055,n644gat,n2406gat,n1188gat,I4000,n1007gat,n1101gat,n1438gat,n264gat,n2750gat,n613gat,n694gat,n160gat,n2790gat,I776,n849gat,n2013gat,n2040gat,n783gat,n2735gat,n251gat,n2948gat,I27,I3300,n1793gat,n746gat,n886gat,n971gat,n2439gat,n2148gat,n739gat,n1482gat,n1051gat,n1301gat,I196,n740gat,I1201,n752gat,n227gat,n792gat,n1116gat,n1330gat,n1440gat,n1088gat,n71gat,n1186gat,I2275,n267gat,n2813gat,n2775gat,n2061gat,n2244gat,n2347gat,n1153gat,n2754gat,n1254gat,n2078gat,n1562gat,I2414,n2687gat,n1097gat,I1698,n1087gat,n3013gat,I609,n576gat,n1917gat,n419gat,n578gat,n2147gat,n2977gat,n2016gat,n1450gat,n1710gat,n2185gat,n2809gat,n1573gat,I461,n1265gat,n563gat,I2731,n1792gat,n2912gat,I4633,I1236,I1833,I963,n1209gat,n720gat,n1071gat,n1472gat,n2850gat,n393gat,n2902gat,I4429,n463gat,n1549gat,n469gat,n1078gat,n789gat,n514gat,n1721gat,n2342gat,I2127,n809gat,n1476gat,n947gat,n140gat,n2199gat,n2558gat,n453gat,I1204,n1363gat,n1353gat,n2861gat,n382gat,n887gat,n461gat,I375,n475gat,n1884gat,n2198gat,n2423gat,n2727gat,I4756,I3754,n326gat,n2893gat,n266gat,n1758gat,n2744gat,I880,I902,I2380,I2148,n1066gat,n456gat,I1783,n2855gat,I1251,I3691,n2562gat,n212gat,I3948,n2319gat,n1029gat,n1469gat,n42gat,n712gat,n2851gat,n2984gat,n3015gat,n1779gat,n412gat,n1762gat,n1648gat,I4432,I4717,n388gat,n2452gat,n2260gat,I2684,n1596gat,n2665gat,n1865gat,n1436gat,n692gat,n2461gat,I227,n951gat,n709gat,n2572gat,n665gat,n321gat,n2836gat,I359,n715gat,n515gat,n1989gat,n1991gat,n1590gat,n2548gat,I2349,n3033gat,n1437gat,n803gat,n1563gat,n2869gat,n3027gat,n283gat,n248gat,n731gat,n478gat,n1578gat,n1303gat,n1008gat,n2792gat,n2108gat,n2488gat,n290gat,n2810gat,I2372,n352gat,n1935gat,n1033gat,n747gat,n921gat,I4452,n252gat,n2795gat,n1249gat,n3043gat,n2962gat,n122gat,n182gat,n2693gat,n1019gat,n790gat,n449gat,n1319gat,n2099gat,n1661gat,I4499,n1529gat,n2567gat,n1398gat,n2048gat,n2930gat,I1481,n2141gat,I4620,n444gat,n993gat,n2132gat,I414,n2130gat,n1409gat,n2667gat,n710gat,n722gat,I4412,n1382gat,n2897gat,n1302gat,n1322gat,n1031gat,n1211gat,n1378gat,n133gat,n911gat,I3235,I1407,n88gat,n1412gat,n2696gat,n1111gat,I1339,n275gat,n1356gat,n2957gat,n1709gat,n446gat,n1898gat,n3006gat,I4762,n1181gat,n2604gat,n14gat,I3211,n558gat,n1896gat,n2581gat,n2285gat,I4145,n2655gat,n2907gat,I4666,n1923gat,n2192gat,n2679gat,I2263,n2466gat,n346gat,n184gat,n2179gat,I2232,n2549gat,n569gat,n2911gat,n271gat,I2736,n2814gat,n347gat,n2621gat,n2708gat,I3941,n1448gat,I4601,n2262gat,n3054gat,I4663,n1825gat,I3914,I1174,I3401,n187gat,n774gat,I264,I1766,I2843,n2730gat,n2937gat,I1230,I23,I3891,I1016,n494gat,n2137gat,n2502gat,n1657gat,I3957,n2644gat,n517gat,n1199gat,I1124,n1700gat,n990gat,I423,I3465,n2987gat,n287gat,I4542,n241gat,n1607gat,I97,n2429gat,n3041gat,I1453,n147gat,n1783gat,n359gat,n1866gat,n794gat,n2685gat,n2251gat,n2743gat,n1251gat,n1586gat,n642gat,n950gat,n2875gat,n1510gat,n2718gat,n773gat,n1629gat,I1155,n2578gat,n1713gat,n1572gat,n270gat,n2489gat,n1920gat,I2376,n443gat,I1947,I646,n2663gat,n53gat,I1348,n268gat,n955gat,n44gat,I4580,n2091gat,n2545gat,n2568gat,n1160gat,n2927gat,n2352gat,I4138,n1722gat,n2904gat,n2922gat,n1921gat,I4216,n1508gat,n2981gat,n1246gat,n2446gat,n1075gat,n318gat,n1954gat,n1321gat,n838gat,n2454gat,n1517gat,n1093gat,n2923gat,I2400,n2188gat,n527gat,n2001gat,n2829gat,I3148,I11,n3000gat,n2530gat,n1860gat,n146gat,n63gat,n1240gat,n2901gat,n1156gat,n1359gat,n892gat,n1052gat,I2319,n1190gat,n1005gat,n1411gat,n2768gat,I837,n356gat,n1365gat,n1706gat,n1736gat,n888gat,n2990gat,n2349gat,n1158gat,n616gat,n2149gat,I2428,I1436,n1919gat,n1025gat,n895gat,n78gat,n1621gat,n2970gat,n2540gat,n1610gat,I320,n3009gat,n1151gat,n714gat,I1516,n612gat,n468gat,n771gat,n1222gat,n1326gat,n1084gat,I4492,n1059gat,I4489,n2546gat,n2982gat,n507gat,n1708gat,n512gat,n2390gat,I4587,n254gat,I4352,I1874,I2248,I3951,I1035,n523gat,n223gat,n2688gat,I4478,n1800gat,n1357gat,n1630gat,n695gat,n2989gat,n663gat,n2803gat,n1134gat,n1840gat,I4684,I1322,n11gat,n956gat,n2607gat,n2331gat,I4449,n706gat,n1684gat,n1273gat,n384gat,n2345gat,n3046gat,n2664gat,n128gat,n369gat,n2283gat,n973gat,n1355gat,n2339gat,n647gat,n2550gat,n2195gat,n1496gat,I4369,n1148gat,n152gat,I3520,n2740gat,n2671gat,n845gat,n1558gat,n2354gat,n181gat,I3312,n344gat,n1666gat,n48gat,n2102gat,I4067,n2980gat,n2239gat,n1777gat,n2337gat,I885,n2388gat,n1183gat,n717gat,I1450,n1973gat,n1256gat,n582gat,I4741,n1377gat,n1635gat,I3412,n2666gat,I1923,n2213gat,n1312gat,n418gat,I4687,n2057gat,n2733gat,n72gat,n2828gat,n1243gat,I4732,n1120gat,n1180gat,n2940gat,n1272gat,I4615,n3031gat,n2458gat,n949gat,n1782gat,n402gat,n1636gat,n2444gat,I1800,n1086gat,I1319,n1863gat,I3174,n1505gat,I368,I4735,I220,n64gat,n2742gat,n41gat,n525gat,n1214gat,n2673gat,n1858gat,n92gat,I1141,I1843,n2798gat,n2991gat,n2009gat,n1561gat,n3047gat,n2394gat,n3019gat,n1442gat,n937gat,n1723gat,n1780gat,n124gat,n1102gat,n1210gat,n2238gat,n1368gat,n767gat,n1177gat,n269gat,n2747gat,n497gat,n1277gat,n50gat,n2291gat,n1499gat,I3457,n1818gat,n2888gat,n2668gat,I2035,I2153,n3004gat,n231gat,n1235gat,n3028gat,n943gat,n772gat,I337,n1293gat,n1786gat,n2969gat,n2914gat,n1839gat,n2259gat,n1796gat,n1516gat,n1546gat,n651gat,n2556gat,I583,n2817gat,n1164gat,I2040,n1238gat,n1423gat,n1787gat,n362gat,I4023,n906gat,n1306gat,n893gat,n258gat,n2042gat,n1588gat,n274gat,I4329,I81,n705gat,n762gat,n61gat,n2777gat,n914gat,n1934gat,I1467,I3587,n1964gat,n2649gat,n896gat,n1000gat,n654gat,n1402gat,n1184gat,n1627gat,n1729gat,n86gat,n1569gat,I709,n579gat,I4651,I4675,n2832gat,I1127,n2661gat,I4020,n2734gat,I4482,n2472gat,n1245gat,n1267gat,n1262gat,n2393gat,I2260,n2464gat,I473,I3306,n260gat,n421gat,n2189gat,n1113gat,I3831,n143gat,I4654,I3808,n1155gat,n1449gat,n2830gat,n846gat,n679gat,n1864gat,n1067gat,I1617,n178gat,n736gat,I2316,n1564gat,n2332gat,n721gat,n1328gat,n1004gat,n730gat,I3483,I420,I3168,n2857gat,n2778gat,n2818gat,n1968gat,n2011gat,n2800gat,n940gat,n1015gat,n46gat,n2975gat,n639gat,n60gat,I2213,n1384gat,n2033gat,n2876gat,n265gat,n459gat,I4122,n286gat,I4642,n2626gat,n1530gat,n2405gat,n1725gat,I2403,I4657,n2121gat,n999gat,n1681gat,n1206gat,I1915,n1500gat,n2220gat,n452gat,n1426gat,I1088,n1098gat,n764gat,n340gat,n2268gat,n2046gat,n156gat,n630gat,n2415gat,n800gat,n828gat,n2791gat,n2988gat,I406,n404gat,n1929gat,n516gat,n1354gat,I4185,I2389,n2385gat,n82gat,n2526gat,I771,I3736,I3016,I4608,I4699,n2580gat,n2421gat,n139gat,n312gat,n529gat,n697gat,n2717gat,n1247gat,n729gat,n2411gat,n1609gat,n1524gat,n1310gat,n397gat,n2915gat,I4157,n2585gat,n2539gat,n976gat,n889gat,n559gat,n291gat,n400gat,I446,n592gat,n2286gat,n1296gat,n596gat,n998gat,n870gat,n2542gat,n3024gat,n1300gat,I572,n1287gat,n2968gat,n47gat,I4392,n2051gat,I2174,n2603gat,n1261gat,I4681,I4696,n2880gat,n2678gat,I4349,n923gat,n1650gat,n277gat,n1781gat,n234gat,n381gat,n1320gat,n832gat,n787gat,I2425,n1399gat,n952gat,n1990gat,n575gat,n806gat,I1891,n1391gat,I3436,n2856gat,n329gat,n1624gat,n2512gat,n439gat,n1092gat,n1677gat,n1513gat,n2012gat,n1433gat,n1692gat,n2543gat,n1022gat,I4594,n1890gat,I683,n1018gat,I3297,I4548,n253gat,n1571gat,n1893gat,n827gat,n1264gat,n2899gat,n1056gat,n2956gat,n1185gat,n490gat,n3044gat,n975gat,I351,n995gat,n1311gat,n1617gat,n477gat,n1397gat,n939gat,n123gat,n938gat,I4711,I1733,n2898gat,n552gat,n221gat,n2704gat,n2510gat,n1861gat,I199,n455gat,n981gat,n1094gat,n2939gat,n2674gat,n2483gat,n2889gat,n526gat,n1969gat,I698,n2712gat,I1305,n249gat,n2993gat,n1647gat,I2926,n1152gat,n2432gat,n1794gat,n142gat,n2015gat,n411gat,n2174gat,n919gat,n440gat,n2216gat,I2720,I2017,n500gat,I3504,I941,I2889,n626gat,I4669,n2582gat,n1754gat,n2725gat,n875gat,n1484gat,n1171gat,I999,n51gat,n3055gat,n1187gat,n2801gat,n699gat,n1955gat,n1566gat,n2692gat,I3558,I2242,I1385,I916,n1250gat,I1464,n68gat,I378,n570gat,n1806gat,n1323gat,n816gat,I2094,n2039gat,n2945gat,n1020gat,n1501gat,n2186gat,n175gat,I1606,n786gat,I1336,n289gat,n2908gat,n813gat,n560gat,n3060gat,n1121gat,I363,n2591gat,n2412gat,I18,n564gat,n2008gat,n2728gat,n860gat,n625gat,I1374,I4795,I3178,n1788gat,n1592gat,n1574gat,I1402,n640gat,n2495gat,n1221gat,n2583gat,n2831gat,n2759gat,n1755gat,I4630,n928gat,n1232gat,n2019gat,n780gat,n594gat,I214,n728gat,n2739gat,n3062gat,I4566,n1897gat,n1757gat,n2392gat,n3036gat,n2397gat,n1234gat,n2153gat,n1560gat,n1726gat,n43gat,n1975gat,n2909gat,n293gat,n2462gat,n371gat,n691gat,n528gat,n688gat,I1360,n2428gat,n1292gat,n1693gat,n1421gat,n2442gat,I384,I672,I1961,n420gat,n2953gat,n2643gat,n2722gat,n1567gat,n850gat,n3039gat,n2594gat,I509,n162gat,n2752gat,n154gat,n633gat,n2576gat,I2032,n245gat,n2711gat,n2047gat,n3021gat,n1504gat,I354,n2840gat,n2398gat,n383gat,n2874gat,n1278gat,n1591gat,n1480gat,n230gat,I4332,n2178gat,I3923,I634,I2268,I4024,I712,n812gat,n2248gat,n953gat,I92,n1738gat,n282gat,n1663gat,I3876,I1472,n2307gat,n196gat,n1922gat,n3058gat,n3035gat,I30,n2206gat,n67gat,I2354,n2210gat,n186gat,n556gat,n353gat,I2832,n1282gat,n246gat,n56gat,I1752,n879gat,n557gat,n2736gat,n2763gat,n638gat,n1103gat,n2554gat,n2811gat,I4389,n244gat,I1416,n2212gat,I3163,n1393gat,I4496,I925,n87gat,n235gat,n1452gat,n1070gat,n942gat,n405gat,n2155gat,n1899gat,n2933gat,n70gat,I1786,n1471gat,n2142gat,n1587gat,I1719,I2281,n2333gat,n1727gat,I3904,n1674gat,n1972gat,n1628gat,n2357gat,I2813,n2023gat,n145gat,I2145,n524gat,n57gat,n1959gat,n150gat,n2605gat,n1212gat,I3801,n1797gat,I253,n1297gat,n872gat,n2154gat,n2683gat,n2960gat,I1538,n55gat,n1759gat,n869gat,n2779gat,n324gat,n506gat,n1255gat,I2225,n2748gat,n1855gat,n1456gat,n969gat,n678gat,n994gat,n693gat,n2670gat,n1743gat,n868gat,n2799gat,n1050gat,n877gat,I4536,n1083gat;
//# 35 inputs
//# 49 outputs
//# 179 D-type flipflops
//# 1775 inverters
//# 1004 gates (0 ANDs + 0 NANDs + 239 ORs + 765 NORs)
//
//
//
  MSFF DFF_0(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n673gat),.DATA(n2897gat));
  MSFF DFF_1(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n398gat),.DATA(n2782gat));
  MSFF DFF_2(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n402gat),.DATA(n2790gat));
  MSFF DFF_3(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n919gat),.DATA(n2670gat));
  MSFF DFF_4(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n846gat),.DATA(n2793gat));
  MSFF DFF_5(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n394gat),.DATA(n2782gat));
  MSFF DFF_6(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n703gat),.DATA(n2790gat));
  MSFF DFF_7(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n722gat),.DATA(n2670gat));
  MSFF DFF_8(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n726gat),.DATA(n2793gat));
  MSFF DFF_9(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2510gat),.DATA(n748gat));
  MSFF DFF_10(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n271gat),.DATA(n2732gat));
  MSFF DFF_11(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n160gat),.DATA(n2776gat));
  MSFF DFF_12(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n337gat),.DATA(n2735gat));
  MSFF DFF_13(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n842gat),.DATA(n2673gat));
  MSFF DFF_14(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n341gat),.DATA(n2779gat));
  MSFF DFF_15(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2522gat),.DATA(n43gat));
  MSFF DFF_16(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2472gat),.DATA(n1620gat));
  MSFF DFF_17(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2319gat),.DATA(n2470gat));
  MSFF DFF_18(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1821gat),.DATA(n1827gat));
  MSFF DFF_19(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1825gat),.DATA(n1827gat));
  MSFF DFF_20(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2029gat),.DATA(n1816gat));
  MSFF DFF_21(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1829gat),.DATA(n2027gat));
  MSFF DFF_22(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n283gat),.DATA(n2732gat));
  MSFF DFF_23(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n165gat),.DATA(n2776gat));
  MSFF DFF_24(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n279gat),.DATA(n2735gat));
  MSFF DFF_25(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1026gat),.DATA(n2673gat));
  MSFF DFF_26(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n275gat),.DATA(n2779gat));
  MSFF DFF_27(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2476gat),.DATA(n55gat));
  MSFF DFF_28(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1068gat),.DATA(n2914gat));
  MSFF DFF_29(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n957gat),.DATA(n2928gat));
  MSFF DFF_30(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n861gat),.DATA(n2927gat));
  MSFF DFF_31(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1294gat),.DATA(n2896gat));
  MSFF DFF_32(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1241gat),.DATA(n2922gat));
  MSFF DFF_33(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1298gat),.DATA(n2897gat));
  MSFF DFF_34(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n865gat),.DATA(n2894gat));
  MSFF DFF_35(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1080gat),.DATA(n2921gat));
  MSFF DFF_36(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1148gat),.DATA(n2895gat));
  MSFF DFF_37(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2468gat),.DATA(n933gat));
  MSFF DFF_38(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n618gat),.DATA(n2790gat));
  MSFF DFF_39(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n491gat),.DATA(n2782gat));
  MSFF DFF_40(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n622gat),.DATA(n2793gat));
  MSFF DFF_41(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n626gat),.DATA(n2670gat));
  MSFF DFF_42(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n834gat),.DATA(n3064gat));
  MSFF DFF_43(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n707gat),.DATA(n3055gat));
  MSFF DFF_44(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n838gat),.DATA(n3063gat));
  MSFF DFF_45(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n830gat),.DATA(n3062gat));
  MSFF DFF_46(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n614gat),.DATA(n3056gat));
  MSFF DFF_47(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2526gat),.DATA(n504gat));
  MSFF DFF_48(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n680gat),.DATA(n2913gat));
  MSFF DFF_49(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n816gat),.DATA(n2920gat));
  MSFF DFF_50(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n580gat),.DATA(n2905gat));
  MSFF DFF_51(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n824gat),.DATA(n3057gat));
  MSFF DFF_52(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n820gat),.DATA(n3059gat));
  MSFF DFF_53(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n883gat),.DATA(n3058gat));
  MSFF DFF_54(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n584gat),.DATA(n2898gat));
  MSFF DFF_55(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n684gat),.DATA(n3060gat));
  MSFF DFF_56(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n699gat),.DATA(n3061gat));
  MSFF DFF_57(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2464gat),.DATA(n567gat));
  MSFF DFF_58(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2399gat),.DATA(n3048gat));
  MSFF DFF_59(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2343gat),.DATA(n3049gat));
  MSFF DFF_60(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2203gat),.DATA(n3051gat));
  MSFF DFF_61(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2562gat),.DATA(n3047gat));
  MSFF DFF_62(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2207gat),.DATA(n3050gat));
  MSFF DFF_63(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2626gat),.DATA(n3040gat));
  MSFF DFF_64(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2490gat),.DATA(n3044gat));
  MSFF DFF_65(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2622gat),.DATA(n3042gat));
  MSFF DFF_66(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2630gat),.DATA(n3037gat));
  MSFF DFF_67(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2543gat),.DATA(n3041gat));
  MSFF DFF_68(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2102gat),.DATA(n1606gat));
  MSFF DFF_69(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1880gat),.DATA(n3052gat));
  MSFF DFF_70(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1763gat),.DATA(n1610gat));
  MSFF DFF_71(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2155gat),.DATA(n1858gat));
  MSFF DFF_72(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1035gat),.DATA(n2918gat));
  MSFF DFF_73(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1121gat),.DATA(n2952gat));
  MSFF DFF_74(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1072gat),.DATA(n2919gat));
  MSFF DFF_75(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1282gat),.DATA(n2910gat));
  MSFF DFF_76(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1226gat),.DATA(n2907gat));
  MSFF DFF_77(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n931gat),.DATA(n2911gat));
  MSFF DFF_78(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1135gat),.DATA(n2912gat));
  MSFF DFF_79(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1045gat),.DATA(n2909gat));
  MSFF DFF_80(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1197gat),.DATA(n2908gat));
  MSFF DFF_81(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2518gat),.DATA(n2971gat));
  MSFF DFF_82(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n667gat),.DATA(n2904gat));
  MSFF DFF_83(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n659gat),.DATA(n2891gat));
  MSFF DFF_84(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n553gat),.DATA(n2903gat));
  MSFF DFF_85(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n777gat),.DATA(n2915gat));
  MSFF DFF_86(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n561gat),.DATA(n2901gat));
  MSFF DFF_87(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n366gat),.DATA(n2890gat));
  MSFF DFF_88(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n322gat),.DATA(n2888gat));
  MSFF DFF_89(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n318gat),.DATA(n2887gat));
  MSFF DFF_90(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n314gat),.DATA(n2886gat));
  MSFF DFF_91(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2599gat),.DATA(n3010gat));
  MSFF DFF_92(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2588gat),.DATA(n3016gat));
  MSFF DFF_93(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2640gat),.DATA(n3054gat));
  MSFF DFF_94(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2658gat),.DATA(n2579gat));
  MSFF DFF_95(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2495gat),.DATA(n3036gat));
  MSFF DFF_96(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2390gat),.DATA(n3034gat));
  MSFF DFF_97(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2270gat),.DATA(n3031gat));
  MSFF DFF_98(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2339gat),.DATA(n3035gat));
  MSFF DFF_99(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2502gat),.DATA(n2646gat));
  MSFF DFF_100(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2634gat),.DATA(n3053gat));
  MSFF DFF_101(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2506gat),.DATA(n2613gat));
  MSFF DFF_102(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1834gat),.DATA(n1625gat));
  MSFF DFF_103(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1767gat),.DATA(n1626gat));
  MSFF DFF_104(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2084gat),.DATA(n1603gat));
  MSFF DFF_105(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2143gat),.DATA(n2541gat));
  MSFF DFF_106(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2061gat),.DATA(n2557gat));
  MSFF DFF_107(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2139gat),.DATA(n2487gat));
  MSFF DFF_108(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1899gat),.DATA(n2532gat));
  MSFF DFF_109(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1850gat),.DATA(n2628gat));
  MSFF DFF_110(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2403gat),.DATA(n2397gat));
  MSFF DFF_111(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2394gat),.DATA(n2341gat));
  MSFF DFF_112(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2440gat),.DATA(n2560gat));
  MSFF DFF_113(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2407gat),.DATA(n2205gat));
  MSFF DFF_114(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2347gat),.DATA(n2201gat));
  MSFF DFF_115(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1389gat),.DATA(n1793gat));
  MSFF DFF_116(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2021gat),.DATA(n1781gat));
  MSFF DFF_117(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1394gat),.DATA(n1516gat));
  MSFF DFF_118(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1496gat),.DATA(n1392gat));
  MSFF DFF_119(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2091gat),.DATA(n1685gat));
  MSFF DFF_120(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1332gat),.DATA(n1565gat));
  MSFF DFF_121(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1740gat),.DATA(n1330gat));
  MSFF DFF_122(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2179gat),.DATA(n1945gat));
  MSFF DFF_123(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2190gat),.DATA(n2268gat));
  MSFF DFF_124(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2135gat),.DATA(n2337gat));
  MSFF DFF_125(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2262gat),.DATA(n2388gat));
  MSFF DFF_126(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2182gat),.DATA(n1836gat));
  MSFF DFF_127(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1433gat),.DATA(n2983gat));
  MSFF DFF_128(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1316gat),.DATA(n1431gat));
  MSFF DFF_129(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1363gat),.DATA(n1314gat));
  MSFF DFF_130(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1312gat),.DATA(n1361gat));
  MSFF DFF_131(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1775gat),.DATA(n1696gat));
  MSFF DFF_132(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1871gat),.DATA(n2009gat));
  MSFF DFF_133(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2592gat),.DATA(n1773gat));
  MSFF DFF_134(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1508gat),.DATA(n1636gat));
  MSFF DFF_135(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1678gat),.DATA(n1712gat));
  MSFF DFF_136(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2309gat),.DATA(n3000gat));
  MSFF DFF_137(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2450gat),.DATA(n2307gat));
  MSFF DFF_138(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2446gat),.DATA(n2661gat));
  MSFF DFF_139(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2095gat),.DATA(n827gat));
  MSFF DFF_140(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2176gat),.DATA(n2093gat));
  MSFF DFF_141(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2169gat),.DATA(n2174gat));
  MSFF DFF_142(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2454gat),.DATA(n2163gat));
  MSFF DFF_143(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2040gat),.DATA(n1777gat));
  MSFF DFF_144(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2044gat),.DATA(n2015gat));
  MSFF DFF_145(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2037gat),.DATA(n2042gat));
  MSFF DFF_146(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2025gat),.DATA(n2017gat));
  MSFF DFF_147(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2099gat),.DATA(n2023gat));
  MSFF DFF_148(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2266gat),.DATA(n2493gat));
  MSFF DFF_149(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2033gat),.DATA(n2035gat));
  MSFF DFF_150(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2110gat),.DATA(n2031gat));
  MSFF DFF_151(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2125gat),.DATA(n2108gat));
  MSFF DFF_152(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2121gat),.DATA(n2123gat));
  MSFF DFF_153(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2117gat),.DATA(n2119gat));
  MSFF DFF_154(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1975gat),.DATA(n2632gat));
  MSFF DFF_155(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2644gat),.DATA(n2638gat));
  MSFF DFF_156(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n156gat),.DATA(n612gat));
  MSFF DFF_157(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n152gat),.DATA(n705gat));
  MSFF DFF_158(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n331gat),.DATA(n822gat));
  MSFF DFF_159(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n388gat),.DATA(n881gat));
  MSFF DFF_160(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n463gat),.DATA(n818gat));
  MSFF DFF_161(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n327gat),.DATA(n682gat));
  MSFF DFF_162(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n384gat),.DATA(n697gat));
  MSFF DFF_163(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n256gat),.DATA(n836gat));
  MSFF DFF_164(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n470gat),.DATA(n828gat));
  MSFF DFF_165(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n148gat),.DATA(n832gat));
  MSFF DFF_166(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2458gat),.DATA(n2590gat));
  MSFF DFF_167(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n2514gat),.DATA(n2456gat));
  MSFF DFF_168(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1771gat),.DATA(n1613gat));
  MSFF DFF_169(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1336gat),.DATA(n1391gat));
  MSFF DFF_170(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1748gat),.DATA(n1927gat));
  MSFF DFF_171(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1675gat),.DATA(n1713gat));
  MSFF DFF_172(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1807gat),.DATA(n1717gat));
  MSFF DFF_173(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1340gat),.DATA(n1567gat));
  MSFF DFF_174(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1456gat),.DATA(n1564gat));
  MSFF DFF_175(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1525gat),.DATA(n1632gat));
  MSFF DFF_176(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1462gat),.DATA(n1915gat));
  MSFF DFF_177(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1596gat),.DATA(n1800gat));
  MSFF DFF_178(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(n1588gat),.DATA(n1593gat));
//
  NOT NOT1_0(.VSS(VSS),.VDD(VDD),.Y(I1),.A(n3088gat));
  NOT NOT1_1(.VSS(VSS),.VDD(VDD),.Y(n2717gat),.A(I1));
  NOT NOT1_2(.VSS(VSS),.VDD(VDD),.Y(n2715gat),.A(n2717gat));
  NOT NOT1_3(.VSS(VSS),.VDD(VDD),.Y(I5),.A(n3087gat));
  NOT NOT1_4(.VSS(VSS),.VDD(VDD),.Y(n2725gat),.A(I5));
  NOT NOT1_5(.VSS(VSS),.VDD(VDD),.Y(n2723gat),.A(n2725gat));
  NOT NOT1_6(.VSS(VSS),.VDD(VDD),.Y(n296gat),.A(n421gat));
  NOT NOT1_7(.VSS(VSS),.VDD(VDD),.Y(I11),.A(n3093gat));
  NOT NOT1_8(.VSS(VSS),.VDD(VDD),.Y(n2768gat),.A(I11));
  NOT NOT1_9(.VSS(VSS),.VDD(VDD),.Y(I14),.A(n2768gat));
  NOT NOT1_10(.VSS(VSS),.VDD(VDD),.Y(n2767gat),.A(I14));
  NOT NOT1_11(.VSS(VSS),.VDD(VDD),.Y(n373gat),.A(n2767gat));
  NOT NOT1_12(.VSS(VSS),.VDD(VDD),.Y(I18),.A(n3072gat));
  NOT NOT1_13(.VSS(VSS),.VDD(VDD),.Y(n2671gat),.A(I18));
  NOT NOT1_14(.VSS(VSS),.VDD(VDD),.Y(n2669gat),.A(n2671gat));
  NOT NOT1_15(.VSS(VSS),.VDD(VDD),.Y(I23),.A(n3081gat));
  NOT NOT1_16(.VSS(VSS),.VDD(VDD),.Y(n2845gat),.A(I23));
  NOT NOT1_17(.VSS(VSS),.VDD(VDD),.Y(n2844gat),.A(n2845gat));
  NOT NOT1_18(.VSS(VSS),.VDD(VDD),.Y(I27),.A(n3095gat));
  NOT NOT1_19(.VSS(VSS),.VDD(VDD),.Y(n2668gat),.A(I27));
  NOT NOT1_20(.VSS(VSS),.VDD(VDD),.Y(I30),.A(n2668gat));
  NOT NOT1_21(.VSS(VSS),.VDD(VDD),.Y(n2667gat),.A(I30));
  NOT NOT1_22(.VSS(VSS),.VDD(VDD),.Y(n856gat),.A(n2667gat));
  NOT NOT1_23(.VSS(VSS),.VDD(VDD),.Y(I44),.A(n673gat));
  NOT NOT1_24(.VSS(VSS),.VDD(VDD),.Y(n672gat),.A(I44));
  NOT NOT1_25(.VSS(VSS),.VDD(VDD),.Y(I47),.A(n3069gat));
  NOT NOT1_26(.VSS(VSS),.VDD(VDD),.Y(n2783gat),.A(I47));
  NOT NOT1_27(.VSS(VSS),.VDD(VDD),.Y(I50),.A(n2783gat));
  NOT NOT1_28(.VSS(VSS),.VDD(VDD),.Y(n2782gat),.A(I50));
  NOT NOT1_29(.VSS(VSS),.VDD(VDD),.Y(n396gat),.A(n398gat));
  NOT NOT1_30(.VSS(VSS),.VDD(VDD),.Y(I62),.A(n3070gat));
  NOT NOT1_31(.VSS(VSS),.VDD(VDD),.Y(n2791gat),.A(I62));
  NOT NOT1_32(.VSS(VSS),.VDD(VDD),.Y(I65),.A(n2791gat));
  NOT NOT1_33(.VSS(VSS),.VDD(VDD),.Y(n2790gat),.A(I65));
  NOT NOT1_34(.VSS(VSS),.VDD(VDD),.Y(I76),.A(n402gat));
  NOT NOT1_35(.VSS(VSS),.VDD(VDD),.Y(n401gat),.A(I76));
  NOT NOT1_36(.VSS(VSS),.VDD(VDD),.Y(n1645gat),.A(n1499gat));
  NOT NOT1_37(.VSS(VSS),.VDD(VDD),.Y(I81),.A(n2671gat));
  NOT NOT1_38(.VSS(VSS),.VDD(VDD),.Y(n2670gat),.A(I81));
  NOT NOT1_39(.VSS(VSS),.VDD(VDD),.Y(I92),.A(n919gat));
  NOT NOT1_40(.VSS(VSS),.VDD(VDD),.Y(n918gat),.A(I92));
  NOT NOT1_41(.VSS(VSS),.VDD(VDD),.Y(n1553gat),.A(n1616gat));
  NOT NOT1_42(.VSS(VSS),.VDD(VDD),.Y(I97),.A(n3071gat));
  NOT NOT1_43(.VSS(VSS),.VDD(VDD),.Y(n2794gat),.A(I97));
  NOT NOT1_44(.VSS(VSS),.VDD(VDD),.Y(I100),.A(n2794gat));
  NOT NOT1_45(.VSS(VSS),.VDD(VDD),.Y(n2793gat),.A(I100));
  NOT NOT1_46(.VSS(VSS),.VDD(VDD),.Y(I111),.A(n846gat));
  NOT NOT1_47(.VSS(VSS),.VDD(VDD),.Y(n845gat),.A(I111));
  NOT NOT1_48(.VSS(VSS),.VDD(VDD),.Y(n1559gat),.A(n1614gat));
  NOT NOT1_49(.VSS(VSS),.VDD(VDD),.Y(n1643gat),.A(n1641gat));
  NOT NOT1_50(.VSS(VSS),.VDD(VDD),.Y(n1651gat),.A(n1642gat));
  NOT NOT1_51(.VSS(VSS),.VDD(VDD),.Y(n1562gat),.A(n1556gat));
  NOT NOT1_52(.VSS(VSS),.VDD(VDD),.Y(n1560gat),.A(n1557gat));
  NOT NOT1_53(.VSS(VSS),.VDD(VDD),.Y(n1640gat),.A(n1639gat));
  NOT NOT1_54(.VSS(VSS),.VDD(VDD),.Y(n1566gat),.A(n1605gat));
  NOT NOT1_55(.VSS(VSS),.VDD(VDD),.Y(n1554gat),.A(n1555gat));
  NOT NOT1_56(.VSS(VSS),.VDD(VDD),.Y(n1722gat),.A(n1558gat));
  NOT NOT1_57(.VSS(VSS),.VDD(VDD),.Y(n392gat),.A(n394gat));
  NOT NOT1_58(.VSS(VSS),.VDD(VDD),.Y(I149),.A(n703gat));
  NOT NOT1_59(.VSS(VSS),.VDD(VDD),.Y(n702gat),.A(I149));
  NOT NOT1_60(.VSS(VSS),.VDD(VDD),.Y(n1319gat),.A(n1256gat));
  NOT NOT1_61(.VSS(VSS),.VDD(VDD),.Y(n720gat),.A(n722gat));
  NOT NOT1_62(.VSS(VSS),.VDD(VDD),.Y(I171),.A(n726gat));
  NOT NOT1_63(.VSS(VSS),.VDD(VDD),.Y(n725gat),.A(I171));
  NOT NOT1_64(.VSS(VSS),.VDD(VDD),.Y(n1447gat),.A(n1117gat));
  NOT NOT1_65(.VSS(VSS),.VDD(VDD),.Y(n1627gat),.A(n1618gat));
  NOT NOT1_66(.VSS(VSS),.VDD(VDD),.Y(I178),.A(n722gat));
  NOT NOT1_67(.VSS(VSS),.VDD(VDD),.Y(n721gat),.A(I178));
  NOT NOT1_68(.VSS(VSS),.VDD(VDD),.Y(n1380gat),.A(n1114gat));
  NOT NOT1_69(.VSS(VSS),.VDD(VDD),.Y(n1628gat),.A(n1621gat));
  NOT NOT1_70(.VSS(VSS),.VDD(VDD),.Y(n701gat),.A(n703gat));
  NOT NOT1_71(.VSS(VSS),.VDD(VDD),.Y(n1446gat),.A(n1318gat));
  NOT NOT1_72(.VSS(VSS),.VDD(VDD),.Y(n1705gat),.A(n1619gat));
  NOT NOT1_73(.VSS(VSS),.VDD(VDD),.Y(n1706gat),.A(n1622gat));
  NOT NOT1_74(.VSS(VSS),.VDD(VDD),.Y(I192),.A(n3083gat));
  NOT NOT1_75(.VSS(VSS),.VDD(VDD),.Y(n2856gat),.A(I192));
  NOT NOT1_76(.VSS(VSS),.VDD(VDD),.Y(n2854gat),.A(n2856gat));
  NOT NOT1_77(.VSS(VSS),.VDD(VDD),.Y(I196),.A(n2854gat));
  NOT NOT1_78(.VSS(VSS),.VDD(VDD),.Y(n1218gat),.A(I196));
  NOT NOT1_79(.VSS(VSS),.VDD(VDD),.Y(I199),.A(n3085gat));
  NOT NOT1_80(.VSS(VSS),.VDD(VDD),.Y(n2861gat),.A(I199));
  NOT NOT1_81(.VSS(VSS),.VDD(VDD),.Y(n2859gat),.A(n2861gat));
  NOT NOT1_82(.VSS(VSS),.VDD(VDD),.Y(I203),.A(n2859gat));
  NOT NOT1_83(.VSS(VSS),.VDD(VDD),.Y(n1219gat),.A(I203));
  NOT NOT1_84(.VSS(VSS),.VDD(VDD),.Y(I206),.A(n3084gat));
  NOT NOT1_85(.VSS(VSS),.VDD(VDD),.Y(n2864gat),.A(I206));
  NOT NOT1_86(.VSS(VSS),.VDD(VDD),.Y(n2862gat),.A(n2864gat));
  NOT NOT1_87(.VSS(VSS),.VDD(VDD),.Y(I210),.A(n2862gat));
  NOT NOT1_88(.VSS(VSS),.VDD(VDD),.Y(n1220gat),.A(I210));
  NOT NOT1_89(.VSS(VSS),.VDD(VDD),.Y(I214),.A(n2861gat));
  NOT NOT1_90(.VSS(VSS),.VDD(VDD),.Y(n2860gat),.A(I214));
  NOT NOT1_91(.VSS(VSS),.VDD(VDD),.Y(I217),.A(n2860gat));
  NOT NOT1_92(.VSS(VSS),.VDD(VDD),.Y(n1221gat),.A(I217));
  NOT NOT1_93(.VSS(VSS),.VDD(VDD),.Y(I220),.A(n2864gat));
  NOT NOT1_94(.VSS(VSS),.VDD(VDD),.Y(n2863gat),.A(I220));
  NOT NOT1_95(.VSS(VSS),.VDD(VDD),.Y(I223),.A(n2863gat));
  NOT NOT1_96(.VSS(VSS),.VDD(VDD),.Y(n1222gat),.A(I223));
  NOT NOT1_97(.VSS(VSS),.VDD(VDD),.Y(I227),.A(n2856gat));
  NOT NOT1_98(.VSS(VSS),.VDD(VDD),.Y(n2855gat),.A(I227));
  NOT NOT1_99(.VSS(VSS),.VDD(VDD),.Y(I230),.A(n2855gat));
  NOT NOT1_100(.VSS(VSS),.VDD(VDD),.Y(n1223gat),.A(I230));
  NOT NOT1_101(.VSS(VSS),.VDD(VDD),.Y(n640gat),.A(n1213gat));
  NOT NOT1_102(.VSS(VSS),.VDD(VDD),.Y(I237),.A(n640gat));
  NOT NOT1_103(.VSS(VSS),.VDD(VDD),.Y(n753gat),.A(I237));
  NOT NOT1_104(.VSS(VSS),.VDD(VDD),.Y(I240),.A(n2717gat));
  NOT NOT1_105(.VSS(VSS),.VDD(VDD),.Y(n2716gat),.A(I240));
  NOT NOT1_106(.VSS(VSS),.VDD(VDD),.Y(I243),.A(n3089gat));
  NOT NOT1_107(.VSS(VSS),.VDD(VDD),.Y(n2869gat),.A(I243));
  NOT NOT1_108(.VSS(VSS),.VDD(VDD),.Y(n2867gat),.A(n2869gat));
  NOT NOT1_109(.VSS(VSS),.VDD(VDD),.Y(I248),.A(n2869gat));
  NOT NOT1_110(.VSS(VSS),.VDD(VDD),.Y(n2868gat),.A(I248));
  NOT NOT1_111(.VSS(VSS),.VDD(VDD),.Y(I253),.A(n2906gat));
  NOT NOT1_112(.VSS(VSS),.VDD(VDD),.Y(n754gat),.A(I253));
  NOT NOT1_113(.VSS(VSS),.VDD(VDD),.Y(I256),.A(n2725gat));
  NOT NOT1_114(.VSS(VSS),.VDD(VDD),.Y(n2724gat),.A(I256));
  NOT NOT1_115(.VSS(VSS),.VDD(VDD),.Y(I259),.A(n3086gat));
  NOT NOT1_116(.VSS(VSS),.VDD(VDD),.Y(n2728gat),.A(I259));
  NOT NOT1_117(.VSS(VSS),.VDD(VDD),.Y(n2726gat),.A(n2728gat));
  NOT NOT1_118(.VSS(VSS),.VDD(VDD),.Y(I264),.A(n2728gat));
  NOT NOT1_119(.VSS(VSS),.VDD(VDD),.Y(n2727gat),.A(I264));
  NOT NOT1_120(.VSS(VSS),.VDD(VDD),.Y(n422gat),.A(n2889gat));
  NOT NOT1_121(.VSS(VSS),.VDD(VDD),.Y(I270),.A(n422gat));
  NOT NOT1_122(.VSS(VSS),.VDD(VDD),.Y(n755gat),.A(I270));
  NOT NOT1_123(.VSS(VSS),.VDD(VDD),.Y(n747gat),.A(n2906gat));
  NOT NOT1_124(.VSS(VSS),.VDD(VDD),.Y(I275),.A(n747gat));
  NOT NOT1_125(.VSS(VSS),.VDD(VDD),.Y(n756gat),.A(I275));
  NOT NOT1_126(.VSS(VSS),.VDD(VDD),.Y(I278),.A(n2889gat));
  NOT NOT1_127(.VSS(VSS),.VDD(VDD),.Y(n757gat),.A(I278));
  NOT NOT1_128(.VSS(VSS),.VDD(VDD),.Y(I282),.A(n1213gat));
  NOT NOT1_129(.VSS(VSS),.VDD(VDD),.Y(n758gat),.A(I282));
  NOT NOT1_130(.VSS(VSS),.VDD(VDD),.Y(n2508gat),.A(n2510gat));
  NOT NOT1_131(.VSS(VSS),.VDD(VDD),.Y(I297),.A(n3065gat));
  NOT NOT1_132(.VSS(VSS),.VDD(VDD),.Y(n2733gat),.A(I297));
  NOT NOT1_133(.VSS(VSS),.VDD(VDD),.Y(I300),.A(n2733gat));
  NOT NOT1_134(.VSS(VSS),.VDD(VDD),.Y(n2732gat),.A(I300));
  NOT NOT1_135(.VSS(VSS),.VDD(VDD),.Y(I311),.A(n271gat));
  NOT NOT1_136(.VSS(VSS),.VDD(VDD),.Y(n270gat),.A(I311));
  NOT NOT1_137(.VSS(VSS),.VDD(VDD),.Y(I314),.A(n270gat));
  NOT NOT1_138(.VSS(VSS),.VDD(VDD),.Y(n263gat),.A(I314));
  NOT NOT1_139(.VSS(VSS),.VDD(VDD),.Y(I317),.A(n3067gat));
  NOT NOT1_140(.VSS(VSS),.VDD(VDD),.Y(n2777gat),.A(I317));
  NOT NOT1_141(.VSS(VSS),.VDD(VDD),.Y(I320),.A(n2777gat));
  NOT NOT1_142(.VSS(VSS),.VDD(VDD),.Y(n2776gat),.A(I320));
  NOT NOT1_143(.VSS(VSS),.VDD(VDD),.Y(I331),.A(n160gat));
  NOT NOT1_144(.VSS(VSS),.VDD(VDD),.Y(n159gat),.A(I331));
  NOT NOT1_145(.VSS(VSS),.VDD(VDD),.Y(I334),.A(n159gat));
  NOT NOT1_146(.VSS(VSS),.VDD(VDD),.Y(n264gat),.A(I334));
  NOT NOT1_147(.VSS(VSS),.VDD(VDD),.Y(I337),.A(n3066gat));
  NOT NOT1_148(.VSS(VSS),.VDD(VDD),.Y(n2736gat),.A(I337));
  NOT NOT1_149(.VSS(VSS),.VDD(VDD),.Y(I340),.A(n2736gat));
  NOT NOT1_150(.VSS(VSS),.VDD(VDD),.Y(n2735gat),.A(I340));
  NOT NOT1_151(.VSS(VSS),.VDD(VDD),.Y(I351),.A(n337gat));
  NOT NOT1_152(.VSS(VSS),.VDD(VDD),.Y(n336gat),.A(I351));
  NOT NOT1_153(.VSS(VSS),.VDD(VDD),.Y(I354),.A(n336gat));
  NOT NOT1_154(.VSS(VSS),.VDD(VDD),.Y(n265gat),.A(I354));
  NOT NOT1_155(.VSS(VSS),.VDD(VDD),.Y(n158gat),.A(n160gat));
  NOT NOT1_156(.VSS(VSS),.VDD(VDD),.Y(I359),.A(n158gat));
  NOT NOT1_157(.VSS(VSS),.VDD(VDD),.Y(n266gat),.A(I359));
  NOT NOT1_158(.VSS(VSS),.VDD(VDD),.Y(n335gat),.A(n337gat));
  NOT NOT1_159(.VSS(VSS),.VDD(VDD),.Y(I363),.A(n335gat));
  NOT NOT1_160(.VSS(VSS),.VDD(VDD),.Y(n267gat),.A(I363));
  NOT NOT1_161(.VSS(VSS),.VDD(VDD),.Y(n269gat),.A(n271gat));
  NOT NOT1_162(.VSS(VSS),.VDD(VDD),.Y(I368),.A(n269gat));
  NOT NOT1_163(.VSS(VSS),.VDD(VDD),.Y(n268gat),.A(I368));
  NOT NOT1_164(.VSS(VSS),.VDD(VDD),.Y(n41gat),.A(n258gat));
  NOT NOT1_165(.VSS(VSS),.VDD(VDD),.Y(I375),.A(n41gat));
  NOT NOT1_166(.VSS(VSS),.VDD(VDD),.Y(n48gat),.A(I375));
  NOT NOT1_167(.VSS(VSS),.VDD(VDD),.Y(I378),.A(n725gat));
  NOT NOT1_168(.VSS(VSS),.VDD(VDD),.Y(n1018gat),.A(I378));
  NOT NOT1_169(.VSS(VSS),.VDD(VDD),.Y(I381),.A(n3073gat));
  NOT NOT1_170(.VSS(VSS),.VDD(VDD),.Y(n2674gat),.A(I381));
  NOT NOT1_171(.VSS(VSS),.VDD(VDD),.Y(I384),.A(n2674gat));
  NOT NOT1_172(.VSS(VSS),.VDD(VDD),.Y(n2673gat),.A(I384));
  NOT NOT1_173(.VSS(VSS),.VDD(VDD),.Y(I395),.A(n842gat));
  NOT NOT1_174(.VSS(VSS),.VDD(VDD),.Y(n841gat),.A(I395));
  NOT NOT1_175(.VSS(VSS),.VDD(VDD),.Y(I398),.A(n841gat));
  NOT NOT1_176(.VSS(VSS),.VDD(VDD),.Y(n1019gat),.A(I398));
  NOT NOT1_177(.VSS(VSS),.VDD(VDD),.Y(I401),.A(n721gat));
  NOT NOT1_178(.VSS(VSS),.VDD(VDD),.Y(n1020gat),.A(I401));
  NOT NOT1_179(.VSS(VSS),.VDD(VDD),.Y(n840gat),.A(n842gat));
  NOT NOT1_180(.VSS(VSS),.VDD(VDD),.Y(I406),.A(n840gat));
  NOT NOT1_181(.VSS(VSS),.VDD(VDD),.Y(n1021gat),.A(I406));
  NOT NOT1_182(.VSS(VSS),.VDD(VDD),.Y(I409),.A(n720gat));
  NOT NOT1_183(.VSS(VSS),.VDD(VDD),.Y(n1022gat),.A(I409));
  NOT NOT1_184(.VSS(VSS),.VDD(VDD),.Y(n724gat),.A(n726gat));
  NOT NOT1_185(.VSS(VSS),.VDD(VDD),.Y(I414),.A(n724gat));
  NOT NOT1_186(.VSS(VSS),.VDD(VDD),.Y(n1023gat),.A(I414));
  NOT NOT1_187(.VSS(VSS),.VDD(VDD),.Y(I420),.A(n1013gat));
  NOT NOT1_188(.VSS(VSS),.VDD(VDD),.Y(n49gat),.A(I420));
  NOT NOT1_189(.VSS(VSS),.VDD(VDD),.Y(I423),.A(n3068gat));
  NOT NOT1_190(.VSS(VSS),.VDD(VDD),.Y(n2780gat),.A(I423));
  NOT NOT1_191(.VSS(VSS),.VDD(VDD),.Y(I426),.A(n2780gat));
  NOT NOT1_192(.VSS(VSS),.VDD(VDD),.Y(n2779gat),.A(I426));
  NOT NOT1_193(.VSS(VSS),.VDD(VDD),.Y(I437),.A(n341gat));
  NOT NOT1_194(.VSS(VSS),.VDD(VDD),.Y(n340gat),.A(I437));
  NOT NOT1_195(.VSS(VSS),.VDD(VDD),.Y(I440),.A(n340gat));
  NOT NOT1_196(.VSS(VSS),.VDD(VDD),.Y(n480gat),.A(I440));
  NOT NOT1_197(.VSS(VSS),.VDD(VDD),.Y(I443),.A(n702gat));
  NOT NOT1_198(.VSS(VSS),.VDD(VDD),.Y(n481gat),.A(I443));
  NOT NOT1_199(.VSS(VSS),.VDD(VDD),.Y(I446),.A(n394gat));
  NOT NOT1_200(.VSS(VSS),.VDD(VDD),.Y(n393gat),.A(I446));
  NOT NOT1_201(.VSS(VSS),.VDD(VDD),.Y(I449),.A(n393gat));
  NOT NOT1_202(.VSS(VSS),.VDD(VDD),.Y(n482gat),.A(I449));
  NOT NOT1_203(.VSS(VSS),.VDD(VDD),.Y(I453),.A(n701gat));
  NOT NOT1_204(.VSS(VSS),.VDD(VDD),.Y(n483gat),.A(I453));
  NOT NOT1_205(.VSS(VSS),.VDD(VDD),.Y(I456),.A(n392gat));
  NOT NOT1_206(.VSS(VSS),.VDD(VDD),.Y(n484gat),.A(I456));
  NOT NOT1_207(.VSS(VSS),.VDD(VDD),.Y(n339gat),.A(n341gat));
  NOT NOT1_208(.VSS(VSS),.VDD(VDD),.Y(I461),.A(n339gat));
  NOT NOT1_209(.VSS(VSS),.VDD(VDD),.Y(n485gat),.A(I461));
  NOT NOT1_210(.VSS(VSS),.VDD(VDD),.Y(n42gat),.A(n475gat));
  NOT NOT1_211(.VSS(VSS),.VDD(VDD),.Y(I468),.A(n42gat));
  NOT NOT1_212(.VSS(VSS),.VDD(VDD),.Y(n50gat),.A(I468));
  NOT NOT1_213(.VSS(VSS),.VDD(VDD),.Y(n162gat),.A(n1013gat));
  NOT NOT1_214(.VSS(VSS),.VDD(VDD),.Y(I473),.A(n162gat));
  NOT NOT1_215(.VSS(VSS),.VDD(VDD),.Y(n51gat),.A(I473));
  NOT NOT1_216(.VSS(VSS),.VDD(VDD),.Y(I476),.A(n475gat));
  NOT NOT1_217(.VSS(VSS),.VDD(VDD),.Y(n52gat),.A(I476));
  NOT NOT1_218(.VSS(VSS),.VDD(VDD),.Y(I480),.A(n258gat));
  NOT NOT1_219(.VSS(VSS),.VDD(VDD),.Y(n53gat),.A(I480));
  NOT NOT1_220(.VSS(VSS),.VDD(VDD),.Y(n2520gat),.A(n2522gat));
  NOT NOT1_221(.VSS(VSS),.VDD(VDD),.Y(n1448gat),.A(n1376gat));
  NOT NOT1_222(.VSS(VSS),.VDD(VDD),.Y(n1701gat),.A(n1617gat));
  NOT NOT1_223(.VSS(VSS),.VDD(VDD),.Y(n1379gat),.A(n1377gat));
  NOT NOT1_224(.VSS(VSS),.VDD(VDD),.Y(n1615gat),.A(n1624gat));
  NOT NOT1_225(.VSS(VSS),.VDD(VDD),.Y(n1500gat),.A(n1113gat));
  NOT NOT1_226(.VSS(VSS),.VDD(VDD),.Y(n1503gat),.A(n1501gat));
  NOT NOT1_227(.VSS(VSS),.VDD(VDD),.Y(n1779gat),.A(n1623gat));
  NOT NOT1_228(.VSS(VSS),.VDD(VDD),.Y(I509),.A(n3099gat));
  NOT NOT1_229(.VSS(VSS),.VDD(VDD),.Y(n2730gat),.A(I509));
  NOT NOT1_230(.VSS(VSS),.VDD(VDD),.Y(I512),.A(n2730gat));
  NOT NOT1_231(.VSS(VSS),.VDD(VDD),.Y(n2729gat),.A(I512));
  NOT NOT1_232(.VSS(VSS),.VDD(VDD),.Y(n2470gat),.A(n2472gat));
  NOT NOT1_233(.VSS(VSS),.VDD(VDD),.Y(n2317gat),.A(n2319gat));
  NOT NOT1_234(.VSS(VSS),.VDD(VDD),.Y(n1819gat),.A(n1821gat));
  NOT NOT1_235(.VSS(VSS),.VDD(VDD),.Y(n1823gat),.A(n1825gat));
  NOT NOT1_236(.VSS(VSS),.VDD(VDD),.Y(n1816gat),.A(n1817gat));
  NOT NOT1_237(.VSS(VSS),.VDD(VDD),.Y(n2027gat),.A(n2029gat));
  NOT NOT1_238(.VSS(VSS),.VDD(VDD),.Y(I572),.A(n1829gat));
  NOT NOT1_239(.VSS(VSS),.VDD(VDD),.Y(n1828gat),.A(I572));
  NOT NOT1_240(.VSS(VSS),.VDD(VDD),.Y(I576),.A(n3100gat));
  NOT NOT1_241(.VSS(VSS),.VDD(VDD),.Y(n2851gat),.A(I576));
  NOT NOT1_242(.VSS(VSS),.VDD(VDD),.Y(I579),.A(n2851gat));
  NOT NOT1_243(.VSS(VSS),.VDD(VDD),.Y(n2850gat),.A(I579));
  NOT NOT1_244(.VSS(VSS),.VDD(VDD),.Y(I583),.A(n2786gat));
  NOT NOT1_245(.VSS(VSS),.VDD(VDD),.Y(n2785gat),.A(I583));
  NOT NOT1_246(.VSS(VSS),.VDD(VDD),.Y(n92gat),.A(n2785gat));
  NOT NOT1_247(.VSS(VSS),.VDD(VDD),.Y(n637gat),.A(n529gat));
  NOT NOT1_248(.VSS(VSS),.VDD(VDD),.Y(n293gat),.A(n361gat));
  NOT NOT1_249(.VSS(VSS),.VDD(VDD),.Y(I591),.A(n3094gat));
  NOT NOT1_250(.VSS(VSS),.VDD(VDD),.Y(n2722gat),.A(I591));
  NOT NOT1_251(.VSS(VSS),.VDD(VDD),.Y(I594),.A(n2722gat));
  NOT NOT1_252(.VSS(VSS),.VDD(VDD),.Y(n2721gat),.A(I594));
  NOT NOT1_253(.VSS(VSS),.VDD(VDD),.Y(n297gat),.A(n2721gat));
  NOT NOT1_254(.VSS(VSS),.VDD(VDD),.Y(I606),.A(n283gat));
  NOT NOT1_255(.VSS(VSS),.VDD(VDD),.Y(n282gat),.A(I606));
  NOT NOT1_256(.VSS(VSS),.VDD(VDD),.Y(I609),.A(n282gat));
  NOT NOT1_257(.VSS(VSS),.VDD(VDD),.Y(n172gat),.A(I609));
  NOT NOT1_258(.VSS(VSS),.VDD(VDD),.Y(I620),.A(n165gat));
  NOT NOT1_259(.VSS(VSS),.VDD(VDD),.Y(n164gat),.A(I620));
  NOT NOT1_260(.VSS(VSS),.VDD(VDD),.Y(I623),.A(n164gat));
  NOT NOT1_261(.VSS(VSS),.VDD(VDD),.Y(n173gat),.A(I623));
  NOT NOT1_262(.VSS(VSS),.VDD(VDD),.Y(I634),.A(n279gat));
  NOT NOT1_263(.VSS(VSS),.VDD(VDD),.Y(n278gat),.A(I634));
  NOT NOT1_264(.VSS(VSS),.VDD(VDD),.Y(I637),.A(n278gat));
  NOT NOT1_265(.VSS(VSS),.VDD(VDD),.Y(n174gat),.A(I637));
  NOT NOT1_266(.VSS(VSS),.VDD(VDD),.Y(n163gat),.A(n165gat));
  NOT NOT1_267(.VSS(VSS),.VDD(VDD),.Y(I642),.A(n163gat));
  NOT NOT1_268(.VSS(VSS),.VDD(VDD),.Y(n175gat),.A(I642));
  NOT NOT1_269(.VSS(VSS),.VDD(VDD),.Y(n277gat),.A(n279gat));
  NOT NOT1_270(.VSS(VSS),.VDD(VDD),.Y(I646),.A(n277gat));
  NOT NOT1_271(.VSS(VSS),.VDD(VDD),.Y(n176gat),.A(I646));
  NOT NOT1_272(.VSS(VSS),.VDD(VDD),.Y(n281gat),.A(n283gat));
  NOT NOT1_273(.VSS(VSS),.VDD(VDD),.Y(I651),.A(n281gat));
  NOT NOT1_274(.VSS(VSS),.VDD(VDD),.Y(n177gat),.A(I651));
  NOT NOT1_275(.VSS(VSS),.VDD(VDD),.Y(n54gat),.A(n167gat));
  NOT NOT1_276(.VSS(VSS),.VDD(VDD),.Y(I658),.A(n54gat));
  NOT NOT1_277(.VSS(VSS),.VDD(VDD),.Y(n60gat),.A(I658));
  NOT NOT1_278(.VSS(VSS),.VDD(VDD),.Y(I661),.A(n845gat));
  NOT NOT1_279(.VSS(VSS),.VDD(VDD),.Y(n911gat),.A(I661));
  NOT NOT1_280(.VSS(VSS),.VDD(VDD),.Y(I672),.A(n1026gat));
  NOT NOT1_281(.VSS(VSS),.VDD(VDD),.Y(n1025gat),.A(I672));
  NOT NOT1_282(.VSS(VSS),.VDD(VDD),.Y(I675),.A(n1025gat));
  NOT NOT1_283(.VSS(VSS),.VDD(VDD),.Y(n912gat),.A(I675));
  NOT NOT1_284(.VSS(VSS),.VDD(VDD),.Y(I678),.A(n918gat));
  NOT NOT1_285(.VSS(VSS),.VDD(VDD),.Y(n913gat),.A(I678));
  NOT NOT1_286(.VSS(VSS),.VDD(VDD),.Y(n1024gat),.A(n1026gat));
  NOT NOT1_287(.VSS(VSS),.VDD(VDD),.Y(I683),.A(n1024gat));
  NOT NOT1_288(.VSS(VSS),.VDD(VDD),.Y(n914gat),.A(I683));
  NOT NOT1_289(.VSS(VSS),.VDD(VDD),.Y(n917gat),.A(n919gat));
  NOT NOT1_290(.VSS(VSS),.VDD(VDD),.Y(I687),.A(n917gat));
  NOT NOT1_291(.VSS(VSS),.VDD(VDD),.Y(n915gat),.A(I687));
  NOT NOT1_292(.VSS(VSS),.VDD(VDD),.Y(n844gat),.A(n846gat));
  NOT NOT1_293(.VSS(VSS),.VDD(VDD),.Y(I692),.A(n844gat));
  NOT NOT1_294(.VSS(VSS),.VDD(VDD),.Y(n916gat),.A(I692));
  NOT NOT1_295(.VSS(VSS),.VDD(VDD),.Y(I698),.A(n906gat));
  NOT NOT1_296(.VSS(VSS),.VDD(VDD),.Y(n61gat),.A(I698));
  NOT NOT1_297(.VSS(VSS),.VDD(VDD),.Y(I709),.A(n275gat));
  NOT NOT1_298(.VSS(VSS),.VDD(VDD),.Y(n274gat),.A(I709));
  NOT NOT1_299(.VSS(VSS),.VDD(VDD),.Y(I712),.A(n274gat));
  NOT NOT1_300(.VSS(VSS),.VDD(VDD),.Y(n348gat),.A(I712));
  NOT NOT1_301(.VSS(VSS),.VDD(VDD),.Y(I715),.A(n401gat));
  NOT NOT1_302(.VSS(VSS),.VDD(VDD),.Y(n349gat),.A(I715));
  NOT NOT1_303(.VSS(VSS),.VDD(VDD),.Y(I718),.A(n398gat));
  NOT NOT1_304(.VSS(VSS),.VDD(VDD),.Y(n397gat),.A(I718));
  NOT NOT1_305(.VSS(VSS),.VDD(VDD),.Y(I721),.A(n397gat));
  NOT NOT1_306(.VSS(VSS),.VDD(VDD),.Y(n350gat),.A(I721));
  NOT NOT1_307(.VSS(VSS),.VDD(VDD),.Y(n400gat),.A(n402gat));
  NOT NOT1_308(.VSS(VSS),.VDD(VDD),.Y(I726),.A(n400gat));
  NOT NOT1_309(.VSS(VSS),.VDD(VDD),.Y(n351gat),.A(I726));
  NOT NOT1_310(.VSS(VSS),.VDD(VDD),.Y(I729),.A(n396gat));
  NOT NOT1_311(.VSS(VSS),.VDD(VDD),.Y(n352gat),.A(I729));
  NOT NOT1_312(.VSS(VSS),.VDD(VDD),.Y(n273gat),.A(n275gat));
  NOT NOT1_313(.VSS(VSS),.VDD(VDD),.Y(I734),.A(n273gat));
  NOT NOT1_314(.VSS(VSS),.VDD(VDD),.Y(n353gat),.A(I734));
  NOT NOT1_315(.VSS(VSS),.VDD(VDD),.Y(n178gat),.A(n343gat));
  NOT NOT1_316(.VSS(VSS),.VDD(VDD),.Y(I741),.A(n178gat));
  NOT NOT1_317(.VSS(VSS),.VDD(VDD),.Y(n62gat),.A(I741));
  NOT NOT1_318(.VSS(VSS),.VDD(VDD),.Y(n66gat),.A(n906gat));
  NOT NOT1_319(.VSS(VSS),.VDD(VDD),.Y(I746),.A(n66gat));
  NOT NOT1_320(.VSS(VSS),.VDD(VDD),.Y(n63gat),.A(I746));
  NOT NOT1_321(.VSS(VSS),.VDD(VDD),.Y(I749),.A(n343gat));
  NOT NOT1_322(.VSS(VSS),.VDD(VDD),.Y(n64gat),.A(I749));
  NOT NOT1_323(.VSS(VSS),.VDD(VDD),.Y(I753),.A(n167gat));
  NOT NOT1_324(.VSS(VSS),.VDD(VDD),.Y(n65gat),.A(I753));
  NOT NOT1_325(.VSS(VSS),.VDD(VDD),.Y(n2474gat),.A(n2476gat));
  NOT NOT1_326(.VSS(VSS),.VDD(VDD),.Y(I768),.A(n3090gat));
  NOT NOT1_327(.VSS(VSS),.VDD(VDD),.Y(n2832gat),.A(I768));
  NOT NOT1_328(.VSS(VSS),.VDD(VDD),.Y(I771),.A(n2832gat));
  NOT NOT1_329(.VSS(VSS),.VDD(VDD),.Y(n2831gat),.A(I771));
  NOT NOT1_330(.VSS(VSS),.VDD(VDD),.Y(n2731gat),.A(n2733gat));
  NOT NOT1_331(.VSS(VSS),.VDD(VDD),.Y(I776),.A(n3074gat));
  NOT NOT1_332(.VSS(VSS),.VDD(VDD),.Y(n2719gat),.A(I776));
  NOT NOT1_333(.VSS(VSS),.VDD(VDD),.Y(n2718gat),.A(n2719gat));
  NOT NOT1_334(.VSS(VSS),.VDD(VDD),.Y(I790),.A(n1068gat));
  NOT NOT1_335(.VSS(VSS),.VDD(VDD),.Y(n1067gat),.A(I790));
  NOT NOT1_336(.VSS(VSS),.VDD(VDD),.Y(I793),.A(n1067gat));
  NOT NOT1_337(.VSS(VSS),.VDD(VDD),.Y(n949gat),.A(I793));
  NOT NOT1_338(.VSS(VSS),.VDD(VDD),.Y(I796),.A(n3076gat));
  NOT NOT1_339(.VSS(VSS),.VDD(VDD),.Y(n2839gat),.A(I796));
  NOT NOT1_340(.VSS(VSS),.VDD(VDD),.Y(n2838gat),.A(n2839gat));
  NOT NOT1_341(.VSS(VSS),.VDD(VDD),.Y(n2775gat),.A(n2777gat));
  NOT NOT1_342(.VSS(VSS),.VDD(VDD),.Y(I812),.A(n957gat));
  NOT NOT1_343(.VSS(VSS),.VDD(VDD),.Y(n956gat),.A(I812));
  NOT NOT1_344(.VSS(VSS),.VDD(VDD),.Y(I815),.A(n956gat));
  NOT NOT1_345(.VSS(VSS),.VDD(VDD),.Y(n950gat),.A(I815));
  NOT NOT1_346(.VSS(VSS),.VDD(VDD),.Y(I818),.A(n3075gat));
  NOT NOT1_347(.VSS(VSS),.VDD(VDD),.Y(n2712gat),.A(I818));
  NOT NOT1_348(.VSS(VSS),.VDD(VDD),.Y(n2711gat),.A(n2712gat));
  NOT NOT1_349(.VSS(VSS),.VDD(VDD),.Y(n2734gat),.A(n2736gat));
  NOT NOT1_350(.VSS(VSS),.VDD(VDD),.Y(I834),.A(n861gat));
  NOT NOT1_351(.VSS(VSS),.VDD(VDD),.Y(n860gat),.A(I834));
  NOT NOT1_352(.VSS(VSS),.VDD(VDD),.Y(I837),.A(n860gat));
  NOT NOT1_353(.VSS(VSS),.VDD(VDD),.Y(n951gat),.A(I837));
  NOT NOT1_354(.VSS(VSS),.VDD(VDD),.Y(n955gat),.A(n957gat));
  NOT NOT1_355(.VSS(VSS),.VDD(VDD),.Y(I842),.A(n955gat));
  NOT NOT1_356(.VSS(VSS),.VDD(VDD),.Y(n952gat),.A(I842));
  NOT NOT1_357(.VSS(VSS),.VDD(VDD),.Y(n859gat),.A(n861gat));
  NOT NOT1_358(.VSS(VSS),.VDD(VDD),.Y(I846),.A(n859gat));
  NOT NOT1_359(.VSS(VSS),.VDD(VDD),.Y(n953gat),.A(I846));
  NOT NOT1_360(.VSS(VSS),.VDD(VDD),.Y(n1066gat),.A(n1068gat));
  NOT NOT1_361(.VSS(VSS),.VDD(VDD),.Y(I851),.A(n1066gat));
  NOT NOT1_362(.VSS(VSS),.VDD(VDD),.Y(n954gat),.A(I851));
  NOT NOT1_363(.VSS(VSS),.VDD(VDD),.Y(n857gat),.A(n944gat));
  NOT NOT1_364(.VSS(VSS),.VDD(VDD),.Y(I858),.A(n857gat));
  NOT NOT1_365(.VSS(VSS),.VDD(VDD),.Y(n938gat),.A(I858));
  NOT NOT1_366(.VSS(VSS),.VDD(VDD),.Y(n2792gat),.A(n2794gat));
  NOT NOT1_367(.VSS(VSS),.VDD(VDD),.Y(I863),.A(n3080gat));
  NOT NOT1_368(.VSS(VSS),.VDD(VDD),.Y(n2847gat),.A(I863));
  NOT NOT1_369(.VSS(VSS),.VDD(VDD),.Y(n2846gat),.A(n2847gat));
  NOT NOT1_370(.VSS(VSS),.VDD(VDD),.Y(I877),.A(n1294gat));
  NOT NOT1_371(.VSS(VSS),.VDD(VDD),.Y(n1293gat),.A(I877));
  NOT NOT1_372(.VSS(VSS),.VDD(VDD),.Y(I880),.A(n1293gat));
  NOT NOT1_373(.VSS(VSS),.VDD(VDD),.Y(n1233gat),.A(I880));
  NOT NOT1_374(.VSS(VSS),.VDD(VDD),.Y(n2672gat),.A(n2674gat));
  NOT NOT1_375(.VSS(VSS),.VDD(VDD),.Y(I885),.A(n3082gat));
  NOT NOT1_376(.VSS(VSS),.VDD(VDD),.Y(n2853gat),.A(I885));
  NOT NOT1_377(.VSS(VSS),.VDD(VDD),.Y(n2852gat),.A(n2853gat));
  NOT NOT1_378(.VSS(VSS),.VDD(VDD),.Y(I899),.A(n1241gat));
  NOT NOT1_379(.VSS(VSS),.VDD(VDD),.Y(n1240gat),.A(I899));
  NOT NOT1_380(.VSS(VSS),.VDD(VDD),.Y(I902),.A(n1240gat));
  NOT NOT1_381(.VSS(VSS),.VDD(VDD),.Y(n1234gat),.A(I902));
  NOT NOT1_382(.VSS(VSS),.VDD(VDD),.Y(I913),.A(n1298gat));
  NOT NOT1_383(.VSS(VSS),.VDD(VDD),.Y(n1297gat),.A(I913));
  NOT NOT1_384(.VSS(VSS),.VDD(VDD),.Y(I916),.A(n1297gat));
  NOT NOT1_385(.VSS(VSS),.VDD(VDD),.Y(n1235gat),.A(I916));
  NOT NOT1_386(.VSS(VSS),.VDD(VDD),.Y(n1239gat),.A(n1241gat));
  NOT NOT1_387(.VSS(VSS),.VDD(VDD),.Y(I921),.A(n1239gat));
  NOT NOT1_388(.VSS(VSS),.VDD(VDD),.Y(n1236gat),.A(I921));
  NOT NOT1_389(.VSS(VSS),.VDD(VDD),.Y(n1296gat),.A(n1298gat));
  NOT NOT1_390(.VSS(VSS),.VDD(VDD),.Y(I925),.A(n1296gat));
  NOT NOT1_391(.VSS(VSS),.VDD(VDD),.Y(n1237gat),.A(I925));
  NOT NOT1_392(.VSS(VSS),.VDD(VDD),.Y(n1292gat),.A(n1294gat));
  NOT NOT1_393(.VSS(VSS),.VDD(VDD),.Y(I930),.A(n1292gat));
  NOT NOT1_394(.VSS(VSS),.VDD(VDD),.Y(n1238gat),.A(I930));
  NOT NOT1_395(.VSS(VSS),.VDD(VDD),.Y(I936),.A(n1228gat));
  NOT NOT1_396(.VSS(VSS),.VDD(VDD),.Y(n939gat),.A(I936));
  NOT NOT1_397(.VSS(VSS),.VDD(VDD),.Y(n2778gat),.A(n2780gat));
  NOT NOT1_398(.VSS(VSS),.VDD(VDD),.Y(I941),.A(n3077gat));
  NOT NOT1_399(.VSS(VSS),.VDD(VDD),.Y(n2837gat),.A(I941));
  NOT NOT1_400(.VSS(VSS),.VDD(VDD),.Y(n2836gat),.A(n2837gat));
  NOT NOT1_401(.VSS(VSS),.VDD(VDD),.Y(I955),.A(n865gat));
  NOT NOT1_402(.VSS(VSS),.VDD(VDD),.Y(n864gat),.A(I955));
  NOT NOT1_403(.VSS(VSS),.VDD(VDD),.Y(I958),.A(n864gat));
  NOT NOT1_404(.VSS(VSS),.VDD(VDD),.Y(n1055gat),.A(I958));
  NOT NOT1_405(.VSS(VSS),.VDD(VDD),.Y(n2789gat),.A(n2791gat));
  NOT NOT1_406(.VSS(VSS),.VDD(VDD),.Y(I963),.A(n3079gat));
  NOT NOT1_407(.VSS(VSS),.VDD(VDD),.Y(n2841gat),.A(I963));
  NOT NOT1_408(.VSS(VSS),.VDD(VDD),.Y(n2840gat),.A(n2841gat));
  NOT NOT1_409(.VSS(VSS),.VDD(VDD),.Y(I977),.A(n1080gat));
  NOT NOT1_410(.VSS(VSS),.VDD(VDD),.Y(n1079gat),.A(I977));
  NOT NOT1_411(.VSS(VSS),.VDD(VDD),.Y(I980),.A(n1079gat));
  NOT NOT1_412(.VSS(VSS),.VDD(VDD),.Y(n1056gat),.A(I980));
  NOT NOT1_413(.VSS(VSS),.VDD(VDD),.Y(n2781gat),.A(n2783gat));
  NOT NOT1_414(.VSS(VSS),.VDD(VDD),.Y(I985),.A(n3078gat));
  NOT NOT1_415(.VSS(VSS),.VDD(VDD),.Y(n2843gat),.A(I985));
  NOT NOT1_416(.VSS(VSS),.VDD(VDD),.Y(n2842gat),.A(n2843gat));
  NOT NOT1_417(.VSS(VSS),.VDD(VDD),.Y(I999),.A(n1148gat));
  NOT NOT1_418(.VSS(VSS),.VDD(VDD),.Y(n1147gat),.A(I999));
  NOT NOT1_419(.VSS(VSS),.VDD(VDD),.Y(I1002),.A(n1147gat));
  NOT NOT1_420(.VSS(VSS),.VDD(VDD),.Y(n1057gat),.A(I1002));
  NOT NOT1_421(.VSS(VSS),.VDD(VDD),.Y(n1078gat),.A(n1080gat));
  NOT NOT1_422(.VSS(VSS),.VDD(VDD),.Y(I1007),.A(n1078gat));
  NOT NOT1_423(.VSS(VSS),.VDD(VDD),.Y(n1058gat),.A(I1007));
  NOT NOT1_424(.VSS(VSS),.VDD(VDD),.Y(n1146gat),.A(n1148gat));
  NOT NOT1_425(.VSS(VSS),.VDD(VDD),.Y(I1011),.A(n1146gat));
  NOT NOT1_426(.VSS(VSS),.VDD(VDD),.Y(n1059gat),.A(I1011));
  NOT NOT1_427(.VSS(VSS),.VDD(VDD),.Y(n863gat),.A(n865gat));
  NOT NOT1_428(.VSS(VSS),.VDD(VDD),.Y(I1016),.A(n863gat));
  NOT NOT1_429(.VSS(VSS),.VDD(VDD),.Y(n1060gat),.A(I1016));
  NOT NOT1_430(.VSS(VSS),.VDD(VDD),.Y(n928gat),.A(n1050gat));
  NOT NOT1_431(.VSS(VSS),.VDD(VDD),.Y(I1023),.A(n928gat));
  NOT NOT1_432(.VSS(VSS),.VDD(VDD),.Y(n940gat),.A(I1023));
  NOT NOT1_433(.VSS(VSS),.VDD(VDD),.Y(n858gat),.A(n1228gat));
  NOT NOT1_434(.VSS(VSS),.VDD(VDD),.Y(I1028),.A(n858gat));
  NOT NOT1_435(.VSS(VSS),.VDD(VDD),.Y(n941gat),.A(I1028));
  NOT NOT1_436(.VSS(VSS),.VDD(VDD),.Y(I1031),.A(n1050gat));
  NOT NOT1_437(.VSS(VSS),.VDD(VDD),.Y(n942gat),.A(I1031));
  NOT NOT1_438(.VSS(VSS),.VDD(VDD),.Y(I1035),.A(n944gat));
  NOT NOT1_439(.VSS(VSS),.VDD(VDD),.Y(n943gat),.A(I1035));
  NOT NOT1_440(.VSS(VSS),.VDD(VDD),.Y(n2466gat),.A(n2468gat));
  NOT NOT1_441(.VSS(VSS),.VDD(VDD),.Y(n2720gat),.A(n2722gat));
  NOT NOT1_442(.VSS(VSS),.VDD(VDD),.Y(n740gat),.A(n2667gat));
  NOT NOT1_443(.VSS(VSS),.VDD(VDD),.Y(n2784gat),.A(n2786gat));
  NOT NOT1_444(.VSS(VSS),.VDD(VDD),.Y(n743gat),.A(n746gat));
  NOT NOT1_445(.VSS(VSS),.VDD(VDD),.Y(n294gat),.A(n360gat));
  NOT NOT1_446(.VSS(VSS),.VDD(VDD),.Y(n374gat),.A(n2767gat));
  NOT NOT1_447(.VSS(VSS),.VDD(VDD),.Y(n616gat),.A(n618gat));
  NOT NOT1_448(.VSS(VSS),.VDD(VDD),.Y(I1067),.A(n616gat));
  NOT NOT1_449(.VSS(VSS),.VDD(VDD),.Y(n501gat),.A(I1067));
  NOT NOT1_450(.VSS(VSS),.VDD(VDD),.Y(n489gat),.A(n491gat));
  NOT NOT1_451(.VSS(VSS),.VDD(VDD),.Y(I1079),.A(n489gat));
  NOT NOT1_452(.VSS(VSS),.VDD(VDD),.Y(n502gat),.A(I1079));
  NOT NOT1_453(.VSS(VSS),.VDD(VDD),.Y(I1082),.A(n618gat));
  NOT NOT1_454(.VSS(VSS),.VDD(VDD),.Y(n617gat),.A(I1082));
  NOT NOT1_455(.VSS(VSS),.VDD(VDD),.Y(I1085),.A(n617gat));
  NOT NOT1_456(.VSS(VSS),.VDD(VDD),.Y(n499gat),.A(I1085));
  NOT NOT1_457(.VSS(VSS),.VDD(VDD),.Y(I1088),.A(n491gat));
  NOT NOT1_458(.VSS(VSS),.VDD(VDD),.Y(n490gat),.A(I1088));
  NOT NOT1_459(.VSS(VSS),.VDD(VDD),.Y(I1091),.A(n490gat));
  NOT NOT1_460(.VSS(VSS),.VDD(VDD),.Y(n500gat),.A(I1091));
  NOT NOT1_461(.VSS(VSS),.VDD(VDD),.Y(n620gat),.A(n622gat));
  NOT NOT1_462(.VSS(VSS),.VDD(VDD),.Y(I1103),.A(n620gat));
  NOT NOT1_463(.VSS(VSS),.VDD(VDD),.Y(n738gat),.A(I1103));
  NOT NOT1_464(.VSS(VSS),.VDD(VDD),.Y(n624gat),.A(n626gat));
  NOT NOT1_465(.VSS(VSS),.VDD(VDD),.Y(I1115),.A(n624gat));
  NOT NOT1_466(.VSS(VSS),.VDD(VDD),.Y(n737gat),.A(I1115));
  NOT NOT1_467(.VSS(VSS),.VDD(VDD),.Y(I1118),.A(n622gat));
  NOT NOT1_468(.VSS(VSS),.VDD(VDD),.Y(n621gat),.A(I1118));
  NOT NOT1_469(.VSS(VSS),.VDD(VDD),.Y(I1121),.A(n621gat));
  NOT NOT1_470(.VSS(VSS),.VDD(VDD),.Y(n733gat),.A(I1121));
  NOT NOT1_471(.VSS(VSS),.VDD(VDD),.Y(I1124),.A(n626gat));
  NOT NOT1_472(.VSS(VSS),.VDD(VDD),.Y(n625gat),.A(I1124));
  NOT NOT1_473(.VSS(VSS),.VDD(VDD),.Y(I1127),.A(n625gat));
  NOT NOT1_474(.VSS(VSS),.VDD(VDD),.Y(n735gat),.A(I1127));
  NOT NOT1_475(.VSS(VSS),.VDD(VDD),.Y(I1138),.A(n834gat));
  NOT NOT1_476(.VSS(VSS),.VDD(VDD),.Y(n833gat),.A(I1138));
  NOT NOT1_477(.VSS(VSS),.VDD(VDD),.Y(I1141),.A(n833gat));
  NOT NOT1_478(.VSS(VSS),.VDD(VDD),.Y(n714gat),.A(I1141));
  NOT NOT1_479(.VSS(VSS),.VDD(VDD),.Y(I1152),.A(n707gat));
  NOT NOT1_480(.VSS(VSS),.VDD(VDD),.Y(n706gat),.A(I1152));
  NOT NOT1_481(.VSS(VSS),.VDD(VDD),.Y(I1155),.A(n706gat));
  NOT NOT1_482(.VSS(VSS),.VDD(VDD),.Y(n715gat),.A(I1155));
  NOT NOT1_483(.VSS(VSS),.VDD(VDD),.Y(I1166),.A(n838gat));
  NOT NOT1_484(.VSS(VSS),.VDD(VDD),.Y(n837gat),.A(I1166));
  NOT NOT1_485(.VSS(VSS),.VDD(VDD),.Y(I1169),.A(n837gat));
  NOT NOT1_486(.VSS(VSS),.VDD(VDD),.Y(n716gat),.A(I1169));
  NOT NOT1_487(.VSS(VSS),.VDD(VDD),.Y(n705gat),.A(n707gat));
  NOT NOT1_488(.VSS(VSS),.VDD(VDD),.Y(I1174),.A(n705gat));
  NOT NOT1_489(.VSS(VSS),.VDD(VDD),.Y(n717gat),.A(I1174));
  NOT NOT1_490(.VSS(VSS),.VDD(VDD),.Y(n836gat),.A(n838gat));
  NOT NOT1_491(.VSS(VSS),.VDD(VDD),.Y(I1178),.A(n836gat));
  NOT NOT1_492(.VSS(VSS),.VDD(VDD),.Y(n718gat),.A(I1178));
  NOT NOT1_493(.VSS(VSS),.VDD(VDD),.Y(n832gat),.A(n834gat));
  NOT NOT1_494(.VSS(VSS),.VDD(VDD),.Y(I1183),.A(n832gat));
  NOT NOT1_495(.VSS(VSS),.VDD(VDD),.Y(n719gat),.A(I1183));
  NOT NOT1_496(.VSS(VSS),.VDD(VDD),.Y(n515gat),.A(n709gat));
  NOT NOT1_497(.VSS(VSS),.VDD(VDD),.Y(I1190),.A(n515gat));
  NOT NOT1_498(.VSS(VSS),.VDD(VDD),.Y(n509gat),.A(I1190));
  NOT NOT1_499(.VSS(VSS),.VDD(VDD),.Y(I1201),.A(n830gat));
  NOT NOT1_500(.VSS(VSS),.VDD(VDD),.Y(n829gat),.A(I1201));
  NOT NOT1_501(.VSS(VSS),.VDD(VDD),.Y(I1204),.A(n829gat));
  NOT NOT1_502(.VSS(VSS),.VDD(VDD),.Y(n734gat),.A(I1204));
  NOT NOT1_503(.VSS(VSS),.VDD(VDD),.Y(n828gat),.A(n830gat));
  NOT NOT1_504(.VSS(VSS),.VDD(VDD),.Y(I1209),.A(n828gat));
  NOT NOT1_505(.VSS(VSS),.VDD(VDD),.Y(n736gat),.A(I1209));
  NOT NOT1_506(.VSS(VSS),.VDD(VDD),.Y(I1216),.A(n728gat));
  NOT NOT1_507(.VSS(VSS),.VDD(VDD),.Y(n510gat),.A(I1216));
  NOT NOT1_508(.VSS(VSS),.VDD(VDD),.Y(I1227),.A(n614gat));
  NOT NOT1_509(.VSS(VSS),.VDD(VDD),.Y(n613gat),.A(I1227));
  NOT NOT1_510(.VSS(VSS),.VDD(VDD),.Y(I1230),.A(n613gat));
  NOT NOT1_511(.VSS(VSS),.VDD(VDD),.Y(n498gat),.A(I1230));
  NOT NOT1_512(.VSS(VSS),.VDD(VDD),.Y(n612gat),.A(n614gat));
  NOT NOT1_513(.VSS(VSS),.VDD(VDD),.Y(I1236),.A(n612gat));
  NOT NOT1_514(.VSS(VSS),.VDD(VDD),.Y(n503gat),.A(I1236));
  NOT NOT1_515(.VSS(VSS),.VDD(VDD),.Y(n404gat),.A(n493gat));
  NOT NOT1_516(.VSS(VSS),.VDD(VDD),.Y(I1243),.A(n404gat));
  NOT NOT1_517(.VSS(VSS),.VDD(VDD),.Y(n511gat),.A(I1243));
  NOT NOT1_518(.VSS(VSS),.VDD(VDD),.Y(n405gat),.A(n728gat));
  NOT NOT1_519(.VSS(VSS),.VDD(VDD),.Y(I1248),.A(n405gat));
  NOT NOT1_520(.VSS(VSS),.VDD(VDD),.Y(n512gat),.A(I1248));
  NOT NOT1_521(.VSS(VSS),.VDD(VDD),.Y(I1251),.A(n493gat));
  NOT NOT1_522(.VSS(VSS),.VDD(VDD),.Y(n513gat),.A(I1251));
  NOT NOT1_523(.VSS(VSS),.VDD(VDD),.Y(I1255),.A(n709gat));
  NOT NOT1_524(.VSS(VSS),.VDD(VDD),.Y(n514gat),.A(I1255));
  NOT NOT1_525(.VSS(VSS),.VDD(VDD),.Y(n2524gat),.A(n2526gat));
  NOT NOT1_526(.VSS(VSS),.VDD(VDD),.Y(n17gat),.A(n564gat));
  NOT NOT1_527(.VSS(VSS),.VDD(VDD),.Y(n79gat),.A(n86gat));
  NOT NOT1_528(.VSS(VSS),.VDD(VDD),.Y(n219gat),.A(n78gat));
  NOT NOT1_529(.VSS(VSS),.VDD(VDD),.Y(n563gat),.A(I1278));
  NOT NOT1_530(.VSS(VSS),.VDD(VDD),.Y(n289gat),.A(n563gat));
  NOT NOT1_531(.VSS(VSS),.VDD(VDD),.Y(n179gat),.A(n287gat));
  NOT NOT1_532(.VSS(VSS),.VDD(VDD),.Y(n188gat),.A(n288gat));
  NOT NOT1_533(.VSS(VSS),.VDD(VDD),.Y(n72gat),.A(n181gat));
  NOT NOT1_534(.VSS(VSS),.VDD(VDD),.Y(n111gat),.A(n182gat));
  NOT NOT1_535(.VSS(VSS),.VDD(VDD),.Y(I1302),.A(n680gat));
  NOT NOT1_536(.VSS(VSS),.VDD(VDD),.Y(n679gat),.A(I1302));
  NOT NOT1_537(.VSS(VSS),.VDD(VDD),.Y(I1305),.A(n679gat));
  NOT NOT1_538(.VSS(VSS),.VDD(VDD),.Y(n808gat),.A(I1305));
  NOT NOT1_539(.VSS(VSS),.VDD(VDD),.Y(I1319),.A(n816gat));
  NOT NOT1_540(.VSS(VSS),.VDD(VDD),.Y(n815gat),.A(I1319));
  NOT NOT1_541(.VSS(VSS),.VDD(VDD),.Y(I1322),.A(n815gat));
  NOT NOT1_542(.VSS(VSS),.VDD(VDD),.Y(n809gat),.A(I1322));
  NOT NOT1_543(.VSS(VSS),.VDD(VDD),.Y(I1336),.A(n580gat));
  NOT NOT1_544(.VSS(VSS),.VDD(VDD),.Y(n579gat),.A(I1336));
  NOT NOT1_545(.VSS(VSS),.VDD(VDD),.Y(I1339),.A(n579gat));
  NOT NOT1_546(.VSS(VSS),.VDD(VDD),.Y(n810gat),.A(I1339));
  NOT NOT1_547(.VSS(VSS),.VDD(VDD),.Y(n814gat),.A(n816gat));
  NOT NOT1_548(.VSS(VSS),.VDD(VDD),.Y(I1344),.A(n814gat));
  NOT NOT1_549(.VSS(VSS),.VDD(VDD),.Y(n811gat),.A(I1344));
  NOT NOT1_550(.VSS(VSS),.VDD(VDD),.Y(n578gat),.A(n580gat));
  NOT NOT1_551(.VSS(VSS),.VDD(VDD),.Y(I1348),.A(n578gat));
  NOT NOT1_552(.VSS(VSS),.VDD(VDD),.Y(n812gat),.A(I1348));
  NOT NOT1_553(.VSS(VSS),.VDD(VDD),.Y(n678gat),.A(n680gat));
  NOT NOT1_554(.VSS(VSS),.VDD(VDD),.Y(I1353),.A(n678gat));
  NOT NOT1_555(.VSS(VSS),.VDD(VDD),.Y(n813gat),.A(I1353));
  NOT NOT1_556(.VSS(VSS),.VDD(VDD),.Y(n677gat),.A(n803gat));
  NOT NOT1_557(.VSS(VSS),.VDD(VDD),.Y(I1360),.A(n677gat));
  NOT NOT1_558(.VSS(VSS),.VDD(VDD),.Y(n572gat),.A(I1360));
  NOT NOT1_559(.VSS(VSS),.VDD(VDD),.Y(I1371),.A(n824gat));
  NOT NOT1_560(.VSS(VSS),.VDD(VDD),.Y(n823gat),.A(I1371));
  NOT NOT1_561(.VSS(VSS),.VDD(VDD),.Y(I1374),.A(n823gat));
  NOT NOT1_562(.VSS(VSS),.VDD(VDD),.Y(n591gat),.A(I1374));
  NOT NOT1_563(.VSS(VSS),.VDD(VDD),.Y(I1385),.A(n820gat));
  NOT NOT1_564(.VSS(VSS),.VDD(VDD),.Y(n819gat),.A(I1385));
  NOT NOT1_565(.VSS(VSS),.VDD(VDD),.Y(I1388),.A(n819gat));
  NOT NOT1_566(.VSS(VSS),.VDD(VDD),.Y(n592gat),.A(I1388));
  NOT NOT1_567(.VSS(VSS),.VDD(VDD),.Y(I1399),.A(n883gat));
  NOT NOT1_568(.VSS(VSS),.VDD(VDD),.Y(n882gat),.A(I1399));
  NOT NOT1_569(.VSS(VSS),.VDD(VDD),.Y(I1402),.A(n882gat));
  NOT NOT1_570(.VSS(VSS),.VDD(VDD),.Y(n593gat),.A(I1402));
  NOT NOT1_571(.VSS(VSS),.VDD(VDD),.Y(n818gat),.A(n820gat));
  NOT NOT1_572(.VSS(VSS),.VDD(VDD),.Y(I1407),.A(n818gat));
  NOT NOT1_573(.VSS(VSS),.VDD(VDD),.Y(n594gat),.A(I1407));
  NOT NOT1_574(.VSS(VSS),.VDD(VDD),.Y(n881gat),.A(n883gat));
  NOT NOT1_575(.VSS(VSS),.VDD(VDD),.Y(I1411),.A(n881gat));
  NOT NOT1_576(.VSS(VSS),.VDD(VDD),.Y(n595gat),.A(I1411));
  NOT NOT1_577(.VSS(VSS),.VDD(VDD),.Y(n822gat),.A(n824gat));
  NOT NOT1_578(.VSS(VSS),.VDD(VDD),.Y(I1416),.A(n822gat));
  NOT NOT1_579(.VSS(VSS),.VDD(VDD),.Y(n596gat),.A(I1416));
  NOT NOT1_580(.VSS(VSS),.VDD(VDD),.Y(I1422),.A(n586gat));
  NOT NOT1_581(.VSS(VSS),.VDD(VDD),.Y(n573gat),.A(I1422));
  NOT NOT1_582(.VSS(VSS),.VDD(VDD),.Y(I1436),.A(n584gat));
  NOT NOT1_583(.VSS(VSS),.VDD(VDD),.Y(n583gat),.A(I1436));
  NOT NOT1_584(.VSS(VSS),.VDD(VDD),.Y(I1439),.A(n583gat));
  NOT NOT1_585(.VSS(VSS),.VDD(VDD),.Y(n691gat),.A(I1439));
  NOT NOT1_586(.VSS(VSS),.VDD(VDD),.Y(I1450),.A(n684gat));
  NOT NOT1_587(.VSS(VSS),.VDD(VDD),.Y(n683gat),.A(I1450));
  NOT NOT1_588(.VSS(VSS),.VDD(VDD),.Y(I1453),.A(n683gat));
  NOT NOT1_589(.VSS(VSS),.VDD(VDD),.Y(n692gat),.A(I1453));
  NOT NOT1_590(.VSS(VSS),.VDD(VDD),.Y(I1464),.A(n699gat));
  NOT NOT1_591(.VSS(VSS),.VDD(VDD),.Y(n698gat),.A(I1464));
  NOT NOT1_592(.VSS(VSS),.VDD(VDD),.Y(I1467),.A(n698gat));
  NOT NOT1_593(.VSS(VSS),.VDD(VDD),.Y(n693gat),.A(I1467));
  NOT NOT1_594(.VSS(VSS),.VDD(VDD),.Y(n682gat),.A(n684gat));
  NOT NOT1_595(.VSS(VSS),.VDD(VDD),.Y(I1472),.A(n682gat));
  NOT NOT1_596(.VSS(VSS),.VDD(VDD),.Y(n694gat),.A(I1472));
  NOT NOT1_597(.VSS(VSS),.VDD(VDD),.Y(n697gat),.A(n699gat));
  NOT NOT1_598(.VSS(VSS),.VDD(VDD),.Y(I1476),.A(n697gat));
  NOT NOT1_599(.VSS(VSS),.VDD(VDD),.Y(n695gat),.A(I1476));
  NOT NOT1_600(.VSS(VSS),.VDD(VDD),.Y(n582gat),.A(n584gat));
  NOT NOT1_601(.VSS(VSS),.VDD(VDD),.Y(I1481),.A(n582gat));
  NOT NOT1_602(.VSS(VSS),.VDD(VDD),.Y(n696gat),.A(I1481));
  NOT NOT1_603(.VSS(VSS),.VDD(VDD),.Y(n456gat),.A(n686gat));
  NOT NOT1_604(.VSS(VSS),.VDD(VDD),.Y(I1488),.A(n456gat));
  NOT NOT1_605(.VSS(VSS),.VDD(VDD),.Y(n574gat),.A(I1488));
  NOT NOT1_606(.VSS(VSS),.VDD(VDD),.Y(n565gat),.A(n586gat));
  NOT NOT1_607(.VSS(VSS),.VDD(VDD),.Y(I1493),.A(n565gat));
  NOT NOT1_608(.VSS(VSS),.VDD(VDD),.Y(n575gat),.A(I1493));
  NOT NOT1_609(.VSS(VSS),.VDD(VDD),.Y(I1496),.A(n686gat));
  NOT NOT1_610(.VSS(VSS),.VDD(VDD),.Y(n576gat),.A(I1496));
  NOT NOT1_611(.VSS(VSS),.VDD(VDD),.Y(I1500),.A(n803gat));
  NOT NOT1_612(.VSS(VSS),.VDD(VDD),.Y(n577gat),.A(I1500));
  NOT NOT1_613(.VSS(VSS),.VDD(VDD),.Y(n2462gat),.A(n2464gat));
  NOT NOT1_614(.VSS(VSS),.VDD(VDD),.Y(n2665gat),.A(I1516));
  NOT NOT1_615(.VSS(VSS),.VDD(VDD),.Y(n2596gat),.A(n2665gat));
  NOT NOT1_616(.VSS(VSS),.VDD(VDD),.Y(n189gat),.A(n286gat));
  NOT NOT1_617(.VSS(VSS),.VDD(VDD),.Y(n194gat),.A(n187gat));
  NOT NOT1_618(.VSS(VSS),.VDD(VDD),.Y(n21gat),.A(n15gat));
  NOT NOT1_619(.VSS(VSS),.VDD(VDD),.Y(I1538),.A(n2399gat));
  NOT NOT1_620(.VSS(VSS),.VDD(VDD),.Y(n2398gat),.A(I1538));
  NOT NOT1_621(.VSS(VSS),.VDD(VDD),.Y(n2353gat),.A(n2398gat));
  NOT NOT1_622(.VSS(VSS),.VDD(VDD),.Y(I1550),.A(n2343gat));
  NOT NOT1_623(.VSS(VSS),.VDD(VDD),.Y(n2342gat),.A(I1550));
  NOT NOT1_624(.VSS(VSS),.VDD(VDD),.Y(n2284gat),.A(n2342gat));
  NOT NOT1_625(.VSS(VSS),.VDD(VDD),.Y(n2201gat),.A(n2203gat));
  NOT NOT1_626(.VSS(VSS),.VDD(VDD),.Y(n2354gat),.A(n2201gat));
  NOT NOT1_627(.VSS(VSS),.VDD(VDD),.Y(n2560gat),.A(n2562gat));
  NOT NOT1_628(.VSS(VSS),.VDD(VDD),.Y(n2356gat),.A(n2560gat));
  NOT NOT1_629(.VSS(VSS),.VDD(VDD),.Y(n2205gat),.A(n2207gat));
  NOT NOT1_630(.VSS(VSS),.VDD(VDD),.Y(n2214gat),.A(n2205gat));
  NOT NOT1_631(.VSS(VSS),.VDD(VDD),.Y(n2286gat),.A(I1585));
  NOT NOT1_632(.VSS(VSS),.VDD(VDD),.Y(n2624gat),.A(n2626gat));
  NOT NOT1_633(.VSS(VSS),.VDD(VDD),.Y(I1606),.A(n2490gat));
  NOT NOT1_634(.VSS(VSS),.VDD(VDD),.Y(n2489gat),.A(I1606));
  NOT NOT1_635(.VSS(VSS),.VDD(VDD),.Y(I1617),.A(n2622gat));
  NOT NOT1_636(.VSS(VSS),.VDD(VDD),.Y(n2621gat),.A(I1617));
  NOT NOT1_637(.VSS(VSS),.VDD(VDD),.Y(n2533gat),.A(n2534gat));
  NOT NOT1_638(.VSS(VSS),.VDD(VDD),.Y(I1630),.A(n2630gat));
  NOT NOT1_639(.VSS(VSS),.VDD(VDD),.Y(n2629gat),.A(I1630));
  NOT NOT1_640(.VSS(VSS),.VDD(VDD),.Y(n2486gat),.A(n2629gat));
  NOT NOT1_641(.VSS(VSS),.VDD(VDD),.Y(n2541gat),.A(n2543gat));
  NOT NOT1_642(.VSS(VSS),.VDD(VDD),.Y(n2429gat),.A(n2541gat));
  NOT NOT1_643(.VSS(VSS),.VDD(VDD),.Y(n2432gat),.A(n2430gat));
  NOT NOT1_644(.VSS(VSS),.VDD(VDD),.Y(I1655),.A(n2102gat));
  NOT NOT1_645(.VSS(VSS),.VDD(VDD),.Y(n2101gat),.A(I1655));
  NOT NOT1_646(.VSS(VSS),.VDD(VDD),.Y(n1693gat),.A(n2101gat));
  NOT NOT1_647(.VSS(VSS),.VDD(VDD),.Y(I1667),.A(n1880gat));
  NOT NOT1_648(.VSS(VSS),.VDD(VDD),.Y(n1879gat),.A(I1667));
  NOT NOT1_649(.VSS(VSS),.VDD(VDD),.Y(n1698gat),.A(n1934gat));
  NOT NOT1_650(.VSS(VSS),.VDD(VDD),.Y(n1543gat),.A(n1606gat));
  NOT NOT1_651(.VSS(VSS),.VDD(VDD),.Y(I1683),.A(n1763gat));
  NOT NOT1_652(.VSS(VSS),.VDD(VDD),.Y(n1762gat),.A(I1683));
  NOT NOT1_653(.VSS(VSS),.VDD(VDD),.Y(n1673gat),.A(n2989gat));
  NOT NOT1_654(.VSS(VSS),.VDD(VDD),.Y(n1858gat),.A(n1673gat));
  NOT NOT1_655(.VSS(VSS),.VDD(VDD),.Y(I1698),.A(n2155gat));
  NOT NOT1_656(.VSS(VSS),.VDD(VDD),.Y(n2154gat),.A(I1698));
  NOT NOT1_657(.VSS(VSS),.VDD(VDD),.Y(n2488gat),.A(n2490gat));
  NOT NOT1_658(.VSS(VSS),.VDD(VDD),.Y(I1703),.A(n2626gat));
  NOT NOT1_659(.VSS(VSS),.VDD(VDD),.Y(n2625gat),.A(I1703));
  NOT NOT1_660(.VSS(VSS),.VDD(VDD),.Y(n2530gat),.A(n2531gat));
  NOT NOT1_661(.VSS(VSS),.VDD(VDD),.Y(I1708),.A(n2543gat));
  NOT NOT1_662(.VSS(VSS),.VDD(VDD),.Y(n2542gat),.A(I1708));
  NOT NOT1_663(.VSS(VSS),.VDD(VDD),.Y(n2482gat),.A(n2542gat));
  NOT NOT1_664(.VSS(VSS),.VDD(VDD),.Y(n2426gat),.A(n2480gat));
  NOT NOT1_665(.VSS(VSS),.VDD(VDD),.Y(n2153gat),.A(n2155gat));
  NOT NOT1_666(.VSS(VSS),.VDD(VDD),.Y(n2341gat),.A(n2343gat));
  NOT NOT1_667(.VSS(VSS),.VDD(VDD),.Y(n2355gat),.A(n2341gat));
  NOT NOT1_668(.VSS(VSS),.VDD(VDD),.Y(I1719),.A(n2562gat));
  NOT NOT1_669(.VSS(VSS),.VDD(VDD),.Y(n2561gat),.A(I1719));
  NOT NOT1_670(.VSS(VSS),.VDD(VDD),.Y(n2443gat),.A(n2561gat));
  NOT NOT1_671(.VSS(VSS),.VDD(VDD),.Y(n2289gat),.A(I1724));
  NOT NOT1_672(.VSS(VSS),.VDD(VDD),.Y(n2148gat),.A(I1734));
  NOT NOT1_673(.VSS(VSS),.VDD(VDD),.Y(n855gat),.A(n2148gat));
  NOT NOT1_674(.VSS(VSS),.VDD(VDD),.Y(n759gat),.A(n855gat));
  NOT NOT1_675(.VSS(VSS),.VDD(VDD),.Y(I1749),.A(n1035gat));
  NOT NOT1_676(.VSS(VSS),.VDD(VDD),.Y(n1034gat),.A(I1749));
  NOT NOT1_677(.VSS(VSS),.VDD(VDD),.Y(I1752),.A(n1034gat));
  NOT NOT1_678(.VSS(VSS),.VDD(VDD),.Y(n1189gat),.A(I1752));
  NOT NOT1_679(.VSS(VSS),.VDD(VDD),.Y(n1075gat),.A(n855gat));
  NOT NOT1_680(.VSS(VSS),.VDD(VDD),.Y(I1766),.A(n1121gat));
  NOT NOT1_681(.VSS(VSS),.VDD(VDD),.Y(n1120gat),.A(I1766));
  NOT NOT1_682(.VSS(VSS),.VDD(VDD),.Y(I1769),.A(n1120gat));
  NOT NOT1_683(.VSS(VSS),.VDD(VDD),.Y(n1190gat),.A(I1769));
  NOT NOT1_684(.VSS(VSS),.VDD(VDD),.Y(n760gat),.A(n855gat));
  NOT NOT1_685(.VSS(VSS),.VDD(VDD),.Y(I1783),.A(n1072gat));
  NOT NOT1_686(.VSS(VSS),.VDD(VDD),.Y(n1071gat),.A(I1783));
  NOT NOT1_687(.VSS(VSS),.VDD(VDD),.Y(I1786),.A(n1071gat));
  NOT NOT1_688(.VSS(VSS),.VDD(VDD),.Y(n1191gat),.A(I1786));
  NOT NOT1_689(.VSS(VSS),.VDD(VDD),.Y(n1119gat),.A(n1121gat));
  NOT NOT1_690(.VSS(VSS),.VDD(VDD),.Y(I1791),.A(n1119gat));
  NOT NOT1_691(.VSS(VSS),.VDD(VDD),.Y(n1192gat),.A(I1791));
  NOT NOT1_692(.VSS(VSS),.VDD(VDD),.Y(n1070gat),.A(n1072gat));
  NOT NOT1_693(.VSS(VSS),.VDD(VDD),.Y(I1795),.A(n1070gat));
  NOT NOT1_694(.VSS(VSS),.VDD(VDD),.Y(n1193gat),.A(I1795));
  NOT NOT1_695(.VSS(VSS),.VDD(VDD),.Y(n1033gat),.A(n1035gat));
  NOT NOT1_696(.VSS(VSS),.VDD(VDD),.Y(I1800),.A(n1033gat));
  NOT NOT1_697(.VSS(VSS),.VDD(VDD),.Y(n1194gat),.A(I1800));
  NOT NOT1_698(.VSS(VSS),.VDD(VDD),.Y(n1183gat),.A(n1184gat));
  NOT NOT1_699(.VSS(VSS),.VDD(VDD),.Y(I1807),.A(n1183gat));
  NOT NOT1_700(.VSS(VSS),.VDD(VDD),.Y(n1274gat),.A(I1807));
  NOT NOT1_701(.VSS(VSS),.VDD(VDD),.Y(n644gat),.A(n855gat));
  NOT NOT1_702(.VSS(VSS),.VDD(VDD),.Y(n1280gat),.A(n1282gat));
  NOT NOT1_703(.VSS(VSS),.VDD(VDD),.Y(n641gat),.A(n855gat));
  NOT NOT1_704(.VSS(VSS),.VDD(VDD),.Y(I1833),.A(n1226gat));
  NOT NOT1_705(.VSS(VSS),.VDD(VDD),.Y(n1225gat),.A(I1833));
  NOT NOT1_706(.VSS(VSS),.VDD(VDD),.Y(I1837),.A(n1282gat));
  NOT NOT1_707(.VSS(VSS),.VDD(VDD),.Y(n1281gat),.A(I1837));
  NOT NOT1_708(.VSS(VSS),.VDD(VDD),.Y(n1224gat),.A(n1226gat));
  NOT NOT1_709(.VSS(VSS),.VDD(VDD),.Y(I1843),.A(n2970gat));
  NOT NOT1_710(.VSS(VSS),.VDD(VDD),.Y(n1275gat),.A(I1843));
  NOT NOT1_711(.VSS(VSS),.VDD(VDD),.Y(n761gat),.A(n855gat));
  NOT NOT1_712(.VSS(VSS),.VDD(VDD),.Y(I1857),.A(n931gat));
  NOT NOT1_713(.VSS(VSS),.VDD(VDD),.Y(n930gat),.A(I1857));
  NOT NOT1_714(.VSS(VSS),.VDD(VDD),.Y(I1860),.A(n930gat));
  NOT NOT1_715(.VSS(VSS),.VDD(VDD),.Y(n1206gat),.A(I1860));
  NOT NOT1_716(.VSS(VSS),.VDD(VDD),.Y(n762gat),.A(n855gat));
  NOT NOT1_717(.VSS(VSS),.VDD(VDD),.Y(I1874),.A(n1135gat));
  NOT NOT1_718(.VSS(VSS),.VDD(VDD),.Y(n1134gat),.A(I1874));
  NOT NOT1_719(.VSS(VSS),.VDD(VDD),.Y(I1877),.A(n1134gat));
  NOT NOT1_720(.VSS(VSS),.VDD(VDD),.Y(n1207gat),.A(I1877));
  NOT NOT1_721(.VSS(VSS),.VDD(VDD),.Y(n643gat),.A(n855gat));
  NOT NOT1_722(.VSS(VSS),.VDD(VDD),.Y(I1891),.A(n1045gat));
  NOT NOT1_723(.VSS(VSS),.VDD(VDD),.Y(n1044gat),.A(I1891));
  NOT NOT1_724(.VSS(VSS),.VDD(VDD),.Y(I1894),.A(n1044gat));
  NOT NOT1_725(.VSS(VSS),.VDD(VDD),.Y(n1208gat),.A(I1894));
  NOT NOT1_726(.VSS(VSS),.VDD(VDD),.Y(n1133gat),.A(n1135gat));
  NOT NOT1_727(.VSS(VSS),.VDD(VDD),.Y(I1899),.A(n1133gat));
  NOT NOT1_728(.VSS(VSS),.VDD(VDD),.Y(n1209gat),.A(I1899));
  NOT NOT1_729(.VSS(VSS),.VDD(VDD),.Y(n1043gat),.A(n1045gat));
  NOT NOT1_730(.VSS(VSS),.VDD(VDD),.Y(I1903),.A(n1043gat));
  NOT NOT1_731(.VSS(VSS),.VDD(VDD),.Y(n1210gat),.A(I1903));
  NOT NOT1_732(.VSS(VSS),.VDD(VDD),.Y(n929gat),.A(n931gat));
  NOT NOT1_733(.VSS(VSS),.VDD(VDD),.Y(I1908),.A(n929gat));
  NOT NOT1_734(.VSS(VSS),.VDD(VDD),.Y(n1211gat),.A(I1908));
  NOT NOT1_735(.VSS(VSS),.VDD(VDD),.Y(n1268gat),.A(n1201gat));
  NOT NOT1_736(.VSS(VSS),.VDD(VDD),.Y(I1915),.A(n1268gat));
  NOT NOT1_737(.VSS(VSS),.VDD(VDD),.Y(n1276gat),.A(I1915));
  NOT NOT1_738(.VSS(VSS),.VDD(VDD),.Y(n1329gat),.A(n2970gat));
  NOT NOT1_739(.VSS(VSS),.VDD(VDD),.Y(I1920),.A(n1329gat));
  NOT NOT1_740(.VSS(VSS),.VDD(VDD),.Y(n1277gat),.A(I1920));
  NOT NOT1_741(.VSS(VSS),.VDD(VDD),.Y(I1923),.A(n1201gat));
  NOT NOT1_742(.VSS(VSS),.VDD(VDD),.Y(n1278gat),.A(I1923));
  NOT NOT1_743(.VSS(VSS),.VDD(VDD),.Y(I1927),.A(n1184gat));
  NOT NOT1_744(.VSS(VSS),.VDD(VDD),.Y(n1279gat),.A(I1927));
  NOT NOT1_745(.VSS(VSS),.VDD(VDD),.Y(n1284gat),.A(n1269gat));
  NOT NOT1_746(.VSS(VSS),.VDD(VDD),.Y(n642gat),.A(n855gat));
  NOT NOT1_747(.VSS(VSS),.VDD(VDD),.Y(n1195gat),.A(n1197gat));
  NOT NOT1_748(.VSS(VSS),.VDD(VDD),.Y(I1947),.A(n1197gat));
  NOT NOT1_749(.VSS(VSS),.VDD(VDD),.Y(n1196gat),.A(I1947));
  NOT NOT1_750(.VSS(VSS),.VDD(VDD),.Y(n2516gat),.A(n2518gat));
  NOT NOT1_751(.VSS(VSS),.VDD(VDD),.Y(I1961),.A(n2516gat));
  NOT NOT1_752(.VSS(VSS),.VDD(VDD),.Y(n3017gat),.A(I1961));
  NOT NOT1_753(.VSS(VSS),.VDD(VDD),.Y(n851gat),.A(n853gat));
  NOT NOT1_754(.VSS(VSS),.VDD(VDD),.Y(n1725gat),.A(n2148gat));
  NOT NOT1_755(.VSS(VSS),.VDD(VDD),.Y(n664gat),.A(n1725gat));
  NOT NOT1_756(.VSS(VSS),.VDD(VDD),.Y(n852gat),.A(n854gat));
  NOT NOT1_757(.VSS(VSS),.VDD(VDD),.Y(I1981),.A(n667gat));
  NOT NOT1_758(.VSS(VSS),.VDD(VDD),.Y(n666gat),.A(I1981));
  NOT NOT1_759(.VSS(VSS),.VDD(VDD),.Y(n368gat),.A(n1725gat));
  NOT NOT1_760(.VSS(VSS),.VDD(VDD),.Y(I1996),.A(n659gat));
  NOT NOT1_761(.VSS(VSS),.VDD(VDD),.Y(n658gat),.A(I1996));
  NOT NOT1_762(.VSS(VSS),.VDD(VDD),.Y(I1999),.A(n658gat));
  NOT NOT1_763(.VSS(VSS),.VDD(VDD),.Y(n784gat),.A(I1999));
  NOT NOT1_764(.VSS(VSS),.VDD(VDD),.Y(n662gat),.A(n1725gat));
  NOT NOT1_765(.VSS(VSS),.VDD(VDD),.Y(I2014),.A(n553gat));
  NOT NOT1_766(.VSS(VSS),.VDD(VDD),.Y(n552gat),.A(I2014));
  NOT NOT1_767(.VSS(VSS),.VDD(VDD),.Y(I2017),.A(n552gat));
  NOT NOT1_768(.VSS(VSS),.VDD(VDD),.Y(n785gat),.A(I2017));
  NOT NOT1_769(.VSS(VSS),.VDD(VDD),.Y(n661gat),.A(n1725gat));
  NOT NOT1_770(.VSS(VSS),.VDD(VDD),.Y(I2032),.A(n777gat));
  NOT NOT1_771(.VSS(VSS),.VDD(VDD),.Y(n776gat),.A(I2032));
  NOT NOT1_772(.VSS(VSS),.VDD(VDD),.Y(I2035),.A(n776gat));
  NOT NOT1_773(.VSS(VSS),.VDD(VDD),.Y(n786gat),.A(I2035));
  NOT NOT1_774(.VSS(VSS),.VDD(VDD),.Y(n551gat),.A(n553gat));
  NOT NOT1_775(.VSS(VSS),.VDD(VDD),.Y(I2040),.A(n551gat));
  NOT NOT1_776(.VSS(VSS),.VDD(VDD),.Y(n787gat),.A(I2040));
  NOT NOT1_777(.VSS(VSS),.VDD(VDD),.Y(n775gat),.A(n777gat));
  NOT NOT1_778(.VSS(VSS),.VDD(VDD),.Y(I2044),.A(n775gat));
  NOT NOT1_779(.VSS(VSS),.VDD(VDD),.Y(n788gat),.A(I2044));
  NOT NOT1_780(.VSS(VSS),.VDD(VDD),.Y(n657gat),.A(n659gat));
  NOT NOT1_781(.VSS(VSS),.VDD(VDD),.Y(I2049),.A(n657gat));
  NOT NOT1_782(.VSS(VSS),.VDD(VDD),.Y(n789gat),.A(I2049));
  NOT NOT1_783(.VSS(VSS),.VDD(VDD),.Y(n35gat),.A(n779gat));
  NOT NOT1_784(.VSS(VSS),.VDD(VDD),.Y(I2056),.A(n35gat));
  NOT NOT1_785(.VSS(VSS),.VDD(VDD),.Y(n125gat),.A(I2056));
  NOT NOT1_786(.VSS(VSS),.VDD(VDD),.Y(n558gat),.A(n1725gat));
  NOT NOT1_787(.VSS(VSS),.VDD(VDD),.Y(n559gat),.A(n561gat));
  NOT NOT1_788(.VSS(VSS),.VDD(VDD),.Y(n371gat),.A(n1725gat));
  NOT NOT1_789(.VSS(VSS),.VDD(VDD),.Y(I2084),.A(n366gat));
  NOT NOT1_790(.VSS(VSS),.VDD(VDD),.Y(n365gat),.A(I2084));
  NOT NOT1_791(.VSS(VSS),.VDD(VDD),.Y(I2088),.A(n561gat));
  NOT NOT1_792(.VSS(VSS),.VDD(VDD),.Y(n560gat),.A(I2088));
  NOT NOT1_793(.VSS(VSS),.VDD(VDD),.Y(n364gat),.A(n366gat));
  NOT NOT1_794(.VSS(VSS),.VDD(VDD),.Y(I2094),.A(n2876gat));
  NOT NOT1_795(.VSS(VSS),.VDD(VDD),.Y(n126gat),.A(I2094));
  NOT NOT1_796(.VSS(VSS),.VDD(VDD),.Y(n663gat),.A(n1725gat));
  NOT NOT1_797(.VSS(VSS),.VDD(VDD),.Y(I2109),.A(n322gat));
  NOT NOT1_798(.VSS(VSS),.VDD(VDD),.Y(n321gat),.A(I2109));
  NOT NOT1_799(.VSS(VSS),.VDD(VDD),.Y(I2112),.A(n321gat));
  NOT NOT1_800(.VSS(VSS),.VDD(VDD),.Y(n226gat),.A(I2112));
  NOT NOT1_801(.VSS(VSS),.VDD(VDD),.Y(n370gat),.A(n1725gat));
  NOT NOT1_802(.VSS(VSS),.VDD(VDD),.Y(I2127),.A(n318gat));
  NOT NOT1_803(.VSS(VSS),.VDD(VDD),.Y(n317gat),.A(I2127));
  NOT NOT1_804(.VSS(VSS),.VDD(VDD),.Y(I2130),.A(n317gat));
  NOT NOT1_805(.VSS(VSS),.VDD(VDD),.Y(n227gat),.A(I2130));
  NOT NOT1_806(.VSS(VSS),.VDD(VDD),.Y(n369gat),.A(n1725gat));
  NOT NOT1_807(.VSS(VSS),.VDD(VDD),.Y(I2145),.A(n314gat));
  NOT NOT1_808(.VSS(VSS),.VDD(VDD),.Y(n313gat),.A(I2145));
  NOT NOT1_809(.VSS(VSS),.VDD(VDD),.Y(I2148),.A(n313gat));
  NOT NOT1_810(.VSS(VSS),.VDD(VDD),.Y(n228gat),.A(I2148));
  NOT NOT1_811(.VSS(VSS),.VDD(VDD),.Y(n316gat),.A(n318gat));
  NOT NOT1_812(.VSS(VSS),.VDD(VDD),.Y(I2153),.A(n316gat));
  NOT NOT1_813(.VSS(VSS),.VDD(VDD),.Y(n229gat),.A(I2153));
  NOT NOT1_814(.VSS(VSS),.VDD(VDD),.Y(n312gat),.A(n314gat));
  NOT NOT1_815(.VSS(VSS),.VDD(VDD),.Y(I2157),.A(n312gat));
  NOT NOT1_816(.VSS(VSS),.VDD(VDD),.Y(n230gat),.A(I2157));
  NOT NOT1_817(.VSS(VSS),.VDD(VDD),.Y(n320gat),.A(n322gat));
  NOT NOT1_818(.VSS(VSS),.VDD(VDD),.Y(I2162),.A(n320gat));
  NOT NOT1_819(.VSS(VSS),.VDD(VDD),.Y(n231gat),.A(I2162));
  NOT NOT1_820(.VSS(VSS),.VDD(VDD),.Y(n34gat),.A(n221gat));
  NOT NOT1_821(.VSS(VSS),.VDD(VDD),.Y(I2169),.A(n34gat));
  NOT NOT1_822(.VSS(VSS),.VDD(VDD),.Y(n127gat),.A(I2169));
  NOT NOT1_823(.VSS(VSS),.VDD(VDD),.Y(n133gat),.A(n2876gat));
  NOT NOT1_824(.VSS(VSS),.VDD(VDD),.Y(I2174),.A(n133gat));
  NOT NOT1_825(.VSS(VSS),.VDD(VDD),.Y(n128gat),.A(I2174));
  NOT NOT1_826(.VSS(VSS),.VDD(VDD),.Y(I2177),.A(n221gat));
  NOT NOT1_827(.VSS(VSS),.VDD(VDD),.Y(n129gat),.A(I2177));
  NOT NOT1_828(.VSS(VSS),.VDD(VDD),.Y(I2181),.A(n779gat));
  NOT NOT1_829(.VSS(VSS),.VDD(VDD),.Y(n130gat),.A(I2181));
  NOT NOT1_830(.VSS(VSS),.VDD(VDD),.Y(n665gat),.A(n667gat));
  NOT NOT1_831(.VSS(VSS),.VDD(VDD),.Y(n1601gat),.A(n120gat));
  NOT NOT1_832(.VSS(VSS),.VDD(VDD),.Y(n2597gat),.A(n2599gat));
  NOT NOT1_833(.VSS(VSS),.VDD(VDD),.Y(n2595gat),.A(n2594gat));
  NOT NOT1_834(.VSS(VSS),.VDD(VDD),.Y(n2586gat),.A(n2588gat));
  NOT NOT1_835(.VSS(VSS),.VDD(VDD),.Y(I2213),.A(n2342gat));
  NOT NOT1_836(.VSS(VSS),.VDD(VDD),.Y(n2573gat),.A(I2213));
  NOT NOT1_837(.VSS(VSS),.VDD(VDD),.Y(n2638gat),.A(n2640gat));
  NOT NOT1_838(.VSS(VSS),.VDD(VDD),.Y(I2225),.A(n2638gat));
  NOT NOT1_839(.VSS(VSS),.VDD(VDD),.Y(n2574gat),.A(I2225));
  NOT NOT1_840(.VSS(VSS),.VDD(VDD),.Y(I2228),.A(n2561gat));
  NOT NOT1_841(.VSS(VSS),.VDD(VDD),.Y(n2575gat),.A(I2228));
  NOT NOT1_842(.VSS(VSS),.VDD(VDD),.Y(I2232),.A(n2640gat));
  NOT NOT1_843(.VSS(VSS),.VDD(VDD),.Y(n2639gat),.A(I2232));
  NOT NOT1_844(.VSS(VSS),.VDD(VDD),.Y(I2235),.A(n2639gat));
  NOT NOT1_845(.VSS(VSS),.VDD(VDD),.Y(n2576gat),.A(I2235));
  NOT NOT1_846(.VSS(VSS),.VDD(VDD),.Y(I2238),.A(n2560gat));
  NOT NOT1_847(.VSS(VSS),.VDD(VDD),.Y(n2577gat),.A(I2238));
  NOT NOT1_848(.VSS(VSS),.VDD(VDD),.Y(I2242),.A(n2341gat));
  NOT NOT1_849(.VSS(VSS),.VDD(VDD),.Y(n2578gat),.A(I2242));
  NOT NOT1_850(.VSS(VSS),.VDD(VDD),.Y(I2248),.A(n2568gat));
  NOT NOT1_851(.VSS(VSS),.VDD(VDD),.Y(n2582gat),.A(I2248));
  NOT NOT1_852(.VSS(VSS),.VDD(VDD),.Y(I2251),.A(n2207gat));
  NOT NOT1_853(.VSS(VSS),.VDD(VDD),.Y(n2206gat),.A(I2251));
  NOT NOT1_854(.VSS(VSS),.VDD(VDD),.Y(I2254),.A(n2206gat));
  NOT NOT1_855(.VSS(VSS),.VDD(VDD),.Y(n2414gat),.A(I2254));
  NOT NOT1_856(.VSS(VSS),.VDD(VDD),.Y(I2257),.A(n2398gat));
  NOT NOT1_857(.VSS(VSS),.VDD(VDD),.Y(n2415gat),.A(I2257));
  NOT NOT1_858(.VSS(VSS),.VDD(VDD),.Y(I2260),.A(n2203gat));
  NOT NOT1_859(.VSS(VSS),.VDD(VDD),.Y(n2202gat),.A(I2260));
  NOT NOT1_860(.VSS(VSS),.VDD(VDD),.Y(I2263),.A(n2202gat));
  NOT NOT1_861(.VSS(VSS),.VDD(VDD),.Y(n2416gat),.A(I2263));
  NOT NOT1_862(.VSS(VSS),.VDD(VDD),.Y(n2397gat),.A(n2399gat));
  NOT NOT1_863(.VSS(VSS),.VDD(VDD),.Y(I2268),.A(n2397gat));
  NOT NOT1_864(.VSS(VSS),.VDD(VDD),.Y(n2417gat),.A(I2268));
  NOT NOT1_865(.VSS(VSS),.VDD(VDD),.Y(I2271),.A(n2201gat));
  NOT NOT1_866(.VSS(VSS),.VDD(VDD),.Y(n2418gat),.A(I2271));
  NOT NOT1_867(.VSS(VSS),.VDD(VDD),.Y(I2275),.A(n2205gat));
  NOT NOT1_868(.VSS(VSS),.VDD(VDD),.Y(n2419gat),.A(I2275));
  NOT NOT1_869(.VSS(VSS),.VDD(VDD),.Y(I2281),.A(n2409gat));
  NOT NOT1_870(.VSS(VSS),.VDD(VDD),.Y(n2585gat),.A(I2281));
  NOT NOT1_871(.VSS(VSS),.VDD(VDD),.Y(n2656gat),.A(n2658gat));
  NOT NOT1_872(.VSS(VSS),.VDD(VDD),.Y(n2493gat),.A(n2495gat));
  NOT NOT1_873(.VSS(VSS),.VDD(VDD),.Y(n2388gat),.A(n2390gat));
  NOT NOT1_874(.VSS(VSS),.VDD(VDD),.Y(I2316),.A(n2390gat));
  NOT NOT1_875(.VSS(VSS),.VDD(VDD),.Y(n2389gat),.A(I2316));
  NOT NOT1_876(.VSS(VSS),.VDD(VDD),.Y(I2319),.A(n2495gat));
  NOT NOT1_877(.VSS(VSS),.VDD(VDD),.Y(n2494gat),.A(I2319));
  NOT NOT1_878(.VSS(VSS),.VDD(VDD),.Y(I2324),.A(n3014gat));
  NOT NOT1_879(.VSS(VSS),.VDD(VDD),.Y(n2649gat),.A(I2324));
  NOT NOT1_880(.VSS(VSS),.VDD(VDD),.Y(n2268gat),.A(n2270gat));
  NOT NOT1_881(.VSS(VSS),.VDD(VDD),.Y(I2344),.A(n2339gat));
  NOT NOT1_882(.VSS(VSS),.VDD(VDD),.Y(n2338gat),.A(I2344));
  NOT NOT1_883(.VSS(VSS),.VDD(VDD),.Y(n2337gat),.A(n2339gat));
  NOT NOT1_884(.VSS(VSS),.VDD(VDD),.Y(I2349),.A(n2270gat));
  NOT NOT1_885(.VSS(VSS),.VDD(VDD),.Y(n2269gat),.A(I2349));
  NOT NOT1_886(.VSS(VSS),.VDD(VDD),.Y(I2354),.A(n2880gat));
  NOT NOT1_887(.VSS(VSS),.VDD(VDD),.Y(n2652gat),.A(I2354));
  NOT NOT1_888(.VSS(VSS),.VDD(VDD),.Y(n2500gat),.A(n2502gat));
  NOT NOT1_889(.VSS(VSS),.VDD(VDD),.Y(n2620gat),.A(n2622gat));
  NOT NOT1_890(.VSS(VSS),.VDD(VDD),.Y(n2612gat),.A(n2620gat));
  NOT NOT1_891(.VSS(VSS),.VDD(VDD),.Y(I2372),.A(n2612gat));
  NOT NOT1_892(.VSS(VSS),.VDD(VDD),.Y(n2606gat),.A(I2372));
  NOT NOT1_893(.VSS(VSS),.VDD(VDD),.Y(n2532gat),.A(n2625gat));
  NOT NOT1_894(.VSS(VSS),.VDD(VDD),.Y(I2376),.A(n2532gat));
  NOT NOT1_895(.VSS(VSS),.VDD(VDD),.Y(n2607gat),.A(I2376));
  NOT NOT1_896(.VSS(VSS),.VDD(VDD),.Y(n2540gat),.A(n2488gat));
  NOT NOT1_897(.VSS(VSS),.VDD(VDD),.Y(I2380),.A(n2540gat));
  NOT NOT1_898(.VSS(VSS),.VDD(VDD),.Y(n2608gat),.A(I2380));
  NOT NOT1_899(.VSS(VSS),.VDD(VDD),.Y(n2536gat),.A(n2624gat));
  NOT NOT1_900(.VSS(VSS),.VDD(VDD),.Y(I2385),.A(n2536gat));
  NOT NOT1_901(.VSS(VSS),.VDD(VDD),.Y(n2609gat),.A(I2385));
  NOT NOT1_902(.VSS(VSS),.VDD(VDD),.Y(n2487gat),.A(n2489gat));
  NOT NOT1_903(.VSS(VSS),.VDD(VDD),.Y(I2389),.A(n2487gat));
  NOT NOT1_904(.VSS(VSS),.VDD(VDD),.Y(n2610gat),.A(I2389));
  NOT NOT1_905(.VSS(VSS),.VDD(VDD),.Y(n2557gat),.A(n2621gat));
  NOT NOT1_906(.VSS(VSS),.VDD(VDD),.Y(I2394),.A(n2557gat));
  NOT NOT1_907(.VSS(VSS),.VDD(VDD),.Y(n2611gat),.A(I2394));
  NOT NOT1_908(.VSS(VSS),.VDD(VDD),.Y(I2400),.A(n2601gat));
  NOT NOT1_909(.VSS(VSS),.VDD(VDD),.Y(n2616gat),.A(I2400));
  NOT NOT1_910(.VSS(VSS),.VDD(VDD),.Y(I2403),.A(n2629gat));
  NOT NOT1_911(.VSS(VSS),.VDD(VDD),.Y(n2550gat),.A(I2403));
  NOT NOT1_912(.VSS(VSS),.VDD(VDD),.Y(I2414),.A(n2634gat));
  NOT NOT1_913(.VSS(VSS),.VDD(VDD),.Y(n2633gat),.A(I2414));
  NOT NOT1_914(.VSS(VSS),.VDD(VDD),.Y(I2417),.A(n2633gat));
  NOT NOT1_915(.VSS(VSS),.VDD(VDD),.Y(n2551gat),.A(I2417));
  NOT NOT1_916(.VSS(VSS),.VDD(VDD),.Y(I2420),.A(n2542gat));
  NOT NOT1_917(.VSS(VSS),.VDD(VDD),.Y(n2552gat),.A(I2420));
  NOT NOT1_918(.VSS(VSS),.VDD(VDD),.Y(n2632gat),.A(n2634gat));
  NOT NOT1_919(.VSS(VSS),.VDD(VDD),.Y(I2425),.A(n2632gat));
  NOT NOT1_920(.VSS(VSS),.VDD(VDD),.Y(n2553gat),.A(I2425));
  NOT NOT1_921(.VSS(VSS),.VDD(VDD),.Y(I2428),.A(n2541gat));
  NOT NOT1_922(.VSS(VSS),.VDD(VDD),.Y(n2554gat),.A(I2428));
  NOT NOT1_923(.VSS(VSS),.VDD(VDD),.Y(n2628gat),.A(n2630gat));
  NOT NOT1_924(.VSS(VSS),.VDD(VDD),.Y(I2433),.A(n2628gat));
  NOT NOT1_925(.VSS(VSS),.VDD(VDD),.Y(n2555gat),.A(I2433));
  NOT NOT1_926(.VSS(VSS),.VDD(VDD),.Y(I2439),.A(n2545gat));
  NOT NOT1_927(.VSS(VSS),.VDD(VDD),.Y(n2619gat),.A(I2439));
  NOT NOT1_928(.VSS(VSS),.VDD(VDD),.Y(n2504gat),.A(n2506gat));
  NOT NOT1_929(.VSS(VSS),.VDD(VDD),.Y(n2660gat),.A(n2655gat));
  NOT NOT1_930(.VSS(VSS),.VDD(VDD),.Y(n1528gat),.A(n2293gat));
  NOT NOT1_931(.VSS(VSS),.VDD(VDD),.Y(n1523gat),.A(n2219gat));
  NOT NOT1_932(.VSS(VSS),.VDD(VDD),.Y(n1592gat),.A(n1529gat));
  NOT NOT1_933(.VSS(VSS),.VDD(VDD),.Y(n2666gat),.A(n1704gat));
  NOT NOT1_934(.VSS(VSS),.VDD(VDD),.Y(n2422gat),.A(n3013gat));
  NOT NOT1_935(.VSS(VSS),.VDD(VDD),.Y(n2290gat),.A(n2202gat));
  NOT NOT1_936(.VSS(VSS),.VDD(VDD),.Y(n2081gat),.A(n2218gat));
  NOT NOT1_937(.VSS(VSS),.VDD(VDD),.Y(n2285gat),.A(n2397gat));
  NOT NOT1_938(.VSS(VSS),.VDD(VDD),.Y(n2359gat),.A(n2358gat));
  NOT NOT1_939(.VSS(VSS),.VDD(VDD),.Y(n1414gat),.A(n1415gat));
  NOT NOT1_940(.VSS(VSS),.VDD(VDD),.Y(n566gat),.A(n364gat));
  NOT NOT1_941(.VSS(VSS),.VDD(VDD),.Y(n1480gat),.A(n2292gat));
  NOT NOT1_942(.VSS(VSS),.VDD(VDD),.Y(n1301gat),.A(n1416gat));
  NOT NOT1_943(.VSS(VSS),.VDD(VDD),.Y(n1150gat),.A(n312gat));
  NOT NOT1_944(.VSS(VSS),.VDD(VDD),.Y(n873gat),.A(n316gat));
  NOT NOT1_945(.VSS(VSS),.VDD(VDD),.Y(n2011gat),.A(n2306gat));
  NOT NOT1_946(.VSS(VSS),.VDD(VDD),.Y(n1478gat),.A(n1481gat));
  NOT NOT1_947(.VSS(VSS),.VDD(VDD),.Y(n875gat),.A(n559gat));
  NOT NOT1_948(.VSS(VSS),.VDD(VDD),.Y(n1410gat),.A(n2357gat));
  NOT NOT1_949(.VSS(VSS),.VDD(VDD),.Y(n876gat),.A(n1347gat));
  NOT NOT1_950(.VSS(VSS),.VDD(VDD),.Y(n1160gat),.A(n1484gat));
  NOT NOT1_951(.VSS(VSS),.VDD(VDD),.Y(n1084gat),.A(n657gat));
  NOT NOT1_952(.VSS(VSS),.VDD(VDD),.Y(n983gat),.A(n320gat));
  NOT NOT1_953(.VSS(VSS),.VDD(VDD),.Y(n1482gat),.A(n2363gat));
  NOT NOT1_954(.VSS(VSS),.VDD(VDD),.Y(n1157gat),.A(n1483gat));
  NOT NOT1_955(.VSS(VSS),.VDD(VDD),.Y(n985gat),.A(n775gat));
  NOT NOT1_956(.VSS(VSS),.VDD(VDD),.Y(n1530gat),.A(n2364gat));
  NOT NOT1_957(.VSS(VSS),.VDD(VDD),.Y(n1307gat),.A(n1308gat));
  NOT NOT1_958(.VSS(VSS),.VDD(VDD),.Y(n1085gat),.A(n551gat));
  NOT NOT1_959(.VSS(VSS),.VDD(VDD),.Y(n1479gat),.A(n2291gat));
  NOT NOT1_960(.VSS(VSS),.VDD(VDD),.Y(n1348gat),.A(n1349gat));
  NOT NOT1_961(.VSS(VSS),.VDD(VDD),.Y(n2217gat),.A(n2206gat));
  NOT NOT1_962(.VSS(VSS),.VDD(VDD),.Y(n1591gat),.A(n2223gat));
  NOT NOT1_963(.VSS(VSS),.VDD(VDD),.Y(n1437gat),.A(n1438gat));
  NOT NOT1_964(.VSS(VSS),.VDD(VDD),.Y(n1832gat),.A(n1834gat));
  NOT NOT1_965(.VSS(VSS),.VDD(VDD),.Y(n1765gat),.A(n1767gat));
  NOT NOT1_966(.VSS(VSS),.VDD(VDD),.Y(n1878gat),.A(n1880gat));
  NOT NOT1_967(.VSS(VSS),.VDD(VDD),.Y(n1442gat),.A(n1831gat));
  NOT NOT1_968(.VSS(VSS),.VDD(VDD),.Y(n1444gat),.A(n1442gat));
  NOT NOT1_969(.VSS(VSS),.VDD(VDD),.Y(n1378gat),.A(n2975gat));
  NOT NOT1_970(.VSS(VSS),.VDD(VDD),.Y(n1322gat),.A(n2974gat));
  NOT NOT1_971(.VSS(VSS),.VDD(VDD),.Y(n1439gat),.A(n1486gat));
  NOT NOT1_972(.VSS(VSS),.VDD(VDD),.Y(n1370gat),.A(n1426gat));
  NOT NOT1_973(.VSS(VSS),.VDD(VDD),.Y(n1369gat),.A(n2966gat));
  NOT NOT1_974(.VSS(VSS),.VDD(VDD),.Y(n1366gat),.A(n1365gat));
  NOT NOT1_975(.VSS(VSS),.VDD(VDD),.Y(n1374gat),.A(n2979gat));
  NOT NOT1_976(.VSS(VSS),.VDD(VDD),.Y(n2162gat),.A(n2220gat));
  NOT NOT1_977(.VSS(VSS),.VDD(VDD),.Y(n1450gat),.A(n1423gat));
  NOT NOT1_978(.VSS(VSS),.VDD(VDD),.Y(n1427gat),.A(n1608gat));
  NOT NOT1_979(.VSS(VSS),.VDD(VDD),.Y(n1603gat),.A(n1831gat));
  NOT NOT1_980(.VSS(VSS),.VDD(VDD),.Y(n2082gat),.A(n2084gat));
  NOT NOT1_981(.VSS(VSS),.VDD(VDD),.Y(n1449gat),.A(n1494gat));
  NOT NOT1_982(.VSS(VSS),.VDD(VDD),.Y(n1590gat),.A(n1603gat));
  NOT NOT1_983(.VSS(VSS),.VDD(VDD),.Y(n1248gat),.A(n2954gat));
  NOT NOT1_984(.VSS(VSS),.VDD(VDD),.Y(n1418gat),.A(n1417gat));
  NOT NOT1_985(.VSS(VSS),.VDD(VDD),.Y(n1306gat),.A(n2964gat));
  NOT NOT1_986(.VSS(VSS),.VDD(VDD),.Y(n1353gat),.A(n1419gat));
  NOT NOT1_987(.VSS(VSS),.VDD(VDD),.Y(n1247gat),.A(n2958gat));
  NOT NOT1_988(.VSS(VSS),.VDD(VDD),.Y(n1355gat),.A(n1422gat));
  NOT NOT1_989(.VSS(VSS),.VDD(VDD),.Y(n1300gat),.A(n2963gat));
  NOT NOT1_990(.VSS(VSS),.VDD(VDD),.Y(n1487gat),.A(n1485gat));
  NOT NOT1_991(.VSS(VSS),.VDD(VDD),.Y(n1164gat),.A(n2953gat));
  NOT NOT1_992(.VSS(VSS),.VDD(VDD),.Y(n1356gat),.A(n1354gat));
  NOT NOT1_993(.VSS(VSS),.VDD(VDD),.Y(n1436gat),.A(n1435gat));
  NOT NOT1_994(.VSS(VSS),.VDD(VDD),.Y(n1106gat),.A(n2949gat));
  NOT NOT1_995(.VSS(VSS),.VDD(VDD),.Y(n1425gat),.A(n1421gat));
  NOT NOT1_996(.VSS(VSS),.VDD(VDD),.Y(n1105gat),.A(n2934gat));
  NOT NOT1_997(.VSS(VSS),.VDD(VDD),.Y(n1424gat),.A(n1420gat));
  NOT NOT1_998(.VSS(VSS),.VDD(VDD),.Y(n1309gat),.A(n2959gat));
  NOT NOT1_999(.VSS(VSS),.VDD(VDD),.Y(I2672),.A(n2143gat));
  NOT NOT1_1000(.VSS(VSS),.VDD(VDD),.Y(n2142gat),.A(I2672));
  NOT NOT1_1001(.VSS(VSS),.VDD(VDD),.Y(n1788gat),.A(n2142gat));
  NOT NOT1_1002(.VSS(VSS),.VDD(VDD),.Y(I2684),.A(n2061gat));
  NOT NOT1_1003(.VSS(VSS),.VDD(VDD),.Y(n2060gat),.A(I2684));
  NOT NOT1_1004(.VSS(VSS),.VDD(VDD),.Y(n1786gat),.A(n2060gat));
  NOT NOT1_1005(.VSS(VSS),.VDD(VDD),.Y(I2696),.A(n2139gat));
  NOT NOT1_1006(.VSS(VSS),.VDD(VDD),.Y(n2138gat),.A(I2696));
  NOT NOT1_1007(.VSS(VSS),.VDD(VDD),.Y(n1839gat),.A(n2138gat));
  NOT NOT1_1008(.VSS(VSS),.VDD(VDD),.Y(n1897gat),.A(n1899gat));
  NOT NOT1_1009(.VSS(VSS),.VDD(VDD),.Y(n1884gat),.A(n1897gat));
  NOT NOT1_1010(.VSS(VSS),.VDD(VDD),.Y(n1848gat),.A(n1850gat));
  NOT NOT1_1011(.VSS(VSS),.VDD(VDD),.Y(n1783gat),.A(n1848gat));
  NOT NOT1_1012(.VSS(VSS),.VDD(VDD),.Y(n1548gat),.A(I2721));
  NOT NOT1_1013(.VSS(VSS),.VDD(VDD),.Y(n1719gat),.A(n1548gat));
  NOT NOT1_1014(.VSS(VSS),.VDD(VDD),.Y(n2137gat),.A(n2139gat));
  NOT NOT1_1015(.VSS(VSS),.VDD(VDD),.Y(n1633gat),.A(n2137gat));
  NOT NOT1_1016(.VSS(VSS),.VDD(VDD),.Y(n2059gat),.A(n2061gat));
  NOT NOT1_1017(.VSS(VSS),.VDD(VDD),.Y(n1785gat),.A(n2059gat));
  NOT NOT1_1018(.VSS(VSS),.VDD(VDD),.Y(I2731),.A(n1850gat));
  NOT NOT1_1019(.VSS(VSS),.VDD(VDD),.Y(n1849gat),.A(I2731));
  NOT NOT1_1020(.VSS(VSS),.VDD(VDD),.Y(n1784gat),.A(n1849gat));
  NOT NOT1_1021(.VSS(VSS),.VDD(VDD),.Y(n1716gat),.A(I2736));
  NOT NOT1_1022(.VSS(VSS),.VDD(VDD),.Y(n1635gat),.A(n1716gat));
  NOT NOT1_1023(.VSS(VSS),.VDD(VDD),.Y(n2401gat),.A(n2403gat));
  NOT NOT1_1024(.VSS(VSS),.VDD(VDD),.Y(n1989gat),.A(n2401gat));
  NOT NOT1_1025(.VSS(VSS),.VDD(VDD),.Y(n2392gat),.A(n2394gat));
  NOT NOT1_1026(.VSS(VSS),.VDD(VDD),.Y(n1918gat),.A(n2392gat));
  NOT NOT1_1027(.VSS(VSS),.VDD(VDD),.Y(I2771),.A(n2440gat));
  NOT NOT1_1028(.VSS(VSS),.VDD(VDD),.Y(n2439gat),.A(I2771));
  NOT NOT1_1029(.VSS(VSS),.VDD(VDD),.Y(n1986gat),.A(n2439gat));
  NOT NOT1_1030(.VSS(VSS),.VDD(VDD),.Y(n1866gat),.A(n1865gat));
  NOT NOT1_1031(.VSS(VSS),.VDD(VDD),.Y(I2785),.A(n2407gat));
  NOT NOT1_1032(.VSS(VSS),.VDD(VDD),.Y(n2406gat),.A(I2785));
  NOT NOT1_1033(.VSS(VSS),.VDD(VDD),.Y(n2216gat),.A(n2406gat));
  NOT NOT1_1034(.VSS(VSS),.VDD(VDD),.Y(n2345gat),.A(n2347gat));
  NOT NOT1_1035(.VSS(VSS),.VDD(VDD),.Y(n1988gat),.A(n2345gat));
  NOT NOT1_1036(.VSS(VSS),.VDD(VDD),.Y(n1735gat),.A(n1861gat));
  NOT NOT1_1037(.VSS(VSS),.VDD(VDD),.Y(n1387gat),.A(n1389gat));
  NOT NOT1_1038(.VSS(VSS),.VDD(VDD),.Y(n1694gat),.A(I2813));
  NOT NOT1_1039(.VSS(VSS),.VDD(VDD),.Y(n1777gat),.A(n1694gat));
  NOT NOT1_1040(.VSS(VSS),.VDD(VDD),.Y(n1781gat),.A(n1780gat));
  NOT NOT1_1041(.VSS(VSS),.VDD(VDD),.Y(n2019gat),.A(n2021gat));
  NOT NOT1_1042(.VSS(VSS),.VDD(VDD),.Y(n1549gat),.A(I2832));
  NOT NOT1_1043(.VSS(VSS),.VDD(VDD),.Y(n1551gat),.A(n1549gat));
  NOT NOT1_1044(.VSS(VSS),.VDD(VDD),.Y(I2837),.A(n2347gat));
  NOT NOT1_1045(.VSS(VSS),.VDD(VDD),.Y(n2346gat),.A(I2837));
  NOT NOT1_1046(.VSS(VSS),.VDD(VDD),.Y(n2152gat),.A(n2346gat));
  NOT NOT1_1047(.VSS(VSS),.VDD(VDD),.Y(n2405gat),.A(n2407gat));
  NOT NOT1_1048(.VSS(VSS),.VDD(VDD),.Y(n2351gat),.A(n2405gat));
  NOT NOT1_1049(.VSS(VSS),.VDD(VDD),.Y(I2843),.A(n2403gat));
  NOT NOT1_1050(.VSS(VSS),.VDD(VDD),.Y(n2402gat),.A(I2843));
  NOT NOT1_1051(.VSS(VSS),.VDD(VDD),.Y(n2212gat),.A(n2402gat));
  NOT NOT1_1052(.VSS(VSS),.VDD(VDD),.Y(I2847),.A(n2394gat));
  NOT NOT1_1053(.VSS(VSS),.VDD(VDD),.Y(n2393gat),.A(I2847));
  NOT NOT1_1054(.VSS(VSS),.VDD(VDD),.Y(n1991gat),.A(n2393gat));
  NOT NOT1_1055(.VSS(VSS),.VDD(VDD),.Y(n1665gat),.A(n1666gat));
  NOT NOT1_1056(.VSS(VSS),.VDD(VDD),.Y(n1517gat),.A(n1578gat));
  NOT NOT1_1057(.VSS(VSS),.VDD(VDD),.Y(n1392gat),.A(n1394gat));
  NOT NOT1_1058(.VSS(VSS),.VDD(VDD),.Y(I2873),.A(n1496gat));
  NOT NOT1_1059(.VSS(VSS),.VDD(VDD),.Y(n1495gat),.A(I2873));
  NOT NOT1_1060(.VSS(VSS),.VDD(VDD),.Y(n1685gat),.A(n1604gat));
  NOT NOT1_1061(.VSS(VSS),.VDD(VDD),.Y(I2885),.A(n2091gat));
  NOT NOT1_1062(.VSS(VSS),.VDD(VDD),.Y(n2090gat),.A(I2885));
  NOT NOT1_1063(.VSS(VSS),.VDD(VDD),.Y(n1550gat),.A(I2890));
  NOT NOT1_1064(.VSS(VSS),.VDD(VDD),.Y(n1552gat),.A(n1550gat));
  NOT NOT1_1065(.VSS(VSS),.VDD(VDD),.Y(n1330gat),.A(n1332gat));
  NOT NOT1_1066(.VSS(VSS),.VDD(VDD),.Y(n1738gat),.A(n1740gat));
  NOT NOT1_1067(.VSS(VSS),.VDD(VDD),.Y(I2915),.A(n1740gat));
  NOT NOT1_1068(.VSS(VSS),.VDD(VDD),.Y(n1739gat),.A(I2915));
  NOT NOT1_1069(.VSS(VSS),.VDD(VDD),.Y(n1925gat),.A(n1920gat));
  NOT NOT1_1070(.VSS(VSS),.VDD(VDD),.Y(n1917gat),.A(n1921gat));
  NOT NOT1_1071(.VSS(VSS),.VDD(VDD),.Y(n2141gat),.A(n2143gat));
  NOT NOT1_1072(.VSS(VSS),.VDD(VDD),.Y(n1787gat),.A(n2141gat));
  NOT NOT1_1073(.VSS(VSS),.VDD(VDD),.Y(n1717gat),.A(I2926));
  NOT NOT1_1074(.VSS(VSS),.VDD(VDD),.Y(n1859gat),.A(n1717gat));
  NOT NOT1_1075(.VSS(VSS),.VDD(VDD),.Y(n1922gat),.A(n1798gat));
  NOT NOT1_1076(.VSS(VSS),.VDD(VDD),.Y(n1713gat),.A(I2935));
  NOT NOT1_1077(.VSS(VSS),.VDD(VDD),.Y(n1743gat),.A(n1713gat));
  NOT NOT1_1078(.VSS(VSS),.VDD(VDD),.Y(n1923gat),.A(n1864gat));
  NOT NOT1_1079(.VSS(VSS),.VDD(VDD),.Y(n1945gat),.A(n1690gat));
  NOT NOT1_1080(.VSS(VSS),.VDD(VDD),.Y(I2953),.A(n2179gat));
  NOT NOT1_1081(.VSS(VSS),.VDD(VDD),.Y(n2178gat),.A(I2953));
  NOT NOT1_1082(.VSS(VSS),.VDD(VDD),.Y(n1661gat),.A(n1660gat));
  NOT NOT1_1083(.VSS(VSS),.VDD(VDD),.Y(n1572gat),.A(n1576gat));
  NOT NOT1_1084(.VSS(VSS),.VDD(VDD),.Y(n2438gat),.A(n2440gat));
  NOT NOT1_1085(.VSS(VSS),.VDD(VDD),.Y(n2283gat),.A(n2438gat));
  NOT NOT1_1086(.VSS(VSS),.VDD(VDD),.Y(n1520gat),.A(n1582gat));
  NOT NOT1_1087(.VSS(VSS),.VDD(VDD),.Y(n1580gat),.A(n1577gat));
  NOT NOT1_1088(.VSS(VSS),.VDD(VDD),.Y(n1990gat),.A(n2988gat));
  NOT NOT1_1089(.VSS(VSS),.VDD(VDD),.Y(I2978),.A(n2190gat));
  NOT NOT1_1090(.VSS(VSS),.VDD(VDD),.Y(n2189gat),.A(I2978));
  NOT NOT1_1091(.VSS(VSS),.VDD(VDD),.Y(I2989),.A(n2135gat));
  NOT NOT1_1092(.VSS(VSS),.VDD(VDD),.Y(n2134gat),.A(I2989));
  NOT NOT1_1093(.VSS(VSS),.VDD(VDD),.Y(I3000),.A(n2262gat));
  NOT NOT1_1094(.VSS(VSS),.VDD(VDD),.Y(n2261gat),.A(I3000));
  NOT NOT1_1095(.VSS(VSS),.VDD(VDD),.Y(n2128gat),.A(n2129gat));
  NOT NOT1_1096(.VSS(VSS),.VDD(VDD),.Y(n1836gat),.A(n1695gat));
  NOT NOT1_1097(.VSS(VSS),.VDD(VDD),.Y(I3016),.A(n2182gat));
  NOT NOT1_1098(.VSS(VSS),.VDD(VDD),.Y(n2181gat),.A(I3016));
  NOT NOT1_1099(.VSS(VSS),.VDD(VDD),.Y(n1431gat),.A(n1433gat));
  NOT NOT1_1100(.VSS(VSS),.VDD(VDD),.Y(n1314gat),.A(n1316gat));
  NOT NOT1_1101(.VSS(VSS),.VDD(VDD),.Y(n1361gat),.A(n1363gat));
  NOT NOT1_1102(.VSS(VSS),.VDD(VDD),.Y(I3056),.A(n1312gat));
  NOT NOT1_1103(.VSS(VSS),.VDD(VDD),.Y(n1311gat),.A(I3056));
  NOT NOT1_1104(.VSS(VSS),.VDD(VDD),.Y(n1707gat),.A(n1626gat));
  NOT NOT1_1105(.VSS(VSS),.VDD(VDD),.Y(n1773gat),.A(n1775gat));
  NOT NOT1_1106(.VSS(VSS),.VDD(VDD),.Y(n1659gat),.A(n2987gat));
  NOT NOT1_1107(.VSS(VSS),.VDD(VDD),.Y(n1515gat),.A(n1521gat));
  NOT NOT1_1108(.VSS(VSS),.VDD(VDD),.Y(n1736gat),.A(n1737gat));
  NOT NOT1_1109(.VSS(VSS),.VDD(VDD),.Y(n1658gat),.A(n2216gat));
  NOT NOT1_1110(.VSS(VSS),.VDD(VDD),.Y(n1724gat),.A(n1732gat));
  NOT NOT1_1111(.VSS(VSS),.VDD(VDD),.Y(n1662gat),.A(n1663gat));
  NOT NOT1_1112(.VSS(VSS),.VDD(VDD),.Y(n1656gat),.A(n1655gat));
  NOT NOT1_1113(.VSS(VSS),.VDD(VDD),.Y(n1670gat),.A(n1667gat));
  NOT NOT1_1114(.VSS(VSS),.VDD(VDD),.Y(n1569gat),.A(n1570gat));
  NOT NOT1_1115(.VSS(VSS),.VDD(VDD),.Y(n1568gat),.A(n1575gat));
  NOT NOT1_1116(.VSS(VSS),.VDD(VDD),.Y(n1727gat),.A(n1728gat));
  NOT NOT1_1117(.VSS(VSS),.VDD(VDD),.Y(n1797gat),.A(n1801gat));
  NOT NOT1_1118(.VSS(VSS),.VDD(VDD),.Y(n1730gat),.A(n1731gat));
  NOT NOT1_1119(.VSS(VSS),.VDD(VDD),.Y(n1561gat),.A(n1571gat));
  NOT NOT1_1120(.VSS(VSS),.VDD(VDD),.Y(n1668gat),.A(n1734gat));
  NOT NOT1_1121(.VSS(VSS),.VDD(VDD),.Y(n1742gat),.A(n2216gat));
  NOT NOT1_1122(.VSS(VSS),.VDD(VDD),.Y(n1671gat),.A(n1669gat));
  NOT NOT1_1123(.VSS(VSS),.VDD(VDD),.Y(n1652gat),.A(n1657gat));
  NOT NOT1_1124(.VSS(VSS),.VDD(VDD),.Y(n1648gat),.A(n1729gat));
  NOT NOT1_1125(.VSS(VSS),.VDD(VDD),.Y(n1790gat),.A(n1726gat));
  NOT NOT1_1126(.VSS(VSS),.VDD(VDD),.Y(n2004gat),.A(n1929gat));
  NOT NOT1_1127(.VSS(VSS),.VDD(VDD),.Y(n1869gat),.A(n1871gat));
  NOT NOT1_1128(.VSS(VSS),.VDD(VDD),.Y(I3143),.A(n2592gat));
  NOT NOT1_1129(.VSS(VSS),.VDD(VDD),.Y(n2591gat),.A(I3143));
  NOT NOT1_1130(.VSS(VSS),.VDD(VDD),.Y(n1584gat),.A(n2989gat));
  NOT NOT1_1131(.VSS(VSS),.VDD(VDD),.Y(n1714gat),.A(I3149));
  NOT NOT1_1132(.VSS(VSS),.VDD(VDD),.Y(n1718gat),.A(n1714gat));
  NOT NOT1_1133(.VSS(VSS),.VDD(VDD),.Y(I3163),.A(n1508gat));
  NOT NOT1_1134(.VSS(VSS),.VDD(VDD),.Y(n1507gat),.A(I3163));
  NOT NOT1_1135(.VSS(VSS),.VDD(VDD),.Y(n1396gat),.A(n1401gat));
  NOT NOT1_1136(.VSS(VSS),.VDD(VDD),.Y(I3168),.A(n1394gat));
  NOT NOT1_1137(.VSS(VSS),.VDD(VDD),.Y(n1393gat),.A(I3168));
  NOT NOT1_1138(.VSS(VSS),.VDD(VDD),.Y(n1409gat),.A(n1476gat));
  NOT NOT1_1139(.VSS(VSS),.VDD(VDD),.Y(I3174),.A(n1899gat));
  NOT NOT1_1140(.VSS(VSS),.VDD(VDD),.Y(n1898gat),.A(I3174));
  NOT NOT1_1141(.VSS(VSS),.VDD(VDD),.Y(n1838gat),.A(n1898gat));
  NOT NOT1_1142(.VSS(VSS),.VDD(VDD),.Y(n1712gat),.A(I3179));
  NOT NOT1_1143(.VSS(VSS),.VDD(VDD),.Y(I3191),.A(n1678gat));
  NOT NOT1_1144(.VSS(VSS),.VDD(VDD),.Y(n1677gat),.A(I3191));
  NOT NOT1_1145(.VSS(VSS),.VDD(VDD),.Y(n2000gat),.A(n1412gat));
  NOT NOT1_1146(.VSS(VSS),.VDD(VDD),.Y(n2001gat),.A(n1412gat));
  NOT NOT1_1147(.VSS(VSS),.VDD(VDD),.Y(n1999gat),.A(n2001gat));
  NOT NOT1_1148(.VSS(VSS),.VDD(VDD),.Y(n2307gat),.A(n2309gat));
  NOT NOT1_1149(.VSS(VSS),.VDD(VDD),.Y(I3211),.A(n2663gat));
  NOT NOT1_1150(.VSS(VSS),.VDD(VDD),.Y(n3018gat),.A(I3211));
  NOT NOT1_1151(.VSS(VSS),.VDD(VDD),.Y(n2448gat),.A(n2450gat));
  NOT NOT1_1152(.VSS(VSS),.VDD(VDD),.Y(n2661gat),.A(n2662gat));
  NOT NOT1_1153(.VSS(VSS),.VDD(VDD),.Y(n2444gat),.A(n2446gat));
  NOT NOT1_1154(.VSS(VSS),.VDD(VDD),.Y(I3235),.A(n2238gat));
  NOT NOT1_1155(.VSS(VSS),.VDD(VDD),.Y(n3019gat),.A(I3235));
  NOT NOT1_1156(.VSS(VSS),.VDD(VDD),.Y(n1310gat),.A(n1312gat));
  NOT NOT1_1157(.VSS(VSS),.VDD(VDD),.Y(n199gat),.A(n87gat));
  NOT NOT1_1158(.VSS(VSS),.VDD(VDD),.Y(n195gat),.A(n184gat));
  NOT NOT1_1159(.VSS(VSS),.VDD(VDD),.Y(n827gat),.A(n204gat));
  NOT NOT1_1160(.VSS(VSS),.VDD(VDD),.Y(n2093gat),.A(n2095gat));
  NOT NOT1_1161(.VSS(VSS),.VDD(VDD),.Y(n2174gat),.A(n2176gat));
  NOT NOT1_1162(.VSS(VSS),.VDD(VDD),.Y(I3273),.A(n2169gat));
  NOT NOT1_1163(.VSS(VSS),.VDD(VDD),.Y(n2168gat),.A(I3273));
  NOT NOT1_1164(.VSS(VSS),.VDD(VDD),.Y(n2452gat),.A(n2454gat));
  NOT NOT1_1165(.VSS(VSS),.VDD(VDD),.Y(n1691gat),.A(n2452gat));
  NOT NOT1_1166(.VSS(VSS),.VDD(VDD),.Y(I3287),.A(n1691gat));
  NOT NOT1_1167(.VSS(VSS),.VDD(VDD),.Y(n3020gat),.A(I3287));
  NOT NOT1_1168(.VSS(VSS),.VDD(VDD),.Y(I3290),.A(n1691gat));
  NOT NOT1_1169(.VSS(VSS),.VDD(VDD),.Y(n3021gat),.A(I3290));
  NOT NOT1_1170(.VSS(VSS),.VDD(VDD),.Y(I3293),.A(n1691gat));
  NOT NOT1_1171(.VSS(VSS),.VDD(VDD),.Y(n3022gat),.A(I3293));
  NOT NOT1_1172(.VSS(VSS),.VDD(VDD),.Y(n1699gat),.A(n2452gat));
  NOT NOT1_1173(.VSS(VSS),.VDD(VDD),.Y(I3297),.A(n1699gat));
  NOT NOT1_1174(.VSS(VSS),.VDD(VDD),.Y(n3023gat),.A(I3297));
  NOT NOT1_1175(.VSS(VSS),.VDD(VDD),.Y(I3300),.A(n1699gat));
  NOT NOT1_1176(.VSS(VSS),.VDD(VDD),.Y(n3024gat),.A(I3300));
  NOT NOT1_1177(.VSS(VSS),.VDD(VDD),.Y(I3303),.A(n1691gat));
  NOT NOT1_1178(.VSS(VSS),.VDD(VDD),.Y(n3025gat),.A(I3303));
  NOT NOT1_1179(.VSS(VSS),.VDD(VDD),.Y(I3306),.A(n1699gat));
  NOT NOT1_1180(.VSS(VSS),.VDD(VDD),.Y(n3026gat),.A(I3306));
  NOT NOT1_1181(.VSS(VSS),.VDD(VDD),.Y(I3309),.A(n1699gat));
  NOT NOT1_1182(.VSS(VSS),.VDD(VDD),.Y(n3027gat),.A(I3309));
  NOT NOT1_1183(.VSS(VSS),.VDD(VDD),.Y(I3312),.A(n1699gat));
  NOT NOT1_1184(.VSS(VSS),.VDD(VDD),.Y(n3028gat),.A(I3312));
  NOT NOT1_1185(.VSS(VSS),.VDD(VDD),.Y(I3315),.A(n1869gat));
  NOT NOT1_1186(.VSS(VSS),.VDD(VDD),.Y(n3029gat),.A(I3315));
  NOT NOT1_1187(.VSS(VSS),.VDD(VDD),.Y(I3318),.A(n1869gat));
  NOT NOT1_1188(.VSS(VSS),.VDD(VDD),.Y(n3030gat),.A(I3318));
  NOT NOT1_1189(.VSS(VSS),.VDD(VDD),.Y(n2260gat),.A(n2262gat));
  NOT NOT1_1190(.VSS(VSS),.VDD(VDD),.Y(n2257gat),.A(n2189gat));
  NOT NOT1_1191(.VSS(VSS),.VDD(VDD),.Y(n2188gat),.A(n2190gat));
  NOT NOT1_1192(.VSS(VSS),.VDD(VDD),.Y(n2187gat),.A(n3004gat));
  NOT NOT1_1193(.VSS(VSS),.VDD(VDD),.Y(I3336),.A(n2040gat));
  NOT NOT1_1194(.VSS(VSS),.VDD(VDD),.Y(n2039gat),.A(I3336));
  NOT NOT1_1195(.VSS(VSS),.VDD(VDD),.Y(I3339),.A(n1775gat));
  NOT NOT1_1196(.VSS(VSS),.VDD(VDD),.Y(n1774gat),.A(I3339));
  NOT NOT1_1197(.VSS(VSS),.VDD(VDD),.Y(I3342),.A(n1316gat));
  NOT NOT1_1198(.VSS(VSS),.VDD(VDD),.Y(n1315gat),.A(I3342));
  NOT NOT1_1199(.VSS(VSS),.VDD(VDD),.Y(n2042gat),.A(n2044gat));
  NOT NOT1_1200(.VSS(VSS),.VDD(VDD),.Y(n2035gat),.A(n2037gat));
  NOT NOT1_1201(.VSS(VSS),.VDD(VDD),.Y(n2023gat),.A(n2025gat));
  NOT NOT1_1202(.VSS(VSS),.VDD(VDD),.Y(n2097gat),.A(n2099gat));
  NOT NOT1_1203(.VSS(VSS),.VDD(VDD),.Y(n1855gat),.A(n2014gat));
  NOT NOT1_1204(.VSS(VSS),.VDD(VDD),.Y(I3387),.A(n2194gat));
  NOT NOT1_1205(.VSS(VSS),.VDD(VDD),.Y(n3031gat),.A(I3387));
  NOT NOT1_1206(.VSS(VSS),.VDD(VDD),.Y(I3390),.A(n2261gat));
  NOT NOT1_1207(.VSS(VSS),.VDD(VDD),.Y(n3032gat),.A(I3390));
  NOT NOT1_1208(.VSS(VSS),.VDD(VDD),.Y(n2256gat),.A(n3032gat));
  NOT NOT1_1209(.VSS(VSS),.VDD(VDD),.Y(I3394),.A(n2260gat));
  NOT NOT1_1210(.VSS(VSS),.VDD(VDD),.Y(n3033gat),.A(I3394));
  NOT NOT1_1211(.VSS(VSS),.VDD(VDD),.Y(n2251gat),.A(n3033gat));
  NOT NOT1_1212(.VSS(VSS),.VDD(VDD),.Y(n2184gat),.A(n3003gat));
  NOT NOT1_1213(.VSS(VSS),.VDD(VDD),.Y(I3401),.A(n2192gat));
  NOT NOT1_1214(.VSS(VSS),.VDD(VDD),.Y(n3034gat),.A(I3401));
  NOT NOT1_1215(.VSS(VSS),.VDD(VDD),.Y(n2133gat),.A(n2135gat));
  NOT NOT1_1216(.VSS(VSS),.VDD(VDD),.Y(n2131gat),.A(n2185gat));
  NOT NOT1_1217(.VSS(VSS),.VDD(VDD),.Y(n2049gat),.A(n3001gat));
  NOT NOT1_1218(.VSS(VSS),.VDD(VDD),.Y(I3412),.A(n2057gat));
  NOT NOT1_1219(.VSS(VSS),.VDD(VDD),.Y(n3035gat),.A(I3412));
  NOT NOT1_1220(.VSS(VSS),.VDD(VDD),.Y(n2253gat),.A(n2189gat));
  NOT NOT1_1221(.VSS(VSS),.VDD(VDD),.Y(n2252gat),.A(n2260gat));
  NOT NOT1_1222(.VSS(VSS),.VDD(VDD),.Y(n2248gat),.A(n3006gat));
  NOT NOT1_1223(.VSS(VSS),.VDD(VDD),.Y(n2264gat),.A(n2266gat));
  NOT NOT1_1224(.VSS(VSS),.VDD(VDD),.Y(I3429),.A(n2266gat));
  NOT NOT1_1225(.VSS(VSS),.VDD(VDD),.Y(n2265gat),.A(I3429));
  NOT NOT1_1226(.VSS(VSS),.VDD(VDD),.Y(n2492gat),.A(n2329gat));
  NOT NOT1_1227(.VSS(VSS),.VDD(VDD),.Y(I3436),.A(n2492gat));
  NOT NOT1_1228(.VSS(VSS),.VDD(VDD),.Y(n3036gat),.A(I3436));
  NOT NOT1_1229(.VSS(VSS),.VDD(VDD),.Y(n1709gat),.A(n1849gat));
  NOT NOT1_1230(.VSS(VSS),.VDD(VDD),.Y(n1845gat),.A(n2141gat));
  NOT NOT1_1231(.VSS(VSS),.VDD(VDD),.Y(n1891gat),.A(n2059gat));
  NOT NOT1_1232(.VSS(VSS),.VDD(VDD),.Y(n1963gat),.A(n2137gat));
  NOT NOT1_1233(.VSS(VSS),.VDD(VDD),.Y(n1886gat),.A(n1897gat));
  NOT NOT1_1234(.VSS(VSS),.VDD(VDD),.Y(n1968gat),.A(n1958gat));
  NOT NOT1_1235(.VSS(VSS),.VDD(VDD),.Y(n1629gat),.A(n1895gat));
  NOT NOT1_1236(.VSS(VSS),.VDD(VDD),.Y(n1631gat),.A(n1848gat));
  NOT NOT1_1237(.VSS(VSS),.VDD(VDD),.Y(n1711gat),.A(n2990gat));
  NOT NOT1_1238(.VSS(VSS),.VDD(VDD),.Y(n2200gat),.A(n2078gat));
  NOT NOT1_1239(.VSS(VSS),.VDD(VDD),.Y(n2437gat),.A(n2195gat));
  NOT NOT1_1240(.VSS(VSS),.VDD(VDD),.Y(I3457),.A(n2556gat));
  NOT NOT1_1241(.VSS(VSS),.VDD(VDD),.Y(n3037gat),.A(I3457));
  NOT NOT1_1242(.VSS(VSS),.VDD(VDD),.Y(n1956gat),.A(n1898gat));
  NOT NOT1_1243(.VSS(VSS),.VDD(VDD),.Y(I3461),.A(n1956gat));
  NOT NOT1_1244(.VSS(VSS),.VDD(VDD),.Y(n3038gat),.A(I3461));
  NOT NOT1_1245(.VSS(VSS),.VDD(VDD),.Y(n1954gat),.A(n3038gat));
  NOT NOT1_1246(.VSS(VSS),.VDD(VDD),.Y(I3465),.A(n1886gat));
  NOT NOT1_1247(.VSS(VSS),.VDD(VDD),.Y(n3039gat),.A(I3465));
  NOT NOT1_1248(.VSS(VSS),.VDD(VDD),.Y(n1888gat),.A(n3039gat));
  NOT NOT1_1249(.VSS(VSS),.VDD(VDD),.Y(n2048gat),.A(n2994gat));
  NOT NOT1_1250(.VSS(VSS),.VDD(VDD),.Y(I3472),.A(n2539gat));
  NOT NOT1_1251(.VSS(VSS),.VDD(VDD),.Y(n3040gat),.A(I3472));
  NOT NOT1_1252(.VSS(VSS),.VDD(VDD),.Y(n1969gat),.A(n2142gat));
  NOT NOT1_1253(.VSS(VSS),.VDD(VDD),.Y(n1893gat),.A(n2060gat));
  NOT NOT1_1254(.VSS(VSS),.VDD(VDD),.Y(n1892gat),.A(n2993gat));
  NOT NOT1_1255(.VSS(VSS),.VDD(VDD),.Y(I3483),.A(n2436gat));
  NOT NOT1_1256(.VSS(VSS),.VDD(VDD),.Y(n3041gat),.A(I3483));
  NOT NOT1_1257(.VSS(VSS),.VDD(VDD),.Y(n2056gat),.A(n2998gat));
  NOT NOT1_1258(.VSS(VSS),.VDD(VDD),.Y(I3491),.A(n2387gat));
  NOT NOT1_1259(.VSS(VSS),.VDD(VDD),.Y(n3042gat),.A(I3491));
  NOT NOT1_1260(.VSS(VSS),.VDD(VDD),.Y(I3494),.A(n1963gat));
  NOT NOT1_1261(.VSS(VSS),.VDD(VDD),.Y(n3043gat),.A(I3494));
  NOT NOT1_1262(.VSS(VSS),.VDD(VDD),.Y(n1960gat),.A(n3043gat));
  NOT NOT1_1263(.VSS(VSS),.VDD(VDD),.Y(n1887gat),.A(n2138gat));
  NOT NOT1_1264(.VSS(VSS),.VDD(VDD),.Y(n1961gat),.A(n2996gat));
  NOT NOT1_1265(.VSS(VSS),.VDD(VDD),.Y(I3504),.A(n2330gat));
  NOT NOT1_1266(.VSS(VSS),.VDD(VDD),.Y(n3044gat),.A(I3504));
  NOT NOT1_1267(.VSS(VSS),.VDD(VDD),.Y(n2199gat),.A(n2147gat));
  NOT NOT1_1268(.VSS(VSS),.VDD(VDD),.Y(I3509),.A(n2438gat));
  NOT NOT1_1269(.VSS(VSS),.VDD(VDD),.Y(n3045gat),.A(I3509));
  NOT NOT1_1270(.VSS(VSS),.VDD(VDD),.Y(n2332gat),.A(n3045gat));
  NOT NOT1_1271(.VSS(VSS),.VDD(VDD),.Y(I3513),.A(n2439gat));
  NOT NOT1_1272(.VSS(VSS),.VDD(VDD),.Y(n3046gat),.A(I3513));
  NOT NOT1_1273(.VSS(VSS),.VDD(VDD),.Y(n2259gat),.A(n3046gat));
  NOT NOT1_1274(.VSS(VSS),.VDD(VDD),.Y(n2328gat),.A(n3008gat));
  NOT NOT1_1275(.VSS(VSS),.VDD(VDD),.Y(I3520),.A(n2498gat));
  NOT NOT1_1276(.VSS(VSS),.VDD(VDD),.Y(n3047gat),.A(I3520));
  NOT NOT1_1277(.VSS(VSS),.VDD(VDD),.Y(n2151gat),.A(n2193gat));
  NOT NOT1_1278(.VSS(VSS),.VDD(VDD),.Y(n2209gat),.A(n3005gat));
  NOT NOT1_1279(.VSS(VSS),.VDD(VDD),.Y(I3530),.A(n2396gat));
  NOT NOT1_1280(.VSS(VSS),.VDD(VDD),.Y(n3048gat),.A(I3530));
  NOT NOT1_1281(.VSS(VSS),.VDD(VDD),.Y(n2052gat),.A(n2393gat));
  NOT NOT1_1282(.VSS(VSS),.VDD(VDD),.Y(n2058gat),.A(n2997gat));
  NOT NOT1_1283(.VSS(VSS),.VDD(VDD),.Y(I3539),.A(n2198gat));
  NOT NOT1_1284(.VSS(VSS),.VDD(VDD),.Y(n3049gat),.A(I3539));
  NOT NOT1_1285(.VSS(VSS),.VDD(VDD),.Y(n2349gat),.A(n2215gat));
  NOT NOT1_1286(.VSS(VSS),.VDD(VDD),.Y(n2281gat),.A(n3009gat));
  NOT NOT1_1287(.VSS(VSS),.VDD(VDD),.Y(I3549),.A(n2197gat));
  NOT NOT1_1288(.VSS(VSS),.VDD(VDD),.Y(n3050gat),.A(I3549));
  NOT NOT1_1289(.VSS(VSS),.VDD(VDD),.Y(n2146gat),.A(n3002gat));
  NOT NOT1_1290(.VSS(VSS),.VDD(VDD),.Y(I3558),.A(n2196gat));
  NOT NOT1_1291(.VSS(VSS),.VDD(VDD),.Y(n3051gat),.A(I3558));
  NOT NOT1_1292(.VSS(VSS),.VDD(VDD),.Y(n2031gat),.A(n2033gat));
  NOT NOT1_1293(.VSS(VSS),.VDD(VDD),.Y(n2108gat),.A(n2110gat));
  NOT NOT1_1294(.VSS(VSS),.VDD(VDD),.Y(I3587),.A(n2125gat));
  NOT NOT1_1295(.VSS(VSS),.VDD(VDD),.Y(n2124gat),.A(I3587));
  NOT NOT1_1296(.VSS(VSS),.VDD(VDD),.Y(n2123gat),.A(n2125gat));
  NOT NOT1_1297(.VSS(VSS),.VDD(VDD),.Y(n2119gat),.A(n2121gat));
  NOT NOT1_1298(.VSS(VSS),.VDD(VDD),.Y(n2115gat),.A(n2117gat));
  NOT NOT1_1299(.VSS(VSS),.VDD(VDD),.Y(I3610),.A(n1882gat));
  NOT NOT1_1300(.VSS(VSS),.VDD(VDD),.Y(n3052gat),.A(I3610));
  NOT NOT1_1301(.VSS(VSS),.VDD(VDD),.Y(I3621),.A(n1975gat));
  NOT NOT1_1302(.VSS(VSS),.VDD(VDD),.Y(n1974gat),.A(I3621));
  NOT NOT1_1303(.VSS(VSS),.VDD(VDD),.Y(n1955gat),.A(n1956gat));
  NOT NOT1_1304(.VSS(VSS),.VDD(VDD),.Y(n1970gat),.A(n1896gat));
  NOT NOT1_1305(.VSS(VSS),.VDD(VDD),.Y(n1973gat),.A(n1975gat));
  NOT NOT1_1306(.VSS(VSS),.VDD(VDD),.Y(n2558gat),.A(n2559gat));
  NOT NOT1_1307(.VSS(VSS),.VDD(VDD),.Y(I3635),.A(n2558gat));
  NOT NOT1_1308(.VSS(VSS),.VDD(VDD),.Y(n3053gat),.A(I3635));
  NOT NOT1_1309(.VSS(VSS),.VDD(VDD),.Y(I3646),.A(n2644gat));
  NOT NOT1_1310(.VSS(VSS),.VDD(VDD),.Y(n2643gat),.A(I3646));
  NOT NOT1_1311(.VSS(VSS),.VDD(VDD),.Y(n2333gat),.A(n2438gat));
  NOT NOT1_1312(.VSS(VSS),.VDD(VDD),.Y(n2564gat),.A(n2352gat));
  NOT NOT1_1313(.VSS(VSS),.VDD(VDD),.Y(n2642gat),.A(n2644gat));
  NOT NOT1_1314(.VSS(VSS),.VDD(VDD),.Y(n2636gat),.A(n2637gat));
  NOT NOT1_1315(.VSS(VSS),.VDD(VDD),.Y(I3660),.A(n2636gat));
  NOT NOT1_1316(.VSS(VSS),.VDD(VDD),.Y(n3054gat),.A(I3660));
  NOT NOT1_1317(.VSS(VSS),.VDD(VDD),.Y(n88gat),.A(n84gat));
  NOT NOT1_1318(.VSS(VSS),.VDD(VDD),.Y(n375gat),.A(n110gat));
  NOT NOT1_1319(.VSS(VSS),.VDD(VDD),.Y(I3677),.A(n156gat));
  NOT NOT1_1320(.VSS(VSS),.VDD(VDD),.Y(n155gat),.A(I3677));
  NOT NOT1_1321(.VSS(VSS),.VDD(VDD),.Y(n253gat),.A(n1702gat));
  NOT NOT1_1322(.VSS(VSS),.VDD(VDD),.Y(n150gat),.A(n152gat));
  NOT NOT1_1323(.VSS(VSS),.VDD(VDD),.Y(I3691),.A(n152gat));
  NOT NOT1_1324(.VSS(VSS),.VDD(VDD),.Y(n151gat),.A(I3691));
  NOT NOT1_1325(.VSS(VSS),.VDD(VDD),.Y(n243gat),.A(n1702gat));
  NOT NOT1_1326(.VSS(VSS),.VDD(VDD),.Y(n233gat),.A(n243gat));
  NOT NOT1_1327(.VSS(VSS),.VDD(VDD),.Y(n154gat),.A(n156gat));
  NOT NOT1_1328(.VSS(VSS),.VDD(VDD),.Y(n800gat),.A(n2874gat));
  NOT NOT1_1329(.VSS(VSS),.VDD(VDD),.Y(I3703),.A(n2917gat));
  NOT NOT1_1330(.VSS(VSS),.VDD(VDD),.Y(n3055gat),.A(I3703));
  NOT NOT1_1331(.VSS(VSS),.VDD(VDD),.Y(n235gat),.A(n2878gat));
  NOT NOT1_1332(.VSS(VSS),.VDD(VDD),.Y(I3713),.A(n2892gat));
  NOT NOT1_1333(.VSS(VSS),.VDD(VDD),.Y(n3056gat),.A(I3713));
  NOT NOT1_1334(.VSS(VSS),.VDD(VDD),.Y(n372gat),.A(n212gat));
  NOT NOT1_1335(.VSS(VSS),.VDD(VDD),.Y(n329gat),.A(n331gat));
  NOT NOT1_1336(.VSS(VSS),.VDD(VDD),.Y(I3736),.A(n388gat));
  NOT NOT1_1337(.VSS(VSS),.VDD(VDD),.Y(n387gat),.A(I3736));
  NOT NOT1_1338(.VSS(VSS),.VDD(VDD),.Y(n334gat),.A(n1700gat));
  NOT NOT1_1339(.VSS(VSS),.VDD(VDD),.Y(n386gat),.A(n388gat));
  NOT NOT1_1340(.VSS(VSS),.VDD(VDD),.Y(I3742),.A(n331gat));
  NOT NOT1_1341(.VSS(VSS),.VDD(VDD),.Y(n330gat),.A(I3742));
  NOT NOT1_1342(.VSS(VSS),.VDD(VDD),.Y(n1430gat),.A(n1700gat));
  NOT NOT1_1343(.VSS(VSS),.VDD(VDD),.Y(n1490gat),.A(n1430gat));
  NOT NOT1_1344(.VSS(VSS),.VDD(VDD),.Y(n452gat),.A(n2885gat));
  NOT NOT1_1345(.VSS(VSS),.VDD(VDD),.Y(I3754),.A(n2900gat));
  NOT NOT1_1346(.VSS(VSS),.VDD(VDD),.Y(n3057gat),.A(I3754));
  NOT NOT1_1347(.VSS(VSS),.VDD(VDD),.Y(n333gat),.A(n2883gat));
  NOT NOT1_1348(.VSS(VSS),.VDD(VDD),.Y(I3765),.A(n2929gat));
  NOT NOT1_1349(.VSS(VSS),.VDD(VDD),.Y(n3058gat),.A(I3765));
  NOT NOT1_1350(.VSS(VSS),.VDD(VDD),.Y(I3777),.A(n463gat));
  NOT NOT1_1351(.VSS(VSS),.VDD(VDD),.Y(n462gat),.A(I3777));
  NOT NOT1_1352(.VSS(VSS),.VDD(VDD),.Y(n325gat),.A(n327gat));
  NOT NOT1_1353(.VSS(VSS),.VDD(VDD),.Y(n457gat),.A(n2884gat));
  NOT NOT1_1354(.VSS(VSS),.VDD(VDD),.Y(n461gat),.A(n463gat));
  NOT NOT1_1355(.VSS(VSS),.VDD(VDD),.Y(n458gat),.A(n2902gat));
  NOT NOT1_1356(.VSS(VSS),.VDD(VDD),.Y(I3801),.A(n2925gat));
  NOT NOT1_1357(.VSS(VSS),.VDD(VDD),.Y(n3059gat),.A(I3801));
  NOT NOT1_1358(.VSS(VSS),.VDD(VDD),.Y(n144gat),.A(n247gat));
  NOT NOT1_1359(.VSS(VSS),.VDD(VDD),.Y(I3808),.A(n327gat));
  NOT NOT1_1360(.VSS(VSS),.VDD(VDD),.Y(n326gat),.A(I3808));
  NOT NOT1_1361(.VSS(VSS),.VDD(VDD),.Y(n878gat),.A(n2879gat));
  NOT NOT1_1362(.VSS(VSS),.VDD(VDD),.Y(I3817),.A(n2916gat));
  NOT NOT1_1363(.VSS(VSS),.VDD(VDD),.Y(n3060gat),.A(I3817));
  NOT NOT1_1364(.VSS(VSS),.VDD(VDD),.Y(n382gat),.A(n384gat));
  NOT NOT1_1365(.VSS(VSS),.VDD(VDD),.Y(I3831),.A(n384gat));
  NOT NOT1_1366(.VSS(VSS),.VDD(VDD),.Y(n383gat),.A(I3831));
  NOT NOT1_1367(.VSS(VSS),.VDD(VDD),.Y(n134gat),.A(n2875gat));
  NOT NOT1_1368(.VSS(VSS),.VDD(VDD),.Y(I3841),.A(n2899gat));
  NOT NOT1_1369(.VSS(VSS),.VDD(VDD),.Y(n3061gat),.A(I3841));
  NOT NOT1_1370(.VSS(VSS),.VDD(VDD),.Y(n254gat),.A(n256gat));
  NOT NOT1_1371(.VSS(VSS),.VDD(VDD),.Y(n252gat),.A(n2877gat));
  NOT NOT1_1372(.VSS(VSS),.VDD(VDD),.Y(n468gat),.A(n470gat));
  NOT NOT1_1373(.VSS(VSS),.VDD(VDD),.Y(I3867),.A(n470gat));
  NOT NOT1_1374(.VSS(VSS),.VDD(VDD),.Y(n469gat),.A(I3867));
  NOT NOT1_1375(.VSS(VSS),.VDD(VDD),.Y(n381gat),.A(n2893gat));
  NOT NOT1_1376(.VSS(VSS),.VDD(VDD),.Y(I3876),.A(n2926gat));
  NOT NOT1_1377(.VSS(VSS),.VDD(VDD),.Y(n3062gat),.A(I3876));
  NOT NOT1_1378(.VSS(VSS),.VDD(VDD),.Y(n241gat),.A(n140gat));
  NOT NOT1_1379(.VSS(VSS),.VDD(VDD),.Y(I3882),.A(n256gat));
  NOT NOT1_1380(.VSS(VSS),.VDD(VDD),.Y(n255gat),.A(I3882));
  NOT NOT1_1381(.VSS(VSS),.VDD(VDD),.Y(n802gat),.A(n2882gat));
  NOT NOT1_1382(.VSS(VSS),.VDD(VDD),.Y(I3891),.A(n2924gat));
  NOT NOT1_1383(.VSS(VSS),.VDD(VDD),.Y(n3063gat),.A(I3891));
  NOT NOT1_1384(.VSS(VSS),.VDD(VDD),.Y(n146gat),.A(n148gat));
  NOT NOT1_1385(.VSS(VSS),.VDD(VDD),.Y(I3904),.A(n148gat));
  NOT NOT1_1386(.VSS(VSS),.VDD(VDD),.Y(n147gat),.A(I3904));
  NOT NOT1_1387(.VSS(VSS),.VDD(VDD),.Y(n380gat),.A(n2881gat));
  NOT NOT1_1388(.VSS(VSS),.VDD(VDD),.Y(I3914),.A(n2923gat));
  NOT NOT1_1389(.VSS(VSS),.VDD(VDD),.Y(n3064gat),.A(I3914));
  NOT NOT1_1390(.VSS(VSS),.VDD(VDD),.Y(n69gat),.A(n68gat));
  NOT NOT1_1391(.VSS(VSS),.VDD(VDD),.Y(n1885gat),.A(n2048gat));
  NOT NOT1_1392(.VSS(VSS),.VDD(VDD),.Y(I3923),.A(n2710gat));
  NOT NOT1_1393(.VSS(VSS),.VDD(VDD),.Y(n2707gat),.A(I3923));
  NOT NOT1_1394(.VSS(VSS),.VDD(VDD),.Y(n16gat),.A(n564gat));
  NOT NOT1_1395(.VSS(VSS),.VDD(VDD),.Y(n295gat),.A(n357gat));
  NOT NOT1_1396(.VSS(VSS),.VDD(VDD),.Y(n11gat),.A(n12gat));
  NOT NOT1_1397(.VSS(VSS),.VDD(VDD),.Y(n1889gat),.A(n1961gat));
  NOT NOT1_1398(.VSS(VSS),.VDD(VDD),.Y(I3935),.A(n2704gat));
  NOT NOT1_1399(.VSS(VSS),.VDD(VDD),.Y(n2700gat),.A(I3935));
  NOT NOT1_1400(.VSS(VSS),.VDD(VDD),.Y(n2051gat),.A(n2056gat));
  NOT NOT1_1401(.VSS(VSS),.VDD(VDD),.Y(I3941),.A(n2684gat));
  NOT NOT1_1402(.VSS(VSS),.VDD(VDD),.Y(n2680gat),.A(I3941));
  NOT NOT1_1403(.VSS(VSS),.VDD(VDD),.Y(n1350gat),.A(n1831gat));
  NOT NOT1_1404(.VSS(VSS),.VDD(VDD),.Y(I3945),.A(n1350gat));
  NOT NOT1_1405(.VSS(VSS),.VDD(VDD),.Y(n2696gat),.A(I3945));
  NOT NOT1_1406(.VSS(VSS),.VDD(VDD),.Y(I3948),.A(n2696gat));
  NOT NOT1_1407(.VSS(VSS),.VDD(VDD),.Y(n2692gat),.A(I3948));
  NOT NOT1_1408(.VSS(VSS),.VDD(VDD),.Y(I3951),.A(n2448gat));
  NOT NOT1_1409(.VSS(VSS),.VDD(VDD),.Y(n2683gat),.A(I3951));
  NOT NOT1_1410(.VSS(VSS),.VDD(VDD),.Y(I3954),.A(n2683gat));
  NOT NOT1_1411(.VSS(VSS),.VDD(VDD),.Y(n2679gat),.A(I3954));
  NOT NOT1_1412(.VSS(VSS),.VDD(VDD),.Y(I3957),.A(n2450gat));
  NOT NOT1_1413(.VSS(VSS),.VDD(VDD),.Y(n2449gat),.A(I3957));
  NOT NOT1_1414(.VSS(VSS),.VDD(VDD),.Y(n1754gat),.A(n2449gat));
  NOT NOT1_1415(.VSS(VSS),.VDD(VDD),.Y(I3962),.A(n2830gat));
  NOT NOT1_1416(.VSS(VSS),.VDD(VDD),.Y(n2827gat),.A(I3962));
  NOT NOT1_1417(.VSS(VSS),.VDD(VDD),.Y(n2590gat),.A(n2592gat));
  NOT NOT1_1418(.VSS(VSS),.VDD(VDD),.Y(n2456gat),.A(n2458gat));
  NOT NOT1_1419(.VSS(VSS),.VDD(VDD),.Y(n2512gat),.A(n2514gat));
  NOT NOT1_1420(.VSS(VSS),.VDD(VDD),.Y(n1544gat),.A(n1625gat));
  NOT NOT1_1421(.VSS(VSS),.VDD(VDD),.Y(n1769gat),.A(n1771gat));
  NOT NOT1_1422(.VSS(VSS),.VDD(VDD),.Y(n1683gat),.A(n1756gat));
  NOT NOT1_1423(.VSS(VSS),.VDD(VDD),.Y(n2167gat),.A(n2169gat));
  NOT NOT1_1424(.VSS(VSS),.VDD(VDD),.Y(n2013gat),.A(I4000));
  NOT NOT1_1425(.VSS(VSS),.VDD(VDD),.Y(n1791gat),.A(n2013gat));
  NOT NOT1_1426(.VSS(VSS),.VDD(VDD),.Y(n2691gat),.A(n2695gat));
  NOT NOT1_1427(.VSS(VSS),.VDD(VDD),.Y(n1518gat),.A(n1694gat));
  NOT NOT1_1428(.VSS(VSS),.VDD(VDD),.Y(n2699gat),.A(n2703gat));
  NOT NOT1_1429(.VSS(VSS),.VDD(VDD),.Y(n2159gat),.A(n1412gat));
  NOT NOT1_1430(.VSS(VSS),.VDD(VDD),.Y(n2478gat),.A(n2579gat));
  NOT NOT1_1431(.VSS(VSS),.VDD(VDD),.Y(I4014),.A(n2744gat));
  NOT NOT1_1432(.VSS(VSS),.VDD(VDD),.Y(n2740gat),.A(I4014));
  NOT NOT1_1433(.VSS(VSS),.VDD(VDD),.Y(n2158gat),.A(n1412gat));
  NOT NOT1_1434(.VSS(VSS),.VDD(VDD),.Y(n2186gat),.A(n2613gat));
  NOT NOT1_1435(.VSS(VSS),.VDD(VDD),.Y(I4020),.A(n2800gat));
  NOT NOT1_1436(.VSS(VSS),.VDD(VDD),.Y(n2797gat),.A(I4020));
  NOT NOT1_1437(.VSS(VSS),.VDD(VDD),.Y(n2288gat),.A(I4024));
  NOT NOT1_1438(.VSS(VSS),.VDD(VDD),.Y(n1513gat),.A(n2288gat));
  NOT NOT1_1439(.VSS(VSS),.VDD(VDD),.Y(n2537gat),.A(n2538gat));
  NOT NOT1_1440(.VSS(VSS),.VDD(VDD),.Y(n2442gat),.A(n2483gat));
  NOT NOT1_1441(.VSS(VSS),.VDD(VDD),.Y(n1334gat),.A(n1336gat));
  NOT NOT1_1442(.VSS(VSS),.VDD(VDD),.Y(I4055),.A(n1748gat));
  NOT NOT1_1443(.VSS(VSS),.VDD(VDD),.Y(n1747gat),.A(I4055));
  NOT NOT1_1444(.VSS(VSS),.VDD(VDD),.Y(I4067),.A(n1675gat));
  NOT NOT1_1445(.VSS(VSS),.VDD(VDD),.Y(n1674gat),.A(I4067));
  NOT NOT1_1446(.VSS(VSS),.VDD(VDD),.Y(n1403gat),.A(n1402gat));
  NOT NOT1_1447(.VSS(VSS),.VDD(VDD),.Y(I4081),.A(n1807gat));
  NOT NOT1_1448(.VSS(VSS),.VDD(VDD),.Y(n1806gat),.A(I4081));
  NOT NOT1_1449(.VSS(VSS),.VDD(VDD),.Y(n1634gat),.A(n1712gat));
  NOT NOT1_1450(.VSS(VSS),.VDD(VDD),.Y(n1338gat),.A(n1340gat));
  NOT NOT1_1451(.VSS(VSS),.VDD(VDD),.Y(I4105),.A(n1456gat));
  NOT NOT1_1452(.VSS(VSS),.VDD(VDD),.Y(n1455gat),.A(I4105));
  NOT NOT1_1453(.VSS(VSS),.VDD(VDD),.Y(I4108),.A(n1340gat));
  NOT NOT1_1454(.VSS(VSS),.VDD(VDD),.Y(n1339gat),.A(I4108));
  NOT NOT1_1455(.VSS(VSS),.VDD(VDD),.Y(n1505gat),.A(n2980gat));
  NOT NOT1_1456(.VSS(VSS),.VDD(VDD),.Y(I4117),.A(n1505gat));
  NOT NOT1_1457(.VSS(VSS),.VDD(VDD),.Y(n2758gat),.A(I4117));
  NOT NOT1_1458(.VSS(VSS),.VDD(VDD),.Y(n2755gat),.A(n2758gat));
  NOT NOT1_1459(.VSS(VSS),.VDD(VDD),.Y(n1546gat),.A(n2980gat));
  NOT NOT1_1460(.VSS(VSS),.VDD(VDD),.Y(I4122),.A(n1546gat));
  NOT NOT1_1461(.VSS(VSS),.VDD(VDD),.Y(n2752gat),.A(I4122));
  NOT NOT1_1462(.VSS(VSS),.VDD(VDD),.Y(n2748gat),.A(n2752gat));
  NOT NOT1_1463(.VSS(VSS),.VDD(VDD),.Y(n2012gat),.A(n2016gat));
  NOT NOT1_1464(.VSS(VSS),.VDD(VDD),.Y(n2002gat),.A(n2008gat));
  NOT NOT1_1465(.VSS(VSS),.VDD(VDD),.Y(I4129),.A(n3097gat));
  NOT NOT1_1466(.VSS(VSS),.VDD(VDD),.Y(n2858gat),.A(I4129));
  NOT NOT1_1467(.VSS(VSS),.VDD(VDD),.Y(n2857gat),.A(n2858gat));
  NOT NOT1_1468(.VSS(VSS),.VDD(VDD),.Y(I4135),.A(n3098gat));
  NOT NOT1_1469(.VSS(VSS),.VDD(VDD),.Y(n2766gat),.A(I4135));
  NOT NOT1_1470(.VSS(VSS),.VDD(VDD),.Y(I4138),.A(n2766gat));
  NOT NOT1_1471(.VSS(VSS),.VDD(VDD),.Y(n2765gat),.A(I4138));
  NOT NOT1_1472(.VSS(VSS),.VDD(VDD),.Y(n1684gat),.A(n1759gat));
  NOT NOT1_1473(.VSS(VSS),.VDD(VDD),.Y(n1632gat),.A(I4145));
  NOT NOT1_1474(.VSS(VSS),.VDD(VDD),.Y(I4157),.A(n1525gat));
  NOT NOT1_1475(.VSS(VSS),.VDD(VDD),.Y(n1524gat),.A(I4157));
  NOT NOT1_1476(.VSS(VSS),.VDD(VDD),.Y(n1862gat),.A(n1863gat));
  NOT NOT1_1477(.VSS(VSS),.VDD(VDD),.Y(n1919gat),.A(n1860gat));
  NOT NOT1_1478(.VSS(VSS),.VDD(VDD),.Y(n1460gat),.A(n1462gat));
  NOT NOT1_1479(.VSS(VSS),.VDD(VDD),.Y(I4185),.A(n1596gat));
  NOT NOT1_1480(.VSS(VSS),.VDD(VDD),.Y(n1595gat),.A(I4185));
  NOT NOT1_1481(.VSS(VSS),.VDD(VDD),.Y(n1454gat),.A(n1469gat));
  NOT NOT1_1482(.VSS(VSS),.VDD(VDD),.Y(n1468gat),.A(n1519gat));
  NOT NOT1_1483(.VSS(VSS),.VDD(VDD),.Y(I4194),.A(n1462gat));
  NOT NOT1_1484(.VSS(VSS),.VDD(VDD),.Y(n1461gat),.A(I4194));
  NOT NOT1_1485(.VSS(VSS),.VDD(VDD),.Y(n1477gat),.A(n2984gat));
  NOT NOT1_1486(.VSS(VSS),.VDD(VDD),.Y(n1594gat),.A(n1596gat));
  NOT NOT1_1487(.VSS(VSS),.VDD(VDD),.Y(I4212),.A(n1588gat));
  NOT NOT1_1488(.VSS(VSS),.VDD(VDD),.Y(n1587gat),.A(I4212));
  NOT NOT1_1489(.VSS(VSS),.VDD(VDD),.Y(n1681gat),.A(I4217));
  NOT NOT1_1490(.VSS(VSS),.VDD(VDD),.Y(I4222),.A(n1761gat));
  NOT NOT1_1491(.VSS(VSS),.VDD(VDD),.Y(n2751gat),.A(I4222));
  NOT NOT1_1492(.VSS(VSS),.VDD(VDD),.Y(n2747gat),.A(n2751gat));
  NOT NOT1_1493(.VSS(VSS),.VDD(VDD),.Y(I4227),.A(n1760gat));
  NOT NOT1_1494(.VSS(VSS),.VDD(VDD),.Y(n2743gat),.A(I4227));
  NOT NOT1_1495(.VSS(VSS),.VDD(VDD),.Y(n2739gat),.A(n2743gat));
  NOT NOT1_1496(.VSS(VSS),.VDD(VDD),.Y(n1978gat),.A(n2286gat));
  NOT NOT1_1497(.VSS(VSS),.VDD(VDD),.Y(I4233),.A(n1721gat));
  NOT NOT1_1498(.VSS(VSS),.VDD(VDD),.Y(n2808gat),.A(I4233));
  NOT NOT1_1499(.VSS(VSS),.VDD(VDD),.Y(I4236),.A(n2808gat));
  NOT NOT1_1500(.VSS(VSS),.VDD(VDD),.Y(n2804gat),.A(I4236));
  NOT NOT1_1501(.VSS(VSS),.VDD(VDD),.Y(n517gat),.A(n518gat));
  NOT NOT1_1502(.VSS(VSS),.VDD(VDD),.Y(n417gat),.A(n418gat));
  NOT NOT1_1503(.VSS(VSS),.VDD(VDD),.Y(n413gat),.A(n411gat));
  NOT NOT1_1504(.VSS(VSS),.VDD(VDD),.Y(n412gat),.A(n522gat));
  NOT NOT1_1505(.VSS(VSS),.VDD(VDD),.Y(n406gat),.A(n516gat));
  NOT NOT1_1506(.VSS(VSS),.VDD(VDD),.Y(n407gat),.A(n355gat));
  NOT NOT1_1507(.VSS(VSS),.VDD(VDD),.Y(n290gat),.A(n525gat));
  NOT NOT1_1508(.VSS(VSS),.VDD(VDD),.Y(n527gat),.A(n356gat));
  NOT NOT1_1509(.VSS(VSS),.VDD(VDD),.Y(n416gat),.A(n415gat));
  NOT NOT1_1510(.VSS(VSS),.VDD(VDD),.Y(n528gat),.A(n521gat));
  NOT NOT1_1511(.VSS(VSS),.VDD(VDD),.Y(n358gat),.A(n532gat));
  NOT NOT1_1512(.VSS(VSS),.VDD(VDD),.Y(n639gat),.A(n523gat));
  NOT NOT1_1513(.VSS(VSS),.VDD(VDD),.Y(n1111gat),.A(n635gat));
  NOT NOT1_1514(.VSS(VSS),.VDD(VDD),.Y(n524gat),.A(n414gat));
  NOT NOT1_1515(.VSS(VSS),.VDD(VDD),.Y(n1112gat),.A(n630gat));
  NOT NOT1_1516(.VSS(VSS),.VDD(VDD),.Y(n741gat),.A(n629gat));
  NOT NOT1_1517(.VSS(VSS),.VDD(VDD),.Y(n633gat),.A(n634gat));
  NOT NOT1_1518(.VSS(VSS),.VDD(VDD),.Y(n926gat),.A(n632gat));
  NOT NOT1_1519(.VSS(VSS),.VDD(VDD),.Y(n670gat),.A(n636gat));
  NOT NOT1_1520(.VSS(VSS),.VDD(VDD),.Y(n1123gat),.A(n632gat));
  NOT NOT1_1521(.VSS(VSS),.VDD(VDD),.Y(n1007gat),.A(n635gat));
  NOT NOT1_1522(.VSS(VSS),.VDD(VDD),.Y(n1006gat),.A(n630gat));
  NOT NOT1_1523(.VSS(VSS),.VDD(VDD),.Y(I4309),.A(n2941gat));
  NOT NOT1_1524(.VSS(VSS),.VDD(VDD),.Y(n2814gat),.A(I4309));
  NOT NOT1_1525(.VSS(VSS),.VDD(VDD),.Y(I4312),.A(n2814gat));
  NOT NOT1_1526(.VSS(VSS),.VDD(VDD),.Y(n2811gat),.A(I4312));
  NOT NOT1_1527(.VSS(VSS),.VDD(VDD),.Y(n1002gat),.A(n2946gat));
  NOT NOT1_1528(.VSS(VSS),.VDD(VDD),.Y(I4329),.A(n2950gat));
  NOT NOT1_1529(.VSS(VSS),.VDD(VDD),.Y(n2813gat),.A(I4329));
  NOT NOT1_1530(.VSS(VSS),.VDD(VDD),.Y(I4332),.A(n2813gat));
  NOT NOT1_1531(.VSS(VSS),.VDD(VDD),.Y(n2810gat),.A(I4332));
  NOT NOT1_1532(.VSS(VSS),.VDD(VDD),.Y(n888gat),.A(n2933gat));
  NOT NOT1_1533(.VSS(VSS),.VDD(VDD),.Y(I4349),.A(n2935gat));
  NOT NOT1_1534(.VSS(VSS),.VDD(VDD),.Y(n2818gat),.A(I4349));
  NOT NOT1_1535(.VSS(VSS),.VDD(VDD),.Y(I4352),.A(n2818gat));
  NOT NOT1_1536(.VSS(VSS),.VDD(VDD),.Y(n2816gat),.A(I4352));
  NOT NOT1_1537(.VSS(VSS),.VDD(VDD),.Y(n898gat),.A(n2940gat));
  NOT NOT1_1538(.VSS(VSS),.VDD(VDD),.Y(I4369),.A(n2937gat));
  NOT NOT1_1539(.VSS(VSS),.VDD(VDD),.Y(n2817gat),.A(I4369));
  NOT NOT1_1540(.VSS(VSS),.VDD(VDD),.Y(I4372),.A(n2817gat));
  NOT NOT1_1541(.VSS(VSS),.VDD(VDD),.Y(n2815gat),.A(I4372));
  NOT NOT1_1542(.VSS(VSS),.VDD(VDD),.Y(n1179gat),.A(n2947gat));
  NOT NOT1_1543(.VSS(VSS),.VDD(VDD),.Y(I4389),.A(n2956gat));
  NOT NOT1_1544(.VSS(VSS),.VDD(VDD),.Y(n2824gat),.A(I4389));
  NOT NOT1_1545(.VSS(VSS),.VDD(VDD),.Y(I4392),.A(n2824gat));
  NOT NOT1_1546(.VSS(VSS),.VDD(VDD),.Y(n2821gat),.A(I4392));
  NOT NOT1_1547(.VSS(VSS),.VDD(VDD),.Y(n897gat),.A(n2939gat));
  NOT NOT1_1548(.VSS(VSS),.VDD(VDD),.Y(I4409),.A(n2938gat));
  NOT NOT1_1549(.VSS(VSS),.VDD(VDD),.Y(n2823gat),.A(I4409));
  NOT NOT1_1550(.VSS(VSS),.VDD(VDD),.Y(I4412),.A(n2823gat));
  NOT NOT1_1551(.VSS(VSS),.VDD(VDD),.Y(n2820gat),.A(I4412));
  NOT NOT1_1552(.VSS(VSS),.VDD(VDD),.Y(n894gat),.A(n2932gat));
  NOT NOT1_1553(.VSS(VSS),.VDD(VDD),.Y(I4429),.A(n2936gat));
  NOT NOT1_1554(.VSS(VSS),.VDD(VDD),.Y(n2829gat),.A(I4429));
  NOT NOT1_1555(.VSS(VSS),.VDD(VDD),.Y(I4432),.A(n2829gat));
  NOT NOT1_1556(.VSS(VSS),.VDD(VDD),.Y(n2826gat),.A(I4432));
  NOT NOT1_1557(.VSS(VSS),.VDD(VDD),.Y(n1180gat),.A(n2948gat));
  NOT NOT1_1558(.VSS(VSS),.VDD(VDD),.Y(I4449),.A(n2955gat));
  NOT NOT1_1559(.VSS(VSS),.VDD(VDD),.Y(n2828gat),.A(I4449));
  NOT NOT1_1560(.VSS(VSS),.VDD(VDD),.Y(I4452),.A(n2828gat));
  NOT NOT1_1561(.VSS(VSS),.VDD(VDD),.Y(n2825gat),.A(I4452));
  NOT NOT1_1562(.VSS(VSS),.VDD(VDD),.Y(n671gat),.A(n673gat));
  NOT NOT1_1563(.VSS(VSS),.VDD(VDD),.Y(n628gat),.A(n631gat));
  NOT NOT1_1564(.VSS(VSS),.VDD(VDD),.Y(n976gat),.A(n628gat));
  NOT NOT1_1565(.VSS(VSS),.VDD(VDD),.Y(I4475),.A(n2951gat));
  NOT NOT1_1566(.VSS(VSS),.VDD(VDD),.Y(n2807gat),.A(I4475));
  NOT NOT1_1567(.VSS(VSS),.VDD(VDD),.Y(I4478),.A(n2807gat));
  NOT NOT1_1568(.VSS(VSS),.VDD(VDD),.Y(n2803gat),.A(I4478));
  NOT NOT1_1569(.VSS(VSS),.VDD(VDD),.Y(n2127gat),.A(n2389gat));
  NOT NOT1_1570(.VSS(VSS),.VDD(VDD),.Y(I4482),.A(n2127gat));
  NOT NOT1_1571(.VSS(VSS),.VDD(VDD),.Y(n2682gat),.A(I4482));
  NOT NOT1_1572(.VSS(VSS),.VDD(VDD),.Y(I4485),.A(n2682gat));
  NOT NOT1_1573(.VSS(VSS),.VDD(VDD),.Y(n2678gat),.A(I4485));
  NOT NOT1_1574(.VSS(VSS),.VDD(VDD),.Y(n2046gat),.A(n2269gat));
  NOT NOT1_1575(.VSS(VSS),.VDD(VDD),.Y(I4489),.A(n2046gat));
  NOT NOT1_1576(.VSS(VSS),.VDD(VDD),.Y(n2681gat),.A(I4489));
  NOT NOT1_1577(.VSS(VSS),.VDD(VDD),.Y(I4492),.A(n2681gat));
  NOT NOT1_1578(.VSS(VSS),.VDD(VDD),.Y(n2677gat),.A(I4492));
  NOT NOT1_1579(.VSS(VSS),.VDD(VDD),.Y(n1708gat),.A(n2338gat));
  NOT NOT1_1580(.VSS(VSS),.VDD(VDD),.Y(I4496),.A(n1708gat));
  NOT NOT1_1581(.VSS(VSS),.VDD(VDD),.Y(n2688gat),.A(I4496));
  NOT NOT1_1582(.VSS(VSS),.VDD(VDD),.Y(I4499),.A(n2688gat));
  NOT NOT1_1583(.VSS(VSS),.VDD(VDD),.Y(n2686gat),.A(I4499));
  NOT NOT1_1584(.VSS(VSS),.VDD(VDD),.Y(n455gat),.A(n291gat));
  NOT NOT1_1585(.VSS(VSS),.VDD(VDD),.Y(n2237gat),.A(n2646gat));
  NOT NOT1_1586(.VSS(VSS),.VDD(VDD),.Y(I4506),.A(n2764gat));
  NOT NOT1_1587(.VSS(VSS),.VDD(VDD),.Y(n2763gat),.A(I4506));
  NOT NOT1_1588(.VSS(VSS),.VDD(VDD),.Y(n1782gat),.A(n2971gat));
  NOT NOT1_1589(.VSS(VSS),.VDD(VDD),.Y(I4512),.A(n2762gat));
  NOT NOT1_1590(.VSS(VSS),.VDD(VDD),.Y(n2760gat),.A(I4512));
  NOT NOT1_1591(.VSS(VSS),.VDD(VDD),.Y(n2325gat),.A(n3010gat));
  NOT NOT1_1592(.VSS(VSS),.VDD(VDD),.Y(I4518),.A(n2761gat));
  NOT NOT1_1593(.VSS(VSS),.VDD(VDD),.Y(n2759gat),.A(I4518));
  NOT NOT1_1594(.VSS(VSS),.VDD(VDD),.Y(n2245gat),.A(n504gat));
  NOT NOT1_1595(.VSS(VSS),.VDD(VDD),.Y(I4524),.A(n2757gat));
  NOT NOT1_1596(.VSS(VSS),.VDD(VDD),.Y(n2754gat),.A(I4524));
  NOT NOT1_1597(.VSS(VSS),.VDD(VDD),.Y(n2244gat),.A(n567gat));
  NOT NOT1_1598(.VSS(VSS),.VDD(VDD),.Y(I4530),.A(n2756gat));
  NOT NOT1_1599(.VSS(VSS),.VDD(VDD),.Y(n2753gat),.A(I4530));
  NOT NOT1_1600(.VSS(VSS),.VDD(VDD),.Y(n2243gat),.A(n55gat));
  NOT NOT1_1601(.VSS(VSS),.VDD(VDD),.Y(I4536),.A(n2750gat));
  NOT NOT1_1602(.VSS(VSS),.VDD(VDD),.Y(n2746gat),.A(I4536));
  NOT NOT1_1603(.VSS(VSS),.VDD(VDD),.Y(n2246gat),.A(n933gat));
  NOT NOT1_1604(.VSS(VSS),.VDD(VDD),.Y(I4542),.A(n2749gat));
  NOT NOT1_1605(.VSS(VSS),.VDD(VDD),.Y(n2745gat),.A(I4542));
  NOT NOT1_1606(.VSS(VSS),.VDD(VDD),.Y(n2384gat),.A(n43gat));
  NOT NOT1_1607(.VSS(VSS),.VDD(VDD),.Y(I4548),.A(n2742gat));
  NOT NOT1_1608(.VSS(VSS),.VDD(VDD),.Y(n2738gat),.A(I4548));
  NOT NOT1_1609(.VSS(VSS),.VDD(VDD),.Y(n2385gat),.A(n748gat));
  NOT NOT1_1610(.VSS(VSS),.VDD(VDD),.Y(I4554),.A(n2741gat));
  NOT NOT1_1611(.VSS(VSS),.VDD(VDD),.Y(n2737gat),.A(I4554));
  NOT NOT1_1612(.VSS(VSS),.VDD(VDD),.Y(n1286gat),.A(n1269gat));
  NOT NOT1_1613(.VSS(VSS),.VDD(VDD),.Y(I4558),.A(n1286gat));
  NOT NOT1_1614(.VSS(VSS),.VDD(VDD),.Y(n2687gat),.A(I4558));
  NOT NOT1_1615(.VSS(VSS),.VDD(VDD),.Y(n2685gat),.A(n2687gat));
  NOT NOT1_1616(.VSS(VSS),.VDD(VDD),.Y(n1328gat),.A(n1224gat));
  NOT NOT1_1617(.VSS(VSS),.VDD(VDD),.Y(n1381gat),.A(n1328gat));
  NOT NOT1_1618(.VSS(VSS),.VDD(VDD),.Y(n1384gat),.A(n2184gat));
  NOT NOT1_1619(.VSS(VSS),.VDD(VDD),.Y(I4566),.A(n2694gat));
  NOT NOT1_1620(.VSS(VSS),.VDD(VDD),.Y(n2690gat),.A(I4566));
  NOT NOT1_1621(.VSS(VSS),.VDD(VDD),.Y(n1382gat),.A(n1280gat));
  NOT NOT1_1622(.VSS(VSS),.VDD(VDD),.Y(n1451gat),.A(n1382gat));
  NOT NOT1_1623(.VSS(VSS),.VDD(VDD),.Y(n1453gat),.A(n2187gat));
  NOT NOT1_1624(.VSS(VSS),.VDD(VDD),.Y(I4573),.A(n2693gat));
  NOT NOT1_1625(.VSS(VSS),.VDD(VDD),.Y(n2689gat),.A(I4573));
  NOT NOT1_1626(.VSS(VSS),.VDD(VDD),.Y(n927gat),.A(n1133gat));
  NOT NOT1_1627(.VSS(VSS),.VDD(VDD),.Y(n925gat),.A(n927gat));
  NOT NOT1_1628(.VSS(VSS),.VDD(VDD),.Y(n1452gat),.A(n2049gat));
  NOT NOT1_1629(.VSS(VSS),.VDD(VDD),.Y(I4580),.A(n2702gat));
  NOT NOT1_1630(.VSS(VSS),.VDD(VDD),.Y(n2698gat),.A(I4580));
  NOT NOT1_1631(.VSS(VSS),.VDD(VDD),.Y(n923gat),.A(n1043gat));
  NOT NOT1_1632(.VSS(VSS),.VDD(VDD),.Y(n921gat),.A(n923gat));
  NOT NOT1_1633(.VSS(VSS),.VDD(VDD),.Y(n1890gat),.A(n2328gat));
  NOT NOT1_1634(.VSS(VSS),.VDD(VDD),.Y(I4587),.A(n2701gat));
  NOT NOT1_1635(.VSS(VSS),.VDD(VDD),.Y(n2697gat),.A(I4587));
  NOT NOT1_1636(.VSS(VSS),.VDD(VDD),.Y(n850gat),.A(n929gat));
  NOT NOT1_1637(.VSS(VSS),.VDD(VDD),.Y(n739gat),.A(n850gat));
  NOT NOT1_1638(.VSS(VSS),.VDD(VDD),.Y(n1841gat),.A(n2058gat));
  NOT NOT1_1639(.VSS(VSS),.VDD(VDD),.Y(I4594),.A(n2709gat));
  NOT NOT1_1640(.VSS(VSS),.VDD(VDD),.Y(n2706gat),.A(I4594));
  NOT NOT1_1641(.VSS(VSS),.VDD(VDD),.Y(n922gat),.A(n1119gat));
  NOT NOT1_1642(.VSS(VSS),.VDD(VDD),.Y(n848gat),.A(n922gat));
  NOT NOT1_1643(.VSS(VSS),.VDD(VDD),.Y(n2047gat),.A(n2209gat));
  NOT NOT1_1644(.VSS(VSS),.VDD(VDD),.Y(I4601),.A(n2708gat));
  NOT NOT1_1645(.VSS(VSS),.VDD(VDD),.Y(n2705gat),.A(I4601));
  NOT NOT1_1646(.VSS(VSS),.VDD(VDD),.Y(n924gat),.A(n1070gat));
  NOT NOT1_1647(.VSS(VSS),.VDD(VDD),.Y(n849gat),.A(n924gat));
  NOT NOT1_1648(.VSS(VSS),.VDD(VDD),.Y(n2050gat),.A(n2146gat));
  NOT NOT1_1649(.VSS(VSS),.VDD(VDD),.Y(I4608),.A(n2799gat));
  NOT NOT1_1650(.VSS(VSS),.VDD(VDD),.Y(n2796gat),.A(I4608));
  NOT NOT1_1651(.VSS(VSS),.VDD(VDD),.Y(n1118gat),.A(n1033gat));
  NOT NOT1_1652(.VSS(VSS),.VDD(VDD),.Y(n1032gat),.A(n1118gat));
  NOT NOT1_1653(.VSS(VSS),.VDD(VDD),.Y(n2054gat),.A(n2281gat));
  NOT NOT1_1654(.VSS(VSS),.VDD(VDD),.Y(I4615),.A(n2798gat));
  NOT NOT1_1655(.VSS(VSS),.VDD(VDD),.Y(n2795gat),.A(I4615));
  NOT NOT1_1656(.VSS(VSS),.VDD(VDD),.Y(I4620),.A(n1745gat));
  NOT NOT1_1657(.VSS(VSS),.VDD(VDD),.Y(n2806gat),.A(I4620));
  NOT NOT1_1658(.VSS(VSS),.VDD(VDD),.Y(I4623),.A(n2806gat));
  NOT NOT1_1659(.VSS(VSS),.VDD(VDD),.Y(n2802gat),.A(I4623));
  NOT NOT1_1660(.VSS(VSS),.VDD(VDD),.Y(I4626),.A(n1871gat));
  NOT NOT1_1661(.VSS(VSS),.VDD(VDD),.Y(n1870gat),.A(I4626));
  NOT NOT1_1662(.VSS(VSS),.VDD(VDD),.Y(n1086gat),.A(n1870gat));
  NOT NOT1_1663(.VSS(VSS),.VDD(VDD),.Y(I4630),.A(n1086gat));
  NOT NOT1_1664(.VSS(VSS),.VDD(VDD),.Y(n2805gat),.A(I4630));
  NOT NOT1_1665(.VSS(VSS),.VDD(VDD),.Y(I4633),.A(n2805gat));
  NOT NOT1_1666(.VSS(VSS),.VDD(VDD),.Y(n2801gat),.A(I4633));
  NOT NOT1_1667(.VSS(VSS),.VDD(VDD),.Y(n67gat),.A(n85gat));
  NOT NOT1_1668(.VSS(VSS),.VDD(VDD),.Y(n71gat),.A(n180gat));
  NOT NOT1_1669(.VSS(VSS),.VDD(VDD),.Y(n1840gat),.A(n1892gat));
  NOT NOT1_1670(.VSS(VSS),.VDD(VDD),.Y(I4642),.A(n2812gat));
  NOT NOT1_1671(.VSS(VSS),.VDD(VDD),.Y(n2809gat),.A(I4642));
  NOT NOT1_1672(.VSS(VSS),.VDD(VDD),.Y(n76gat),.A(n82gat));
  NOT NOT1_1673(.VSS(VSS),.VDD(VDD),.Y(n14gat),.A(n186gat));
  NOT NOT1_1674(.VSS(VSS),.VDD(VDD),.Y(n1842gat),.A(n1711gat));
  NOT NOT1_1675(.VSS(VSS),.VDD(VDD),.Y(I4651),.A(n2822gat));
  NOT NOT1_1676(.VSS(VSS),.VDD(VDD),.Y(n2819gat),.A(I4651));
  NOT NOT1_1677(.VSS(VSS),.VDD(VDD),.Y(I4654),.A(n2819gat));
  NOT NOT1_1678(.VSS(VSS),.VDD(VDD),.Y(n3104gat),.A(I4654));
  NOT NOT1_1679(.VSS(VSS),.VDD(VDD),.Y(I4657),.A(n2809gat));
  NOT NOT1_1680(.VSS(VSS),.VDD(VDD),.Y(n3105gat),.A(I4657));
  NOT NOT1_1681(.VSS(VSS),.VDD(VDD),.Y(I4660),.A(n2801gat));
  NOT NOT1_1682(.VSS(VSS),.VDD(VDD),.Y(n3106gat),.A(I4660));
  NOT NOT1_1683(.VSS(VSS),.VDD(VDD),.Y(I4663),.A(n2802gat));
  NOT NOT1_1684(.VSS(VSS),.VDD(VDD),.Y(n3107gat),.A(I4663));
  NOT NOT1_1685(.VSS(VSS),.VDD(VDD),.Y(I4666),.A(n2795gat));
  NOT NOT1_1686(.VSS(VSS),.VDD(VDD),.Y(n3108gat),.A(I4666));
  NOT NOT1_1687(.VSS(VSS),.VDD(VDD),.Y(I4669),.A(n2796gat));
  NOT NOT1_1688(.VSS(VSS),.VDD(VDD),.Y(n3109gat),.A(I4669));
  NOT NOT1_1689(.VSS(VSS),.VDD(VDD),.Y(I4672),.A(n2705gat));
  NOT NOT1_1690(.VSS(VSS),.VDD(VDD),.Y(n3110gat),.A(I4672));
  NOT NOT1_1691(.VSS(VSS),.VDD(VDD),.Y(I4675),.A(n2706gat));
  NOT NOT1_1692(.VSS(VSS),.VDD(VDD),.Y(n3111gat),.A(I4675));
  NOT NOT1_1693(.VSS(VSS),.VDD(VDD),.Y(I4678),.A(n2697gat));
  NOT NOT1_1694(.VSS(VSS),.VDD(VDD),.Y(n3112gat),.A(I4678));
  NOT NOT1_1695(.VSS(VSS),.VDD(VDD),.Y(I4681),.A(n2698gat));
  NOT NOT1_1696(.VSS(VSS),.VDD(VDD),.Y(n3113gat),.A(I4681));
  NOT NOT1_1697(.VSS(VSS),.VDD(VDD),.Y(I4684),.A(n2689gat));
  NOT NOT1_1698(.VSS(VSS),.VDD(VDD),.Y(n3114gat),.A(I4684));
  NOT NOT1_1699(.VSS(VSS),.VDD(VDD),.Y(I4687),.A(n2690gat));
  NOT NOT1_1700(.VSS(VSS),.VDD(VDD),.Y(n3115gat),.A(I4687));
  NOT NOT1_1701(.VSS(VSS),.VDD(VDD),.Y(I4690),.A(n2685gat));
  NOT NOT1_1702(.VSS(VSS),.VDD(VDD),.Y(n3116gat),.A(I4690));
  NOT NOT1_1703(.VSS(VSS),.VDD(VDD),.Y(I4693),.A(n2737gat));
  NOT NOT1_1704(.VSS(VSS),.VDD(VDD),.Y(n3117gat),.A(I4693));
  NOT NOT1_1705(.VSS(VSS),.VDD(VDD),.Y(I4696),.A(n2738gat));
  NOT NOT1_1706(.VSS(VSS),.VDD(VDD),.Y(n3118gat),.A(I4696));
  NOT NOT1_1707(.VSS(VSS),.VDD(VDD),.Y(I4699),.A(n2745gat));
  NOT NOT1_1708(.VSS(VSS),.VDD(VDD),.Y(n3119gat),.A(I4699));
  NOT NOT1_1709(.VSS(VSS),.VDD(VDD),.Y(I4702),.A(n2746gat));
  NOT NOT1_1710(.VSS(VSS),.VDD(VDD),.Y(n3120gat),.A(I4702));
  NOT NOT1_1711(.VSS(VSS),.VDD(VDD),.Y(I4705),.A(n2753gat));
  NOT NOT1_1712(.VSS(VSS),.VDD(VDD),.Y(n3121gat),.A(I4705));
  NOT NOT1_1713(.VSS(VSS),.VDD(VDD),.Y(I4708),.A(n2754gat));
  NOT NOT1_1714(.VSS(VSS),.VDD(VDD),.Y(n3122gat),.A(I4708));
  NOT NOT1_1715(.VSS(VSS),.VDD(VDD),.Y(I4711),.A(n2759gat));
  NOT NOT1_1716(.VSS(VSS),.VDD(VDD),.Y(n3123gat),.A(I4711));
  NOT NOT1_1717(.VSS(VSS),.VDD(VDD),.Y(I4714),.A(n2760gat));
  NOT NOT1_1718(.VSS(VSS),.VDD(VDD),.Y(n3124gat),.A(I4714));
  NOT NOT1_1719(.VSS(VSS),.VDD(VDD),.Y(I4717),.A(n2763gat));
  NOT NOT1_1720(.VSS(VSS),.VDD(VDD),.Y(n3125gat),.A(I4717));
  NOT NOT1_1721(.VSS(VSS),.VDD(VDD),.Y(I4720),.A(n2686gat));
  NOT NOT1_1722(.VSS(VSS),.VDD(VDD),.Y(n3126gat),.A(I4720));
  NOT NOT1_1723(.VSS(VSS),.VDD(VDD),.Y(I4723),.A(n2677gat));
  NOT NOT1_1724(.VSS(VSS),.VDD(VDD),.Y(n3127gat),.A(I4723));
  NOT NOT1_1725(.VSS(VSS),.VDD(VDD),.Y(I4726),.A(n2678gat));
  NOT NOT1_1726(.VSS(VSS),.VDD(VDD),.Y(n3128gat),.A(I4726));
  NOT NOT1_1727(.VSS(VSS),.VDD(VDD),.Y(I4729),.A(n2803gat));
  NOT NOT1_1728(.VSS(VSS),.VDD(VDD),.Y(n3129gat),.A(I4729));
  NOT NOT1_1729(.VSS(VSS),.VDD(VDD),.Y(I4732),.A(n2825gat));
  NOT NOT1_1730(.VSS(VSS),.VDD(VDD),.Y(n3130gat),.A(I4732));
  NOT NOT1_1731(.VSS(VSS),.VDD(VDD),.Y(I4735),.A(n2826gat));
  NOT NOT1_1732(.VSS(VSS),.VDD(VDD),.Y(n3131gat),.A(I4735));
  NOT NOT1_1733(.VSS(VSS),.VDD(VDD),.Y(I4738),.A(n2820gat));
  NOT NOT1_1734(.VSS(VSS),.VDD(VDD),.Y(n3132gat),.A(I4738));
  NOT NOT1_1735(.VSS(VSS),.VDD(VDD),.Y(I4741),.A(n2821gat));
  NOT NOT1_1736(.VSS(VSS),.VDD(VDD),.Y(n3133gat),.A(I4741));
  NOT NOT1_1737(.VSS(VSS),.VDD(VDD),.Y(I4744),.A(n2815gat));
  NOT NOT1_1738(.VSS(VSS),.VDD(VDD),.Y(n3134gat),.A(I4744));
  NOT NOT1_1739(.VSS(VSS),.VDD(VDD),.Y(I4747),.A(n2816gat));
  NOT NOT1_1740(.VSS(VSS),.VDD(VDD),.Y(n3135gat),.A(I4747));
  NOT NOT1_1741(.VSS(VSS),.VDD(VDD),.Y(I4750),.A(n2810gat));
  NOT NOT1_1742(.VSS(VSS),.VDD(VDD),.Y(n3136gat),.A(I4750));
  NOT NOT1_1743(.VSS(VSS),.VDD(VDD),.Y(I4753),.A(n2811gat));
  NOT NOT1_1744(.VSS(VSS),.VDD(VDD),.Y(n3137gat),.A(I4753));
  NOT NOT1_1745(.VSS(VSS),.VDD(VDD),.Y(I4756),.A(n2804gat));
  NOT NOT1_1746(.VSS(VSS),.VDD(VDD),.Y(n3138gat),.A(I4756));
  NOT NOT1_1747(.VSS(VSS),.VDD(VDD),.Y(I4759),.A(n2739gat));
  NOT NOT1_1748(.VSS(VSS),.VDD(VDD),.Y(n3139gat),.A(I4759));
  NOT NOT1_1749(.VSS(VSS),.VDD(VDD),.Y(I4762),.A(n2747gat));
  NOT NOT1_1750(.VSS(VSS),.VDD(VDD),.Y(n3140gat),.A(I4762));
  NOT NOT1_1751(.VSS(VSS),.VDD(VDD),.Y(I4765),.A(n2748gat));
  NOT NOT1_1752(.VSS(VSS),.VDD(VDD),.Y(n3141gat),.A(I4765));
  NOT NOT1_1753(.VSS(VSS),.VDD(VDD),.Y(I4768),.A(n2755gat));
  NOT NOT1_1754(.VSS(VSS),.VDD(VDD),.Y(n3142gat),.A(I4768));
  NOT NOT1_1755(.VSS(VSS),.VDD(VDD),.Y(I4771),.A(n2797gat));
  NOT NOT1_1756(.VSS(VSS),.VDD(VDD),.Y(n3143gat),.A(I4771));
  NOT NOT1_1757(.VSS(VSS),.VDD(VDD),.Y(I4774),.A(n2740gat));
  NOT NOT1_1758(.VSS(VSS),.VDD(VDD),.Y(n3144gat),.A(I4774));
  NOT NOT1_1759(.VSS(VSS),.VDD(VDD),.Y(I4777),.A(n2699gat));
  NOT NOT1_1760(.VSS(VSS),.VDD(VDD),.Y(n3145gat),.A(I4777));
  NOT NOT1_1761(.VSS(VSS),.VDD(VDD),.Y(I4780),.A(n2691gat));
  NOT NOT1_1762(.VSS(VSS),.VDD(VDD),.Y(n3146gat),.A(I4780));
  NOT NOT1_1763(.VSS(VSS),.VDD(VDD),.Y(I4783),.A(n2827gat));
  NOT NOT1_1764(.VSS(VSS),.VDD(VDD),.Y(n3147gat),.A(I4783));
  NOT NOT1_1765(.VSS(VSS),.VDD(VDD),.Y(I4786),.A(n2679gat));
  NOT NOT1_1766(.VSS(VSS),.VDD(VDD),.Y(n3148gat),.A(I4786));
  NOT NOT1_1767(.VSS(VSS),.VDD(VDD),.Y(I4789),.A(n2692gat));
  NOT NOT1_1768(.VSS(VSS),.VDD(VDD),.Y(n3149gat),.A(I4789));
  NOT NOT1_1769(.VSS(VSS),.VDD(VDD),.Y(I4792),.A(n2680gat));
  NOT NOT1_1770(.VSS(VSS),.VDD(VDD),.Y(n3150gat),.A(I4792));
  NOT NOT1_1771(.VSS(VSS),.VDD(VDD),.Y(I4795),.A(n2700gat));
  NOT NOT1_1772(.VSS(VSS),.VDD(VDD),.Y(n3151gat),.A(I4795));
  NOT NOT1_1773(.VSS(VSS),.VDD(VDD),.Y(I4798),.A(n2707gat));
  NOT NOT1_1774(.VSS(VSS),.VDD(VDD),.Y(n3152gat),.A(I4798));
//
  OR2 OR2_0(.VSS(VSS),.VDD(VDD),.Y(n2897gat),.A(n648gat),.B(n442gat));
  OR4 OR4_0(.VSS(VSS),.VDD(VDD),.Y(n1213gat),.A(n1214gat),.B(n1215gat),.C(n1216gat),.D(n1217gat));
  OR2 OR2_1(.VSS(VSS),.VDD(VDD),.Y(n2906gat),.A(n745gat),.B(n638gat));
  OR2 OR2_2(.VSS(VSS),.VDD(VDD),.Y(n2889gat),.A(n423gat),.B(n362gat));
  OR4 OR4_1(.VSS(VSS),.VDD(VDD),.Y(n748gat),.A(n749gat),.B(n750gat),.C(n751gat),.D(n752gat));
  OR4 OR4_2(.VSS(VSS),.VDD(VDD),.Y(n258gat),.A(n259gat),.B(n260gat),.C(n261gat),.D(n262gat));
  OR4 OR4_3(.VSS(VSS),.VDD(VDD),.Y(n1013gat),.A(n1014gat),.B(n1015gat),.C(n1016gat),.D(n1017gat));
  OR4 OR4_4(.VSS(VSS),.VDD(VDD),.Y(n475gat),.A(n476gat),.B(n477gat),.C(n478gat),.D(n479gat));
  OR4 OR4_5(.VSS(VSS),.VDD(VDD),.Y(n43gat),.A(n44gat),.B(n45gat),.C(n46gat),.D(n47gat));
  OR2 OR2_3(.VSS(VSS),.VDD(VDD),.Y(n2786gat),.A(n3091gat),.B(n3092gat));
  OR4 OR4_6(.VSS(VSS),.VDD(VDD),.Y(n167gat),.A(n168gat),.B(n169gat),.C(n170gat),.D(n171gat));
  OR4 OR4_7(.VSS(VSS),.VDD(VDD),.Y(n906gat),.A(n907gat),.B(n908gat),.C(n909gat),.D(n910gat));
  OR4 OR4_8(.VSS(VSS),.VDD(VDD),.Y(n343gat),.A(n344gat),.B(n345gat),.C(n346gat),.D(n347gat));
  OR4 OR4_9(.VSS(VSS),.VDD(VDD),.Y(n55gat),.A(n56gat),.B(n57gat),.C(n58gat),.D(n59gat));
  OR2 OR2_4(.VSS(VSS),.VDD(VDD),.Y(n2914gat),.A(n768gat),.B(n655gat));
  OR2 OR2_5(.VSS(VSS),.VDD(VDD),.Y(n2928gat),.A(n963gat),.B(n868gat));
  OR2 OR2_6(.VSS(VSS),.VDD(VDD),.Y(n2927gat),.A(n962gat),.B(n959gat));
  OR4 OR4_10(.VSS(VSS),.VDD(VDD),.Y(n944gat),.A(n945gat),.B(n946gat),.C(n947gat),.D(n948gat));
  OR2 OR2_7(.VSS(VSS),.VDD(VDD),.Y(n2896gat),.A(n647gat),.B(n441gat));
  OR2 OR2_8(.VSS(VSS),.VDD(VDD),.Y(n2922gat),.A(n967gat),.B(n792gat));
  OR4 OR4_11(.VSS(VSS),.VDD(VDD),.Y(n1228gat),.A(n1229gat),.B(n1230gat),.C(n1231gat),.D(n1232gat));
  OR2 OR2_9(.VSS(VSS),.VDD(VDD),.Y(n2894gat),.A(n443gat),.B(n439gat));
  OR2 OR2_10(.VSS(VSS),.VDD(VDD),.Y(n2921gat),.A(n966gat),.B(n790gat));
  OR2 OR2_11(.VSS(VSS),.VDD(VDD),.Y(n2895gat),.A(n444gat),.B(n440gat));
  OR4 OR4_12(.VSS(VSS),.VDD(VDD),.Y(n1050gat),.A(n1051gat),.B(n1052gat),.C(n1053gat),.D(n1054gat));
  OR4 OR4_13(.VSS(VSS),.VDD(VDD),.Y(n933gat),.A(n934gat),.B(n935gat),.C(n936gat),.D(n937gat));
  OR4 OR4_14(.VSS(VSS),.VDD(VDD),.Y(n709gat),.A(n710gat),.B(n711gat),.C(n712gat),.D(n713gat));
  OR4 OR4_15(.VSS(VSS),.VDD(VDD),.Y(n728gat),.A(n729gat),.B(n730gat),.C(n731gat),.D(n732gat));
  OR4 OR4_16(.VSS(VSS),.VDD(VDD),.Y(n493gat),.A(n494gat),.B(n495gat),.C(n496gat),.D(n497gat));
  OR4 OR4_17(.VSS(VSS),.VDD(VDD),.Y(n504gat),.A(n505gat),.B(n506gat),.C(n507gat),.D(n508gat));
  OR3 OR3_0(.VSS(VSS),.VDD(VDD),.Y(I1277),.A(n2860gat),.B(n2855gat),.C(n2863gat));
  OR3 OR3_1(.VSS(VSS),.VDD(VDD),.Y(I1278),.A(n740gat),.B(n3030gat),.C(I1277));
  OR2 OR2_12(.VSS(VSS),.VDD(VDD),.Y(n2913gat),.A(n767gat),.B(n653gat));
  OR2 OR2_13(.VSS(VSS),.VDD(VDD),.Y(n2920gat),.A(n867gat),.B(n771gat));
  OR2 OR2_14(.VSS(VSS),.VDD(VDD),.Y(n2905gat),.A(n964gat),.B(n961gat));
  OR4 OR4_18(.VSS(VSS),.VDD(VDD),.Y(n803gat),.A(n804gat),.B(n805gat),.C(n806gat),.D(n807gat));
  OR4 OR4_19(.VSS(VSS),.VDD(VDD),.Y(n586gat),.A(n587gat),.B(n588gat),.C(n589gat),.D(n590gat));
  OR2 OR2_15(.VSS(VSS),.VDD(VDD),.Y(n2898gat),.A(n447gat),.B(n445gat));
  OR4 OR4_20(.VSS(VSS),.VDD(VDD),.Y(n686gat),.A(n687gat),.B(n688gat),.C(n689gat),.D(n690gat));
  OR4 OR4_21(.VSS(VSS),.VDD(VDD),.Y(n567gat),.A(n568gat),.B(n569gat),.C(n570gat),.D(n571gat));
  OR3 OR3_2(.VSS(VSS),.VDD(VDD),.Y(I1515),.A(n2474gat),.B(n2524gat),.C(n2831gat));
  OR3 OR3_3(.VSS(VSS),.VDD(VDD),.Y(I1516),.A(n2466gat),.B(n2462gat),.C(I1515));
  OR3 OR3_4(.VSS(VSS),.VDD(VDD),.Y(I1584),.A(n2353gat),.B(n2284gat),.C(n2354gat));
  OR3 OR3_5(.VSS(VSS),.VDD(VDD),.Y(I1585),.A(n2356gat),.B(n2214gat),.C(I1584));
  OR2 OR2_16(.VSS(VSS),.VDD(VDD),.Y(n2989gat),.A(n1693gat),.B(n1692gat));
  OR3 OR3_6(.VSS(VSS),.VDD(VDD),.Y(I1723),.A(n2354gat),.B(n2353gat),.C(n2214gat));
  OR3 OR3_7(.VSS(VSS),.VDD(VDD),.Y(I1724),.A(n2355gat),.B(n2443gat),.C(I1723));
  OR3 OR3_8(.VSS(VSS),.VDD(VDD),.Y(I1733),.A(n2286gat),.B(n2428gat),.C(n2289gat));
  OR3 OR3_9(.VSS(VSS),.VDD(VDD),.Y(I1734),.A(n1604gat),.B(n2214gat),.C(I1733));
  OR2 OR2_17(.VSS(VSS),.VDD(VDD),.Y(n2918gat),.A(n769gat),.B(n759gat));
  OR2 OR2_18(.VSS(VSS),.VDD(VDD),.Y(n2952gat),.A(n1076gat),.B(n1075gat));
  OR2 OR2_19(.VSS(VSS),.VDD(VDD),.Y(n2919gat),.A(n766gat),.B(n760gat));
  OR4 OR4_22(.VSS(VSS),.VDD(VDD),.Y(n1184gat),.A(n1185gat),.B(n1186gat),.C(n1187gat),.D(n1188gat));
  OR2 OR2_20(.VSS(VSS),.VDD(VDD),.Y(n2910gat),.A(n645gat),.B(n644gat));
  OR2 OR2_21(.VSS(VSS),.VDD(VDD),.Y(n2907gat),.A(n646gat),.B(n641gat));
  OR2 OR2_22(.VSS(VSS),.VDD(VDD),.Y(n2970gat),.A(n1383gat),.B(n1327gat));
  OR2 OR2_23(.VSS(VSS),.VDD(VDD),.Y(n2911gat),.A(n761gat),.B(n651gat));
  OR2 OR2_24(.VSS(VSS),.VDD(VDD),.Y(n2912gat),.A(n762gat),.B(n652gat));
  OR2 OR2_25(.VSS(VSS),.VDD(VDD),.Y(n2909gat),.A(n765gat),.B(n643gat));
  OR4 OR4_23(.VSS(VSS),.VDD(VDD),.Y(n1201gat),.A(n1202gat),.B(n1203gat),.C(n1204gat),.D(n1205gat));
  OR4 OR4_24(.VSS(VSS),.VDD(VDD),.Y(n1269gat),.A(n1270gat),.B(n1271gat),.C(n1272gat),.D(n1273gat));
  OR2 OR2_26(.VSS(VSS),.VDD(VDD),.Y(n2908gat),.A(n763gat),.B(n642gat));
  OR2 OR2_27(.VSS(VSS),.VDD(VDD),.Y(n2971gat),.A(n1287gat),.B(n1285gat));
  OR3 OR3_10(.VSS(VSS),.VDD(VDD),.Y(n2904gat),.A(n793gat),.B(n664gat),.C(n556gat));
  OR3 OR3_11(.VSS(VSS),.VDD(VDD),.Y(n2891gat),.A(n795gat),.B(n656gat),.C(n368gat));
  OR3 OR3_12(.VSS(VSS),.VDD(VDD),.Y(n2903gat),.A(n794gat),.B(n773gat),.C(n662gat));
  OR3 OR3_13(.VSS(VSS),.VDD(VDD),.Y(n2915gat),.A(n965gat),.B(n960gat),.C(n661gat));
  OR4 OR4_25(.VSS(VSS),.VDD(VDD),.Y(n779gat),.A(n780gat),.B(n781gat),.C(n782gat),.D(n783gat));
  OR3 OR3_14(.VSS(VSS),.VDD(VDD),.Y(n2901gat),.A(n558gat),.B(n555gat),.C(n450gat));
  OR3 OR3_15(.VSS(VSS),.VDD(VDD),.Y(n2890gat),.A(n654gat),.B(n557gat),.C(n371gat));
  OR2 OR2_28(.VSS(VSS),.VDD(VDD),.Y(n2876gat),.A(n874gat),.B(n132gat));
  OR3 OR3_16(.VSS(VSS),.VDD(VDD),.Y(n2888gat),.A(n663gat),.B(n649gat),.C(n449gat));
  OR3 OR3_17(.VSS(VSS),.VDD(VDD),.Y(n2887gat),.A(n791gat),.B(n650gat),.C(n370gat));
  OR3 OR3_18(.VSS(VSS),.VDD(VDD),.Y(n2886gat),.A(n774gat),.B(n764gat),.C(n369gat));
  OR4 OR4_26(.VSS(VSS),.VDD(VDD),.Y(n221gat),.A(n222gat),.B(n223gat),.C(n224gat),.D(n225gat));
  OR4 OR4_27(.VSS(VSS),.VDD(VDD),.Y(n120gat),.A(n121gat),.B(n122gat),.C(n123gat),.D(n124gat));
  OR2 OR2_29(.VSS(VSS),.VDD(VDD),.Y(n3010gat),.A(n2460gat),.B(n2423gat));
  OR2 OR2_30(.VSS(VSS),.VDD(VDD),.Y(n3016gat),.A(n2596gat),.B(n2595gat));
  OR4 OR4_28(.VSS(VSS),.VDD(VDD),.Y(n2568gat),.A(n2569gat),.B(n2570gat),.C(n2571gat),.D(n2572gat));
  OR4 OR4_29(.VSS(VSS),.VDD(VDD),.Y(n2409gat),.A(n2410gat),.B(n2411gat),.C(n2412gat),.D(n2413gat));
  OR2 OR2_31(.VSS(VSS),.VDD(VDD),.Y(n2579gat),.A(n2580gat),.B(n2581gat));
  OR2 OR2_32(.VSS(VSS),.VDD(VDD),.Y(n3014gat),.A(n2567gat),.B(n2499gat));
  OR2 OR2_33(.VSS(VSS),.VDD(VDD),.Y(n2880gat),.A(n299gat),.B(n207gat));
  OR2 OR2_34(.VSS(VSS),.VDD(VDD),.Y(n2646gat),.A(n2647gat),.B(n2648gat));
  OR4 OR4_30(.VSS(VSS),.VDD(VDD),.Y(n2601gat),.A(n2602gat),.B(n2603gat),.C(n2604gat),.D(n2605gat));
  OR4 OR4_31(.VSS(VSS),.VDD(VDD),.Y(n2545gat),.A(n2546gat),.B(n2547gat),.C(n2548gat),.D(n2549gat));
  OR2 OR2_35(.VSS(VSS),.VDD(VDD),.Y(n2613gat),.A(n2614gat),.B(n2615gat));
  OR2 OR2_36(.VSS(VSS),.VDD(VDD),.Y(n3013gat),.A(n2461gat),.B(n2421gat));
  OR4 OR4_32(.VSS(VSS),.VDD(VDD),.Y(n2930gat),.A(n1153gat),.B(n1151gat),.C(n982gat),.D(n877gat));
  OR4 OR4_33(.VSS(VSS),.VDD(VDD),.Y(n2957gat),.A(n1159gat),.B(n1158gat),.C(n1156gat),.D(n1155gat));
  OR2 OR2_37(.VSS(VSS),.VDD(VDD),.Y(n2975gat),.A(n1443gat),.B(n1325gat));
  OR2 OR2_38(.VSS(VSS),.VDD(VDD),.Y(n2974gat),.A(n1321gat),.B(n1320gat));
  OR2 OR2_39(.VSS(VSS),.VDD(VDD),.Y(n2966gat),.A(n1368gat),.B(n1258gat));
  OR2 OR2_40(.VSS(VSS),.VDD(VDD),.Y(n2979gat),.A(n1373gat),.B(n1372gat));
  OR4 OR4_34(.VSS(VSS),.VDD(VDD),.Y(n2978gat),.A(n1441gat),.B(n1440gat),.C(n1371gat),.D(n1367gat));
  OR2 OR2_41(.VSS(VSS),.VDD(VDD),.Y(n2982gat),.A(n1504gat),.B(n1502gat));
  OR2 OR2_42(.VSS(VSS),.VDD(VDD),.Y(n2954gat),.A(n1250gat),.B(n1103gat));
  OR2 OR2_43(.VSS(VSS),.VDD(VDD),.Y(n2964gat),.A(n1304gat),.B(n1249gat));
  OR2 OR2_44(.VSS(VSS),.VDD(VDD),.Y(n2958gat),.A(n1246gat),.B(n1161gat));
  OR2 OR2_45(.VSS(VSS),.VDD(VDD),.Y(n2963gat),.A(n1291gat),.B(n1245gat));
  OR4 OR4_35(.VSS(VSS),.VDD(VDD),.Y(n2973gat),.A(n1352gat),.B(n1351gat),.C(n1303gat),.D(n1302gat));
  OR2 OR2_46(.VSS(VSS),.VDD(VDD),.Y(n2953gat),.A(n1163gat),.B(n1102gat));
  OR2 OR2_47(.VSS(VSS),.VDD(VDD),.Y(n2949gat),.A(n1101gat),.B(n996gat));
  OR2 OR2_48(.VSS(VSS),.VDD(VDD),.Y(n2934gat),.A(n1104gat),.B(n887gat));
  OR2 OR2_49(.VSS(VSS),.VDD(VDD),.Y(n2959gat),.A(n1305gat),.B(n1162gat));
  OR4 OR4_36(.VSS(VSS),.VDD(VDD),.Y(n2977gat),.A(n1360gat),.B(n1359gat),.C(n1358gat),.D(n1357gat));
  OR3 OR3_19(.VSS(VSS),.VDD(VDD),.Y(I2720),.A(n1788gat),.B(n1786gat),.C(n1839gat));
  OR3 OR3_20(.VSS(VSS),.VDD(VDD),.Y(I2721),.A(n1884gat),.B(n1783gat),.C(I2720));
  OR3 OR3_21(.VSS(VSS),.VDD(VDD),.Y(I2735),.A(n1788gat),.B(n1884gat),.C(n1633gat));
  OR3 OR3_22(.VSS(VSS),.VDD(VDD),.Y(I2736),.A(n1785gat),.B(n1784gat),.C(I2735));
  OR3 OR3_23(.VSS(VSS),.VDD(VDD),.Y(I2812),.A(n1703gat),.B(n1704gat),.C(n1778gat));
  OR4 OR4_37(.VSS(VSS),.VDD(VDD),.Y(I2813),.A(n1609gat),.B(n1702gat),.C(n1700gat),.D(I2812));
  OR3 OR3_24(.VSS(VSS),.VDD(VDD),.Y(I2831),.A(n1839gat),.B(n1786gat),.C(n1788gat));
  OR3 OR3_25(.VSS(VSS),.VDD(VDD),.Y(I2832),.A(n1884gat),.B(n1784gat),.C(I2831));
  OR3 OR3_26(.VSS(VSS),.VDD(VDD),.Y(I2889),.A(n1784gat),.B(n1633gat),.C(n1884gat));
  OR3 OR3_27(.VSS(VSS),.VDD(VDD),.Y(I2890),.A(n1788gat),.B(n1786gat),.C(I2889));
  OR3 OR3_28(.VSS(VSS),.VDD(VDD),.Y(I2925),.A(n1784gat),.B(n1785gat),.C(n1633gat));
  OR3 OR3_29(.VSS(VSS),.VDD(VDD),.Y(I2926),.A(n1884gat),.B(n1787gat),.C(I2925));
  OR3 OR3_30(.VSS(VSS),.VDD(VDD),.Y(I2934),.A(n1784gat),.B(n1839gat),.C(n1788gat));
  OR3 OR3_31(.VSS(VSS),.VDD(VDD),.Y(I2935),.A(n1785gat),.B(n1884gat),.C(I2934));
  OR2 OR2_50(.VSS(VSS),.VDD(VDD),.Y(n2988gat),.A(n1733gat),.B(n1581gat));
  OR2 OR2_51(.VSS(VSS),.VDD(VDD),.Y(n2983gat),.A(n2079gat),.B(n2073gat));
  OR2 OR2_52(.VSS(VSS),.VDD(VDD),.Y(n2987gat),.A(n1574gat),.B(n1573gat));
  OR3 OR3_32(.VSS(VSS),.VDD(VDD),.Y(n2992gat),.A(n1723gat),.B(n1647gat),.C(n1646gat));
  OR3 OR3_33(.VSS(VSS),.VDD(VDD),.Y(n2986gat),.A(n1650gat),.B(n1649gat),.C(n1563gat));
  OR3 OR3_34(.VSS(VSS),.VDD(VDD),.Y(n2991gat),.A(n1654gat),.B(n1653gat),.C(n1644gat));
  OR3 OR3_35(.VSS(VSS),.VDD(VDD),.Y(I3148),.A(n1839gat),.B(n1884gat),.C(n1784gat));
  OR3 OR3_36(.VSS(VSS),.VDD(VDD),.Y(I3149),.A(n1786gat),.B(n1787gat),.C(I3148));
  OR3 OR3_37(.VSS(VSS),.VDD(VDD),.Y(I3178),.A(n1838gat),.B(n1785gat),.C(n1788gat));
  OR3 OR3_38(.VSS(VSS),.VDD(VDD),.Y(I3179),.A(n1839gat),.B(n1784gat),.C(I3178));
  OR3 OR3_39(.VSS(VSS),.VDD(VDD),.Y(n2981gat),.A(n1413gat),.B(n1408gat),.C(n1407gat));
  OR2 OR2_53(.VSS(VSS),.VDD(VDD),.Y(n3000gat),.A(n2000gat),.B(n1999gat));
  OR3 OR3_40(.VSS(VSS),.VDD(VDD),.Y(n3004gat),.A(n2258gat),.B(n2257gat),.C(n2255gat));
  OR2 OR2_54(.VSS(VSS),.VDD(VDD),.Y(n3003gat),.A(n2256gat),.B(n2251gat));
  OR2 OR2_55(.VSS(VSS),.VDD(VDD),.Y(n3001gat),.A(n2132gat),.B(n2130gat));
  OR2 OR2_56(.VSS(VSS),.VDD(VDD),.Y(n3006gat),.A(n2253gat),.B(n2252gat));
  OR2 OR2_57(.VSS(VSS),.VDD(VDD),.Y(n3007gat),.A(n2250gat),.B(n2249gat));
  OR2 OR2_58(.VSS(VSS),.VDD(VDD),.Y(n2990gat),.A(n1710gat),.B(n1630gat));
  OR2 OR2_59(.VSS(VSS),.VDD(VDD),.Y(n2994gat),.A(n1954gat),.B(n1888gat));
  OR3 OR3_41(.VSS(VSS),.VDD(VDD),.Y(n2993gat),.A(n1894gat),.B(n1847gat),.C(n1846gat));
  OR2 OR2_60(.VSS(VSS),.VDD(VDD),.Y(n2998gat),.A(n2055gat),.B(n1967gat));
  OR3 OR3_42(.VSS(VSS),.VDD(VDD),.Y(n2996gat),.A(n1960gat),.B(n1959gat),.C(n1957gat));
  OR2 OR2_61(.VSS(VSS),.VDD(VDD),.Y(n3008gat),.A(n2332gat),.B(n2259gat));
  OR2 OR2_62(.VSS(VSS),.VDD(VDD),.Y(n3005gat),.A(n2211gat),.B(n2210gat));
  OR3 OR3_43(.VSS(VSS),.VDD(VDD),.Y(n2997gat),.A(n2053gat),.B(n2052gat),.C(n1964gat));
  OR2 OR2_63(.VSS(VSS),.VDD(VDD),.Y(n3009gat),.A(n2350gat),.B(n2282gat));
  OR3 OR3_44(.VSS(VSS),.VDD(VDD),.Y(n3002gat),.A(n2213gat),.B(n2150gat),.C(n2149gat));
  OR2 OR2_64(.VSS(VSS),.VDD(VDD),.Y(n2995gat),.A(n1962gat),.B(n1955gat));
  OR2 OR2_65(.VSS(VSS),.VDD(VDD),.Y(n2999gat),.A(n1972gat),.B(n1971gat));
  OR2 OR2_66(.VSS(VSS),.VDD(VDD),.Y(n3011gat),.A(n2333gat),.B(n2331gat));
  OR2 OR2_67(.VSS(VSS),.VDD(VDD),.Y(n3015gat),.A(n2566gat),.B(n2565gat));
  OR3 OR3_45(.VSS(VSS),.VDD(VDD),.Y(n2874gat),.A(n141gat),.B(n38gat),.C(n37gat));
  OR2 OR2_68(.VSS(VSS),.VDD(VDD),.Y(n2917gat),.A(n1074gat),.B(n872gat));
  OR2 OR2_69(.VSS(VSS),.VDD(VDD),.Y(n2878gat),.A(n234gat),.B(n137gat));
  OR2 OR2_70(.VSS(VSS),.VDD(VDD),.Y(n2892gat),.A(n378gat),.B(n377gat));
  OR3 OR3_46(.VSS(VSS),.VDD(VDD),.Y(n2885gat),.A(n250gat),.B(n249gat),.C(n248gat));
  OR3 OR3_47(.VSS(VSS),.VDD(VDD),.Y(n2900gat),.A(n869gat),.B(n453gat),.C(n448gat));
  OR2 OR2_71(.VSS(VSS),.VDD(VDD),.Y(n2883gat),.A(n251gat),.B(n244gat));
  OR3 OR3_48(.VSS(VSS),.VDD(VDD),.Y(n2929gat),.A(n974gat),.B(n973gat),.C(n870gat));
  OR2 OR2_72(.VSS(VSS),.VDD(VDD),.Y(n2884gat),.A(n246gat),.B(n245gat));
  OR2 OR2_73(.VSS(VSS),.VDD(VDD),.Y(n2902gat),.A(n460gat),.B(n459gat));
  OR3 OR3_49(.VSS(VSS),.VDD(VDD),.Y(n2925gat),.A(n975gat),.B(n972gat),.C(n969gat));
  OR2 OR2_74(.VSS(VSS),.VDD(VDD),.Y(n2879gat),.A(n145gat),.B(n143gat));
  OR3 OR3_50(.VSS(VSS),.VDD(VDD),.Y(n2916gat),.A(n971gat),.B(n970gat),.C(n968gat));
  OR3 OR3_51(.VSS(VSS),.VDD(VDD),.Y(n2875gat),.A(n142gat),.B(n40gat),.C(n39gat));
  OR3 OR3_52(.VSS(VSS),.VDD(VDD),.Y(n2899gat),.A(n772gat),.B(n451gat),.C(n446gat));
  OR2 OR2_75(.VSS(VSS),.VDD(VDD),.Y(n2877gat),.A(n139gat),.B(n136gat));
  OR2 OR2_76(.VSS(VSS),.VDD(VDD),.Y(n2893gat),.A(n391gat),.B(n390gat));
  OR2 OR2_77(.VSS(VSS),.VDD(VDD),.Y(n2926gat),.A(n1083gat),.B(n1077gat));
  OR2 OR2_78(.VSS(VSS),.VDD(VDD),.Y(n2882gat),.A(n242gat),.B(n240gat));
  OR2 OR2_79(.VSS(VSS),.VDD(VDD),.Y(n2924gat),.A(n871gat),.B(n797gat));
  OR3 OR3_53(.VSS(VSS),.VDD(VDD),.Y(n2881gat),.A(n324gat),.B(n238gat),.C(n237gat));
  OR2 OR2_80(.VSS(VSS),.VDD(VDD),.Y(n2923gat),.A(n1082gat),.B(n796gat));
  OR2 OR2_81(.VSS(VSS),.VDD(VDD),.Y(n2710gat),.A(n69gat),.B(n1885gat));
  OR2 OR2_82(.VSS(VSS),.VDD(VDD),.Y(n2704gat),.A(n11gat),.B(n1889gat));
  OR2 OR2_83(.VSS(VSS),.VDD(VDD),.Y(n2684gat),.A(n1599gat),.B(n2051gat));
  OR2 OR2_84(.VSS(VSS),.VDD(VDD),.Y(n2830gat),.A(n2444gat),.B(n1754gat));
  OR3 OR3_54(.VSS(VSS),.VDD(VDD),.Y(I3999),.A(n2167gat),.B(n2031gat),.C(n2174gat));
  OR4 OR4_38(.VSS(VSS),.VDD(VDD),.Y(I4000),.A(n2108gat),.B(n2093gat),.C(n2035gat),.D(I3999));
  OR2 OR2_85(.VSS(VSS),.VDD(VDD),.Y(n2695gat),.A(n1586gat),.B(n1791gat));
  OR2 OR2_86(.VSS(VSS),.VDD(VDD),.Y(n2703gat),.A(n1755gat),.B(n1518gat));
  OR2 OR2_87(.VSS(VSS),.VDD(VDD),.Y(n2744gat),.A(n2159gat),.B(n2478gat));
  OR2 OR2_88(.VSS(VSS),.VDD(VDD),.Y(n2800gat),.A(n2158gat),.B(n2186gat));
  OR3 OR3_55(.VSS(VSS),.VDD(VDD),.Y(I4023),.A(n2443gat),.B(n2290gat),.C(n2214gat));
  OR3 OR3_56(.VSS(VSS),.VDD(VDD),.Y(I4024),.A(n2353gat),.B(n2284gat),.C(I4023));
  OR4 OR4_39(.VSS(VSS),.VDD(VDD),.Y(n2980gat),.A(n1470gat),.B(n1400gat),.C(n1399gat),.D(n1398gat));
  OR3 OR3_57(.VSS(VSS),.VDD(VDD),.Y(I4144),.A(n1633gat),.B(n1838gat),.C(n1786gat));
  OR3 OR3_58(.VSS(VSS),.VDD(VDD),.Y(I4145),.A(n1788gat),.B(n1784gat),.C(I4144));
  OR2 OR2_89(.VSS(VSS),.VDD(VDD),.Y(n2984gat),.A(n1467gat),.B(n1466gat));
  OR4 OR4_40(.VSS(VSS),.VDD(VDD),.Y(n2985gat),.A(n1686gat),.B(n1533gat),.C(n1532gat),.D(n1531gat));
  OR3 OR3_59(.VSS(VSS),.VDD(VDD),.Y(I4216),.A(n1427gat),.B(n1595gat),.C(n1677gat));
  OR3 OR3_60(.VSS(VSS),.VDD(VDD),.Y(I4217),.A(n1392gat),.B(n2989gat),.C(I4216));
  OR4 OR4_41(.VSS(VSS),.VDD(VDD),.Y(n2931gat),.A(n1100gat),.B(n994gat),.C(n989gat),.D(n880gat));
  OR2 OR2_90(.VSS(VSS),.VDD(VDD),.Y(n2943gat),.A(n1012gat),.B(n905gat));
  OR2 OR2_91(.VSS(VSS),.VDD(VDD),.Y(n2941gat),.A(n1003gat),.B(n902gat));
  OR4 OR4_42(.VSS(VSS),.VDD(VDD),.Y(n2946gat),.A(n1099gat),.B(n998gat),.C(n995gat),.D(n980gat));
  OR2 OR2_92(.VSS(VSS),.VDD(VDD),.Y(n2960gat),.A(n1175gat),.B(n1174gat));
  OR2 OR2_93(.VSS(VSS),.VDD(VDD),.Y(n2950gat),.A(n1001gat),.B(n999gat));
  OR2 OR2_94(.VSS(VSS),.VDD(VDD),.Y(n2969gat),.A(n1323gat),.B(n1264gat));
  OR4 OR4_43(.VSS(VSS),.VDD(VDD),.Y(n2933gat),.A(n981gat),.B(n890gat),.C(n889gat),.D(n886gat));
  OR2 OR2_95(.VSS(VSS),.VDD(VDD),.Y(n2935gat),.A(n892gat),.B(n891gat));
  OR2 OR2_96(.VSS(VSS),.VDD(VDD),.Y(n2942gat),.A(n904gat),.B(n903gat));
  OR4 OR4_44(.VSS(VSS),.VDD(VDD),.Y(n2940gat),.A(n1152gat),.B(n1092gat),.C(n997gat),.D(n993gat));
  OR2 OR2_97(.VSS(VSS),.VDD(VDD),.Y(n2937gat),.A(n900gat),.B(n895gat));
  OR4 OR4_45(.VSS(VSS),.VDD(VDD),.Y(n2947gat),.A(n1094gat),.B(n1093gat),.C(n988gat),.D(n984gat));
  OR2 OR2_98(.VSS(VSS),.VDD(VDD),.Y(n2965gat),.A(n1267gat),.B(n1257gat));
  OR2 OR2_99(.VSS(VSS),.VDD(VDD),.Y(n2956gat),.A(n1178gat),.B(n1116gat));
  OR2 OR2_100(.VSS(VSS),.VDD(VDD),.Y(n2961gat),.A(n1375gat),.B(n1324gat));
  OR4 OR4_46(.VSS(VSS),.VDD(VDD),.Y(n2939gat),.A(n1091gat),.B(n1088gat),.C(n992gat),.D(n987gat));
  OR2 OR2_101(.VSS(VSS),.VDD(VDD),.Y(n2938gat),.A(n899gat),.B(n896gat));
  OR2 OR2_102(.VSS(VSS),.VDD(VDD),.Y(n2967gat),.A(n1262gat),.B(n1260gat));
  OR4 OR4_47(.VSS(VSS),.VDD(VDD),.Y(n2932gat),.A(n1098gat),.B(n1090gat),.C(n986gat),.D(n885gat));
  OR2 OR2_103(.VSS(VSS),.VDD(VDD),.Y(n2936gat),.A(n901gat),.B(n893gat));
  OR4 OR4_48(.VSS(VSS),.VDD(VDD),.Y(n2948gat),.A(n1097gat),.B(n1089gat),.C(n1087gat),.D(n991gat));
  OR2 OR2_104(.VSS(VSS),.VDD(VDD),.Y(n2968gat),.A(n1326gat),.B(n1261gat));
  OR2 OR2_105(.VSS(VSS),.VDD(VDD),.Y(n2955gat),.A(n1177gat),.B(n1115gat));
  OR2 OR2_106(.VSS(VSS),.VDD(VDD),.Y(n2944gat),.A(n977gat),.B(n976gat));
  OR4 OR4_49(.VSS(VSS),.VDD(VDD),.Y(n2945gat),.A(n1096gat),.B(n1095gat),.C(n990gat),.D(n979gat));
  OR2 OR2_107(.VSS(VSS),.VDD(VDD),.Y(n2962gat),.A(n1176gat),.B(n1173gat));
  OR2 OR2_108(.VSS(VSS),.VDD(VDD),.Y(n2951gat),.A(n1004gat),.B(n1000gat));
  OR2 OR2_109(.VSS(VSS),.VDD(VDD),.Y(n2764gat),.A(n1029gat),.B(n2237gat));
  OR2 OR2_110(.VSS(VSS),.VDD(VDD),.Y(n2762gat),.A(n1028gat),.B(n1782gat));
  OR2 OR2_111(.VSS(VSS),.VDD(VDD),.Y(n2761gat),.A(n1031gat),.B(n2325gat));
  OR2 OR2_112(.VSS(VSS),.VDD(VDD),.Y(n2757gat),.A(n1030gat),.B(n2245gat));
  OR2 OR2_113(.VSS(VSS),.VDD(VDD),.Y(n2756gat),.A(n1011gat),.B(n2244gat));
  OR2 OR2_114(.VSS(VSS),.VDD(VDD),.Y(n2750gat),.A(n1181gat),.B(n2243gat));
  OR2 OR2_115(.VSS(VSS),.VDD(VDD),.Y(n2749gat),.A(n1010gat),.B(n2246gat));
  OR2 OR2_116(.VSS(VSS),.VDD(VDD),.Y(n2742gat),.A(n1005gat),.B(n2384gat));
  OR2 OR2_117(.VSS(VSS),.VDD(VDD),.Y(n2741gat),.A(n1182gat),.B(n2385gat));
  OR2 OR2_118(.VSS(VSS),.VDD(VDD),.Y(n2694gat),.A(n1381gat),.B(n1384gat));
  OR2 OR2_119(.VSS(VSS),.VDD(VDD),.Y(n2693gat),.A(n1451gat),.B(n1453gat));
  OR2 OR2_120(.VSS(VSS),.VDD(VDD),.Y(n2702gat),.A(n925gat),.B(n1452gat));
  OR2 OR2_121(.VSS(VSS),.VDD(VDD),.Y(n2701gat),.A(n921gat),.B(n1890gat));
  OR2 OR2_122(.VSS(VSS),.VDD(VDD),.Y(n2709gat),.A(n739gat),.B(n1841gat));
  OR2 OR2_123(.VSS(VSS),.VDD(VDD),.Y(n2708gat),.A(n848gat),.B(n2047gat));
  OR2 OR2_124(.VSS(VSS),.VDD(VDD),.Y(n2799gat),.A(n849gat),.B(n2050gat));
  OR2 OR2_125(.VSS(VSS),.VDD(VDD),.Y(n2798gat),.A(n1032gat),.B(n2054gat));
  OR3 OR3_61(.VSS(VSS),.VDD(VDD),.Y(n2812gat),.A(n73gat),.B(n70gat),.C(n1840gat));
  OR3 OR3_62(.VSS(VSS),.VDD(VDD),.Y(n2822gat),.A(n77gat),.B(n13gat),.C(n1842gat));
//
  NOR2 NOR2_0(.VSS(VSS),.VDD(VDD),.Y(n421gat),.A(n2715gat),.B(n2723gat));
  NOR2 NOR2_1(.VSS(VSS),.VDD(VDD),.Y(n648gat),.A(n373gat),.B(n2669gat));
  NOR2 NOR2_2(.VSS(VSS),.VDD(VDD),.Y(n442gat),.A(n2844gat),.B(n856gat));
  NOR2 NOR2_3(.VSS(VSS),.VDD(VDD),.Y(n1499gat),.A(n396gat),.B(n401gat));
  NOR2 NOR2_4(.VSS(VSS),.VDD(VDD),.Y(n1616gat),.A(n918gat),.B(n396gat));
  NOR2 NOR2_5(.VSS(VSS),.VDD(VDD),.Y(n1614gat),.A(n396gat),.B(n845gat));
  NOR3 NOR3_0(.VSS(VSS),.VDD(VDD),.Y(n1641gat),.A(n1645gat),.B(n1553gat),.C(n1559gat));
  NOR3 NOR3_1(.VSS(VSS),.VDD(VDD),.Y(n1642gat),.A(n1559gat),.B(n1616gat),.C(n1645gat));
  NOR3 NOR3_2(.VSS(VSS),.VDD(VDD),.Y(n1556gat),.A(n1614gat),.B(n1645gat),.C(n1616gat));
  NOR3 NOR3_3(.VSS(VSS),.VDD(VDD),.Y(n1557gat),.A(n1553gat),.B(n1645gat),.C(n1614gat));
  NOR3 NOR3_4(.VSS(VSS),.VDD(VDD),.Y(n1639gat),.A(n1499gat),.B(n1559gat),.C(n1553gat));
  NOR4 NOR4_0(.VSS(VSS),.VDD(VDD),.Y(n1605gat),.A(n1614gat),.B(n1616gat),.C(n1499gat),.D(n396gat));
  NOR3 NOR3_5(.VSS(VSS),.VDD(VDD),.Y(n1555gat),.A(n1616gat),.B(n1559gat),.C(n1499gat));
  NOR3 NOR3_6(.VSS(VSS),.VDD(VDD),.Y(n1558gat),.A(n1614gat),.B(n1553gat),.C(n1499gat));
  NOR2 NOR2_6(.VSS(VSS),.VDD(VDD),.Y(n1256gat),.A(n392gat),.B(n702gat));
  NOR2 NOR2_7(.VSS(VSS),.VDD(VDD),.Y(n1117gat),.A(n720gat),.B(n725gat));
  NOR2 NOR2_8(.VSS(VSS),.VDD(VDD),.Y(n1618gat),.A(n1319gat),.B(n1447gat));
  NOR2 NOR2_9(.VSS(VSS),.VDD(VDD),.Y(n1114gat),.A(n725gat),.B(n721gat));
  NOR2 NOR2_10(.VSS(VSS),.VDD(VDD),.Y(n1621gat),.A(n1319gat),.B(n1380gat));
  NOR2 NOR2_11(.VSS(VSS),.VDD(VDD),.Y(n1318gat),.A(n392gat),.B(n701gat));
  NOR2 NOR2_12(.VSS(VSS),.VDD(VDD),.Y(n1619gat),.A(n1447gat),.B(n1446gat));
  NOR2 NOR2_13(.VSS(VSS),.VDD(VDD),.Y(n1622gat),.A(n1380gat),.B(n1446gat));
  NOR3 NOR3_7(.VSS(VSS),.VDD(VDD),.Y(n1214gat),.A(n1218gat),.B(n1219gat),.C(n1220gat));
  NOR3 NOR3_8(.VSS(VSS),.VDD(VDD),.Y(n1215gat),.A(n1218gat),.B(n1221gat),.C(n1222gat));
  NOR3 NOR3_9(.VSS(VSS),.VDD(VDD),.Y(n1216gat),.A(n1223gat),.B(n1219gat),.C(n1222gat));
  NOR3 NOR3_10(.VSS(VSS),.VDD(VDD),.Y(n1217gat),.A(n1223gat),.B(n1221gat),.C(n1220gat));
  NOR2 NOR2_14(.VSS(VSS),.VDD(VDD),.Y(n745gat),.A(n2716gat),.B(n2867gat));
  NOR2 NOR2_15(.VSS(VSS),.VDD(VDD),.Y(n638gat),.A(n2715gat),.B(n2868gat));
  NOR2 NOR2_16(.VSS(VSS),.VDD(VDD),.Y(n423gat),.A(n2724gat),.B(n2726gat));
  NOR2 NOR2_17(.VSS(VSS),.VDD(VDD),.Y(n362gat),.A(n2723gat),.B(n2727gat));
  NOR3 NOR3_11(.VSS(VSS),.VDD(VDD),.Y(n749gat),.A(n753gat),.B(n754gat),.C(n755gat));
  NOR3 NOR3_12(.VSS(VSS),.VDD(VDD),.Y(n750gat),.A(n753gat),.B(n756gat),.C(n757gat));
  NOR3 NOR3_13(.VSS(VSS),.VDD(VDD),.Y(n751gat),.A(n758gat),.B(n754gat),.C(n757gat));
  NOR3 NOR3_14(.VSS(VSS),.VDD(VDD),.Y(n752gat),.A(n758gat),.B(n756gat),.C(n755gat));
  NOR3 NOR3_15(.VSS(VSS),.VDD(VDD),.Y(n259gat),.A(n263gat),.B(n264gat),.C(n265gat));
  NOR3 NOR3_16(.VSS(VSS),.VDD(VDD),.Y(n260gat),.A(n263gat),.B(n266gat),.C(n267gat));
  NOR3 NOR3_17(.VSS(VSS),.VDD(VDD),.Y(n261gat),.A(n268gat),.B(n264gat),.C(n267gat));
  NOR3 NOR3_18(.VSS(VSS),.VDD(VDD),.Y(n262gat),.A(n268gat),.B(n266gat),.C(n265gat));
  NOR3 NOR3_19(.VSS(VSS),.VDD(VDD),.Y(n1014gat),.A(n1018gat),.B(n1019gat),.C(n1020gat));
  NOR3 NOR3_20(.VSS(VSS),.VDD(VDD),.Y(n1015gat),.A(n1018gat),.B(n1021gat),.C(n1022gat));
  NOR3 NOR3_21(.VSS(VSS),.VDD(VDD),.Y(n1016gat),.A(n1023gat),.B(n1019gat),.C(n1022gat));
  NOR3 NOR3_22(.VSS(VSS),.VDD(VDD),.Y(n1017gat),.A(n1023gat),.B(n1021gat),.C(n1020gat));
  NOR3 NOR3_23(.VSS(VSS),.VDD(VDD),.Y(n476gat),.A(n480gat),.B(n481gat),.C(n482gat));
  NOR3 NOR3_24(.VSS(VSS),.VDD(VDD),.Y(n477gat),.A(n480gat),.B(n483gat),.C(n484gat));
  NOR3 NOR3_25(.VSS(VSS),.VDD(VDD),.Y(n478gat),.A(n485gat),.B(n481gat),.C(n484gat));
  NOR3 NOR3_26(.VSS(VSS),.VDD(VDD),.Y(n479gat),.A(n485gat),.B(n483gat),.C(n482gat));
  NOR3 NOR3_27(.VSS(VSS),.VDD(VDD),.Y(n44gat),.A(n48gat),.B(n49gat),.C(n50gat));
  NOR3 NOR3_28(.VSS(VSS),.VDD(VDD),.Y(n45gat),.A(n48gat),.B(n51gat),.C(n52gat));
  NOR3 NOR3_29(.VSS(VSS),.VDD(VDD),.Y(n46gat),.A(n53gat),.B(n49gat),.C(n52gat));
  NOR3 NOR3_30(.VSS(VSS),.VDD(VDD),.Y(n47gat),.A(n53gat),.B(n51gat),.C(n50gat));
  NOR2 NOR2_18(.VSS(VSS),.VDD(VDD),.Y(n1376gat),.A(n724gat),.B(n720gat));
  NOR2 NOR2_19(.VSS(VSS),.VDD(VDD),.Y(n1617gat),.A(n1319gat),.B(n1448gat));
  NOR2 NOR2_20(.VSS(VSS),.VDD(VDD),.Y(n1377gat),.A(n724gat),.B(n721gat));
  NOR2 NOR2_21(.VSS(VSS),.VDD(VDD),.Y(n1624gat),.A(n1319gat),.B(n1379gat));
  NOR2 NOR2_22(.VSS(VSS),.VDD(VDD),.Y(n1113gat),.A(n393gat),.B(n701gat));
  NOR2 NOR2_23(.VSS(VSS),.VDD(VDD),.Y(n1501gat),.A(n1448gat),.B(n1500gat));
  NOR2 NOR2_24(.VSS(VSS),.VDD(VDD),.Y(n1623gat),.A(n1379gat),.B(n1446gat));
  NOR2 NOR2_25(.VSS(VSS),.VDD(VDD),.Y(n1620gat),.A(n1448gat),.B(n1446gat));
  NOR2 NOR2_26(.VSS(VSS),.VDD(VDD),.Y(n1827gat),.A(n2729gat),.B(n2317gat));
  NOR2 NOR2_27(.VSS(VSS),.VDD(VDD),.Y(n1817gat),.A(n1819gat),.B(n1823gat));
  NOR2 NOR2_28(.VSS(VSS),.VDD(VDD),.Y(n1935gat),.A(n1816gat),.B(n1828gat));
  NOR2 NOR2_29(.VSS(VSS),.VDD(VDD),.Y(n529gat),.A(n2724gat),.B(n2715gat));
  NOR2 NOR2_30(.VSS(VSS),.VDD(VDD),.Y(n361gat),.A(n2859gat),.B(n2726gat));
  NOR3 NOR3_31(.VSS(VSS),.VDD(VDD),.Y(n168gat),.A(n172gat),.B(n173gat),.C(n174gat));
  NOR3 NOR3_32(.VSS(VSS),.VDD(VDD),.Y(n169gat),.A(n172gat),.B(n175gat),.C(n176gat));
  NOR3 NOR3_33(.VSS(VSS),.VDD(VDD),.Y(n170gat),.A(n177gat),.B(n173gat),.C(n176gat));
  NOR3 NOR3_34(.VSS(VSS),.VDD(VDD),.Y(n171gat),.A(n177gat),.B(n175gat),.C(n174gat));
  NOR3 NOR3_35(.VSS(VSS),.VDD(VDD),.Y(n907gat),.A(n911gat),.B(n912gat),.C(n913gat));
  NOR3 NOR3_36(.VSS(VSS),.VDD(VDD),.Y(n908gat),.A(n911gat),.B(n914gat),.C(n915gat));
  NOR3 NOR3_37(.VSS(VSS),.VDD(VDD),.Y(n909gat),.A(n916gat),.B(n912gat),.C(n915gat));
  NOR3 NOR3_38(.VSS(VSS),.VDD(VDD),.Y(n910gat),.A(n916gat),.B(n914gat),.C(n913gat));
  NOR3 NOR3_39(.VSS(VSS),.VDD(VDD),.Y(n344gat),.A(n348gat),.B(n349gat),.C(n350gat));
  NOR3 NOR3_40(.VSS(VSS),.VDD(VDD),.Y(n345gat),.A(n348gat),.B(n351gat),.C(n352gat));
  NOR3 NOR3_41(.VSS(VSS),.VDD(VDD),.Y(n346gat),.A(n353gat),.B(n349gat),.C(n352gat));
  NOR3 NOR3_42(.VSS(VSS),.VDD(VDD),.Y(n347gat),.A(n353gat),.B(n351gat),.C(n350gat));
  NOR3 NOR3_43(.VSS(VSS),.VDD(VDD),.Y(n56gat),.A(n60gat),.B(n61gat),.C(n62gat));
  NOR3 NOR3_44(.VSS(VSS),.VDD(VDD),.Y(n57gat),.A(n60gat),.B(n63gat),.C(n64gat));
  NOR3 NOR3_45(.VSS(VSS),.VDD(VDD),.Y(n58gat),.A(n65gat),.B(n61gat),.C(n64gat));
  NOR3 NOR3_46(.VSS(VSS),.VDD(VDD),.Y(n59gat),.A(n65gat),.B(n63gat),.C(n62gat));
  NOR2 NOR2_31(.VSS(VSS),.VDD(VDD),.Y(n768gat),.A(n373gat),.B(n2731gat));
  NOR2 NOR2_32(.VSS(VSS),.VDD(VDD),.Y(n655gat),.A(n856gat),.B(n2718gat));
  NOR2 NOR2_33(.VSS(VSS),.VDD(VDD),.Y(n963gat),.A(n856gat),.B(n2838gat));
  NOR2 NOR2_34(.VSS(VSS),.VDD(VDD),.Y(n868gat),.A(n2775gat),.B(n373gat));
  NOR2 NOR2_35(.VSS(VSS),.VDD(VDD),.Y(n962gat),.A(n856gat),.B(n2711gat));
  NOR2 NOR2_36(.VSS(VSS),.VDD(VDD),.Y(n959gat),.A(n373gat),.B(n2734gat));
  NOR3 NOR3_47(.VSS(VSS),.VDD(VDD),.Y(n945gat),.A(n949gat),.B(n950gat),.C(n951gat));
  NOR3 NOR3_48(.VSS(VSS),.VDD(VDD),.Y(n946gat),.A(n949gat),.B(n952gat),.C(n953gat));
  NOR3 NOR3_49(.VSS(VSS),.VDD(VDD),.Y(n947gat),.A(n954gat),.B(n950gat),.C(n953gat));
  NOR3 NOR3_50(.VSS(VSS),.VDD(VDD),.Y(n948gat),.A(n954gat),.B(n952gat),.C(n951gat));
  NOR2 NOR2_37(.VSS(VSS),.VDD(VDD),.Y(n647gat),.A(n2792gat),.B(n373gat));
  NOR2 NOR2_38(.VSS(VSS),.VDD(VDD),.Y(n441gat),.A(n856gat),.B(n2846gat));
  NOR2 NOR2_39(.VSS(VSS),.VDD(VDD),.Y(n967gat),.A(n373gat),.B(n2672gat));
  NOR2 NOR2_40(.VSS(VSS),.VDD(VDD),.Y(n792gat),.A(n2852gat),.B(n856gat));
  NOR3 NOR3_51(.VSS(VSS),.VDD(VDD),.Y(n1229gat),.A(n1233gat),.B(n1234gat),.C(n1235gat));
  NOR3 NOR3_52(.VSS(VSS),.VDD(VDD),.Y(n1230gat),.A(n1233gat),.B(n1236gat),.C(n1237gat));
  NOR3 NOR3_53(.VSS(VSS),.VDD(VDD),.Y(n1231gat),.A(n1238gat),.B(n1234gat),.C(n1237gat));
  NOR3 NOR3_54(.VSS(VSS),.VDD(VDD),.Y(n1232gat),.A(n1238gat),.B(n1236gat),.C(n1235gat));
  NOR2 NOR2_41(.VSS(VSS),.VDD(VDD),.Y(n443gat),.A(n2778gat),.B(n373gat));
  NOR2 NOR2_42(.VSS(VSS),.VDD(VDD),.Y(n439gat),.A(n856gat),.B(n2836gat));
  NOR2 NOR2_43(.VSS(VSS),.VDD(VDD),.Y(n966gat),.A(n2789gat),.B(n373gat));
  NOR2 NOR2_44(.VSS(VSS),.VDD(VDD),.Y(n790gat),.A(n856gat),.B(n2840gat));
  NOR2 NOR2_45(.VSS(VSS),.VDD(VDD),.Y(n444gat),.A(n373gat),.B(n2781gat));
  NOR2 NOR2_46(.VSS(VSS),.VDD(VDD),.Y(n440gat),.A(n856gat),.B(n2842gat));
  NOR3 NOR3_55(.VSS(VSS),.VDD(VDD),.Y(n1051gat),.A(n1055gat),.B(n1056gat),.C(n1057gat));
  NOR3 NOR3_56(.VSS(VSS),.VDD(VDD),.Y(n1052gat),.A(n1055gat),.B(n1058gat),.C(n1059gat));
  NOR3 NOR3_57(.VSS(VSS),.VDD(VDD),.Y(n1053gat),.A(n1060gat),.B(n1056gat),.C(n1059gat));
  NOR3 NOR3_58(.VSS(VSS),.VDD(VDD),.Y(n1054gat),.A(n1060gat),.B(n1058gat),.C(n1057gat));
  NOR3 NOR3_59(.VSS(VSS),.VDD(VDD),.Y(n934gat),.A(n938gat),.B(n939gat),.C(n940gat));
  NOR3 NOR3_60(.VSS(VSS),.VDD(VDD),.Y(n935gat),.A(n938gat),.B(n941gat),.C(n942gat));
  NOR3 NOR3_61(.VSS(VSS),.VDD(VDD),.Y(n936gat),.A(n943gat),.B(n939gat),.C(n942gat));
  NOR3 NOR3_62(.VSS(VSS),.VDD(VDD),.Y(n937gat),.A(n943gat),.B(n941gat),.C(n940gat));
  NOR2 NOR2_47(.VSS(VSS),.VDD(VDD),.Y(n746gat),.A(n2716gat),.B(n2723gat));
  NOR2 NOR2_48(.VSS(VSS),.VDD(VDD),.Y(n360gat),.A(n2859gat),.B(n2727gat));
  NOR3 NOR3_63(.VSS(VSS),.VDD(VDD),.Y(n710gat),.A(n714gat),.B(n715gat),.C(n716gat));
  NOR3 NOR3_64(.VSS(VSS),.VDD(VDD),.Y(n711gat),.A(n714gat),.B(n717gat),.C(n718gat));
  NOR3 NOR3_65(.VSS(VSS),.VDD(VDD),.Y(n712gat),.A(n719gat),.B(n715gat),.C(n718gat));
  NOR3 NOR3_66(.VSS(VSS),.VDD(VDD),.Y(n713gat),.A(n719gat),.B(n717gat),.C(n716gat));
  NOR3 NOR3_67(.VSS(VSS),.VDD(VDD),.Y(n729gat),.A(n733gat),.B(n734gat),.C(n735gat));
  NOR3 NOR3_68(.VSS(VSS),.VDD(VDD),.Y(n730gat),.A(n733gat),.B(n736gat),.C(n737gat));
  NOR3 NOR3_69(.VSS(VSS),.VDD(VDD),.Y(n731gat),.A(n738gat),.B(n734gat),.C(n737gat));
  NOR3 NOR3_70(.VSS(VSS),.VDD(VDD),.Y(n732gat),.A(n738gat),.B(n736gat),.C(n735gat));
  NOR3 NOR3_71(.VSS(VSS),.VDD(VDD),.Y(n494gat),.A(n498gat),.B(n499gat),.C(n500gat));
  NOR3 NOR3_72(.VSS(VSS),.VDD(VDD),.Y(n495gat),.A(n498gat),.B(n501gat),.C(n502gat));
  NOR3 NOR3_73(.VSS(VSS),.VDD(VDD),.Y(n496gat),.A(n503gat),.B(n499gat),.C(n502gat));
  NOR3 NOR3_74(.VSS(VSS),.VDD(VDD),.Y(n497gat),.A(n503gat),.B(n501gat),.C(n500gat));
  NOR3 NOR3_75(.VSS(VSS),.VDD(VDD),.Y(n505gat),.A(n509gat),.B(n510gat),.C(n511gat));
  NOR3 NOR3_76(.VSS(VSS),.VDD(VDD),.Y(n506gat),.A(n509gat),.B(n512gat),.C(n513gat));
  NOR3 NOR3_77(.VSS(VSS),.VDD(VDD),.Y(n507gat),.A(n514gat),.B(n510gat),.C(n513gat));
  NOR3 NOR3_78(.VSS(VSS),.VDD(VDD),.Y(n508gat),.A(n514gat),.B(n512gat),.C(n511gat));
  NOR4 NOR4_1(.VSS(VSS),.VDD(VDD),.Y(n564gat),.A(n3029gat),.B(n2863gat),.C(n2855gat),.D(n374gat));
  NOR3 NOR3_79(.VSS(VSS),.VDD(VDD),.Y(n86gat),.A(n743gat),.B(n294gat),.C(n17gat));
  NOR2 NOR2_49(.VSS(VSS),.VDD(VDD),.Y(n78gat),.A(n2784gat),.B(n79gat));
  NOR2 NOR2_50(.VSS(VSS),.VDD(VDD),.Y(n767gat),.A(n219gat),.B(n2731gat));
  NOR2 NOR2_51(.VSS(VSS),.VDD(VDD),.Y(n286gat),.A(n289gat),.B(n2723gat));
  NOR2 NOR2_52(.VSS(VSS),.VDD(VDD),.Y(n287gat),.A(n289gat),.B(n2715gat));
  NOR2 NOR2_53(.VSS(VSS),.VDD(VDD),.Y(n288gat),.A(n289gat),.B(n2726gat));
  NOR3 NOR3_80(.VSS(VSS),.VDD(VDD),.Y(n181gat),.A(n286gat),.B(n179gat),.C(n188gat));
  NOR2 NOR2_54(.VSS(VSS),.VDD(VDD),.Y(n182gat),.A(n72gat),.B(n2720gat));
  NOR2 NOR2_55(.VSS(VSS),.VDD(VDD),.Y(n653gat),.A(n2718gat),.B(n111gat));
  NOR2 NOR2_56(.VSS(VSS),.VDD(VDD),.Y(n867gat),.A(n219gat),.B(n2775gat));
  NOR2 NOR2_57(.VSS(VSS),.VDD(VDD),.Y(n771gat),.A(n2838gat),.B(n111gat));
  NOR2 NOR2_58(.VSS(VSS),.VDD(VDD),.Y(n964gat),.A(n111gat),.B(n2711gat));
  NOR2 NOR2_59(.VSS(VSS),.VDD(VDD),.Y(n961gat),.A(n219gat),.B(n2734gat));
  NOR3 NOR3_81(.VSS(VSS),.VDD(VDD),.Y(n804gat),.A(n808gat),.B(n809gat),.C(n810gat));
  NOR3 NOR3_82(.VSS(VSS),.VDD(VDD),.Y(n805gat),.A(n808gat),.B(n811gat),.C(n812gat));
  NOR3 NOR3_83(.VSS(VSS),.VDD(VDD),.Y(n806gat),.A(n813gat),.B(n809gat),.C(n812gat));
  NOR3 NOR3_84(.VSS(VSS),.VDD(VDD),.Y(n807gat),.A(n813gat),.B(n811gat),.C(n810gat));
  NOR3 NOR3_85(.VSS(VSS),.VDD(VDD),.Y(n587gat),.A(n591gat),.B(n592gat),.C(n593gat));
  NOR3 NOR3_86(.VSS(VSS),.VDD(VDD),.Y(n588gat),.A(n591gat),.B(n594gat),.C(n595gat));
  NOR3 NOR3_87(.VSS(VSS),.VDD(VDD),.Y(n589gat),.A(n596gat),.B(n592gat),.C(n595gat));
  NOR3 NOR3_88(.VSS(VSS),.VDD(VDD),.Y(n590gat),.A(n596gat),.B(n594gat),.C(n593gat));
  NOR2 NOR2_60(.VSS(VSS),.VDD(VDD),.Y(n447gat),.A(n2836gat),.B(n111gat));
  NOR2 NOR2_61(.VSS(VSS),.VDD(VDD),.Y(n445gat),.A(n2778gat),.B(n219gat));
  NOR3 NOR3_89(.VSS(VSS),.VDD(VDD),.Y(n687gat),.A(n691gat),.B(n692gat),.C(n693gat));
  NOR3 NOR3_90(.VSS(VSS),.VDD(VDD),.Y(n688gat),.A(n691gat),.B(n694gat),.C(n695gat));
  NOR3 NOR3_91(.VSS(VSS),.VDD(VDD),.Y(n689gat),.A(n696gat),.B(n692gat),.C(n695gat));
  NOR3 NOR3_92(.VSS(VSS),.VDD(VDD),.Y(n690gat),.A(n696gat),.B(n694gat),.C(n693gat));
  NOR3 NOR3_93(.VSS(VSS),.VDD(VDD),.Y(n568gat),.A(n572gat),.B(n573gat),.C(n574gat));
  NOR3 NOR3_94(.VSS(VSS),.VDD(VDD),.Y(n569gat),.A(n572gat),.B(n575gat),.C(n576gat));
  NOR3 NOR3_95(.VSS(VSS),.VDD(VDD),.Y(n570gat),.A(n577gat),.B(n573gat),.C(n576gat));
  NOR3 NOR3_96(.VSS(VSS),.VDD(VDD),.Y(n571gat),.A(n577gat),.B(n575gat),.C(n574gat));
  NOR3 NOR3_97(.VSS(VSS),.VDD(VDD),.Y(n187gat),.A(n189gat),.B(n287gat),.C(n188gat));
  NOR2 NOR2_62(.VSS(VSS),.VDD(VDD),.Y(n197gat),.A(n194gat),.B(n297gat));
  NOR3 NOR3_98(.VSS(VSS),.VDD(VDD),.Y(n15gat),.A(n637gat),.B(n17gat),.C(n293gat));
  NOR2 NOR2_63(.VSS(VSS),.VDD(VDD),.Y(n22gat),.A(n92gat),.B(n21gat));
  NOR2 NOR2_64(.VSS(VSS),.VDD(VDD),.Y(n93gat),.A(n197gat),.B(n22gat));
  NOR2 NOR2_65(.VSS(VSS),.VDD(VDD),.Y(n769gat),.A(n93gat),.B(n2731gat));
  NOR3 NOR3_99(.VSS(VSS),.VDD(VDD),.Y(n2534gat),.A(n2624gat),.B(n2489gat),.C(n2621gat));
  NOR3 NOR3_100(.VSS(VSS),.VDD(VDD),.Y(n2430gat),.A(n2533gat),.B(n2486gat),.C(n2429gat));
  NOR2 NOR2_66(.VSS(VSS),.VDD(VDD),.Y(n1606gat),.A(n3020gat),.B(n270gat));
  NOR2 NOR2_67(.VSS(VSS),.VDD(VDD),.Y(n2239gat),.A(n2850gat),.B(n3019gat));
  NOR3 NOR3_101(.VSS(VSS),.VDD(VDD),.Y(n1934gat),.A(n2470gat),.B(n1935gat),.C(n2239gat));
  NOR2 NOR2_68(.VSS(VSS),.VDD(VDD),.Y(n1610gat),.A(n1698gat),.B(n1543gat));
  NOR2 NOR2_69(.VSS(VSS),.VDD(VDD),.Y(n1692gat),.A(n1879gat),.B(n1762gat));
  NOR2 NOR2_70(.VSS(VSS),.VDD(VDD),.Y(n2433gat),.A(n2432gat),.B(n2154gat));
  NOR3 NOR3_102(.VSS(VSS),.VDD(VDD),.Y(n2531gat),.A(n2488gat),.B(n2625gat),.C(n2621gat));
  NOR3 NOR3_103(.VSS(VSS),.VDD(VDD),.Y(n2480gat),.A(n2530gat),.B(n2482gat),.C(n2486gat));
  NOR2 NOR2_71(.VSS(VSS),.VDD(VDD),.Y(n2427gat),.A(n2426gat),.B(n2153gat));
  NOR2 NOR2_72(.VSS(VSS),.VDD(VDD),.Y(n2428gat),.A(n2433gat),.B(n2427gat));
  NOR2 NOR2_73(.VSS(VSS),.VDD(VDD),.Y(n1778gat),.A(n3026gat),.B(n1779gat));
  NOR2 NOR2_74(.VSS(VSS),.VDD(VDD),.Y(n1609gat),.A(n1503gat),.B(n3025gat));
  NOR2 NOR2_75(.VSS(VSS),.VDD(VDD),.Y(n1702gat),.A(n3024gat),.B(n1615gat));
  NOR2 NOR2_76(.VSS(VSS),.VDD(VDD),.Y(n1700gat),.A(n1701gat),.B(n3023gat));
  NOR4 NOR4_2(.VSS(VSS),.VDD(VDD),.Y(n1604gat),.A(n1778gat),.B(n1609gat),.C(n1702gat),.D(n1700gat));
  NOR2 NOR2_77(.VSS(VSS),.VDD(VDD),.Y(n1076gat),.A(n93gat),.B(n2775gat));
  NOR2 NOR2_78(.VSS(VSS),.VDD(VDD),.Y(n766gat),.A(n93gat),.B(n2734gat));
  NOR3 NOR3_104(.VSS(VSS),.VDD(VDD),.Y(n1185gat),.A(n1189gat),.B(n1190gat),.C(n1191gat));
  NOR3 NOR3_105(.VSS(VSS),.VDD(VDD),.Y(n1186gat),.A(n1189gat),.B(n1192gat),.C(n1193gat));
  NOR3 NOR3_106(.VSS(VSS),.VDD(VDD),.Y(n1187gat),.A(n1194gat),.B(n1190gat),.C(n1193gat));
  NOR3 NOR3_107(.VSS(VSS),.VDD(VDD),.Y(n1188gat),.A(n1194gat),.B(n1192gat),.C(n1191gat));
  NOR2 NOR2_79(.VSS(VSS),.VDD(VDD),.Y(n645gat),.A(n2792gat),.B(n93gat));
  NOR2 NOR2_80(.VSS(VSS),.VDD(VDD),.Y(n646gat),.A(n93gat),.B(n2669gat));
  NOR2 NOR2_81(.VSS(VSS),.VDD(VDD),.Y(n1383gat),.A(n1280gat),.B(n1225gat));
  NOR2 NOR2_82(.VSS(VSS),.VDD(VDD),.Y(n1327gat),.A(n1281gat),.B(n1224gat));
  NOR2 NOR2_83(.VSS(VSS),.VDD(VDD),.Y(n651gat),.A(n93gat),.B(n2778gat));
  NOR2 NOR2_84(.VSS(VSS),.VDD(VDD),.Y(n652gat),.A(n2789gat),.B(n93gat));
  NOR2 NOR2_85(.VSS(VSS),.VDD(VDD),.Y(n765gat),.A(n2781gat),.B(n93gat));
  NOR3 NOR3_108(.VSS(VSS),.VDD(VDD),.Y(n1202gat),.A(n1206gat),.B(n1207gat),.C(n1208gat));
  NOR3 NOR3_109(.VSS(VSS),.VDD(VDD),.Y(n1203gat),.A(n1206gat),.B(n1209gat),.C(n1210gat));
  NOR3 NOR3_110(.VSS(VSS),.VDD(VDD),.Y(n1204gat),.A(n1211gat),.B(n1207gat),.C(n1210gat));
  NOR3 NOR3_111(.VSS(VSS),.VDD(VDD),.Y(n1205gat),.A(n1211gat),.B(n1209gat),.C(n1208gat));
  NOR3 NOR3_112(.VSS(VSS),.VDD(VDD),.Y(n1270gat),.A(n1274gat),.B(n1275gat),.C(n1276gat));
  NOR3 NOR3_113(.VSS(VSS),.VDD(VDD),.Y(n1271gat),.A(n1274gat),.B(n1277gat),.C(n1278gat));
  NOR3 NOR3_114(.VSS(VSS),.VDD(VDD),.Y(n1272gat),.A(n1279gat),.B(n1275gat),.C(n1278gat));
  NOR3 NOR3_115(.VSS(VSS),.VDD(VDD),.Y(n1273gat),.A(n1279gat),.B(n1277gat),.C(n1276gat));
  NOR2 NOR2_86(.VSS(VSS),.VDD(VDD),.Y(n763gat),.A(n2672gat),.B(n93gat));
  NOR2 NOR2_87(.VSS(VSS),.VDD(VDD),.Y(n1287gat),.A(n1284gat),.B(n1195gat));
  NOR2 NOR2_88(.VSS(VSS),.VDD(VDD),.Y(n1285gat),.A(n1196gat),.B(n1269gat));
  NOR2 NOR2_89(.VSS(VSS),.VDD(VDD),.Y(n853gat),.A(n740gat),.B(n2148gat));
  NOR2 NOR2_90(.VSS(VSS),.VDD(VDD),.Y(n793gat),.A(n2852gat),.B(n851gat));
  NOR2 NOR2_91(.VSS(VSS),.VDD(VDD),.Y(n854gat),.A(n2148gat),.B(n374gat));
  NOR2 NOR2_92(.VSS(VSS),.VDD(VDD),.Y(n556gat),.A(n2672gat),.B(n852gat));
  NOR2 NOR2_93(.VSS(VSS),.VDD(VDD),.Y(n795gat),.A(n2731gat),.B(n852gat));
  NOR2 NOR2_94(.VSS(VSS),.VDD(VDD),.Y(n656gat),.A(n851gat),.B(n2718gat));
  NOR2 NOR2_95(.VSS(VSS),.VDD(VDD),.Y(n794gat),.A(n852gat),.B(n2775gat));
  NOR2 NOR2_96(.VSS(VSS),.VDD(VDD),.Y(n773gat),.A(n851gat),.B(n2838gat));
  NOR2 NOR2_97(.VSS(VSS),.VDD(VDD),.Y(n965gat),.A(n2711gat),.B(n851gat));
  NOR2 NOR2_98(.VSS(VSS),.VDD(VDD),.Y(n960gat),.A(n2734gat),.B(n852gat));
  NOR3 NOR3_116(.VSS(VSS),.VDD(VDD),.Y(n780gat),.A(n784gat),.B(n785gat),.C(n786gat));
  NOR3 NOR3_117(.VSS(VSS),.VDD(VDD),.Y(n781gat),.A(n784gat),.B(n787gat),.C(n788gat));
  NOR3 NOR3_118(.VSS(VSS),.VDD(VDD),.Y(n782gat),.A(n789gat),.B(n785gat),.C(n788gat));
  NOR3 NOR3_119(.VSS(VSS),.VDD(VDD),.Y(n783gat),.A(n789gat),.B(n787gat),.C(n786gat));
  NOR2 NOR2_99(.VSS(VSS),.VDD(VDD),.Y(n555gat),.A(n852gat),.B(n2792gat));
  NOR2 NOR2_100(.VSS(VSS),.VDD(VDD),.Y(n450gat),.A(n851gat),.B(n2846gat));
  NOR2 NOR2_101(.VSS(VSS),.VDD(VDD),.Y(n654gat),.A(n851gat),.B(n2844gat));
  NOR2 NOR2_102(.VSS(VSS),.VDD(VDD),.Y(n557gat),.A(n2669gat),.B(n852gat));
  NOR2 NOR2_103(.VSS(VSS),.VDD(VDD),.Y(n874gat),.A(n559gat),.B(n365gat));
  NOR2 NOR2_104(.VSS(VSS),.VDD(VDD),.Y(n132gat),.A(n560gat),.B(n364gat));
  NOR2 NOR2_105(.VSS(VSS),.VDD(VDD),.Y(n649gat),.A(n2778gat),.B(n852gat));
  NOR2 NOR2_106(.VSS(VSS),.VDD(VDD),.Y(n449gat),.A(n2836gat),.B(n851gat));
  NOR2 NOR2_107(.VSS(VSS),.VDD(VDD),.Y(n791gat),.A(n851gat),.B(n2840gat));
  NOR2 NOR2_108(.VSS(VSS),.VDD(VDD),.Y(n650gat),.A(n852gat),.B(n2789gat));
  NOR2 NOR2_109(.VSS(VSS),.VDD(VDD),.Y(n774gat),.A(n2842gat),.B(n851gat));
  NOR2 NOR2_110(.VSS(VSS),.VDD(VDD),.Y(n764gat),.A(n852gat),.B(n2781gat));
  NOR3 NOR3_120(.VSS(VSS),.VDD(VDD),.Y(n222gat),.A(n226gat),.B(n227gat),.C(n228gat));
  NOR3 NOR3_121(.VSS(VSS),.VDD(VDD),.Y(n223gat),.A(n226gat),.B(n229gat),.C(n230gat));
  NOR3 NOR3_122(.VSS(VSS),.VDD(VDD),.Y(n224gat),.A(n231gat),.B(n227gat),.C(n230gat));
  NOR3 NOR3_123(.VSS(VSS),.VDD(VDD),.Y(n225gat),.A(n231gat),.B(n229gat),.C(n228gat));
  NOR3 NOR3_124(.VSS(VSS),.VDD(VDD),.Y(n121gat),.A(n125gat),.B(n126gat),.C(n127gat));
  NOR3 NOR3_125(.VSS(VSS),.VDD(VDD),.Y(n122gat),.A(n125gat),.B(n128gat),.C(n129gat));
  NOR3 NOR3_126(.VSS(VSS),.VDD(VDD),.Y(n123gat),.A(n130gat),.B(n126gat),.C(n129gat));
  NOR3 NOR3_127(.VSS(VSS),.VDD(VDD),.Y(n124gat),.A(n130gat),.B(n128gat),.C(n127gat));
  NOR2 NOR2_111(.VSS(VSS),.VDD(VDD),.Y(n2460gat),.A(n666gat),.B(n120gat));
  NOR2 NOR2_112(.VSS(VSS),.VDD(VDD),.Y(n2423gat),.A(n665gat),.B(n1601gat));
  NOR3 NOR3_128(.VSS(VSS),.VDD(VDD),.Y(n2594gat),.A(n3017gat),.B(n2520gat),.C(n2597gat));
  NOR3 NOR3_129(.VSS(VSS),.VDD(VDD),.Y(n2569gat),.A(n2573gat),.B(n2574gat),.C(n2575gat));
  NOR3 NOR3_130(.VSS(VSS),.VDD(VDD),.Y(n2570gat),.A(n2573gat),.B(n2576gat),.C(n2577gat));
  NOR3 NOR3_131(.VSS(VSS),.VDD(VDD),.Y(n2571gat),.A(n2578gat),.B(n2574gat),.C(n2577gat));
  NOR3 NOR3_132(.VSS(VSS),.VDD(VDD),.Y(n2572gat),.A(n2578gat),.B(n2576gat),.C(n2575gat));
  NOR3 NOR3_133(.VSS(VSS),.VDD(VDD),.Y(n2410gat),.A(n2414gat),.B(n2415gat),.C(n2416gat));
  NOR3 NOR3_134(.VSS(VSS),.VDD(VDD),.Y(n2411gat),.A(n2414gat),.B(n2417gat),.C(n2418gat));
  NOR3 NOR3_135(.VSS(VSS),.VDD(VDD),.Y(n2412gat),.A(n2419gat),.B(n2415gat),.C(n2418gat));
  NOR3 NOR3_136(.VSS(VSS),.VDD(VDD),.Y(n2413gat),.A(n2419gat),.B(n2417gat),.C(n2416gat));
  NOR2 NOR2_113(.VSS(VSS),.VDD(VDD),.Y(n2583gat),.A(n2582gat),.B(n2585gat));
  NOR2 NOR2_114(.VSS(VSS),.VDD(VDD),.Y(n2580gat),.A(n2582gat),.B(n2583gat));
  NOR2 NOR2_115(.VSS(VSS),.VDD(VDD),.Y(n2581gat),.A(n2583gat),.B(n2585gat));
  NOR2 NOR2_116(.VSS(VSS),.VDD(VDD),.Y(n2567gat),.A(n2493gat),.B(n2388gat));
  NOR2 NOR2_117(.VSS(VSS),.VDD(VDD),.Y(n2499gat),.A(n2389gat),.B(n2494gat));
  NOR2 NOR2_118(.VSS(VSS),.VDD(VDD),.Y(n299gat),.A(n2268gat),.B(n2338gat));
  NOR2 NOR2_119(.VSS(VSS),.VDD(VDD),.Y(n207gat),.A(n2337gat),.B(n2269gat));
  NOR2 NOR2_120(.VSS(VSS),.VDD(VDD),.Y(n2650gat),.A(n2649gat),.B(n2652gat));
  NOR2 NOR2_121(.VSS(VSS),.VDD(VDD),.Y(n2647gat),.A(n2649gat),.B(n2650gat));
  NOR2 NOR2_122(.VSS(VSS),.VDD(VDD),.Y(n2648gat),.A(n2650gat),.B(n2652gat));
  NOR3 NOR3_137(.VSS(VSS),.VDD(VDD),.Y(n2602gat),.A(n2606gat),.B(n2607gat),.C(n2608gat));
  NOR3 NOR3_138(.VSS(VSS),.VDD(VDD),.Y(n2603gat),.A(n2606gat),.B(n2609gat),.C(n2610gat));
  NOR3 NOR3_139(.VSS(VSS),.VDD(VDD),.Y(n2604gat),.A(n2611gat),.B(n2607gat),.C(n2610gat));
  NOR3 NOR3_140(.VSS(VSS),.VDD(VDD),.Y(n2605gat),.A(n2611gat),.B(n2609gat),.C(n2608gat));
  NOR3 NOR3_141(.VSS(VSS),.VDD(VDD),.Y(n2546gat),.A(n2550gat),.B(n2551gat),.C(n2552gat));
  NOR3 NOR3_142(.VSS(VSS),.VDD(VDD),.Y(n2547gat),.A(n2550gat),.B(n2553gat),.C(n2554gat));
  NOR3 NOR3_143(.VSS(VSS),.VDD(VDD),.Y(n2548gat),.A(n2555gat),.B(n2551gat),.C(n2554gat));
  NOR3 NOR3_144(.VSS(VSS),.VDD(VDD),.Y(n2549gat),.A(n2555gat),.B(n2553gat),.C(n2552gat));
  NOR2 NOR2_123(.VSS(VSS),.VDD(VDD),.Y(n2617gat),.A(n2616gat),.B(n2619gat));
  NOR2 NOR2_124(.VSS(VSS),.VDD(VDD),.Y(n2614gat),.A(n2616gat),.B(n2617gat));
  NOR2 NOR2_125(.VSS(VSS),.VDD(VDD),.Y(n2615gat),.A(n2617gat),.B(n2619gat));
  NOR4 NOR4_3(.VSS(VSS),.VDD(VDD),.Y(n2655gat),.A(n2508gat),.B(n2656gat),.C(n2500gat),.D(n2504gat));
  NOR3 NOR3_145(.VSS(VSS),.VDD(VDD),.Y(n2293gat),.A(n2353gat),.B(n2284gat),.C(n2443gat));
  NOR2 NOR2_126(.VSS(VSS),.VDD(VDD),.Y(n2219gat),.A(n2354gat),.B(n2214gat));
  NOR2 NOR2_127(.VSS(VSS),.VDD(VDD),.Y(n1529gat),.A(n1528gat),.B(n1523gat));
  NOR2 NOR2_128(.VSS(VSS),.VDD(VDD),.Y(n1704gat),.A(n3027gat),.B(n1706gat));
  NOR2 NOR2_129(.VSS(VSS),.VDD(VDD),.Y(n2461gat),.A(n120gat),.B(n2666gat));
  NOR2 NOR2_130(.VSS(VSS),.VDD(VDD),.Y(n2421gat),.A(n1601gat),.B(n1704gat));
  NOR2 NOR2_131(.VSS(VSS),.VDD(VDD),.Y(n1598gat),.A(n1592gat),.B(n2422gat));
  NOR2 NOR2_132(.VSS(VSS),.VDD(VDD),.Y(n2218gat),.A(n2214gat),.B(n2290gat));
  NOR3 NOR3_146(.VSS(VSS),.VDD(VDD),.Y(n2358gat),.A(n2285gat),.B(n2356gat),.C(n2355gat));
  NOR2 NOR2_133(.VSS(VSS),.VDD(VDD),.Y(n1415gat),.A(n2081gat),.B(n2359gat));
  NOR2 NOR2_134(.VSS(VSS),.VDD(VDD),.Y(n1153gat),.A(n1414gat),.B(n566gat));
  NOR3 NOR3_147(.VSS(VSS),.VDD(VDD),.Y(n2292gat),.A(n2443gat),.B(n2284gat),.C(n2285gat));
  NOR2 NOR2_135(.VSS(VSS),.VDD(VDD),.Y(n1416gat),.A(n2081gat),.B(n1480gat));
  NOR2 NOR2_136(.VSS(VSS),.VDD(VDD),.Y(n1151gat),.A(n1301gat),.B(n1150gat));
  NOR3 NOR3_148(.VSS(VSS),.VDD(VDD),.Y(n2306gat),.A(n2356gat),.B(n2284gat),.C(n2285gat));
  NOR2 NOR2_137(.VSS(VSS),.VDD(VDD),.Y(n1481gat),.A(n2081gat),.B(n2011gat));
  NOR2 NOR2_138(.VSS(VSS),.VDD(VDD),.Y(n982gat),.A(n873gat),.B(n1478gat));
  NOR3 NOR3_149(.VSS(VSS),.VDD(VDD),.Y(n2357gat),.A(n2285gat),.B(n2355gat),.C(n2443gat));
  NOR2 NOR2_139(.VSS(VSS),.VDD(VDD),.Y(n1347gat),.A(n2081gat),.B(n1410gat));
  NOR2 NOR2_140(.VSS(VSS),.VDD(VDD),.Y(n877gat),.A(n875gat),.B(n876gat));
  NOR2 NOR2_141(.VSS(VSS),.VDD(VDD),.Y(n1484gat),.A(n2081gat),.B(n1528gat));
  NOR2 NOR2_142(.VSS(VSS),.VDD(VDD),.Y(n1159gat),.A(n1160gat),.B(n1084gat));
  NOR3 NOR3_150(.VSS(VSS),.VDD(VDD),.Y(n2363gat),.A(n2353gat),.B(n2356gat),.C(n2355gat));
  NOR2 NOR2_143(.VSS(VSS),.VDD(VDD),.Y(n1483gat),.A(n2081gat),.B(n1482gat));
  NOR2 NOR2_144(.VSS(VSS),.VDD(VDD),.Y(n1158gat),.A(n983gat),.B(n1157gat));
  NOR3 NOR3_151(.VSS(VSS),.VDD(VDD),.Y(n2364gat),.A(n2353gat),.B(n2284gat),.C(n2356gat));
  NOR2 NOR2_145(.VSS(VSS),.VDD(VDD),.Y(n1308gat),.A(n2081gat),.B(n1530gat));
  NOR2 NOR2_146(.VSS(VSS),.VDD(VDD),.Y(n1156gat),.A(n985gat),.B(n1307gat));
  NOR3 NOR3_152(.VSS(VSS),.VDD(VDD),.Y(n2291gat),.A(n2353gat),.B(n2355gat),.C(n2443gat));
  NOR2 NOR2_147(.VSS(VSS),.VDD(VDD),.Y(n1349gat),.A(n1479gat),.B(n2081gat));
  NOR2 NOR2_148(.VSS(VSS),.VDD(VDD),.Y(n1155gat),.A(n1085gat),.B(n1348gat));
  NOR3 NOR3_153(.VSS(VSS),.VDD(VDD),.Y(n1154gat),.A(n1598gat),.B(n2930gat),.C(n2957gat));
  NOR2 NOR2_149(.VSS(VSS),.VDD(VDD),.Y(n1703gat),.A(n1705gat),.B(n3028gat));
  NOR2 NOR2_150(.VSS(VSS),.VDD(VDD),.Y(n1608gat),.A(n1704gat),.B(n1703gat));
  NOR2 NOR2_151(.VSS(VSS),.VDD(VDD),.Y(n1411gat),.A(n1154gat),.B(n1608gat));
  NOR2 NOR2_152(.VSS(VSS),.VDD(VDD),.Y(n2223gat),.A(n2354gat),.B(n2217gat));
  NOR2 NOR2_153(.VSS(VSS),.VDD(VDD),.Y(n1438gat),.A(n1591gat),.B(n1480gat));
  NOR2 NOR2_154(.VSS(VSS),.VDD(VDD),.Y(n1625gat),.A(n3021gat),.B(n1628gat));
  NOR2 NOR2_155(.VSS(VSS),.VDD(VDD),.Y(n1626gat),.A(n1627gat),.B(n3022gat));
  NOR3 NOR3_154(.VSS(VSS),.VDD(VDD),.Y(n1831gat),.A(n1832gat),.B(n1765gat),.C(n1878gat));
  NOR2 NOR2_156(.VSS(VSS),.VDD(VDD),.Y(n1443gat),.A(n1442gat),.B(n706gat));
  NOR2 NOR2_157(.VSS(VSS),.VDD(VDD),.Y(n1325gat),.A(n1444gat),.B(n164gat));
  NOR2 NOR2_158(.VSS(VSS),.VDD(VDD),.Y(n1441gat),.A(n1437gat),.B(n1378gat));
  NOR2 NOR2_159(.VSS(VSS),.VDD(VDD),.Y(n1321gat),.A(n1442gat),.B(n837gat));
  NOR2 NOR2_160(.VSS(VSS),.VDD(VDD),.Y(n1320gat),.A(n1444gat),.B(n278gat));
  NOR2 NOR2_161(.VSS(VSS),.VDD(VDD),.Y(n1486gat),.A(n1482gat),.B(n1591gat));
  NOR2 NOR2_162(.VSS(VSS),.VDD(VDD),.Y(n1440gat),.A(n1322gat),.B(n1439gat));
  NOR2 NOR2_163(.VSS(VSS),.VDD(VDD),.Y(n1426gat),.A(n2011gat),.B(n1591gat));
  NOR2 NOR2_164(.VSS(VSS),.VDD(VDD),.Y(n1368gat),.A(n1442gat),.B(n613gat));
  NOR2 NOR2_165(.VSS(VSS),.VDD(VDD),.Y(n1258gat),.A(n274gat),.B(n1444gat));
  NOR2 NOR2_166(.VSS(VSS),.VDD(VDD),.Y(n1371gat),.A(n1370gat),.B(n1369gat));
  NOR2 NOR2_167(.VSS(VSS),.VDD(VDD),.Y(n1365gat),.A(n1479gat),.B(n1591gat));
  NOR2 NOR2_168(.VSS(VSS),.VDD(VDD),.Y(n1373gat),.A(n833gat),.B(n1442gat));
  NOR2 NOR2_169(.VSS(VSS),.VDD(VDD),.Y(n1372gat),.A(n282gat),.B(n1444gat));
  NOR2 NOR2_170(.VSS(VSS),.VDD(VDD),.Y(n1367gat),.A(n1366gat),.B(n1374gat));
  NOR2 NOR2_171(.VSS(VSS),.VDD(VDD),.Y(n2220gat),.A(n2290gat),.B(n2217gat));
  NOR2 NOR2_172(.VSS(VSS),.VDD(VDD),.Y(n1423gat),.A(n2162gat),.B(n1530gat));
  NOR2 NOR2_173(.VSS(VSS),.VDD(VDD),.Y(n1498gat),.A(n1609gat),.B(n1427gat));
  NOR2 NOR2_174(.VSS(VSS),.VDD(VDD),.Y(n1504gat),.A(n1450gat),.B(n1498gat));
  NOR2 NOR2_175(.VSS(VSS),.VDD(VDD),.Y(n1607gat),.A(n2082gat),.B(n1609gat));
  NOR2 NOR2_176(.VSS(VSS),.VDD(VDD),.Y(n1494gat),.A(n1528gat),.B(n2162gat));
  NOR2 NOR2_177(.VSS(VSS),.VDD(VDD),.Y(n1502gat),.A(n1607gat),.B(n1449gat));
  NOR2 NOR2_178(.VSS(VSS),.VDD(VDD),.Y(n1250gat),.A(n1603gat),.B(n815gat));
  NOR2 NOR2_179(.VSS(VSS),.VDD(VDD),.Y(n1103gat),.A(n956gat),.B(n1590gat));
  NOR2 NOR2_180(.VSS(VSS),.VDD(VDD),.Y(n1417gat),.A(n2162gat),.B(n1480gat));
  NOR2 NOR2_181(.VSS(VSS),.VDD(VDD),.Y(n1352gat),.A(n1248gat),.B(n1418gat));
  NOR2 NOR2_182(.VSS(VSS),.VDD(VDD),.Y(n1304gat),.A(n1590gat),.B(n1067gat));
  NOR2 NOR2_183(.VSS(VSS),.VDD(VDD),.Y(n1249gat),.A(n679gat),.B(n1603gat));
  NOR2 NOR2_184(.VSS(VSS),.VDD(VDD),.Y(n1419gat),.A(n2162gat),.B(n1479gat));
  NOR2 NOR2_185(.VSS(VSS),.VDD(VDD),.Y(n1351gat),.A(n1306gat),.B(n1353gat));
  NOR2 NOR2_186(.VSS(VSS),.VDD(VDD),.Y(n1246gat),.A(n864gat),.B(n1590gat));
  NOR2 NOR2_187(.VSS(VSS),.VDD(VDD),.Y(n1161gat),.A(n583gat),.B(n1603gat));
  NOR2 NOR2_188(.VSS(VSS),.VDD(VDD),.Y(n1422gat),.A(n2011gat),.B(n2162gat));
  NOR2 NOR2_189(.VSS(VSS),.VDD(VDD),.Y(n1303gat),.A(n1247gat),.B(n1355gat));
  NOR2 NOR2_190(.VSS(VSS),.VDD(VDD),.Y(n1291gat),.A(n1603gat),.B(n579gat));
  NOR2 NOR2_191(.VSS(VSS),.VDD(VDD),.Y(n1245gat),.A(n1590gat),.B(n860gat));
  NOR2 NOR2_192(.VSS(VSS),.VDD(VDD),.Y(n1485gat),.A(n1482gat),.B(n2162gat));
  NOR2 NOR2_193(.VSS(VSS),.VDD(VDD),.Y(n1302gat),.A(n1300gat),.B(n1487gat));
  NOR2 NOR2_194(.VSS(VSS),.VDD(VDD),.Y(n1163gat),.A(n882gat),.B(n1603gat));
  NOR2 NOR2_195(.VSS(VSS),.VDD(VDD),.Y(n1102gat),.A(n1297gat),.B(n1590gat));
  NOR2 NOR2_196(.VSS(VSS),.VDD(VDD),.Y(n1354gat),.A(n1591gat),.B(n1530gat));
  NOR2 NOR2_197(.VSS(VSS),.VDD(VDD),.Y(n1360gat),.A(n1164gat),.B(n1356gat));
  NOR2 NOR2_198(.VSS(VSS),.VDD(VDD),.Y(n1435gat),.A(n1591gat),.B(n1528gat));
  NOR2 NOR2_199(.VSS(VSS),.VDD(VDD),.Y(n1101gat),.A(n1590gat),.B(n1293gat));
  NOR2 NOR2_200(.VSS(VSS),.VDD(VDD),.Y(n996gat),.A(n1603gat),.B(n823gat));
  NOR2 NOR2_201(.VSS(VSS),.VDD(VDD),.Y(n1359gat),.A(n1436gat),.B(n1106gat));
  NOR2 NOR2_202(.VSS(VSS),.VDD(VDD),.Y(n1421gat),.A(n2162gat),.B(n2359gat));
  NOR2 NOR2_203(.VSS(VSS),.VDD(VDD),.Y(n1104gat),.A(n1079gat),.B(n1590gat));
  NOR2 NOR2_204(.VSS(VSS),.VDD(VDD),.Y(n887gat),.A(n1603gat),.B(n683gat));
  NOR2 NOR2_205(.VSS(VSS),.VDD(VDD),.Y(n1358gat),.A(n1425gat),.B(n1105gat));
  NOR2 NOR2_206(.VSS(VSS),.VDD(VDD),.Y(n1420gat),.A(n1410gat),.B(n2162gat));
  NOR2 NOR2_207(.VSS(VSS),.VDD(VDD),.Y(n1305gat),.A(n1147gat),.B(n1590gat));
  NOR2 NOR2_208(.VSS(VSS),.VDD(VDD),.Y(n1162gat),.A(n698gat),.B(n1603gat));
  NOR2 NOR2_209(.VSS(VSS),.VDD(VDD),.Y(n1357gat),.A(n1424gat),.B(n1309gat));
  NOR4 NOR4_4(.VSS(VSS),.VDD(VDD),.Y(n1428gat),.A(n2978gat),.B(n2982gat),.C(n2973gat),.D(n2977gat));
  NOR2 NOR2_210(.VSS(VSS),.VDD(VDD),.Y(n1794gat),.A(n1673gat),.B(n1719gat));
  NOR2 NOR2_211(.VSS(VSS),.VDD(VDD),.Y(n1796gat),.A(n1858gat),.B(n1635gat));
  NOR2 NOR2_212(.VSS(VSS),.VDD(VDD),.Y(n1792gat),.A(n1794gat),.B(n1796gat));
  NOR3 NOR3_155(.VSS(VSS),.VDD(VDD),.Y(n1865gat),.A(n1989gat),.B(n1918gat),.C(n1986gat));
  NOR3 NOR3_156(.VSS(VSS),.VDD(VDD),.Y(n1861gat),.A(n1866gat),.B(n2216gat),.C(n1988gat));
  NOR2 NOR2_213(.VSS(VSS),.VDD(VDD),.Y(n1793gat),.A(n1792gat),.B(n1735gat));
  NOR2 NOR2_214(.VSS(VSS),.VDD(VDD),.Y(n1406gat),.A(n1428gat),.B(n1387gat));
  NOR3 NOR3_157(.VSS(VSS),.VDD(VDD),.Y(n1780gat),.A(n1777gat),.B(n1625gat),.C(n1626gat));
  NOR2 NOR2_215(.VSS(VSS),.VDD(VDD),.Y(n2016gat),.A(n2019gat),.B(n1878gat));
  NOR2 NOR2_216(.VSS(VSS),.VDD(VDD),.Y(n2664gat),.A(n2850gat),.B(n3018gat));
  NOR3 NOR3_158(.VSS(VSS),.VDD(VDD),.Y(n1666gat),.A(n1986gat),.B(n2212gat),.C(n1991gat));
  NOR3 NOR3_159(.VSS(VSS),.VDD(VDD),.Y(n1578gat),.A(n2152gat),.B(n2351gat),.C(n1665gat));
  NOR2 NOR2_217(.VSS(VSS),.VDD(VDD),.Y(n1516gat),.A(n1551gat),.B(n1517gat));
  NOR3 NOR3_160(.VSS(VSS),.VDD(VDD),.Y(n1864gat),.A(n1858gat),.B(n1495gat),.C(n2090gat));
  NOR2 NOR2_218(.VSS(VSS),.VDD(VDD),.Y(n1565gat),.A(n1735gat),.B(n1552gat));
  NOR2 NOR2_219(.VSS(VSS),.VDD(VDD),.Y(n1921gat),.A(n1738gat),.B(n1673gat));
  NOR2 NOR2_220(.VSS(VSS),.VDD(VDD),.Y(n1798gat),.A(n1739gat),.B(n1673gat));
  NOR3 NOR3_161(.VSS(VSS),.VDD(VDD),.Y(n1920gat),.A(n1864gat),.B(n1921gat),.C(n1798gat));
  NOR2 NOR2_221(.VSS(VSS),.VDD(VDD),.Y(n1926gat),.A(n1925gat),.B(n1635gat));
  NOR2 NOR2_222(.VSS(VSS),.VDD(VDD),.Y(n1916gat),.A(n1917gat),.B(n1859gat));
  NOR2 NOR2_223(.VSS(VSS),.VDD(VDD),.Y(n1994gat),.A(n1719gat),.B(n1922gat));
  NOR2 NOR2_224(.VSS(VSS),.VDD(VDD),.Y(n1924gat),.A(n1743gat),.B(n1923gat));
  NOR4 NOR4_5(.VSS(VSS),.VDD(VDD),.Y(n2078gat),.A(n1926gat),.B(n1916gat),.C(n1994gat),.D(n1924gat));
  NOR2 NOR2_225(.VSS(VSS),.VDD(VDD),.Y(n1690gat),.A(n1700gat),.B(n1702gat));
  NOR3 NOR3_162(.VSS(VSS),.VDD(VDD),.Y(n1660gat),.A(n1918gat),.B(n1986gat),.C(n2212gat));
  NOR3 NOR3_163(.VSS(VSS),.VDD(VDD),.Y(n1576gat),.A(n2351gat),.B(n1988gat),.C(n1661gat));
  NOR2 NOR2_226(.VSS(VSS),.VDD(VDD),.Y(n1733gat),.A(n1673gat),.B(n1572gat));
  NOR3 NOR3_164(.VSS(VSS),.VDD(VDD),.Y(n1582gat),.A(n2283gat),.B(n1991gat),.C(n2212gat));
  NOR3 NOR3_165(.VSS(VSS),.VDD(VDD),.Y(n1577gat),.A(n1520gat),.B(n2351gat),.C(n1988gat));
  NOR2 NOR2_227(.VSS(VSS),.VDD(VDD),.Y(n1581gat),.A(n1858gat),.B(n1580gat));
  NOR3 NOR3_166(.VSS(VSS),.VDD(VDD),.Y(n2129gat),.A(n2189gat),.B(n2134gat),.C(n2261gat));
  NOR4 NOR4_6(.VSS(VSS),.VDD(VDD),.Y(n2079gat),.A(n2078gat),.B(n2178gat),.C(n1990gat),.D(n2128gat));
  NOR4 NOR4_7(.VSS(VSS),.VDD(VDD),.Y(n1695gat),.A(n1609gat),.B(n1778gat),.C(n1704gat),.D(n1703gat));
  NOR3 NOR3_167(.VSS(VSS),.VDD(VDD),.Y(n2073gat),.A(n2078gat),.B(n1990gat),.C(n2181gat));
  NOR2 NOR2_228(.VSS(VSS),.VDD(VDD),.Y(n1696gat),.A(n1707gat),.B(n1698gat));
  NOR2 NOR2_229(.VSS(VSS),.VDD(VDD),.Y(n1758gat),.A(n1311gat),.B(n1773gat));
  NOR3 NOR3_168(.VSS(VSS),.VDD(VDD),.Y(n1574gat),.A(n1719gat),.B(n1673gat),.C(n1444gat));
  NOR3 NOR3_169(.VSS(VSS),.VDD(VDD),.Y(n1573gat),.A(n1444gat),.B(n1858gat),.C(n1635gat));
  NOR2 NOR2_230(.VSS(VSS),.VDD(VDD),.Y(n1521gat),.A(n2283gat),.B(n1991gat));
  NOR2 NOR2_231(.VSS(VSS),.VDD(VDD),.Y(n1737gat),.A(n2212gat),.B(n2152gat));
  NOR3 NOR3_170(.VSS(VSS),.VDD(VDD),.Y(n1732gat),.A(n1515gat),.B(n1736gat),.C(n1658gat));
  NOR3 NOR3_171(.VSS(VSS),.VDD(VDD),.Y(n1723gat),.A(n1659gat),.B(n1722gat),.C(n1724gat));
  NOR2 NOR2_232(.VSS(VSS),.VDD(VDD),.Y(n1663gat),.A(n1986gat),.B(n1918gat));
  NOR3 NOR3_172(.VSS(VSS),.VDD(VDD),.Y(n1655gat),.A(n1736gat),.B(n1662gat),.C(n1658gat));
  NOR3 NOR3_173(.VSS(VSS),.VDD(VDD),.Y(n1647gat),.A(n1656gat),.B(n1659gat),.C(n1554gat));
  NOR2 NOR2_233(.VSS(VSS),.VDD(VDD),.Y(n1667gat),.A(n1991gat),.B(n1986gat));
  NOR3 NOR3_174(.VSS(VSS),.VDD(VDD),.Y(n1570gat),.A(n1736gat),.B(n1658gat),.C(n1670gat));
  NOR3 NOR3_175(.VSS(VSS),.VDD(VDD),.Y(n1646gat),.A(n1569gat),.B(n1659gat),.C(n1566gat));
  NOR2 NOR2_234(.VSS(VSS),.VDD(VDD),.Y(n1575gat),.A(n1918gat),.B(n2283gat));
  NOR3 NOR3_176(.VSS(VSS),.VDD(VDD),.Y(n1728gat),.A(n1568gat),.B(n1736gat),.C(n1658gat));
  NOR3 NOR3_177(.VSS(VSS),.VDD(VDD),.Y(n1650gat),.A(n1727gat),.B(n1659gat),.C(n1640gat));
  NOR2 NOR2_235(.VSS(VSS),.VDD(VDD),.Y(n1801gat),.A(n2152gat),.B(n1989gat));
  NOR3 NOR3_178(.VSS(VSS),.VDD(VDD),.Y(n1731gat),.A(n1658gat),.B(n1515gat),.C(n1797gat));
  NOR3 NOR3_179(.VSS(VSS),.VDD(VDD),.Y(n1649gat),.A(n1560gat),.B(n1659gat),.C(n1730gat));
  NOR3 NOR3_180(.VSS(VSS),.VDD(VDD),.Y(n1571gat),.A(n1670gat),.B(n1658gat),.C(n1797gat));
  NOR3 NOR3_181(.VSS(VSS),.VDD(VDD),.Y(n1563gat),.A(n1561gat),.B(n1562gat),.C(n1659gat));
  NOR2 NOR2_236(.VSS(VSS),.VDD(VDD),.Y(n1734gat),.A(n1988gat),.B(n2212gat));
  NOR3 NOR3_182(.VSS(VSS),.VDD(VDD),.Y(n1669gat),.A(n1668gat),.B(n1742gat),.C(n1670gat));
  NOR2 NOR2_237(.VSS(VSS),.VDD(VDD),.Y(n1654gat),.A(n1671gat),.B(n1659gat));
  NOR3 NOR3_183(.VSS(VSS),.VDD(VDD),.Y(n1657gat),.A(n1662gat),.B(n1797gat),.C(n1658gat));
  NOR3 NOR3_184(.VSS(VSS),.VDD(VDD),.Y(n1653gat),.A(n1651gat),.B(n1652gat),.C(n1659gat));
  NOR3 NOR3_185(.VSS(VSS),.VDD(VDD),.Y(n1729gat),.A(n1658gat),.B(n1797gat),.C(n1568gat));
  NOR3 NOR3_186(.VSS(VSS),.VDD(VDD),.Y(n1644gat),.A(n1643gat),.B(n1648gat),.C(n1659gat));
  NOR3 NOR3_187(.VSS(VSS),.VDD(VDD),.Y(n1726gat),.A(n2992gat),.B(n2986gat),.C(n2991gat));
  NOR2 NOR2_238(.VSS(VSS),.VDD(VDD),.Y(n1929gat),.A(n1758gat),.B(n1790gat));
  NOR3 NOR3_188(.VSS(VSS),.VDD(VDD),.Y(n2009gat),.A(n2016gat),.B(n2664gat),.C(n2004gat));
  NOR3 NOR3_189(.VSS(VSS),.VDD(VDD),.Y(n1413gat),.A(n1869gat),.B(n672gat),.C(n2591gat));
  NOR2 NOR2_239(.VSS(VSS),.VDD(VDD),.Y(n1636gat),.A(n1584gat),.B(n1718gat));
  NOR2 NOR2_240(.VSS(VSS),.VDD(VDD),.Y(n1401gat),.A(n1584gat),.B(n1590gat));
  NOR3 NOR3_190(.VSS(VSS),.VDD(VDD),.Y(n1408gat),.A(n1507gat),.B(n1396gat),.C(n1393gat));
  NOR2 NOR2_241(.VSS(VSS),.VDD(VDD),.Y(n1476gat),.A(n1858gat),.B(n1590gat));
  NOR3 NOR3_191(.VSS(VSS),.VDD(VDD),.Y(n1407gat),.A(n1393gat),.B(n1409gat),.C(n1677gat));
  NOR3 NOR3_192(.VSS(VSS),.VDD(VDD),.Y(n1412gat),.A(n1411gat),.B(n1406gat),.C(n2981gat));
  NOR3 NOR3_193(.VSS(VSS),.VDD(VDD),.Y(n2663gat),.A(n2586gat),.B(n2660gat),.C(n2307gat));
  NOR2 NOR2_242(.VSS(VSS),.VDD(VDD),.Y(n2662gat),.A(n2660gat),.B(n2586gat));
  NOR2 NOR2_243(.VSS(VSS),.VDD(VDD),.Y(n2238gat),.A(n2448gat),.B(n2444gat));
  NOR3 NOR3_194(.VSS(VSS),.VDD(VDD),.Y(n87gat),.A(n743gat),.B(n17gat),.C(n293gat));
  NOR2 NOR2_244(.VSS(VSS),.VDD(VDD),.Y(n200gat),.A(n199gat),.B(n92gat));
  NOR3 NOR3_195(.VSS(VSS),.VDD(VDD),.Y(n184gat),.A(n189gat),.B(n188gat),.C(n179gat));
  NOR2 NOR2_245(.VSS(VSS),.VDD(VDD),.Y(n196gat),.A(n297gat),.B(n195gat));
  NOR2 NOR2_246(.VSS(VSS),.VDD(VDD),.Y(n204gat),.A(n200gat),.B(n196gat));
  NOR4 NOR4_8(.VSS(VSS),.VDD(VDD),.Y(n2163gat),.A(n1790gat),.B(n1310gat),.C(n2664gat),.D(n2168gat));
  NOR2 NOR2_247(.VSS(VSS),.VDD(VDD),.Y(n2258gat),.A(n2260gat),.B(n2189gat));
  NOR2 NOR2_248(.VSS(VSS),.VDD(VDD),.Y(n2255gat),.A(n2261gat),.B(n2188gat));
  NOR3 NOR3_196(.VSS(VSS),.VDD(VDD),.Y(n2015gat),.A(n2039gat),.B(n1774gat),.C(n1315gat));
  NOR2 NOR2_249(.VSS(VSS),.VDD(VDD),.Y(n2017gat),.A(n1790gat),.B(n2016gat));
  NOR2 NOR2_250(.VSS(VSS),.VDD(VDD),.Y(n2018gat),.A(n2016gat),.B(n2097gat));
  NOR4 NOR4_9(.VSS(VSS),.VDD(VDD),.Y(n2014gat),.A(n2035gat),.B(n2093gat),.C(n2018gat),.D(n2664gat));
  NOR2 NOR2_251(.VSS(VSS),.VDD(VDD),.Y(n2194gat),.A(n2187gat),.B(n1855gat));
  NOR2 NOR2_252(.VSS(VSS),.VDD(VDD),.Y(n2192gat),.A(n2184gat),.B(n1855gat));
  NOR2 NOR2_253(.VSS(VSS),.VDD(VDD),.Y(n2185gat),.A(n2261gat),.B(n2189gat));
  NOR2 NOR2_254(.VSS(VSS),.VDD(VDD),.Y(n2132gat),.A(n2133gat),.B(n2131gat));
  NOR2 NOR2_255(.VSS(VSS),.VDD(VDD),.Y(n2130gat),.A(n2134gat),.B(n2185gat));
  NOR2 NOR2_256(.VSS(VSS),.VDD(VDD),.Y(n2057gat),.A(n2049gat),.B(n1855gat));
  NOR2 NOR2_257(.VSS(VSS),.VDD(VDD),.Y(n2250gat),.A(n2248gat),.B(n2264gat));
  NOR2 NOR2_258(.VSS(VSS),.VDD(VDD),.Y(n2249gat),.A(n2265gat),.B(n3006gat));
  NOR2 NOR2_259(.VSS(VSS),.VDD(VDD),.Y(n2329gat),.A(n1855gat),.B(n3007gat));
  NOR2 NOR2_260(.VSS(VSS),.VDD(VDD),.Y(n1958gat),.A(n1963gat),.B(n1886gat));
  NOR3 NOR3_197(.VSS(VSS),.VDD(VDD),.Y(n1895gat),.A(n1845gat),.B(n1891gat),.C(n1968gat));
  NOR2 NOR2_261(.VSS(VSS),.VDD(VDD),.Y(n1710gat),.A(n1709gat),.B(n1629gat));
  NOR2 NOR2_262(.VSS(VSS),.VDD(VDD),.Y(n1630gat),.A(n1895gat),.B(n1631gat));
  NOR2 NOR2_263(.VSS(VSS),.VDD(VDD),.Y(n2195gat),.A(n2200gat),.B(n1855gat));
  NOR2 NOR2_264(.VSS(VSS),.VDD(VDD),.Y(n2556gat),.A(n1711gat),.B(n2437gat));
  NOR2 NOR2_265(.VSS(VSS),.VDD(VDD),.Y(n2539gat),.A(n2048gat),.B(n2437gat));
  NOR3 NOR3_198(.VSS(VSS),.VDD(VDD),.Y(n1894gat),.A(n1968gat),.B(n1891gat),.C(n1969gat));
  NOR2 NOR2_266(.VSS(VSS),.VDD(VDD),.Y(n1847gat),.A(n1958gat),.B(n1845gat));
  NOR2 NOR2_267(.VSS(VSS),.VDD(VDD),.Y(n1846gat),.A(n1845gat),.B(n1893gat));
  NOR2 NOR2_268(.VSS(VSS),.VDD(VDD),.Y(n2436gat),.A(n2437gat),.B(n1892gat));
  NOR2 NOR2_269(.VSS(VSS),.VDD(VDD),.Y(n2055gat),.A(n1891gat),.B(n1958gat));
  NOR2 NOR2_270(.VSS(VSS),.VDD(VDD),.Y(n1967gat),.A(n1893gat),.B(n1968gat));
  NOR2 NOR2_271(.VSS(VSS),.VDD(VDD),.Y(n2387gat),.A(n2056gat),.B(n2437gat));
  NOR2 NOR2_272(.VSS(VSS),.VDD(VDD),.Y(n1959gat),.A(n1956gat),.B(n1963gat));
  NOR2 NOR2_273(.VSS(VSS),.VDD(VDD),.Y(n1957gat),.A(n1886gat),.B(n1887gat));
  NOR2 NOR2_274(.VSS(VSS),.VDD(VDD),.Y(n2330gat),.A(n2437gat),.B(n1961gat));
  NOR2 NOR2_275(.VSS(VSS),.VDD(VDD),.Y(n2147gat),.A(n2988gat),.B(n1855gat));
  NOR2 NOR2_276(.VSS(VSS),.VDD(VDD),.Y(n2498gat),.A(n2199gat),.B(n2328gat));
  NOR2 NOR2_277(.VSS(VSS),.VDD(VDD),.Y(n2193gat),.A(n2393gat),.B(n2439gat));
  NOR2 NOR2_278(.VSS(VSS),.VDD(VDD),.Y(n2211gat),.A(n2193gat),.B(n2402gat));
  NOR2 NOR2_279(.VSS(VSS),.VDD(VDD),.Y(n2210gat),.A(n2401gat),.B(n2151gat));
  NOR2 NOR2_280(.VSS(VSS),.VDD(VDD),.Y(n2396gat),.A(n2199gat),.B(n2209gat));
  NOR2 NOR2_281(.VSS(VSS),.VDD(VDD),.Y(n2053gat),.A(n2393gat),.B(n2438gat));
  NOR2 NOR2_282(.VSS(VSS),.VDD(VDD),.Y(n1964gat),.A(n2392gat),.B(n2439gat));
  NOR2 NOR2_283(.VSS(VSS),.VDD(VDD),.Y(n2198gat),.A(n2199gat),.B(n2058gat));
  NOR3 NOR3_199(.VSS(VSS),.VDD(VDD),.Y(n2215gat),.A(n2346gat),.B(n2151gat),.C(n2402gat));
  NOR2 NOR2_284(.VSS(VSS),.VDD(VDD),.Y(n2350gat),.A(n2405gat),.B(n2349gat));
  NOR2 NOR2_285(.VSS(VSS),.VDD(VDD),.Y(n2282gat),.A(n2406gat),.B(n2215gat));
  NOR2 NOR2_286(.VSS(VSS),.VDD(VDD),.Y(n2197gat),.A(n2199gat),.B(n2281gat));
  NOR3 NOR3_200(.VSS(VSS),.VDD(VDD),.Y(n2213gat),.A(n2402gat),.B(n2151gat),.C(n2345gat));
  NOR2 NOR2_287(.VSS(VSS),.VDD(VDD),.Y(n2150gat),.A(n2401gat),.B(n2346gat));
  NOR2 NOR2_288(.VSS(VSS),.VDD(VDD),.Y(n2149gat),.A(n2193gat),.B(n2346gat));
  NOR2 NOR2_289(.VSS(VSS),.VDD(VDD),.Y(n2196gat),.A(n2199gat),.B(n2146gat));
  NOR3 NOR3_201(.VSS(VSS),.VDD(VDD),.Y(n1882gat),.A(n2124gat),.B(n2115gat),.C(n2239gat));
  NOR2 NOR2_290(.VSS(VSS),.VDD(VDD),.Y(n1962gat),.A(n1963gat),.B(n1893gat));
  NOR2 NOR2_291(.VSS(VSS),.VDD(VDD),.Y(n1896gat),.A(n2995gat),.B(n1895gat));
  NOR2 NOR2_292(.VSS(VSS),.VDD(VDD),.Y(n1972gat),.A(n1974gat),.B(n1970gat));
  NOR2 NOR2_293(.VSS(VSS),.VDD(VDD),.Y(n1971gat),.A(n1896gat),.B(n1973gat));
  NOR2 NOR2_294(.VSS(VSS),.VDD(VDD),.Y(n2559gat),.A(n2999gat),.B(n2437gat));
  NOR2 NOR2_295(.VSS(VSS),.VDD(VDD),.Y(n2331gat),.A(n2393gat),.B(n2401gat));
  NOR2 NOR2_296(.VSS(VSS),.VDD(VDD),.Y(n2352gat),.A(n3011gat),.B(n2215gat));
  NOR2 NOR2_297(.VSS(VSS),.VDD(VDD),.Y(n2566gat),.A(n2643gat),.B(n2564gat));
  NOR2 NOR2_298(.VSS(VSS),.VDD(VDD),.Y(n2565gat),.A(n2352gat),.B(n2642gat));
  NOR2 NOR2_299(.VSS(VSS),.VDD(VDD),.Y(n2637gat),.A(n3015gat),.B(n2199gat));
  NOR3 NOR3_202(.VSS(VSS),.VDD(VDD),.Y(n84gat),.A(n296gat),.B(n17gat),.C(n294gat));
  NOR2 NOR2_300(.VSS(VSS),.VDD(VDD),.Y(n89gat),.A(n88gat),.B(n2784gat));
  NOR2 NOR2_301(.VSS(VSS),.VDD(VDD),.Y(n110gat),.A(n182gat),.B(n89gat));
  NOR2 NOR2_302(.VSS(VSS),.VDD(VDD),.Y(n1074gat),.A(n2775gat),.B(n110gat));
  NOR3 NOR3_203(.VSS(VSS),.VDD(VDD),.Y(n141gat),.A(n155gat),.B(n253gat),.C(n150gat));
  NOR2 NOR2_303(.VSS(VSS),.VDD(VDD),.Y(n38gat),.A(n151gat),.B(n233gat));
  NOR2 NOR2_304(.VSS(VSS),.VDD(VDD),.Y(n37gat),.A(n151gat),.B(n154gat));
  NOR2 NOR2_305(.VSS(VSS),.VDD(VDD),.Y(n872gat),.A(n375gat),.B(n800gat));
  NOR2 NOR2_306(.VSS(VSS),.VDD(VDD),.Y(n234gat),.A(n155gat),.B(n233gat));
  NOR2 NOR2_307(.VSS(VSS),.VDD(VDD),.Y(n137gat),.A(n154gat),.B(n253gat));
  NOR2 NOR2_308(.VSS(VSS),.VDD(VDD),.Y(n378gat),.A(n375gat),.B(n235gat));
  NOR2 NOR2_309(.VSS(VSS),.VDD(VDD),.Y(n377gat),.A(n110gat),.B(n2778gat));
  NOR2 NOR2_310(.VSS(VSS),.VDD(VDD),.Y(n869gat),.A(n219gat),.B(n2792gat));
  NOR2 NOR2_311(.VSS(VSS),.VDD(VDD),.Y(n212gat),.A(n182gat),.B(n78gat));
  NOR3 NOR3_204(.VSS(VSS),.VDD(VDD),.Y(n250gat),.A(n329gat),.B(n387gat),.C(n334gat));
  NOR2 NOR2_312(.VSS(VSS),.VDD(VDD),.Y(n249gat),.A(n386gat),.B(n330gat));
  NOR2 NOR2_313(.VSS(VSS),.VDD(VDD),.Y(n248gat),.A(n330gat),.B(n1490gat));
  NOR2 NOR2_314(.VSS(VSS),.VDD(VDD),.Y(n453gat),.A(n372gat),.B(n452gat));
  NOR2 NOR2_315(.VSS(VSS),.VDD(VDD),.Y(n448gat),.A(n111gat),.B(n2846gat));
  NOR2 NOR2_316(.VSS(VSS),.VDD(VDD),.Y(n974gat),.A(n2844gat),.B(n111gat));
  NOR2 NOR2_317(.VSS(VSS),.VDD(VDD),.Y(n251gat),.A(n1490gat),.B(n387gat));
  NOR2 NOR2_318(.VSS(VSS),.VDD(VDD),.Y(n244gat),.A(n334gat),.B(n386gat));
  NOR2 NOR2_319(.VSS(VSS),.VDD(VDD),.Y(n973gat),.A(n372gat),.B(n333gat));
  NOR2 NOR2_320(.VSS(VSS),.VDD(VDD),.Y(n870gat),.A(n2669gat),.B(n219gat));
  NOR2 NOR2_321(.VSS(VSS),.VDD(VDD),.Y(n975gat),.A(n111gat),.B(n2852gat));
  NOR3 NOR3_205(.VSS(VSS),.VDD(VDD),.Y(n246gat),.A(n330gat),.B(n325gat),.C(n334gat));
  NOR2 NOR2_322(.VSS(VSS),.VDD(VDD),.Y(n245gat),.A(n386gat),.B(n334gat));
  NOR2 NOR2_323(.VSS(VSS),.VDD(VDD),.Y(n460gat),.A(n462gat),.B(n2884gat));
  NOR2 NOR2_324(.VSS(VSS),.VDD(VDD),.Y(n459gat),.A(n457gat),.B(n461gat));
  NOR2 NOR2_325(.VSS(VSS),.VDD(VDD),.Y(n972gat),.A(n372gat),.B(n458gat));
  NOR2 NOR2_326(.VSS(VSS),.VDD(VDD),.Y(n969gat),.A(n219gat),.B(n2672gat));
  NOR2 NOR2_327(.VSS(VSS),.VDD(VDD),.Y(n971gat),.A(n111gat),.B(n2840gat));
  NOR3 NOR3_206(.VSS(VSS),.VDD(VDD),.Y(n247gat),.A(n334gat),.B(n387gat),.C(n330gat));
  NOR2 NOR2_328(.VSS(VSS),.VDD(VDD),.Y(n145gat),.A(n144gat),.B(n325gat));
  NOR2 NOR2_329(.VSS(VSS),.VDD(VDD),.Y(n143gat),.A(n326gat),.B(n247gat));
  NOR2 NOR2_330(.VSS(VSS),.VDD(VDD),.Y(n970gat),.A(n372gat),.B(n878gat));
  NOR2 NOR2_331(.VSS(VSS),.VDD(VDD),.Y(n968gat),.A(n2789gat),.B(n219gat));
  NOR2 NOR2_332(.VSS(VSS),.VDD(VDD),.Y(n772gat),.A(n111gat),.B(n2842gat));
  NOR3 NOR3_207(.VSS(VSS),.VDD(VDD),.Y(n142gat),.A(n382gat),.B(n326gat),.C(n144gat));
  NOR2 NOR2_333(.VSS(VSS),.VDD(VDD),.Y(n40gat),.A(n325gat),.B(n383gat));
  NOR2 NOR2_334(.VSS(VSS),.VDD(VDD),.Y(n39gat),.A(n383gat),.B(n247gat));
  NOR2 NOR2_335(.VSS(VSS),.VDD(VDD),.Y(n451gat),.A(n134gat),.B(n372gat));
  NOR2 NOR2_336(.VSS(VSS),.VDD(VDD),.Y(n446gat),.A(n219gat),.B(n2781gat));
  NOR3 NOR3_208(.VSS(VSS),.VDD(VDD),.Y(n139gat),.A(n253gat),.B(n151gat),.C(n254gat));
  NOR2 NOR2_337(.VSS(VSS),.VDD(VDD),.Y(n136gat),.A(n253gat),.B(n154gat));
  NOR2 NOR2_338(.VSS(VSS),.VDD(VDD),.Y(n391gat),.A(n252gat),.B(n468gat));
  NOR2 NOR2_339(.VSS(VSS),.VDD(VDD),.Y(n390gat),.A(n469gat),.B(n2877gat));
  NOR2 NOR2_340(.VSS(VSS),.VDD(VDD),.Y(n1083gat),.A(n381gat),.B(n375gat));
  NOR2 NOR2_341(.VSS(VSS),.VDD(VDD),.Y(n1077gat),.A(n110gat),.B(n2672gat));
  NOR3 NOR3_209(.VSS(VSS),.VDD(VDD),.Y(n140gat),.A(n151gat),.B(n253gat),.C(n155gat));
  NOR2 NOR2_342(.VSS(VSS),.VDD(VDD),.Y(n242gat),.A(n254gat),.B(n241gat));
  NOR2 NOR2_343(.VSS(VSS),.VDD(VDD),.Y(n240gat),.A(n255gat),.B(n140gat));
  NOR2 NOR2_344(.VSS(VSS),.VDD(VDD),.Y(n871gat),.A(n802gat),.B(n375gat));
  NOR2 NOR2_345(.VSS(VSS),.VDD(VDD),.Y(n797gat),.A(n110gat),.B(n2734gat));
  NOR3 NOR3_210(.VSS(VSS),.VDD(VDD),.Y(n324gat),.A(n255gat),.B(n146gat),.C(n241gat));
  NOR2 NOR2_346(.VSS(VSS),.VDD(VDD),.Y(n238gat),.A(n147gat),.B(n254gat));
  NOR2 NOR2_347(.VSS(VSS),.VDD(VDD),.Y(n237gat),.A(n140gat),.B(n147gat));
  NOR2 NOR2_348(.VSS(VSS),.VDD(VDD),.Y(n1082gat),.A(n375gat),.B(n380gat));
  NOR2 NOR2_349(.VSS(VSS),.VDD(VDD),.Y(n796gat),.A(n2731gat),.B(n110gat));
  NOR3 NOR3_211(.VSS(VSS),.VDD(VDD),.Y(n85gat),.A(n17gat),.B(n294gat),.C(n637gat));
  NOR3 NOR3_212(.VSS(VSS),.VDD(VDD),.Y(n180gat),.A(n286gat),.B(n188gat),.C(n287gat));
  NOR2 NOR2_350(.VSS(VSS),.VDD(VDD),.Y(n68gat),.A(n85gat),.B(n180gat));
  NOR3 NOR3_213(.VSS(VSS),.VDD(VDD),.Y(n186gat),.A(n189gat),.B(n287gat),.C(n288gat));
  NOR2 NOR2_351(.VSS(VSS),.VDD(VDD),.Y(n357gat),.A(n2726gat),.B(n2860gat));
  NOR3 NOR3_214(.VSS(VSS),.VDD(VDD),.Y(n82gat),.A(n16gat),.B(n295gat),.C(n637gat));
  NOR2 NOR2_352(.VSS(VSS),.VDD(VDD),.Y(n12gat),.A(n186gat),.B(n82gat));
  NOR2 NOR2_353(.VSS(VSS),.VDD(VDD),.Y(n1599gat),.A(n1691gat),.B(n336gat));
  NOR2 NOR2_354(.VSS(VSS),.VDD(VDD),.Y(n1613gat),.A(n1544gat),.B(n1698gat));
  NOR3 NOR3_215(.VSS(VSS),.VDD(VDD),.Y(n1756gat),.A(n2512gat),.B(n1769gat),.C(n1773gat));
  NOR2 NOR2_355(.VSS(VSS),.VDD(VDD),.Y(n1586gat),.A(n1869gat),.B(n1683gat));
  NOR3 NOR3_216(.VSS(VSS),.VDD(VDD),.Y(n1755gat),.A(n1769gat),.B(n1773gat),.C(n2512gat));
  NOR3 NOR3_217(.VSS(VSS),.VDD(VDD),.Y(n2538gat),.A(n2620gat),.B(n2625gat),.C(n2488gat));
  NOR3 NOR3_218(.VSS(VSS),.VDD(VDD),.Y(n2483gat),.A(n2537gat),.B(n2482gat),.C(n2486gat));
  NOR2 NOR2_356(.VSS(VSS),.VDD(VDD),.Y(n1391gat),.A(n1513gat),.B(n2442gat));
  NOR3 NOR3_219(.VSS(VSS),.VDD(VDD),.Y(n1471gat),.A(n1334gat),.B(n1858gat),.C(n1604gat));
  NOR2 NOR2_357(.VSS(VSS),.VDD(VDD),.Y(n1469gat),.A(n1858gat),.B(n1608gat));
  NOR3 NOR3_220(.VSS(VSS),.VDD(VDD),.Y(n1472gat),.A(n1476gat),.B(n1471gat),.C(n1469gat));
  NOR2 NOR2_358(.VSS(VSS),.VDD(VDD),.Y(n1927gat),.A(n1790gat),.B(n1635gat));
  NOR2 NOR2_359(.VSS(VSS),.VDD(VDD),.Y(n1470gat),.A(n1472gat),.B(n1747gat));
  NOR3 NOR3_221(.VSS(VSS),.VDD(VDD),.Y(n1402gat),.A(n1858gat),.B(n1393gat),.C(n1604gat));
  NOR2 NOR2_360(.VSS(VSS),.VDD(VDD),.Y(n1400gat),.A(n1674gat),.B(n1403gat));
  NOR2 NOR2_361(.VSS(VSS),.VDD(VDD),.Y(n1567gat),.A(n1634gat),.B(n1735gat));
  NOR3 NOR3_222(.VSS(VSS),.VDD(VDD),.Y(n1399gat),.A(n1806gat),.B(n1338gat),.C(n1584gat));
  NOR4 NOR4_10(.VSS(VSS),.VDD(VDD),.Y(n1564gat),.A(n1584gat),.B(n1719gat),.C(n1790gat),.D(n1576gat));
  NOR2 NOR2_362(.VSS(VSS),.VDD(VDD),.Y(n1600gat),.A(n1685gat),.B(n1427gat));
  NOR3 NOR3_223(.VSS(VSS),.VDD(VDD),.Y(n1519gat),.A(n1584gat),.B(n1339gat),.C(n1600gat));
  NOR2 NOR2_363(.VSS(VSS),.VDD(VDD),.Y(n1397gat),.A(n1519gat),.B(n1401gat));
  NOR2 NOR2_364(.VSS(VSS),.VDD(VDD),.Y(n1398gat),.A(n1455gat),.B(n1397gat));
  NOR2 NOR2_365(.VSS(VSS),.VDD(VDD),.Y(n2008gat),.A(n2012gat),.B(n1774gat));
  NOR2 NOR2_366(.VSS(VSS),.VDD(VDD),.Y(n2005gat),.A(n2002gat),.B(n2857gat));
  NOR2 NOR2_367(.VSS(VSS),.VDD(VDD),.Y(n1818gat),.A(n1823gat),.B(n2005gat));
  NOR3 NOR3_224(.VSS(VSS),.VDD(VDD),.Y(n1759gat),.A(n1818gat),.B(n1935gat),.C(n2765gat));
  NOR3 NOR3_225(.VSS(VSS),.VDD(VDD),.Y(n1686gat),.A(n1774gat),.B(n1869gat),.C(n1684gat));
  NOR2 NOR2_368(.VSS(VSS),.VDD(VDD),.Y(n1533gat),.A(n1524gat),.B(n1403gat));
  NOR3 NOR3_226(.VSS(VSS),.VDD(VDD),.Y(n1863gat),.A(n1991gat),.B(n2283gat),.C(n1989gat));
  NOR3 NOR3_227(.VSS(VSS),.VDD(VDD),.Y(n1860gat),.A(n1988gat),.B(n2216gat),.C(n1862gat));
  NOR2 NOR2_369(.VSS(VSS),.VDD(VDD),.Y(n1915gat),.A(n1859gat),.B(n1919gat));
  NOR2 NOR2_370(.VSS(VSS),.VDD(VDD),.Y(n1510gat),.A(n1584gat),.B(n1460gat));
  NOR2 NOR2_371(.VSS(VSS),.VDD(VDD),.Y(n1800gat),.A(n1635gat),.B(n1919gat));
  NOR2 NOR2_372(.VSS(VSS),.VDD(VDD),.Y(n1459gat),.A(n1595gat),.B(n1454gat));
  NOR2 NOR2_373(.VSS(VSS),.VDD(VDD),.Y(n1458gat),.A(n1510gat),.B(n1459gat));
  NOR2 NOR2_374(.VSS(VSS),.VDD(VDD),.Y(n1532gat),.A(n1677gat),.B(n1458gat));
  NOR2 NOR2_375(.VSS(VSS),.VDD(VDD),.Y(n1467gat),.A(n2289gat),.B(n1468gat));
  NOR3 NOR3_228(.VSS(VSS),.VDD(VDD),.Y(n1466gat),.A(n1392gat),.B(n1461gat),.C(n1396gat));
  NOR2 NOR2_376(.VSS(VSS),.VDD(VDD),.Y(n1531gat),.A(n1507gat),.B(n1477gat));
  NOR2 NOR2_377(.VSS(VSS),.VDD(VDD),.Y(n1593gat),.A(n1551gat),.B(n1310gat));
  NOR3 NOR3_229(.VSS(VSS),.VDD(VDD),.Y(n1602gat),.A(n1594gat),.B(n1587gat),.C(n2989gat));
  NOR3 NOR3_230(.VSS(VSS),.VDD(VDD),.Y(n1761gat),.A(n2985gat),.B(n1602gat),.C(n1681gat));
  NOR3 NOR3_231(.VSS(VSS),.VDD(VDD),.Y(n1760gat),.A(n1681gat),.B(n1602gat),.C(n2985gat));
  NOR3 NOR3_232(.VSS(VSS),.VDD(VDD),.Y(n1721gat),.A(n2442gat),.B(n1690gat),.C(n1978gat));
  NOR2 NOR2_378(.VSS(VSS),.VDD(VDD),.Y(n520gat),.A(n374gat),.B(n2862gat));
  NOR2 NOR2_379(.VSS(VSS),.VDD(VDD),.Y(n519gat),.A(n2854gat),.B(n374gat));
  NOR2 NOR2_380(.VSS(VSS),.VDD(VDD),.Y(n518gat),.A(n520gat),.B(n519gat));
  NOR2 NOR2_381(.VSS(VSS),.VDD(VDD),.Y(n418gat),.A(n374gat),.B(n2723gat));
  NOR2 NOR2_382(.VSS(VSS),.VDD(VDD),.Y(n411gat),.A(n374gat),.B(n2726gat));
  NOR2 NOR2_383(.VSS(VSS),.VDD(VDD),.Y(n522gat),.A(n374gat),.B(n2859gat));
  NOR2 NOR2_384(.VSS(VSS),.VDD(VDD),.Y(n516gat),.A(n374gat),.B(n2715gat));
  NOR4 NOR4_11(.VSS(VSS),.VDD(VDD),.Y(n410gat),.A(n417gat),.B(n413gat),.C(n412gat),.D(n406gat));
  NOR2 NOR2_385(.VSS(VSS),.VDD(VDD),.Y(n354gat),.A(n411gat),.B(n522gat));
  NOR3 NOR3_233(.VSS(VSS),.VDD(VDD),.Y(n355gat),.A(n517gat),.B(n410gat),.C(n354gat));
  NOR2 NOR2_386(.VSS(VSS),.VDD(VDD),.Y(n408gat),.A(n516gat),.B(n407gat));
  NOR2 NOR2_387(.VSS(VSS),.VDD(VDD),.Y(n526gat),.A(n2859gat),.B(n740gat));
  NOR2 NOR2_388(.VSS(VSS),.VDD(VDD),.Y(n531gat),.A(n740gat),.B(n2854gat));
  NOR2 NOR2_389(.VSS(VSS),.VDD(VDD),.Y(n530gat),.A(n2862gat),.B(n740gat));
  NOR3 NOR3_234(.VSS(VSS),.VDD(VDD),.Y(n525gat),.A(n526gat),.B(n531gat),.C(n530gat));
  NOR2 NOR2_390(.VSS(VSS),.VDD(VDD),.Y(n356gat),.A(n2726gat),.B(n740gat));
  NOR2 NOR2_391(.VSS(VSS),.VDD(VDD),.Y(n415gat),.A(n2723gat),.B(n740gat));
  NOR2 NOR2_392(.VSS(VSS),.VDD(VDD),.Y(n521gat),.A(n740gat),.B(n2715gat));
  NOR3 NOR3_235(.VSS(VSS),.VDD(VDD),.Y(n532gat),.A(n527gat),.B(n416gat),.C(n528gat));
  NOR2 NOR2_393(.VSS(VSS),.VDD(VDD),.Y(n359gat),.A(n290gat),.B(n358gat));
  NOR2 NOR2_394(.VSS(VSS),.VDD(VDD),.Y(n420gat),.A(n408gat),.B(n359gat));
  NOR2 NOR2_395(.VSS(VSS),.VDD(VDD),.Y(n523gat),.A(n522gat),.B(n356gat));
  NOR2 NOR2_396(.VSS(VSS),.VDD(VDD),.Y(n634gat),.A(n418gat),.B(n521gat));
  NOR2 NOR2_397(.VSS(VSS),.VDD(VDD),.Y(n414gat),.A(n411gat),.B(n415gat));
  NOR3 NOR3_236(.VSS(VSS),.VDD(VDD),.Y(n635gat),.A(n639gat),.B(n634gat),.C(n414gat));
  NOR2 NOR2_398(.VSS(VSS),.VDD(VDD),.Y(n1100gat),.A(n1297gat),.B(n1111gat));
  NOR3 NOR3_237(.VSS(VSS),.VDD(VDD),.Y(n630gat),.A(n634gat),.B(n523gat),.C(n524gat));
  NOR2 NOR2_399(.VSS(VSS),.VDD(VDD),.Y(n994gat),.A(n1112gat),.B(n882gat));
  NOR3 NOR3_238(.VSS(VSS),.VDD(VDD),.Y(n629gat),.A(n414gat),.B(n634gat),.C(n523gat));
  NOR2 NOR2_400(.VSS(VSS),.VDD(VDD),.Y(n989gat),.A(n721gat),.B(n741gat));
  NOR3 NOR3_239(.VSS(VSS),.VDD(VDD),.Y(n632gat),.A(n414gat),.B(n523gat),.C(n633gat));
  NOR2 NOR2_401(.VSS(VSS),.VDD(VDD),.Y(n880gat),.A(n926gat),.B(n566gat));
  NOR3 NOR3_240(.VSS(VSS),.VDD(VDD),.Y(n636gat),.A(n414gat),.B(n633gat),.C(n639gat));
  NOR2 NOR2_402(.VSS(VSS),.VDD(VDD),.Y(n801gat),.A(n672gat),.B(n670gat));
  NOR2 NOR2_403(.VSS(VSS),.VDD(VDD),.Y(n879gat),.A(n2931gat),.B(n801gat));
  NOR2 NOR2_404(.VSS(VSS),.VDD(VDD),.Y(n1003gat),.A(n420gat),.B(n879gat));
  NOR2 NOR2_405(.VSS(VSS),.VDD(VDD),.Y(n1255gat),.A(n1123gat),.B(n1225gat));
  NOR2 NOR2_406(.VSS(VSS),.VDD(VDD),.Y(n1012gat),.A(n1007gat),.B(n918gat));
  NOR2 NOR2_407(.VSS(VSS),.VDD(VDD),.Y(n905gat),.A(n625gat),.B(n1006gat));
  NOR2 NOR2_408(.VSS(VSS),.VDD(VDD),.Y(n1009gat),.A(n1255gat),.B(n2943gat));
  NOR2 NOR2_409(.VSS(VSS),.VDD(VDD),.Y(n409gat),.A(n406gat),.B(n407gat));
  NOR2 NOR2_410(.VSS(VSS),.VDD(VDD),.Y(n292gat),.A(n415gat),.B(n356gat));
  NOR2 NOR2_411(.VSS(VSS),.VDD(VDD),.Y(n291gat),.A(n290gat),.B(n292gat));
  NOR2 NOR2_412(.VSS(VSS),.VDD(VDD),.Y(n419gat),.A(n409gat),.B(n291gat));
  NOR2 NOR2_413(.VSS(VSS),.VDD(VDD),.Y(n902gat),.A(n1009gat),.B(n419gat));
  NOR2 NOR2_414(.VSS(VSS),.VDD(VDD),.Y(n1099gat),.A(n1111gat),.B(n1293gat));
  NOR2 NOR2_415(.VSS(VSS),.VDD(VDD),.Y(n998gat),.A(n725gat),.B(n741gat));
  NOR2 NOR2_416(.VSS(VSS),.VDD(VDD),.Y(n995gat),.A(n823gat),.B(n1112gat));
  NOR2 NOR2_417(.VSS(VSS),.VDD(VDD),.Y(n980gat),.A(n875gat),.B(n926gat));
  NOR2 NOR2_418(.VSS(VSS),.VDD(VDD),.Y(n1001gat),.A(n420gat),.B(n1002gat));
  NOR2 NOR2_419(.VSS(VSS),.VDD(VDD),.Y(n1175gat),.A(n621gat),.B(n1006gat));
  NOR2 NOR2_420(.VSS(VSS),.VDD(VDD),.Y(n1174gat),.A(n845gat),.B(n1007gat));
  NOR2 NOR2_421(.VSS(VSS),.VDD(VDD),.Y(n1243gat),.A(n1281gat),.B(n1123gat));
  NOR2 NOR2_422(.VSS(VSS),.VDD(VDD),.Y(n1171gat),.A(n2960gat),.B(n1243gat));
  NOR2 NOR2_423(.VSS(VSS),.VDD(VDD),.Y(n999gat),.A(n419gat),.B(n1171gat));
  NOR2 NOR2_424(.VSS(VSS),.VDD(VDD),.Y(n1244gat),.A(n1123gat),.B(n1134gat));
  NOR2 NOR2_425(.VSS(VSS),.VDD(VDD),.Y(n1323gat),.A(n1007gat),.B(n401gat));
  NOR2 NOR2_426(.VSS(VSS),.VDD(VDD),.Y(n1264gat),.A(n1006gat),.B(n617gat));
  NOR2 NOR2_427(.VSS(VSS),.VDD(VDD),.Y(n1265gat),.A(n1244gat),.B(n2969gat));
  NOR2 NOR2_428(.VSS(VSS),.VDD(VDD),.Y(n892gat),.A(n419gat),.B(n1265gat));
  NOR2 NOR2_429(.VSS(VSS),.VDD(VDD),.Y(n981gat),.A(n926gat),.B(n873gat));
  NOR2 NOR2_430(.VSS(VSS),.VDD(VDD),.Y(n890gat),.A(n741gat),.B(n702gat));
  NOR2 NOR2_431(.VSS(VSS),.VDD(VDD),.Y(n889gat),.A(n1111gat),.B(n1079gat));
  NOR2 NOR2_432(.VSS(VSS),.VDD(VDD),.Y(n886gat),.A(n683gat),.B(n1112gat));
  NOR2 NOR2_433(.VSS(VSS),.VDD(VDD),.Y(n891gat),.A(n420gat),.B(n888gat));
  NOR2 NOR2_434(.VSS(VSS),.VDD(VDD),.Y(n904gat),.A(n1006gat),.B(n490gat));
  NOR2 NOR2_435(.VSS(VSS),.VDD(VDD),.Y(n903gat),.A(n1007gat),.B(n397gat));
  NOR2 NOR2_436(.VSS(VSS),.VDD(VDD),.Y(n1254gat),.A(n1123gat),.B(n1044gat));
  NOR2 NOR2_437(.VSS(VSS),.VDD(VDD),.Y(n1008gat),.A(n2942gat),.B(n1254gat));
  NOR2 NOR2_438(.VSS(VSS),.VDD(VDD),.Y(n900gat),.A(n419gat),.B(n1008gat));
  NOR2 NOR2_439(.VSS(VSS),.VDD(VDD),.Y(n1152gat),.A(n926gat),.B(n1150gat));
  NOR2 NOR2_440(.VSS(VSS),.VDD(VDD),.Y(n1092gat),.A(n1147gat),.B(n1111gat));
  NOR2 NOR2_441(.VSS(VSS),.VDD(VDD),.Y(n997gat),.A(n741gat),.B(n393gat));
  NOR2 NOR2_442(.VSS(VSS),.VDD(VDD),.Y(n993gat),.A(n1112gat),.B(n698gat));
  NOR2 NOR2_443(.VSS(VSS),.VDD(VDD),.Y(n895gat),.A(n420gat),.B(n898gat));
  NOR2 NOR2_444(.VSS(VSS),.VDD(VDD),.Y(n1094gat),.A(n1112gat),.B(n583gat));
  NOR2 NOR2_445(.VSS(VSS),.VDD(VDD),.Y(n1093gat),.A(n1111gat),.B(n864gat));
  NOR2 NOR2_446(.VSS(VSS),.VDD(VDD),.Y(n988gat),.A(n340gat),.B(n741gat));
  NOR2 NOR2_447(.VSS(VSS),.VDD(VDD),.Y(n984gat),.A(n926gat),.B(n983gat));
  NOR2 NOR2_448(.VSS(VSS),.VDD(VDD),.Y(n1178gat),.A(n420gat),.B(n1179gat));
  NOR2 NOR2_449(.VSS(VSS),.VDD(VDD),.Y(n1267gat),.A(n613gat),.B(n1006gat));
  NOR2 NOR2_450(.VSS(VSS),.VDD(VDD),.Y(n1257gat),.A(n1007gat),.B(n274gat));
  NOR2 NOR2_451(.VSS(VSS),.VDD(VDD),.Y(n1253gat),.A(n930gat),.B(n1123gat));
  NOR2 NOR2_452(.VSS(VSS),.VDD(VDD),.Y(n1266gat),.A(n2965gat),.B(n1253gat));
  NOR2 NOR2_453(.VSS(VSS),.VDD(VDD),.Y(n1116gat),.A(n419gat),.B(n1266gat));
  NOR2 NOR2_454(.VSS(VSS),.VDD(VDD),.Y(n1375gat),.A(n1006gat),.B(n706gat));
  NOR2 NOR2_455(.VSS(VSS),.VDD(VDD),.Y(n1324gat),.A(n164gat),.B(n1007gat));
  NOR2 NOR2_456(.VSS(VSS),.VDD(VDD),.Y(n1200gat),.A(n1120gat),.B(n1123gat));
  NOR2 NOR2_457(.VSS(VSS),.VDD(VDD),.Y(n1172gat),.A(n2961gat),.B(n1200gat));
  NOR2 NOR2_458(.VSS(VSS),.VDD(VDD),.Y(n899gat),.A(n419gat),.B(n1172gat));
  NOR2 NOR2_459(.VSS(VSS),.VDD(VDD),.Y(n1091gat),.A(n1111gat),.B(n956gat));
  NOR2 NOR2_460(.VSS(VSS),.VDD(VDD),.Y(n1088gat),.A(n1085gat),.B(n926gat));
  NOR2 NOR2_461(.VSS(VSS),.VDD(VDD),.Y(n992gat),.A(n815gat),.B(n1112gat));
  NOR2 NOR2_462(.VSS(VSS),.VDD(VDD),.Y(n987gat),.A(n741gat),.B(n159gat));
  NOR2 NOR2_463(.VSS(VSS),.VDD(VDD),.Y(n896gat),.A(n897gat),.B(n420gat));
  NOR2 NOR2_464(.VSS(VSS),.VDD(VDD),.Y(n1262gat),.A(n837gat),.B(n1006gat));
  NOR2 NOR2_465(.VSS(VSS),.VDD(VDD),.Y(n1260gat),.A(n1007gat),.B(n278gat));
  NOR2 NOR2_466(.VSS(VSS),.VDD(VDD),.Y(n1251gat),.A(n1123gat),.B(n1071gat));
  NOR2 NOR2_467(.VSS(VSS),.VDD(VDD),.Y(n1259gat),.A(n2967gat),.B(n1251gat));
  NOR2 NOR2_468(.VSS(VSS),.VDD(VDD),.Y(n901gat),.A(n419gat),.B(n1259gat));
  NOR2 NOR2_469(.VSS(VSS),.VDD(VDD),.Y(n1098gat),.A(n336gat),.B(n741gat));
  NOR2 NOR2_470(.VSS(VSS),.VDD(VDD),.Y(n1090gat),.A(n1111gat),.B(n860gat));
  NOR2 NOR2_471(.VSS(VSS),.VDD(VDD),.Y(n986gat),.A(n985gat),.B(n926gat));
  NOR2 NOR2_472(.VSS(VSS),.VDD(VDD),.Y(n885gat),.A(n579gat),.B(n1112gat));
  NOR2 NOR2_473(.VSS(VSS),.VDD(VDD),.Y(n893gat),.A(n894gat),.B(n420gat));
  NOR2 NOR2_474(.VSS(VSS),.VDD(VDD),.Y(n1097gat),.A(n270gat),.B(n741gat));
  NOR2 NOR2_475(.VSS(VSS),.VDD(VDD),.Y(n1089gat),.A(n1067gat),.B(n1111gat));
  NOR2 NOR2_476(.VSS(VSS),.VDD(VDD),.Y(n1087gat),.A(n926gat),.B(n1084gat));
  NOR2 NOR2_477(.VSS(VSS),.VDD(VDD),.Y(n991gat),.A(n1112gat),.B(n679gat));
  NOR2 NOR2_478(.VSS(VSS),.VDD(VDD),.Y(n1177gat),.A(n1180gat),.B(n420gat));
  NOR2 NOR2_479(.VSS(VSS),.VDD(VDD),.Y(n1212gat),.A(n1123gat),.B(n1034gat));
  NOR2 NOR2_480(.VSS(VSS),.VDD(VDD),.Y(n1326gat),.A(n1007gat),.B(n282gat));
  NOR2 NOR2_481(.VSS(VSS),.VDD(VDD),.Y(n1261gat),.A(n833gat),.B(n1006gat));
  NOR2 NOR2_482(.VSS(VSS),.VDD(VDD),.Y(n1263gat),.A(n1212gat),.B(n2968gat));
  NOR2 NOR2_483(.VSS(VSS),.VDD(VDD),.Y(n1115gat),.A(n1263gat),.B(n419gat));
  NOR2 NOR2_484(.VSS(VSS),.VDD(VDD),.Y(n977gat),.A(n670gat),.B(n671gat));
  NOR3 NOR3_241(.VSS(VSS),.VDD(VDD),.Y(n631gat),.A(n523gat),.B(n633gat),.C(n524gat));
  NOR2 NOR2_485(.VSS(VSS),.VDD(VDD),.Y(n1096gat),.A(n819gat),.B(n1112gat));
  NOR2 NOR2_486(.VSS(VSS),.VDD(VDD),.Y(n1095gat),.A(n1240gat),.B(n1111gat));
  NOR2 NOR2_487(.VSS(VSS),.VDD(VDD),.Y(n990gat),.A(n841gat),.B(n741gat));
  NOR2 NOR2_488(.VSS(VSS),.VDD(VDD),.Y(n979gat),.A(n1601gat),.B(n926gat));
  NOR2 NOR2_489(.VSS(VSS),.VDD(VDD),.Y(n978gat),.A(n2944gat),.B(n2945gat));
  NOR2 NOR2_490(.VSS(VSS),.VDD(VDD),.Y(n1004gat),.A(n978gat),.B(n420gat));
  NOR2 NOR2_491(.VSS(VSS),.VDD(VDD),.Y(n1199gat),.A(n1123gat),.B(n1284gat));
  NOR2 NOR2_492(.VSS(VSS),.VDD(VDD),.Y(n1176gat),.A(n829gat),.B(n1006gat));
  NOR2 NOR2_493(.VSS(VSS),.VDD(VDD),.Y(n1173gat),.A(n1007gat),.B(n1025gat));
  NOR2 NOR2_494(.VSS(VSS),.VDD(VDD),.Y(n1252gat),.A(n1199gat),.B(n2962gat));
  NOR2 NOR2_495(.VSS(VSS),.VDD(VDD),.Y(n1000gat),.A(n419gat),.B(n1252gat));
  NOR2 NOR2_496(.VSS(VSS),.VDD(VDD),.Y(n1029gat),.A(n978gat),.B(n455gat));
  NOR2 NOR2_497(.VSS(VSS),.VDD(VDD),.Y(n1028gat),.A(n455gat),.B(n879gat));
  NOR2 NOR2_498(.VSS(VSS),.VDD(VDD),.Y(n1031gat),.A(n1002gat),.B(n455gat));
  NOR2 NOR2_499(.VSS(VSS),.VDD(VDD),.Y(n1030gat),.A(n455gat),.B(n888gat));
  NOR2 NOR2_500(.VSS(VSS),.VDD(VDD),.Y(n1011gat),.A(n455gat),.B(n898gat));
  NOR2 NOR2_501(.VSS(VSS),.VDD(VDD),.Y(n1181gat),.A(n455gat),.B(n1179gat));
  NOR2 NOR2_502(.VSS(VSS),.VDD(VDD),.Y(n1010gat),.A(n897gat),.B(n455gat));
  NOR2 NOR2_503(.VSS(VSS),.VDD(VDD),.Y(n1005gat),.A(n894gat),.B(n455gat));
  NOR2 NOR2_504(.VSS(VSS),.VDD(VDD),.Y(n1182gat),.A(n1180gat),.B(n455gat));
  NOR2 NOR2_505(.VSS(VSS),.VDD(VDD),.Y(n1757gat),.A(n1773gat),.B(n1769gat));
  NOR2 NOR2_506(.VSS(VSS),.VDD(VDD),.Y(n1745gat),.A(n1869gat),.B(n1757gat));
  NOR2 NOR2_507(.VSS(VSS),.VDD(VDD),.Y(n73gat),.A(n67gat),.B(n2784gat));
  NOR2 NOR2_508(.VSS(VSS),.VDD(VDD),.Y(n70gat),.A(n71gat),.B(n2720gat));
  NOR2 NOR2_509(.VSS(VSS),.VDD(VDD),.Y(n77gat),.A(n76gat),.B(n2784gat));
  NOR2 NOR2_510(.VSS(VSS),.VDD(VDD),.Y(n13gat),.A(n2720gat),.B(n14gat));

endmodule