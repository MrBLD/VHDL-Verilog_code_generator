module s3858(g20763,g17845,g31861,g8215,g34237,g6752,g24184,g33079,g16686,g16659,g12470,g25583,g9680,g17678,g8416,g10527,g18099,g9743,g114,g13272,g14518,g34915,g25219,g5,g16722,g16748,g33947,g14147,g9555,g24166,g13259,g29215,g8915,g25259,g134,g24167,g92,g8719,g36,g17688,g17580,g17739,g34927,g21270,g29221,g14189,g34437,g12184,g11388,g18100,g126,g33894,g25589,g24185,g8839,g16718,g24164,g6745,g14779,g26876,g8353,g9251,g33959,g8475,g13906,g17646,g13895,g32975,g24180,g34925,g33935,g8785,g24179,g7243,g13085,g24163,g12833,g8918,g21727,g14451,g28041,g34921,g34383,g13039,g6751,g20899,g35,g34233,g17577,g12300,g34923,g16955,g20654,g34425,g14828,g24173,g29210,g8291,g34956,g56,g34919,g28753,g116,g9617,g54,g33948,g14217,g100,g7946,g14421,g20652,g8786,g33636,g13865,g18092,g28042,g16603,g17674,g6747,g10306,g12923,g14705,g84,g23683,g24177,g17778,g24169,g9048,g44,g14635,g90,g12422,g9741,g32429,g13881,g12350,g24181,g24168,g10500,g11770,g8919,g31793,g24162,g33950,g7257,g9817,g11678,g31863,g124,g18098,g30327,g34917,g24178,g17711,g19334,g18096,g25588,g24171,g18097,g16775,g17607,g29213,g25586,g17400,g11447,g31521,g23612,g57,g33533,g26875,g13068,g17649,g34240,g28030,g24165,g29214,g16874,g32454,g8870,g17722,g25582,g9553,g30332,g29212,g13966,g17316,g31656,g34221,g18101,g8920,VDD,g135,g34234,g21292,g34235,g6749,g25114,g33659,g8403,g24170,g7260,g21176,g7245,g24161,g24175,g29220,g12368,g13926,g14662,g10122,g120,g7540,g23002,g16624,g6750,g11349,g8916,g127,g24172,g17291,g25590,g34788,g16744,g8789,g11418,g17639,g17423,g18094,g30329,g8344,g34201,g34232,g21245,g14096,g8277,g17787,g14167,g8787,g12919,g6746,g17871,g14201,g23190,g26801,g8235,g16656,g30331,g113,g34435,g72,g73,g8788,g34972,g18095,g23759,g8279,g8358,g12238,g33435,g8784,g25587,g29219,g33945,g16924,g17760,g6753,g32185,g31860,g34839,g16627,g24183,g125,g20049,g7916,g17819,g29211,g8342,g9497,g34913,g24174,g6744,g33949,g8132,g99,g24182,g13049,g17743,g14597,g14738,g34239,g26877,g34436,g17764,g9682,g21698,g8783,g14125,g25585,g8283,g115,g17320,g29218,g17715,g33874,g23652,g17404,g19357,g17813,g8398,g17604,g64,g24151,g25167,g27831,g16693,g34238,g29216,g13099,g33946,g8917,g91,g20901,g8178,g9615,g14694,g30330,g29217,g17519,g31862,g34597,g24176,g18881,g20557,VSS,g25584,g6748,g12832,g14673,g14749,g9019,CLOCK,g17685,g31665,g34236,g53);
input g57,g6751,g115,g127,g35,g44,g6752,g90,g6753,g64,g126,g56,g72,g116,g91,g54,g125,g114,g6745,VDD,g5,g100,g135,g124,g6749,g6744,g6746,g6747,g99,VSS,g134,g6748,g113,g84,CLOCK,g92,g36,g120,g73,g53,g6750;
output g20763,g31521,g23612,g17845,g33533,g26875,g8215,g31861,g13068,g17649,g34237,g34240,g24184,g33079,g16686,g28030,g16659,g24165,g29214,g25583,g16874,g32454,g8870,g9680,g17722,g17678,g25582,g9553,g8416,g10527,g18099,g29212,g30332,g9743,g13966,g17316,g31656,g34221,g13272,g14518,g18101,g8920,g25219,g34915,g16722,g16748,g34234,g21292,g34235,g25114,g33947,g33659,g8403,g14147,g24170,g7260,g9555,g21176,g24166,g13259,g29215,g8915,g7245,g25259,g24161,g24167,g24175,g29220,g12368,g13926,g8719,g14662,g10122,g7540,g17688,g23002,g16624,g11349,g17580,g17739,g8916,g24172,g17291,g25590,g34788,g34927,g21270,g16744,g29221,g8789,g11418,g14189,g17639,g34437,g17423,g12184,g11388,g18100,g18094,g30329,g8344,g33894,g25589,g34201,g34232,g21245,g8839,g24185,g16718,g24164,g14096,g14779,g26876,g8277,g8353,g9251,g33959,g8475,g13906,g17787,g14167,g17646,g13895,g8787,g12919,g32975,g24180,g17871,g34925,g33935,g8785,g14201,g23190,g26801,g8235,g16656,g7243,g13085,g24179,g24163,g30331,g12833,g34435,g8918,g21727,g14451,g8788,g28041,g18095,g23759,g8279,g34383,g34921,g8358,g12238,g13039,g34972,g20899,g33435,g8784,g25587,g29219,g34233,g33945,g17577,g12300,g16924,g34923,g16955,g17760,g20654,g32185,g34425,g14828,g24173,g29210,g8291,g31860,g34956,g34839,g16627,g28753,g34919,g24183,g9617,g20049,g33948,g7916,g14217,g17819,g29211,g8342,g9497,g34913,g24174,g7946,g14421,g20652,g8786,g33636,g13865,g18092,g28042,g16603,g8132,g17674,g33949,g24182,g10306,g13049,g17743,g12923,g14705,g14597,g14738,g34239,g26877,g34436,g34236,g17764,g23683,g9682,g24177,g17778,g21698,g8783,g14125,g9048,g8283,g25585,g17320,g29218,g24169,g17715,g14635,g33874,g23652,g12422,g17404,g17813,g8398,g9741,g17604,g19357,g24151,g25167,g16693,g27831,g32429,g29216,g13881,g12350,g13099,g33946,g24181,g8917,g10500,g24168,g11770,g8919,g20901,g8178,g31793,g24162,g9615,g14694,g25586,g30330,g7257,g9817,g33950,g11678,g31863,g18098,g30327,g29217,g17519,g34917,g31862,g34597,g24178,g17711,g18881,g19334,g24176,g20557,g25584,g12832,g14673,g14749,g25588,g18097,g9019,g16775,g17607,g29213,g24171,g17685,g34238,g31665,g12470,g18096,g17400,g11447;

  wire g14407,g10200,g9070,g3333,g32541,g26388,g7535,g27306,I20412,g12950,g13910,g3462,g7153,g17693,I15263,g5637,g28343,g8002,I16969,g30003,I17114,g8812,g27416,g22176,g24112,g6462,g13393,g23884,g31930,g24843,g7593,g29852,g28295,g19479,g16164,g14807,g33263,g25876,g24631,g22519,g9177,g4392,I18307,g33449,g2652,g21187,g28585,g34657,g8139,g18325,g9935,g29865,g10390,I31171,g30921,I21258,g15162,g6704,g26784,g33279,g22078,g18394,I18813,g29792,g31252,g31185,g14753,g8792,g7632,I12927,g30102,g21381,I12270,g34276,g17575,g1992,g25087,g27720,g28885,g21988,g17503,g32808,g25148,g22018,g9958,g23984,g19677,g6997,g34938,g22051,g24802,g30092,g26713,g12361,g25848,g30457,g16489,g18826,g20269,I20910,g27371,g14537,g21765,g28374,g14255,g34292,g28602,g1576,g34371,g32507,g13266,g10044,I28349,g13486,g23505,g33791,g12399,g9792,I13744,g11753,g8851,g31969,g30097,I11701,g29008,g23415,g23129,g24892,g23408,g32356,g23985,I14257,g25647,g24748,g32304,g24571,g29736,g23374,g29270,g17189,g21990,g11323,g34029,g18417,g29512,g31069,g25721,g2514,g13221,g11389,I12631,I18205,I30971,g15707,g16162,g31658,g17152,g21823,g27041,g18127,I14630,g25654,I21234,g14838,g32190,g34987,g18751,g18498,g34159,g21163,g33017,g13156,g32321,g10709,g28340,g27528,g27045,g16629,g25577,g25119,I33103,g3219,I16512,g31478,g20182,g31834,g10081,g23905,g29344,g10199,g26268,g9747,I15287,g17419,g11183,g23291,g28158,g14386,g32072,g20036,g32864,g15063,g33858,g20552,g32301,g29857,g9752,g18223,g8201,g33560,g22154,I18568,I32161,g18438,g25180,g6073,g29150,g7513,g8239,g27350,g17706,g17145,g3805,g27149,g28369,I16855,I16695,g14625,g24347,g21709,g4258,g26851,I20165,g16729,g29310,g18170,g29982,g25660,g11917,g28493,g4966,g24098,g34806,g19768,g17365,g33295,g29077,g25322,I12314,g34940,g13912,g33238,g16826,g24406,g24916,g18659,g16674,I31222,g17586,g28163,g12589,g24353,g4801,g10571,I26676,g23857,g13963,g32714,I24674,g9848,g13574,g17183,g19376,g24635,I18398,g25209,g5052,g34134,g31855,g32316,g28482,g21189,g21800,g6837,g9269,g19962,g12651,g32153,g34790,g33551,g32352,g2970,g23478,g34749,g32674,I16821,g23458,g11224,I32613,I18897,g18284,g12523,g23655,g8889,g28321,g32702,g9892,g26900,g20556,g12259,g29793,g33460,g182,g13334,I18280,g11107,g26548,g34014,g27881,g14233,g11046,I12618,g12113,g19480,I22965,g5413,g9499,I14957,g10418,g34786,g19852,g21792,g24679,g22157,g33344,g24058,g28306,g33837,g15483,g28228,g31239,g25618,g29892,g29641,g34819,I18364,g21779,I29285,g19578,g8154,g17290,g26960,g25689,g18883,I32794,g30008,g33499,g25189,g17429,g28538,g21940,g18735,g33583,g7964,I15987,g17531,g10086,I32449,g19394,g19488,g18287,g18706,g30594,g19714,g13761,g2547,g30598,g20027,g18506,g28568,g21845,g13933,g26670,g16764,g12029,g10416,I14033,g25553,g18134,g2927,g25968,g12159,g28113,g8795,I15080,g5037,g23079,g15613,g33721,g22306,g13336,g33080,g19516,g32736,g29615,g11194,g33141,g8515,g18310,g6177,g32565,g33553,I31751,g17513,g30227,g8301,g30190,g28552,g29572,g29740,g31324,g33638,I32195,g13853,g22936,g10323,g27334,g32830,g33382,I26925,g31211,g4492,g20587,g5148,g31646,g7779,g6653,I22353,g11735,g8373,I12577,g22038,g6601,g23938,I26072,I22267,g24649,I12061,g24237,g32601,g17748,g28643,I23119,g18347,g6027,g28734,g6466,g30731,g23543,g30056,g7567,g13024,g29955,I14370,g30735,g17432,I14365,g29184,I23384,g812,g14000,g24685,g34287,g26840,g27650,g10337,g32536,g28048,g27390,g13287,g29519,g13251,g14188,I20819,I22622,g34141,g27435,g17467,g27562,g30609,g17752,g24637,g10366,I32391,g22531,I22380,g16731,g16047,I23372,g33291,g17389,g7985,g24981,g2864,g7196,g33401,g22122,g21182,g12971,g28267,g33071,g33725,g29195,g18658,g11127,g34261,g4242,g28718,g25356,g20522,g19611,g2675,g31839,g23982,g17756,g15110,g16795,g8808,g29486,g25953,g34492,g30730,I14475,g22522,g51,g28648,g24572,g12118,g3085,g19800,g2208,g13027,g23900,g21895,I24709,g34593,g11771,g33896,g17723,g25481,g32055,g24547,g27328,g34516,g14706,g27591,g18391,g32942,g2283,g25530,g15860,g34850,g12204,g8087,g34859,g12074,g17781,g12639,g20057,g33846,g34037,I32690,g10998,g33243,g33660,g28126,g18797,g26398,g33786,g18633,g28562,g32497,g14871,g10883,g21773,g5467,g17093,g25628,g2246,g13846,g28711,g31209,g28860,g20202,g24115,g33456,g20096,g7259,g28624,g25627,g29045,g28353,g1399,g24657,I32617,g31150,g31933,g26733,I12779,g21139,g30361,g34949,g4950,g9771,g3937,I26451,g4785,g10022,g19878,g33121,I31022,g25570,g17193,I22760,g15969,g28942,g20597,g34863,g23789,g24900,g28703,g8691,g30251,I21815,g34646,g28994,g29893,I12545,g13664,g28201,I26936,g14697,I31500,g12953,g26847,g10030,g21886,g34395,g21066,g16853,g15877,g12790,g11032,g24285,I13694,g32018,g25971,g10569,g12904,g11468,g33955,g32118,g27372,g31309,g10655,g31943,g33103,g23066,I25327,g3594,g34478,g12839,g14336,g34984,g24662,g14221,I18633,g9214,g33518,g22173,g23198,g28293,g14813,g31874,g30276,g18595,g30510,g13378,g24952,I32204,g31888,g30437,g31254,g10318,g34352,g11430,g27577,g17618,g7939,I17405,g34535,I23396,g22864,g28444,I29981,g28443,g16777,g10794,g14582,g18933,g24626,g16259,g19353,g25033,g20767,g3578,g15857,g22071,g24088,g24224,g2491,g6990,g20569,g32898,g26093,I32675,g33750,g11977,I25750,g3869,g19903,g14833,g24131,g7845,g33677,g31884,g28414,g21995,g14445,g15861,g5929,g19857,I30468,g19656,g18349,g21791,g13242,g3512,g8280,g14145,I31221,g34683,I15705,I32173,g15829,g23210,g28053,g24464,g30339,g23386,g6715,g23571,g24560,g34703,g27044,g11414,g28965,g18687,g32030,g34599,g34424,g5990,I28838,I18536,g29716,g34926,g15652,g31968,g32016,g30315,g16239,g32918,g23263,g20072,g13941,I22286,g22108,I15831,g27670,g25340,g24303,I17476,g16626,g11372,g14190,g18115,g14218,g13737,g19801,g9653,g23656,g33623,g32410,g4552,g26393,g11419,g20553,I14532,g19652,g8238,g2890,g17811,g246,g21361,I14932,g18830,g32706,g11192,g21398,g33606,g26634,g27336,g29627,g11024,g29954,g23300,g6500,g7344,g34999,g4229,g33637,g14816,I32929,g14768,g18526,g25782,g9828,g22128,I21181,g18501,g21769,g31503,g11234,g18648,g12864,g9602,g25105,g23483,g32849,g21831,I31286,g33104,g34099,g10756,g23544,g17092,I31306,g12882,g34203,g32753,g4515,g6593,g17301,g5587,g11991,g27063,g8362,I12709,I16231,g23639,g5527,g22407,I18758,g15135,g13070,g13976,g11249,g30518,g8106,I26972,g20595,g20386,g25894,g24758,g9280,g4449,g59,I21019,I27738,g30088,I14187,g19333,g31985,I12046,g10925,g21143,g32271,g14121,g29752,g15655,g34427,g24730,g16430,g24774,g11411,g29297,g24701,g3207,I18560,g9072,g6415,g19689,g22497,g33475,g29278,g5813,g15138,g28150,g16163,g17757,g14936,g33778,g26814,g20247,g9831,g18478,g7340,g12571,g1779,g15841,g18359,g26230,g32710,g28339,g18800,I32956,I14955,g586,g19554,g14912,I32752,g18192,g8492,g14793,I31181,g25337,g11360,g5401,I29139,g32631,g33821,g31949,g15843,g28359,g27329,g33911,g23802,g10206,g7615,g23487,I31092,g30030,g32742,g15024,g28592,g21410,I32433,g2685,g22024,I31539,g29164,I18634,g31513,g34856,g21358,g3949,g23204,g27215,g23880,g27254,g8195,I29351,g30205,g16515,g16869,g14993,g33484,g13097,g13545,g28285,g15715,I18131,g12887,g29601,g24925,g8240,g24047,g20585,g30673,g6992,g28596,g15743,g34054,g10732,g6849,g12344,g23531,g34733,g4854,g13241,I32461,g31147,g31302,g1070,g33021,g5377,g9689,g5644,g6982,I14992,g24713,g17686,I11879,g13189,g30203,g34929,g34742,g23076,g28494,g12027,g13306,g5406,I23755,g12151,g23499,g24967,g18166,g10799,g16696,g26809,g7617,g25556,g28086,g24439,g14088,g12189,g32838,I25380,g20109,g6069,g17762,g29527,g24980,g11924,g34655,I21483,g18237,I14046,g5069,g30263,g29273,g19780,g5953,I13335,g31784,g34064,g10272,g25446,g34081,g33510,g13173,I31006,I16160,g11471,g24345,g34463,g16136,g31623,g4907,g3119,I26440,g7522,g33733,g28722,g33270,g32666,g29521,I22718,g9258,I12217,I14690,g9852,g26931,g21894,g26330,g33419,g26890,g32148,g23462,g27627,I15295,g34654,g33394,g14222,g13345,g13176,I14006,g24101,I30644,g10504,g28755,g15838,I31187,g5817,g24252,g6128,g6887,I14939,g28484,g29782,g33479,g31810,g25681,g33364,g30080,I15542,g32010,g34277,g12861,I14705,g22144,g24215,g7092,g10274,I25514,g31275,g34336,g4456,g33812,g18992,g18179,g14343,g8977,g28700,I32991,g23193,g22009,g32426,g24085,I15650,g24308,g32166,g6215,I22958,I13847,I18411,g2051,g1996,g7717,g18387,g18318,g16967,g24453,g15653,g8583,I18529,g29725,g33865,g14431,g6209,g19752,I16289,g34167,I16755,g21603,g3263,g32332,g12429,g11986,g10736,g30563,g29330,g14987,g29484,g13782,I20650,g32145,g33004,g22983,g13772,g18305,g34440,g15082,g17181,g28149,g4871,g2815,g9212,g26920,g17178,I14905,g29943,g22409,g32345,g29593,g15164,g27409,I13751,g33915,g23472,g16261,g20527,g11929,g3171,g33434,g25272,g18990,g13797,g15782,g8734,I17780,g16602,g3719,g8010,g13491,I17140,g34928,g16519,g31815,I24075,g11709,I15633,g30269,g1740,g25973,I27543,g28417,g21359,g25777,g9501,g32045,g20200,g28650,g20149,g12866,g16845,g13289,g18698,I14896,g27439,g19742,g15127,g33469,I33246,I14884,g23503,g32173,g26844,g26157,g25702,g18245,g20236,g24023,g28111,g27430,g29206,g15054,I24616,g28258,g23847,g33356,g25637,g31828,g30026,g13623,I12991,g21817,I14816,g12080,g30007,g9989,g30732,g18566,g14146,g13518,g1585,g13528,g12317,I13057,g15852,g5046,g12884,g12218,g24160,g18427,g34113,g26146,g24430,g5703,g32999,g22759,g7405,g34982,g20193,g33044,I24787,I31686,I18734,g10664,g1211,I17456,g19400,g30240,g2575,g32579,g15008,g13223,g10136,g31143,g22518,g22991,g32349,g7592,g16539,g20554,g32737,g10085,g8228,g29808,g24146,g24707,g14120,g14220,g6741,g10120,g30110,g15056,g29731,I29961,I12530,g27098,g17572,g26571,g30532,g20582,g25271,g6336,g30512,g19697,g14078,g21432,g14914,I14346,g33506,g28241,g27654,g33330,g34461,g23975,g12752,g27930,g24506,g7051,g32131,g11245,g33013,g23870,g34933,g20739,g17324,g32909,g29109,g20568,g30379,g9158,g29640,g4308,g16644,g10490,g20167,I15937,g24021,g3179,g33839,g21884,g31877,I29936,g25214,g24417,g25552,g10805,g17139,g11990,g29876,g8290,g10488,g34445,I29986,g15633,g22058,g31638,I19238,g5767,I31276,g19531,g33566,g34019,g30202,g33804,g33585,I14054,g12921,g9755,g19568,g3925,g8858,I14773,g209,g632,g23246,g34205,g25130,g18639,I17675,g17634,g6395,g26672,I14481,I11835,g9379,g30516,g31848,I12074,g14804,g31250,g34431,g22159,g33092,g29777,I30992,g7004,I12172,g6019,g10530,g18911,g27960,g25880,g34042,g28706,g34909,I14424,g26932,g34190,g19440,g19145,g23342,g32238,g13131,g15030,g32965,g23292,g21124,I12764,g25410,g6113,g12182,g9460,g13255,g25620,g27628,g11957,g8575,g30298,g18610,I17128,g29174,g29148,g20838,g19694,g12246,g24650,g622,g6976,g34138,g24795,g28254,g32912,g21051,g17393,g30672,g24817,g14405,I18614,g32326,I13402,g33466,g15104,g22758,g27501,g32167,g13341,g22708,g11217,g19882,g33815,g21924,g34114,g12435,g28096,I19484,g8872,g18532,g8608,g16514,g30368,g29241,g12186,g22643,g18251,g23936,g15734,g31145,g9489,g25221,g21812,g29813,g12466,g15813,g8587,I20188,g7675,g12795,g15033,g32934,g15171,g20447,g13011,g33755,g18336,g9772,g32544,g18441,g32775,g26777,g14902,g16633,g26343,g18479,g4571,g10118,g20555,I29985,g21382,g392,g16963,g8951,g34961,g4575,I14455,I27401,g18555,g13511,g22865,g24099,g31492,g8957,g34462,g31270,I16688,g34944,g32085,g18723,g10165,g28626,g10793,g11958,g20720,g34295,I21029,g12478,g24962,g1311,g14947,g28676,g27601,g12834,g32470,g7519,g20681,g30270,g3385,g28532,g13330,g13983,g25011,g8681,g21956,g7018,g13000,g32636,g26873,g14251,g23393,g11972,g32861,g23244,g24478,g28512,I17606,I12218,g28565,g18335,g5152,g14708,I31167,g25672,g9311,g25166,g17468,g31904,g14785,g30325,g34490,g10472,g7209,I33235,g7157,g20550,g22982,g14513,g30418,g18777,g34076,g17497,g34199,g5821,g29382,g19710,g10520,g12907,g29985,g34482,I15824,g21395,g24051,g18204,I15176,g21890,g21656,g6283,I13044,g11215,g20073,g19364,g29746,g2012,g29115,g12219,g10893,g9995,g13898,I29965,g33008,g22513,g23008,g33923,g15072,g30259,g19273,g25020,I31983,g18583,g13948,g20713,g30072,I20982,g33536,g2066,g30167,g15153,g14510,g27997,g30136,g29758,g25213,g11470,g20708,I13079,g27008,g17510,g32331,g94,g34060,g16212,g15853,g24309,g34448,g9909,g34253,I27508,g23280,g13115,g30357,g21925,g17058,g27347,I24690,g32733,g25907,g23724,g15747,g2984,g26907,I24600,g29949,g34571,g29197,g28167,g3255,g11951,g25965,g8229,g33415,g25283,g13625,g17523,g29564,g31502,g17654,g30071,g32462,g28815,g1636,I24383,g20055,g34567,g10665,g20371,g12601,g33808,g32758,g32763,g20268,g20380,g29978,g34763,g21407,g25879,I15600,I31782,I18894,g8718,I22692,g11740,g30499,I13597,g34387,g32746,I15043,g9613,I12418,g24951,I15079,I17879,g12853,g12086,g34690,g6621,g31066,g2671,g33710,g19756,g22995,g30311,g21809,g6888,g13485,g29964,g15803,g34729,g21694,g31222,g7972,g7528,g29966,g27651,g10487,I13444,g23507,g26993,I14277,g24338,g14555,g32806,g31886,g27285,g21123,g32335,g9282,g17624,g23305,g16676,g33512,g33567,g32656,g11273,g25183,g18624,g11160,g33349,g26896,g18419,g6299,g28260,g23957,g7780,g27038,g26328,g26968,g30274,g18366,g12512,g11970,g14888,g17616,I21254,g29264,g16522,g25774,I13511,g3376,I27549,I18341,g10620,I15340,g8434,g6818,I22936,g3259,g32568,g24194,g5559,g24447,g30387,g28560,g32387,g23338,I27492,g26944,g19963,g3003,I18373,g17153,I30330,I12878,g21846,g33001,g13302,g18372,g24239,g9021,g13947,g14015,I14351,g23610,g19671,g26842,g29364,g25193,I20957,g27658,g34617,g7296,g28731,g24855,g22107,g7115,g28165,g27228,g7867,g11987,g24293,g17784,g28638,g30430,I18151,I31207,g34963,g26255,g3913,g19560,g13663,g25873,g1189,g10922,g29990,g25657,g31895,g15832,g4277,g9416,g24092,g3451,g23887,g24495,g28327,g25952,g5204,I17355,I32671,g8138,g11147,g25039,g16743,g11932,g34466,g18642,g6295,g10184,g32486,g34922,g24423,g20237,g7520,g26820,g11165,g34077,g22589,g29796,g18983,g17682,g8170,g25009,g27222,g18502,g9300,g9152,g18511,g518,g26957,g2036,g20147,g30226,g23916,I26417,g32221,g14612,I28434,I30741,g28768,g17673,g23769,g9861,g27460,g26314,I30124,I18906,g29742,g17384,I12823,g21362,g21252,g34865,g21276,g31893,g21832,g24648,g9414,I14497,I32874,g4146,g25819,g10685,g15871,g23546,I31477,g18660,g25018,g30193,g13902,g14261,g30363,g23380,g31759,g20070,g4760,g7335,g1564,g9730,g25791,g31908,g29570,g9808,g9305,g34500,g26278,g29606,g23650,g14686,g10684,g23538,g11981,g24527,g14516,g33732,g29284,I31327,g22045,g34498,g26545,g32383,g25537,g18224,I15205,g32708,g20697,g31206,g17747,g20913,g19146,g12888,g18630,g29878,g12995,g21728,I27253,g24313,g19541,g30090,g3672,g12667,g30060,g10653,I16452,g8751,I14923,g16100,g22037,g3921,g23813,g28799,I32791,g3443,g19632,g33684,I13321,g27587,g12538,I11740,g19504,g32050,g25958,g34192,g2579,g34112,g23413,g33097,g19620,g8899,g18416,g18243,I17741,g26636,g24311,g2169,g9890,g32947,g18123,I14291,I27513,g18217,g32600,g22714,g28910,g24008,g23485,g18426,I13336,g16159,g13513,g10528,g28091,g48,g7926,g28110,g25970,g3203,g20383,g1744,g34722,g8046,g18663,g8021,g20381,g8807,g14116,g34073,g21964,g24302,g12191,g32791,I21802,g11815,g29980,g14864,g25533,g25425,g25986,I25736,g12577,g27508,g20601,g16483,g10387,g23970,g34698,g33706,g14185,g10111,g33612,g9750,g1242,g33144,g17679,g15150,g16077,g20528,g23547,g31272,g32259,g27107,g29117,g28139,g31977,g16191,g27454,g19454,g23908,g9040,I17314,g28492,g29335,g862,g18065,g20717,g23401,g4495,g22182,g33991,g20785,g34513,g29685,g9013,g29246,g31779,g21756,g28399,g28657,g23816,g28566,g26892,g1454,g14921,g16630,g28305,g28919,g34756,g14614,g32878,g15912,g19950,g23894,g20498,g28313,g22077,g22084,I23318,g27456,g34080,g26937,g9902,g34836,g17417,g20551,g25748,g24972,g22688,g29151,g4608,I27941,g21155,g26128,g22898,g23748,g27095,I13850,g32789,g31266,g30364,g33334,g33090,g34343,g13114,g6803,g17773,g24609,g12840,g23278,g6545,g18729,g27230,g18367,g34023,g13523,I17852,g10106,g25215,g18258,g6974,g1249,g9511,g6373,g20008,g943,I33106,I15051,g17502,g28683,g8531,g32665,g6645,g14317,g15796,g20775,g3957,g27253,g10213,g13671,g20107,I14593,I13141,g22871,g20132,g3590,g25164,g12093,g11679,g6994,g26305,g22085,g20385,g19571,g26934,g2327,g24509,g22938,g10073,g3698,g10176,g28563,g33855,g26510,g29321,g33402,g26612,g19630,g11189,g27432,g11934,g27349,g3338,g5005,g31887,g28590,g25334,g3161,g22689,g23346,g25661,g18695,g20145,g19961,g27113,g33856,g10307,g18741,g13729,g27235,g10121,g7975,I14016,I17471,g26126,g34994,g2868,g5774,g24310,g20642,g13082,g32434,g18148,g16593,I17401,g25655,g329,g8644,I14660,I14185,g29015,g23929,g19373,g32353,g12121,I12861,g34793,g22079,g34279,g24072,g16321,g572,g21776,g10311,g32605,g24403,g29749,g20695,g2712,g8441,g13257,g23322,g27073,g34000,g12640,g24048,g28421,g27932,g26940,g31117,g16192,g16236,g24554,g194,g28032,I21189,g21788,g3057,g23882,g33459,g15141,g16580,g32977,g26271,g26793,g23574,g8155,g32157,I17125,g24083,g32870,g9049,g21405,g23306,g33488,g17758,g25563,g28483,g8092,g30373,g32408,g30066,g15902,I26460,g11142,g25083,g15632,g15695,g30580,g22520,I32782,I11753,g24316,g10365,g29234,g10042,g32677,g24982,g12558,g30552,g19527,g12980,I13979,g32958,I22180,I12890,g9523,g17792,g25994,g23690,g6109,g19763,g25575,g27564,I14537,g30300,g34100,g13872,g29276,g25961,g34249,g14654,g446,g28344,g9527,g16841,g25411,g14978,g33076,I31132,g10625,g23534,g7886,g4116,g19618,g13065,g19782,g8179,I15148,g11483,g33075,g962,g11357,g18279,g24516,I17639,g16968,g11891,I19917,g4927,g918,g4849,g18404,g22854,g32619,I18360,I28851,I31873,g26177,g2779,I20753,g34025,g23691,g11797,g4564,g30268,g29361,g34694,g31140,g19678,g34317,g34662,g30354,g23619,g2361,g16449,g20902,g29902,g7582,g13059,I14499,g23983,g19486,I16489,g31320,g32455,g34808,g28182,g11017,g34632,g30579,g21294,g14204,g30284,g32105,g8757,I15130,I12355,g21904,g11404,g10057,g24880,g24120,I14967,g23375,g18745,g13104,g24488,g24923,g32738,I30717,g7471,g24142,g20778,g34528,g32970,g32720,I22601,I27567,g33436,g20196,g31997,g2922,g25614,g33036,g21510,g23449,g7496,g23948,I33214,g30346,g24587,g21826,g28162,g34726,g34365,I32824,g7474,g29841,g26574,g4818,g13798,I19837,g28517,g30301,I18875,g32284,g28194,g19613,g18467,g32420,g25939,g33099,g19911,g8273,g10762,g19919,g3791,g32697,g16207,g12914,g24084,g7132,g14028,I17633,g34906,g20994,g23424,g32983,g33186,g20628,g22515,g9687,g5763,g30040,g16591,g10503,g27147,g32626,g18386,I26418,g34622,g5945,g31857,g24087,g23523,g23017,g33845,g33873,g34283,g1648,I12572,g27201,g13709,g27536,g16198,g21951,g12708,g424,g17247,g30210,g25599,g34320,I15306,I15333,g31950,g30257,g23050,g28037,I32517,g34635,g14165,g18878,g1395,I29204,g28580,g15140,g32040,g16179,I17104,g34206,g32625,g18611,g14691,g30345,g20063,g18411,g10553,g30400,g25200,g21918,g33543,g24728,I15448,g27516,g25605,g1379,g7854,g11279,g18331,g28550,g29110,g17929,g28491,g34264,g34878,g34204,g30265,g3941,g34770,g22133,g27153,g27434,g8567,g30256,g14337,g25501,g31902,g18982,g25188,g19522,I22931,g26269,I22754,g28056,g13246,I16471,I31786,g32611,g5373,g23373,g25424,g1955,g24992,g22937,I15089,g33498,g18472,g11172,g13098,g34595,g27120,g20593,g4732,g32655,I12930,g7627,g16760,g6279,g22213,g25983,g16183,g3752,g14382,g33149,g24017,g13564,I26368,g8609,g33315,g23586,g18750,g18483,g12112,I15004,g15608,I25243,g26703,g26652,g10087,g19427,g25560,I28832,g25568,I14650,g19683,g32886,g25573,g22325,I23399,g23502,g25803,I31868,g17491,g33597,g32698,g2338,g3689,g10099,g29928,g13277,g31375,g12526,g30063,g29106,g16249,I31581,g18813,g27013,g9601,g34634,I18504,g25883,I29207,g29208,I18620,g7170,g142,g29976,g16583,g14565,g12868,g28749,g31490,g28518,g32467,g10090,g29883,g9484,g10349,g20217,g33890,g15787,I14935,g23247,g30111,g15779,g32456,g31520,g33341,I18625,I28241,g13980,g31974,g13993,g30416,g11435,g8769,g23105,g34422,g10405,g9568,g10615,I18320,I15214,g32506,I31863,g577,g12867,g15045,I16357,g27507,g26099,g21781,g14521,g7674,g33487,g676,g34784,g18275,I31241,g22369,g34720,g28708,g31758,g16226,g2902,g29805,g30002,g26233,g17411,g19475,I31311,g21850,g12846,g21665,g23184,g32224,g7750,g21178,g33990,g23187,g18874,g21722,g23359,g14630,g24304,I22640,g13008,g31978,I18382,g21610,g1312,g34998,I11665,I21922,g29236,g1322,g28813,g13350,g31911,I23366,g30085,g18147,g15647,g22194,g3352,g6953,g7518,g15567,I32051,I14369,I25692,g21302,g10289,g28824,g23202,g14981,g18495,g32121,g9776,g21982,g34775,g18247,g6035,g12824,g16423,g50,g12546,g9966,g21460,g14176,g30914,g24433,g25751,I12000,I27504,g12022,I26448,g7511,g28207,g34160,g1484,g22047,g13211,g18280,g18587,g12416,g18424,g20079,g14519,g7765,I32243,g32905,g29573,g2084,g20326,g19263,g23551,g4207,g16619,g32567,g29229,g31963,g17809,g15742,g24103,g22070,I12013,g22338,I14505,I27558,g19573,I18716,g14168,g25207,g30466,g34179,g15122,g29768,g32035,g22223,g25300,g22126,g31291,g93,g21424,g14254,g2950,g23238,g305,g13670,g10231,g30568,g10155,g30204,g24949,g10999,g12066,g12886,g8032,g29257,g7228,g14505,g28747,g30115,g30134,g3770,g3068,g5503,g24763,g29649,g32114,g14589,g23811,g10510,g9806,g24996,I18350,g19275,g24097,I31874,g18886,I13276,g32442,g31805,g18191,g22298,g9648,g10544,g14424,g16672,g27524,g28982,g13913,g26863,g8631,g22869,g30138,g34266,g31249,g16723,g16204,g21369,g31153,g22090,g21388,g21246,g8442,g23873,g16701,g33881,g23990,g16219,g12925,g11513,g11029,g34527,g10614,g4411,I24030,g18551,g25722,g12968,g10295,g22718,g24013,g26802,g626,g21434,g3480,g9534,g9480,g13019,I31607,I15308,g26927,g30472,g34840,g32445,g8341,I31791,I14429,g32017,I33020,g34766,g18430,g20191,g4741,g16740,g21935,g18560,g24591,g28547,g2016,g24020,g25289,g6105,g25307,g20165,g30414,g27181,g21557,g34645,g6052,g23993,g16805,g32311,g27937,g24936,g13884,g23285,g14437,g18825,g8651,g1030,g30187,g30076,I32834,g33406,g18809,g18929,g29232,g34135,I27503,g8791,g30125,g12645,g34522,g12016,g781,g29900,g27976,g26575,g26484,g25977,g5160,g33554,g14610,g7766,g29605,g24238,g29520,g19984,g23615,g34739,g6439,I18518,g3187,g4543,g26894,g14334,g12351,g14296,g22842,g27276,g11510,g32228,g27136,I13066,g24392,g17653,I11793,g23760,g20144,I31321,g32675,g34476,g11790,g18748,g32863,g28511,g5787,g32575,I30641,g32108,g16855,g16182,g20324,g10061,I12903,g17148,I16713,g20606,g18705,g2759,g20515,g27990,g34641,g29226,g18604,g26750,g1116,I12463,I18370,g19593,g24312,g31519,g29348,g29228,g33648,g23389,g32027,g32032,g34423,I18842,g25856,g32495,g23997,g6617,g25070,g33298,g33493,g28669,g11780,g17408,g30142,g23569,g4200,g29755,g25174,g18373,g23962,g25044,g32836,g23394,g11772,g4483,g2873,g13656,g15581,I25680,g26148,g10887,g24332,g24678,g34950,g21256,g25788,g17190,g17328,g16486,I27481,g29609,I12402,g32043,g16875,g23171,g32216,g23447,g9904,g25374,g32925,g1974,g22225,g8873,g14316,g11676,g18713,g21250,g18116,g21857,g19434,g16600,g25608,I33255,g9883,g32466,g22687,I17425,g30520,g31787,g28583,g8236,g14157,g20323,g20275,I32843,I32452,g34848,g19208,g26897,g34328,g22011,g33383,g14490,g8364,g31768,g18409,g25097,g14271,g23860,I12411,g9843,g30479,g9900,g27963,g8921,g33558,g27018,g19207,g32896,g30982,g32367,g24517,g24890,g33392,g8538,g6398,I15846,g19698,g13870,g3355,g29202,g11255,g30501,g20670,g34566,g18549,g22682,g33871,g13494,I32815,I24759,g19472,g32571,g17226,g32543,g21052,g23281,g10273,g21873,g14591,g30496,g21933,I15569,g32034,g33011,g20700,g28954,g13778,g31799,g30514,g21711,g21816,g26616,g18906,g14844,I13990,g22016,g34174,g22537,g30448,g26250,g34624,g28075,g33829,I12493,g17755,g30322,g11213,g23614,g27096,g14908,g31528,g27708,g15566,g27722,g14223,g24263,g15735,g30341,g28104,g27346,g26306,g30159,g28571,g16578,g27410,g21984,g34242,g27039,g19478,g32547,g32124,g25662,g23418,g23234,g6474,g26158,g9488,g28395,g27635,g13033,g18499,g17763,g33131,g4939,g5124,g9729,g33789,g19139,g14443,g33323,g13742,g3235,I27429,g23391,g24744,g1171,g8669,g34666,g5759,g27796,g11012,g19693,g26085,I16596,g14701,g16776,I25562,g20588,I12729,g23444,g13047,g28187,g25064,g32973,g30171,g25099,g19384,g27355,g2541,g24658,g25574,g20078,g8912,I13140,g31913,g13632,g723,g23265,g5607,g32893,g10399,g14063,g34523,I17924,g27566,g29901,g33647,g8381,g29963,g34144,g28060,I29228,g27089,g22669,g7392,g32293,I31262,g25974,g26829,g33259,g10652,g20328,g20544,g16987,I32185,g17390,I32699,g24393,g30074,g27246,g7393,g32670,g34968,g32276,g17087,g33828,g21748,g32399,g19411,g26947,g16840,g16751,g26782,g11890,g9203,g32411,g33724,g25677,g31822,g22191,g7836,g26724,g29360,g18597,g33801,g6154,g25760,g7647,g640,I12277,g30432,g32046,g16928,g18540,g14568,g26147,g25249,g3416,g33256,g17224,g24515,g20064,g31116,g19749,g24526,g10072,I15893,g18111,g20774,g19521,g23440,g29555,I16564,g6996,g20903,I14350,g33599,g20028,g32872,g18205,g21983,g21397,g14794,g12288,g33735,g34118,g7149,g33204,g29354,g2555,g20531,g16527,g32847,g14817,g9564,g10704,g34983,g14093,g26206,g20676,g28033,I12849,I33053,g26810,I31212,I32535,g1682,g33574,g18820,g15823,g26954,g33081,g34459,g28660,g28302,g21763,g18893,g30382,g30004,g30469,g27980,g24258,g27520,g8480,I15106,g28332,g24958,g28282,g29867,g12672,g25893,g3484,g26866,g23404,g30192,g20238,g33610,g25591,g17767,g29042,g9760,g32871,g32281,g12306,I28585,g32282,g22980,g33332,g34015,I17801,g20583,g30997,g46,g11571,g25268,g28215,g24016,I14267,g25734,g16637,g1367,g1874,g29907,g14089,I20461,g26162,g17120,g16090,g32846,g32757,g7087,g24908,g12144,g30411,g28361,g28914,g24618,I31101,g969,I31066,g27247,g13030,g1890,g33340,g18736,g27211,g30280,g23876,g18563,g13346,g32155,g13134,g21941,g19657,g6873,g26859,g22310,g7563,I16626,g9672,g29033,g16868,g7222,g24749,g13975,g33897,g14868,g30537,g34953,g18805,g7840,g8037,g26390,g27025,g15780,g25429,g27988,g21975,g24582,g12419,I23684,g9829,g6692,g10795,g3802,g24654,g25110,g25502,g34117,g32019,g33483,I24365,I15300,g19609,I12219,g32835,g12863,g31255,g14347,g5752,g30990,g30392,g25688,g8632,g32263,g33454,g26651,g23958,g28509,g11402,g21892,I31252,g32798,g4567,g23902,g15372,g12543,g8778,g24226,g8476,g19699,g6291,g18776,g23764,g31253,I22589,g31771,g33474,I31600,g34058,g28050,g29979,I13077,I14761,g23893,g20904,g24619,g25514,g24022,g6801,g12018,g18592,g27493,g25184,g5208,g29259,I26710,g34660,g19904,g8124,g11144,g34544,g16303,g25388,I32150,g6900,g10804,g28732,g1706,g30604,I15556,g7715,g8790,g8133,g25613,g25638,g20009,g33058,I22823,g31811,g21556,g27241,g33082,g29948,g28130,g16222,g32995,g20495,I31316,I13762,g33877,g17482,g17176,g14262,g1536,g26718,g14545,I25244,g29509,g19577,g4912,I20433,g28907,g21868,g30470,g24861,g32393,g21385,g23152,g24583,g23998,g33378,g28618,g34418,g11968,g21996,g21848,g30144,g32269,g25712,g11237,I21250,I15299,g26277,g34693,g18650,I22930,I32775,g13831,I18333,g4176,g32534,g25924,g33910,g18109,g23988,g26754,g17284,g12849,g10822,I15474,g34404,g18686,I21033,g16622,g18786,g33683,g34,g32322,g18798,g1291,g24567,g27558,g13411,g3649,g28179,g33803,g33124,I19786,g23138,g30592,g29941,g24259,g32952,g6928,g21409,I29969,g34062,g18693,g10565,g3431,g24496,g33464,g10519,g22841,g34954,g24940,g32650,g33809,I31031,g31501,g8016,g1600,g16237,g22062,g31210,g33785,g30199,g13414,g18384,g27693,g29884,g11527,g33526,g19612,I13759,g32672,g1830,I15834,g7394,g24746,g22082,g7971,g23103,g14055,g11607,g29248,I14714,g14154,g11225,g9805,g34582,g12632,g28840,g11950,g13190,g23216,g3736,g23681,g12772,g5073,g5396,g29924,g18739,g15107,g24305,g7623,g12412,g25467,g11019,g33918,g33061,g9250,g18645,g25488,g18225,g28319,g33412,g34491,I12132,g32098,g21874,g33535,g33040,g19791,g18938,g30338,g29860,g24054,g11936,g20086,I26508,g23909,g29097,g19491,g15757,g8836,g28652,g15678,g23528,g18788,I31016,g14735,g6809,g27116,g14752,g29299,g34209,g24959,g14535,g24603,g24933,g7,g25778,g4245,g9664,g26154,g27974,g14082,g10666,g27487,g27585,g34665,g14130,g24798,I12261,g20000,g17783,g19398,g854,g24934,g33136,g24314,g16628,I25391,I21934,g14959,g3506,g27832,g19452,g2932,g11326,I18574,g32009,g32476,g18594,g27551,g20011,g20183,g11677,g32071,g16689,g13335,I16028,g27146,g21938,g23788,g29811,g20682,g26573,g33872,g16873,g25834,g15070,g17590,g22881,g30593,g9797,I31097,g26165,I31106,g18466,g6040,g8334,g5029,g24941,g22866,g33973,g23794,g25022,g29355,g16957,I26050,g29171,g24946,g15165,g15112,g24865,g11920,g30198,g10116,g30917,g3251,I15190,g26248,g30139,g28178,I15363,I28913,g26182,g26023,g3897,I17814,g31928,g16125,g18700,g29553,g33622,g23275,g5264,g29243,g20782,g10566,g33690,g32667,g25673,g19595,g24639,g22830,g16581,g12909,g29209,g28853,g772,g28420,g29638,g22979,g7387,g23590,g31276,g18752,g33063,g11841,g32651,g29532,g32624,g19865,g29004,g27283,g4273,g20559,g30096,g24050,g34075,g29839,I25541,g26334,g14714,g30920,g13416,g29591,g27102,g18578,g8440,g32154,I31107,g29956,g11038,g20185,g4153,g18569,g27972,g34018,g21707,g22536,g4704,g8859,g25545,g10363,g17742,I19756,g10656,g26380,g17315,g20921,g12978,g28707,g15595,g10408,I27552,g14758,g23609,g23083,g16258,g34536,I13634,g14971,g18593,g32402,g23293,g23388,g31240,g19764,g27249,g25007,g32487,g30238,g26888,g18256,g22833,g32865,g26633,g15795,g4253,g16534,g13124,g30589,g17487,g32524,g2537,g27305,g30350,g13857,I30962,g32306,g26286,g34947,g29797,g19070,g7139,g26377,g32232,g18613,g34438,g15744,g22384,g34150,I33173,g5698,g479,I12963,g24134,g29154,g10882,I24576,g29744,I11878,g34202,g13437,g29319,I14516,g33003,g23658,g28152,g12347,g24064,g3199,g7626,g27387,g7936,I27954,g20189,I18912,I31077,g20113,g23242,g8595,I31151,I31141,g14030,I19012,g27437,g18991,I22844,I24334,g14442,g32639,g12117,I29302,g30149,g29318,g568,g12110,g8069,g3530,g5507,g30079,g22876,g19996,I24680,g2791,g28141,g9742,g17085,g24604,I23321,g29353,g17712,g18726,g20709,g18803,g9490,g18892,I30750,I16024,g31845,g32964,g10812,I26430,g29309,g11897,g27462,g32559,g26280,g32730,g34670,g10218,g9339,I31297,g15724,g23409,g8579,g30536,g32400,g34460,g11384,I20469,g25725,g28140,g11560,g17791,g16326,g18676,g5736,g11395,g31940,g13680,g26351,g26830,g15081,I23363,I22945,g14940,g30460,g23350,g27563,g32572,g13869,g20106,g9586,g15039,g23414,g30447,g9704,g32384,g7655,g18444,I14619,I17615,g7345,g10233,g20641,g8592,g10031,g10529,g31488,g4581,g13706,g27367,g32227,g21736,g18949,g15058,g18326,g1083,g32606,I23369,g18544,g30425,g4219,g34339,g28945,g23778,g8958,g29373,g12881,g23052,g26808,I26682,g21069,I16111,g22063,g34401,g20887,g11345,g21730,g12169,g2741,g21733,g10119,g18880,g23490,g15156,g13739,g28077,g16747,g29951,g26946,g896,I12373,g34569,g34104,I31111,g12440,g21156,g5041,g19375,g8944,g24869,I26638,g13539,g681,g20266,g30024,g18778,g28227,g20664,g25685,g16533,g30194,g21455,g13516,g5583,g25990,g27766,g10043,g29146,g33073,I31291,I13240,g2223,g2151,g22114,g29987,I18006,g21973,g15102,g23192,g5547,g25870,g14572,g28330,g3343,g17619,g28357,g20636,g34614,I33056,g25768,g2145,g29085,I17658,I23099,g15078,g7003,g28479,g5252,g22179,g12228,g28098,g25197,g18504,I21994,g11480,g20065,g278,g21949,g8457,I18446,g19416,g27040,g9055,g29372,g31207,g11763,g25078,g23799,g5889,g33864,g11669,g22625,I32473,g32325,g27151,I23303,g31824,g29778,I25882,I31057,g11769,g22049,I31332,g33417,g24245,g27335,g32700,g1152,g13119,g32288,g13078,g9483,g6984,g22975,g33759,g301,g29800,g25262,I18626,g17780,I12437,g27221,g30033,g25698,g21379,g34225,g18588,g28877,g1932,g6227,g34783,g15125,g25991,g32679,g22130,g31504,g30334,g33969,g26344,g26395,g20633,g19619,g33060,g34415,g25290,g2783,g24514,g22653,g25001,g28545,g4369,g26645,g32143,g33709,g16812,g28144,g1426,g21057,g5348,g936,g10212,g12588,I14833,g28950,g13106,g3893,g32338,g255,g23314,g32250,g30560,g28093,g24935,g29898,g8591,g11383,g17125,I23980,g5232,g28656,g27360,g33552,g22098,g31508,g13540,g3034,g33128,I32305,g20026,g20007,g86,g9779,g25076,g33069,g11584,g29530,g13622,g164,g6369,I33270,g28331,g32540,g19716,g239,g33827,g23540,g9554,g9644,g33912,g15371,g32810,g32123,g21281,g10654,g20211,g25703,g33448,g22523,g20995,I13392,g16765,g8187,g9684,g20737,g18512,g12482,g11706,g25830,g11442,g32703,g19998,g33471,I20166,g16925,g15872,g28946,g33014,g29338,g30355,I13462,I31494,g18605,I11721,g21801,g13132,g21720,g15850,g32804,g14182,I17590,g14247,g33932,g15805,g8984,g18429,g12155,g29807,g22219,g22902,g32109,I33158,I26381,g34007,g3310,g28525,g14556,g23405,g17727,g1002,g25108,g3808,g18199,I15255,g33720,g25756,g31804,g16774,g30378,g15145,I22745,g29802,g11945,g29734,g20168,g18944,g31897,g33132,g33478,I24393,g12970,g6597,g34074,I15862,g18606,g23518,g21908,g27374,g8350,g23022,g15836,g30542,g34781,g847,g11966,I14610,g23729,g21282,I20204,g4332,g32198,g13315,g9804,I11824,g29502,g13431,g17675,g10578,g15111,g6444,g27265,g23649,g29082,g33264,g32068,g25473,g15344,g7289,g14547,g17271,I18066,I12159,g22101,g6267,g18446,g19783,g20875,g30108,I14192,g12972,g25058,g30234,g17512,g9537,g30610,g24508,g33046,g33557,g33564,g29929,g32885,g1270,g9777,g25541,g4983,g34538,g27020,g27876,g18142,g25349,g20586,g13250,g23445,g34930,g28252,g26396,g23890,g12234,g13498,g33995,g17694,g23937,g15704,g18754,g23183,g18810,g29069,g13728,I21115,g26942,g24484,g14192,g12019,g24036,g11425,g2449,g33027,g34980,g269,g25316,g27532,g22516,g19735,g34426,g4000,g28312,g14037,g4408,g34194,g30164,g20734,g11118,g6377,I18903,g32247,g32309,I19348,g19633,g19754,g27534,g23235,I31357,g26156,g7704,g17746,g21937,g9477,g29683,g32206,g20441,g31608,g26803,g22053,g20536,g33602,g34211,g14615,g21012,g30059,g28796,I30469,g20379,g18172,g26303,g17716,g6840,g20871,g25903,g23452,g25693,g17496,g1882,g28279,g11998,g34321,g16187,g11639,g21822,g34125,g24057,I28582,g25607,g32732,g30605,g29741,g19787,g18721,g25124,g32488,g21693,g28324,g14398,g23822,g22847,I13329,I28540,g26615,g24778,g27438,g13526,g24260,g31295,g34543,g20248,g34789,g33491,g27309,g28261,g28469,g32599,g23497,g21378,g16069,g17327,g24295,g16821,g18151,g29585,I17661,g19431,g33346,g26753,g26879,g30337,g6581,g33146,g8558,g30258,g29625,g3562,g10501,g2689,g7549,g29632,g29851,g24218,g12848,g8216,g7163,g20154,g7764,g13794,g18410,g6991,g7252,I22211,g30075,g34773,g21058,g22853,g5551,g9964,g10139,g11023,g15914,g31245,I14381,g33458,g30006,I13124,g22014,g25324,g16025,g32634,I22547,g32573,I31281,g34764,g33114,g25225,g2619,g31317,g3849,g5909,g19408,g20857,g21304,g25452,g20271,g11692,g20212,g33675,g18758,g33550,g7446,I18434,I31694,g25945,g23996,I29013,g18458,g23923,g26234,g22667,g27363,g25984,g33274,I18034,g29383,g33646,g34846,g13138,g32229,I22769,g22113,g30422,g15507,g25581,g29961,g27373,g31495,g27661,g32986,I20882,g34374,g29363,g23849,g24670,g34289,g23986,g12896,g16609,g14830,g33372,g33605,g19422,g14680,g18218,g32712,g31995,g25106,I16090,g8989,g18319,g31474,g10001,I24555,I33047,g27019,g11592,g32015,g33107,g4859,g27106,I16135,g27032,g28729,g12662,g34507,g6137,g8458,I26427,g21915,g21878,g6203,g28758,g7928,g25911,g33900,g34101,g4664,g2273,g8741,g32481,g34393,g13544,g20607,I11866,g29025,g34618,g32825,g32097,g31900,g33790,g9569,I22901,g19545,g29595,g34254,g34246,g13595,g19415,g29535,g15788,g33736,g27366,g16814,g7620,I15241,g27488,g21408,g32629,g32218,I15254,g23041,g18617,g34052,g29349,g34338,g18323,g26933,g27280,g24153,g20095,g7805,g29594,g4185,g26769,g30215,g18523,g5706,g28653,g9887,g33047,I13805,g17770,g31671,g18423,g14383,g28244,I18469,g29999,g8679,g28181,g16124,g17656,g7110,g19338,g10172,g32020,g16772,g31168,I18523,g15784,g13508,g33408,g22202,g34162,g21453,g29079,g21710,g23194,g34687,g24361,g28440,g30459,I18487,g32761,g32292,g1472,g16808,g13509,g33212,g16023,g22654,g2704,g24586,g18740,g24732,g30047,I30734,g13055,g26766,g9932,g23573,g34874,g29903,g13118,I33276,g15166,g27130,g4249,g27090,g11834,g27242,g12878,g29661,g15108,g18943,g16275,g23575,I32446,g16506,g18781,g18453,g25956,g27505,g21787,g33042,g10946,g20372,I27192,g4366,g25867,g25921,g18679,g34521,g23436,I32056,g24330,g34493,g28415,g10918,g31228,g13209,g27561,g11403,g14656,g9856,g27612,g15725,g1280,g30305,g18522,g34910,g23525,I26395,g27058,g25972,g34390,g33018,g10917,g30321,g7631,g29621,g10491,g8764,g30476,g32709,g18932,g7117,g25479,g13510,g16093,g11010,g18749,I12346,g14950,g12656,g28793,g30314,g18559,g14314,g27403,g24606,g33389,g15880,g24102,g30244,g24236,g22993,g7178,g20771,g26605,I27235,g9360,g30919,g4226,g15065,g11705,g15611,g32891,g3821,g18490,g32686,g15673,I20167,g33719,g29227,g15870,g33059,I17692,g28641,g7594,I32518,g2093,g13384,g14515,g29516,g22015,g11498,g31283,g32823,I15129,g8630,g8324,g10348,g19861,g28125,g23283,g18685,g21454,g33810,g9619,g17409,g25126,I14854,g34579,g25156,g10582,g21957,g10380,g22023,g24240,I24699,g28990,g23654,g16876,g29263,g22637,g29568,g28386,g26103,g18447,g14937,I31216,g28255,g23548,g30146,g20540,g29771,g1467,g776,g4210,g29279,g10362,g34619,g13409,g20534,g24396,g3853,g2465,g14127,g24721,g7187,g21560,g24556,g24771,g31883,g5654,g34570,g20910,g1945,g26378,g27298,g9071,g13116,g33035,g14933,g12939,g28664,g3817,g22873,g21882,g15910,g15014,g20157,g14414,g11026,g23334,g33129,g19335,g14227,g28625,g29336,g34429,g24786,g11912,g47,g23869,g15966,g7246,g24405,g13305,g11906,I15843,g11686,g33742,g22080,g21406,g16854,g32715,g17499,g4072,g28088,g2331,g23166,g17242,g14782,g24904,I17143,g11316,g21714,g32254,I27271,g11729,g12040,g17926,g24523,g6537,g11707,I18589,g10191,g22028,g31918,g29056,g32067,g26120,g20153,g34590,g34585,g6799,g25949,g28389,g18380,g2476,I26530,g5164,g4438,g34686,g16216,g16749,g31776,g6697,g5881,g10047,g18329,I23339,g25026,g16161,g31885,g32265,I11629,g7596,g20192,g9833,g33112,g30478,g12188,g21298,g20152,g31293,g31244,g27957,g31002,I33131,g14339,g17521,g27599,g30450,g25325,g16811,g25543,I26406,g31907,I15536,g34762,g12859,g15563,g32613,g32997,g25032,I25579,I13453,I23336,g27365,g30533,g31128,g6804,g26183,g9281,g29308,g11443,g29525,g19597,g28300,g12598,g23111,g22487,g32751,g16312,g31152,g5272,g7566,g27258,g34307,g31115,g20187,g25651,g25935,g27928,I22711,g26948,g27699,g18124,g31282,g24903,g6509,g22121,g32818,g19461,g17414,g34914,g30054,g24998,I24505,g14541,g18978,g30348,g8507,I16646,g23331,g33687,g29233,g31579,g15571,g17690,g23874,g19532,g29838,g23372,g18696,g27105,g23063,g15651,g11988,g25836,g27767,g10411,g28635,g20151,g33977,g26915,g16752,g33994,g26186,g26973,g22180,g34040,g29529,g9558,g22897,g32883,g23006,g32770,g19587,I20399,g32840,g19965,g24979,I18114,g33116,g26870,g27499,g27304,g13141,g10400,g20634,g24669,g1913,g20513,g11737,g22752,g28490,g10410,g18249,g33381,g14538,I17302,g3239,g12223,g26104,I18849,g24919,g13177,g22008,g30105,g16688,I32645,g29712,g30239,g19399,g3668,g26364,g32762,g13333,g28105,g29180,g18338,g21875,g16484,g32504,I15365,g18476,g18644,g25175,g9391,g12415,g18817,g7379,g11312,g21795,g26916,g18285,g14095,g24038,g24743,g4455,g24710,g15859,g17010,g33066,g32633,g21794,g18486,g18737,I24700,g23419,g33617,I18344,g32503,g21393,g30360,g14822,g29774,g6999,g8113,g26721,I24524,g10587,g14511,g22659,g29769,g25067,g29254,g11566,g17777,g30253,g13050,g11232,g33427,g32994,g33299,g2886,g34353,g20543,g9217,g10156,g29945,g25529,g27357,g34145,g31313,g32314,g14206,g6847,I13045,I23348,g29586,g22525,g29977,g8891,g3570,g22115,g32463,g19437,g27050,g24235,g11511,g30061,g29584,g20659,g31975,g18769,g16594,g18608,g16631,I19772,g10554,I12735,I29909,g7947,g28693,g7512,g20108,g24286,g33524,g29189,g14027,g26290,g13105,g18114,g26339,g33928,I13699,g9024,g16422,g24625,g9705,I27546,I22972,I23602,g25139,g34991,g23922,g24031,g32644,g26951,g30600,g20783,g10775,g12035,g2375,g8955,I32464,g34178,g9744,g18515,g33235,g355,g26254,g32029,g24624,g19736,I21978,g30065,g25535,g2860,g28148,g12356,g24333,g34333,g655,I14450,g2975,g22868,g32766,I17475,g33966,g26962,g25604,g15738,I17923,g17056,g22052,g24791,g2807,g18732,g25675,g6483,g23361,g25557,g19401,g32117,g34752,g30335,g2441,I33143,g14198,g13554,g34471,g35002,I15033,g26919,g22896,g32275,g33163,g30534,g23861,g27545,g19687,g12119,g14004,g14044,g33712,g9972,g19960,g17583,g4112,g1300,g20083,g34562,g29554,g1870,g4507,g25288,g9860,g34247,g11849,g32315,g14290,g25539,g6815,g28524,I12848,g2399,g30037,g20777,I22580,g19581,g22312,g34900,g23473,g21916,g16537,I14222,g7803,g27291,g4064,g16292,g29534,g1306,g20525,g30463,g2509,g15170,g24600,g28320,g32654,g28743,g23708,g17140,g18183,g30023,g29143,g31308,g29305,g15731,g34315,g21818,g29293,g23646,g18529,I14290,g22224,g15992,I16779,g23209,g6116,g10124,g10586,g8803,g11561,g12609,g23032,g31070,g20618,g33072,g17239,g20625,g17137,I16671,g18266,g18904,g21872,g31601,g29238,g23792,g9285,g17597,g11119,g14644,g10884,g18981,g24655,g15884,g16601,g24533,g17182,g33889,g33142,g17608,I15364,g33835,g20915,g19061,g739,g33503,I22604,g25407,g31631,g26828,g23855,I31491,g34379,g15105,g18675,g13290,g10429,g25059,g33254,g9934,I20954,g27571,g7994,I20999,g17268,g18554,g19455,g29847,g21228,g26845,g2625,g17612,I29233,g30057,g10838,g32368,g25817,g11153,g18895,g27327,g33843,I14331,g16810,g30465,g4452,I21226,I16775,g27676,g23255,g19206,g16604,I22852,g33556,g12467,g34245,I24414,g27660,g13832,g30230,g33355,g5077,g4480,g31310,g8011,g13699,g21611,g31258,g23745,I31545,g18572,g23850,g22843,I14510,g33571,g25602,g27522,I26880,g19362,g26878,g13079,I30959,g13256,g18346,I21976,g30483,g6428,g9832,g14170,g9373,g27311,g23243,g25505,g24825,g31624,g28679,g32564,g29528,g9591,I14482,g15612,g24907,g15789,g32614,g17528,g1384,g29018,I31191,I31036,I14827,g29080,I32840,g9559,g17144,g22360,g23589,g30250,g2299,g23341,g11268,g20869,g26778,g22994,g26731,g31469,g18233,I22799,g29602,I16733,g15098,g12975,I13065,g15883,g31,g18677,g27383,g33030,g6875,g22118,g12217,g6479,g20162,g6235,g18957,g16290,g13029,g29795,g33162,g18585,g13004,g25203,g28309,g24306,g26078,g25308,g27480,g11618,g28114,g19363,g9819,g25724,g18270,g11852,g25567,I14399,g31869,g29249,g29247,g32985,g20090,g33530,g13525,I14925,g32499,g23989,g23486,g26953,I20130,I11734,g26054,I22845,g2787,g25569,g18619,g29307,g18261,g17873,g31807,g10027,g31852,g33601,g23067,g13036,g32253,g33758,g18361,g25107,g25326,I31156,g34633,g24534,g33844,g26302,g7266,g28094,g17724,g30174,g2852,I33232,g22060,g25656,g11185,g9245,g30010,g13323,g27734,g32052,g4681,I27742,I31616,g33722,I14563,g20198,I21486,g27015,g8745,g16867,g26685,I17883,g27677,g24821,g12333,g32933,g8542,g14596,g32747,g22535,I24625,g5471,I15003,g29862,g26123,I14765,g19659,g20104,g34771,g10110,I18071,g11872,g31853,g20174,g6386,g30283,g34488,g23302,g14707,g28803,g26338,I22114,g28675,g24522,I29585,g17846,g19397,g11409,g18885,g28466,g16260,g24281,g13911,g25510,g686,g19880,g18649,g9660,g32494,g6585,g30031,g33029,g25127,g27468,I20830,g23907,g5016,g25506,g10947,g24367,g23939,g29129,g24715,g34785,I24278,g23378,g24643,g25170,g24541,g21798,g15808,g14626,g11336,g31880,g11126,g21804,g13871,g24082,I24497,g24189,g18718,I15078,g24210,g17638,I12519,g32529,g11994,I32225,g28888,g20133,g24568,g14885,g20703,g21782,g4659,g4628,I28594,g32274,g11993,g30103,g13551,g18715,g20563,g19368,g16861,I32096,g25639,I30761,g34157,g11804,g32464,g7542,g24705,g20616,g34816,I29255,g33342,g6159,I32071,g18155,g30391,I12083,g14248,g28694,g29646,g2648,g24030,g26485,g23552,g10623,I33067,g27031,g351,g11293,g13061,I31242,g30094,g18221,g17617,g22099,g30567,g19686,g13282,g33041,g16487,g25036,g18370,g22074,I30746,g31882,g18712,g25910,g34169,g32170,g28183,g33906,g33866,g26264,g34675,g13460,g34510,g18062,g32280,g30293,I19775,g1752,I33146,g27596,g8895,I14275,g28092,g9698,g9479,g22935,g19462,g6351,g11916,g18138,g15579,g33875,I23585,g5723,g32516,g18103,g5142,g27407,g27402,g25728,g31131,g23139,g29643,g30266,g24422,g19907,g30591,g10427,I19235,g31710,g10677,g17699,g7224,g12154,g18254,I32800,g16712,g8876,g12042,g22882,g11878,g30162,g19653,g34499,g13303,g28372,g32257,g34484,g22207,g18131,g17515,g7868,g24220,g11928,I32651,g24043,g24049,g24731,g22086,g21706,g25674,I26654,g23925,g8357,g22496,g27970,g22939,I14326,g4388,g12014,g28142,g34020,g34761,g31261,g15737,I15981,g33276,g28191,g17593,g18452,g32014,I21831,g21986,g33327,g26275,g28702,g20037,g27467,g17735,g13727,g29517,g18701,g25980,g27985,g9542,g25093,g23565,g22652,g31905,g10585,g13129,g25120,g16126,g29483,g14377,g11037,g32179,g4639,g19935,g24005,g14075,g34097,g31851,g28495,g7236,g6381,g8964,I25105,g25955,I33291,g203,g16651,g9638,g15057,g19600,g28594,g33718,g9982,g26423,g13851,g24380,g15103,g23429,g33477,I20205,g27502,g7138,g28308,g29993,g24457,g23494,g28615,g9478,g23011,g28328,g16181,g19395,g10388,g33303,g25396,I28128,g15748,g19414,g18450,I15811,I12214,g27343,g18104,I27730,g22861,g25202,g16476,g32110,g30336,g21221,g34453,g19747,I18092,g28063,g5835,g24035,g4031,g22091,g33361,g2610,g19760,g13805,I12183,g24145,g32126,g13700,I12278,g30464,g28336,g9415,g32662,g16155,I25846,g20604,g25820,g11035,g16287,g6960,g30308,g31859,g608,I14567,g21183,g23618,g28667,g8080,g32618,g17610,g24248,g10421,g12459,g27271,I23586,g31220,g18297,g31948,g12811,g13130,g32788,g16199,g12855,g14562,g26744,g25038,I13637,I27784,g8805,g8744,g33979,g19762,g5659,g468,g19614,g3494,g12195,g32337,g6303,g14412,g24107,g33863,g23513,g25629,g22073,I14332,g32180,g31666,g31778,g24917,g13627,g18455,g7557,g15815,I20816,g23446,g24331,g24350,g31942,g33120,g7268,g15568,g24630,g12891,g20040,g25447,I13007,g33360,g18684,I33189,g33984,g17505,g11736,g6732,g8504,g11829,I11620,g33600,I20793,g22104,g2445,g26614,g18189,g29637,g28045,g22998,g5901,g12729,g20435,g29669,g32535,g14873,g13915,g11173,g14166,g33273,g14504,g34747,g24337,g4584,g28061,g24961,I21074,g12183,g33420,g19446,g18533,g14180,I29571,g8359,g4991,g11370,g21289,g12294,g31878,g34072,g26725,g21413,g7903,g18235,g28095,g12843,I32297,g21463,g27428,g27084,g16704,I23694,g22158,g29912,g18156,g18727,g17736,g14988,g34255,g8281,g17243,g15720,g34297,g21286,g25045,g33901,I18526,g28613,g16843,g34541,g21351,g23231,g23313,g30016,g33249,g32711,g27225,g34685,I30262,g33934,g24841,g32868,g13216,g23854,g33997,g3368,g4420,g9714,I31474,g17765,g9946,g17509,g24918,g12192,I14352,g32587,g14058,g24269,g33242,g27459,g18989,g30527,g34441,g25080,g31964,g28242,g28036,g26833,g33850,g30127,I28872,I32758,g29743,g17821,g34514,g12890,g22088,g29345,g34701,g6167,g17606,g13280,g32542,g27709,g21772,g14943,g32090,g22160,g12735,g21821,g7666,g11955,g34228,g12100,g31280,g23162,g14892,g10383,I29242,g26835,g33952,g27440,g3490,g24983,I20562,g9528,g34301,g32490,g20784,g15129,I32187,I25242,g20159,g19651,g27087,g20092,g32376,g13660,I21787,g7499,g16702,I32093,g9246,I32985,g6736,g24773,g22359,I17381,I13623,g22973,g14956,g22997,g15074,g33442,g21993,g24010,g16680,g34226,g13215,g33269,g32992,g27617,g7869,g30168,I22425,g10080,g16098,g22923,g22432,g29578,g33705,g32373,g27602,g30535,g31780,g33561,g21365,g31183,g19879,g2089,g12895,g4132,g7541,g30211,g32295,g18316,g30180,g324,g33019,g28705,g14590,g14638,g34031,g19501,I18530,g16741,g29613,g14786,g14627,g29668,g27576,g12590,g33039,I31800,g29887,I32756,I18083,g28085,g22490,g19715,g5681,g15915,g28159,g19953,I17529,I14186,I18861,g26912,g31745,I24705,g28690,g19209,I28572,g9517,g32902,g23475,g12311,g27400,g25019,g3723,g8635,g16800,g17870,I25220,g11953,g25002,g32920,g29252,g16234,g29495,g27251,g19421,g23749,g21754,g26800,I17839,g15746,g20578,g23492,g19330,g5290,g23131,g30564,g16733,g33868,g21716,g27633,g34967,I26531,g18789,g9678,g32721,g10602,g24754,g6957,g2303,g9223,g6955,I31748,g11493,g28136,g13568,g34182,g31325,g24074,I18285,g1287,g7564,g21749,g32640,g30511,g13291,g24645,g25233,g29587,g4382,g21740,I26071,g31524,g27742,g5128,g32750,g4546,g26701,g29190,g33547,g26382,g28673,g32360,I22264,I17173,g29872,g28623,g14045,g6649,g31018,g10649,g17641,g5105,g11030,g21942,I11726,g8626,g28084,g18580,g17779,g9100,g15062,I31878,g25121,g7050,g27338,g31230,g24379,g21674,g19544,g4087,I27539,g32539,g26051,g19649,I23393,g26895,g31831,g18461,g26295,g33293,I13684,g33999,g13876,g23333,I18819,g13600,g10583,g25243,g7888,g18118,g29664,g23510,I18865,g18110,g28498,g24292,g18682,g24544,g6358,g33678,g17672,g21967,g24634,g25593,g28678,g21301,g33703,I31810,g31251,g22863,g19757,I18367,g25735,g7523,g34281,g2417,g30446,g2960,g16190,I21230,g9899,g23010,g33920,g23482,g24125,g8540,I12128,g16681,g7297,g21893,g20509,g8725,g28101,I13183,g34795,g11653,I17653,g34985,I27385,g32453,I32693,g8439,g27362,I27533,g32286,g18918,g17524,g24428,g18510,g18909,g25015,g20541,g16611,I29199,g33603,g23779,g17642,g11303,g33086,g10948,g33368,g30009,g24688,g32859,g7689,g32175,g19534,g27030,g14566,g31916,g33996,g2433,g11269,g28681,g5694,g29302,g27385,g9815,g27091,g33674,g33304,g28066,g18694,g17490,g4311,g26161,g33005,g5357,g15163,g14333,g790,g32469,g12220,g12255,g25088,g599,I32982,g17188,g24681,g18135,g23862,I22822,g20160,I32763,g22150,g1906,I16057,g32748,g5138,I27534,g10182,g25236,g18546,g26049,g34323,g27714,g24317,g24029,g30474,g17364,g20134,g33976,g24789,g32696,g22541,g17213,g29623,g13015,g11039,g2116,g18823,g9618,g9594,I23978,g25381,g21803,g13377,g33262,g20598,g9954,g16272,g5200,g7960,g29869,g26906,g33676,g6903,g16771,g27969,g26543,g19912,g23233,g33135,g27652,g29923,g6497,I12583,g22885,g13304,g31898,g19576,g31554,g34730,I29315,g28827,g4057,g22178,g25874,g23814,I21222,g21731,g10355,g19731,g9822,g16235,g34122,g14841,g16099,g34753,g31541,g10386,I14170,g25527,g28658,g18239,g30089,g30413,g15002,g23252,g14601,g9077,g20612,I13078,g29191,g29583,g11974,g12462,g25231,g1373,g14574,g12049,I23688,g33942,I17636,g34969,g24978,g21876,g12933,g27539,g17096,g13937,g6012,g28814,g1157,g19792,g29477,g25895,I29444,g17600,g16221,g8830,g19266,g33376,g29717,g28645,g27326,g27557,g34995,g10096,g29072,g27315,g4235,I26466,g33713,g31154,g16284,g32057,g18328,g21356,g9616,g25223,g22201,I15223,g20199,g22940,g16685,g31229,g22299,g17476,g17147,g24383,g25267,g16577,g28775,g34887,g14895,g16870,g13175,g11350,I24508,I31342,g5109,g9091,g24343,g32054,g18626,g34986,g8470,g33446,g17151,g25227,g32342,g15154,I27576,g30312,g25034,I19802,g12321,g14741,g20673,g20605,g32317,g31489,g23003,g24364,g27886,g27011,I22665,g23237,g23864,g2661,g23498,g18352,g7835,g19644,I19831,g28851,g25285,g33787,g27457,g28079,g10741,g20384,g2936,g19445,g16177,g31507,g28997,g31923,I13110,g33495,g32774,g7017,g17246,g30559,g34960,g10725,g11122,g19513,g11793,g18102,g2161,g14810,g21747,g7635,g15819,g29028,g13885,g8411,g26218,g22069,g33422,g21789,I25909,g23495,g24943,g21725,g33160,g23517,g30122,g13970,g191,g20922,g559,g29786,I31146,g22622,g2060,I13497,g15806,g34678,g32120,g5770,g9450,g27260,g23433,g17953,g19778,g28911,g13822,g30148,g13174,g24675,g30569,g20506,I26512,g15825,g18242,g30169,g32160,g14675,g11964,g8620,g23299,g9834,I28908,g24559,I24363,g16587,g28670,g34124,g23423,g7806,g18910,I23601,g8840,g29904,g18602,g18669,g4294,g31945,g18710,g25237,g29804,g4473,g7948,g29896,g29359,g7526,g28289,I16502,I32467,g11762,I14764,g25089,I30901,g12644,g21204,g2287,g20610,g9206,g32350,g20179,g34219,g29837,g11563,g12173,g10102,g7167,g18207,g21513,g6255,g15995,g1917,g27289,g25260,g2643,g8177,g28218,I14708,g29973,I18485,g25727,I16829,g14358,g6144,g17180,g27515,g817,g11938,g30328,g16213,g24018,g1825,I21849,g21451,g24718,I31047,g27590,g32412,g4558,I25695,g20322,g33987,g18556,g17264,g29939,g31119,g6187,g18762,g22634,g31827,g23530,g18146,g32531,I16479,g18784,g32645,I13382,g24460,g21160,g22849,g21420,g20594,g18527,g33520,g34877,I17108,g18108,g13986,g18159,g8541,g25775,I28925,g8365,g34876,g14450,g13858,g24297,I20486,g17677,g20626,g10934,g28049,g22640,g11489,g25852,g32370,g23839,g33989,g26309,g32211,g27270,g18897,g2108,g17681,g27342,g17501,g20675,g29068,g24342,g16671,g3167,g18562,g25682,I22499,g16803,g14150,g13060,g13458,g14219,g11130,g1478,I20870,g17952,g32574,I14924,g16768,g9691,g7851,g32086,g23396,g23020,g30277,g12149,g23360,g13716,g13265,g8466,g24760,g30386,g7244,g9830,g24251,g21414,g24385,g6404,g10407,g10726,g27996,g10039,g7624,g32222,I32458,g22836,g22646,g30186,g21403,g22132,g22341,g26899,g29666,g25143,I31869,g9166,g13010,g23230,g1018,g5571,g10570,g17717,I31037,g23422,g28970,I23971,g21770,g11203,g15509,g23841,g33961,g17647,g22543,I25359,g32694,g27653,I26664,g13074,g19794,g7993,I32455,g4427,g20523,I12189,g5327,I12374,g20674,g28263,I23315,g12527,g32718,g24835,g29705,g22102,g21963,g21511,g14238,g16927,g32094,g21251,g9153,I20750,g7158,g25503,I32059,g33359,g34981,g15588,g30021,g13697,g9692,g28051,g16536,g4322,g30264,I11860,g33546,g33975,g24468,g14119,I17783,g24274,g18196,g8508,g13989,g29346,g34224,g1854,g1052,g24270,g9679,g25055,g28239,g24727,g14542,g25648,g20450,g26516,g10737,g24536,g21738,g18481,g33604,g28704,g14397,g33351,g26105,g27875,I17989,g3211,g25633,g16172,g18407,g23881,g5957,g30083,g27281,g28271,g26298,g26913,g28058,g23558,g24532,I15921,g30440,g16286,g31931,g21396,g26079,g26336,I15174,g11615,g24116,g29478,g27292,g13006,g34193,g11537,g28250,g28065,g13032,g11980,g29350,g33450,g14186,g29631,g8680,g12905,g23506,g30543,g21847,g14452,g4054,I16575,g26925,g18290,g30983,I33075,g28733,g21976,g32894,g23885,g34592,g23451,I15042,g19068,g27510,g34351,g30015,g27458,I12858,g15862,I20216,g22680,g8112,g2894,g26327,g10143,g13856,g14432,g30163,g29203,g13580,g30369,g26205,g33248,g18492,I31659,g21339,g24808,g31856,g14946,g24485,I22024,g34867,g9780,g34530,g19885,g32816,g29225,g17427,g27521,g33730,g19738,g20914,I13552,g20627,g11111,I22710,g10414,g21778,g21992,g14395,g22716,g10489,g12129,g29577,g12873,g23398,g13672,g21285,g21987,g11385,g21989,g27685,g15807,g1700,g6988,g26261,g11640,g8282,g33410,g29888,g14911,g136,g29250,g12465,g12823,I14158,g25328,g33840,g22143,g11445,g23395,g10391,g12045,g31271,g12587,g8700,g31763,g14528,g10392,I32973,g18299,g29933,g12075,I11688,g9337,g34198,g1604,g25073,g28966,g20665,g28598,g9639,g5535,g33363,g29920,g31990,I29149,g29169,I24695,g13018,g19748,g32359,g14613,g25885,g10521,g28710,g26576,g31797,g24156,g12314,g34755,g30408,g9338,g34110,g22544,g25449,g33239,g3436,g32407,I15736,g18369,g21759,g29579,g12147,g32182,g25196,g30176,g14755,g24872,g30220,g11996,g21431,I17249,I12544,g31516,g28151,g34311,I31046,I16780,g12806,g24004,g10130,g30173,g33983,g25551,g12793,g18814,I14999,g11204,g24374,g29856,g32839,g15634,g14496,g7827,g24027,g34385,g16268,g21206,g12163,I31727,g28197,g32955,g16662,g7397,g28010,g24660,g22317,I16770,g23251,g34767,I14883,I18245,g30036,g21307,g16473,I15168,g21911,g5731,g19140,g27829,g31146,g14184,g1664,g20649,g20088,g25737,g30421,g25100,g12374,g32841,g27509,g14695,g14033,g12109,g21732,g28290,g10618,g9731,I23756,I17787,I12056,g2357,I26679,g4527,g21686,g32386,g34568,g20581,g25964,g25357,I13802,g14503,g25622,g33834,g28080,g21336,g22852,g26956,g12550,g23377,g9827,g15373,I31147,g23763,g11231,g13329,g15962,g32759,g28078,g12,g16227,g28185,g34186,g7183,g13279,g10166,g17720,g28998,g6549,g22636,g25152,I31814,g34710,g33331,I23987,I18048,g13474,g26911,I29891,g12903,g28164,I12360,g17179,g3742,g29665,I30054,g25150,g27376,g28719,I28480,g17199,g22976,g11992,g13321,g15143,g26765,g24301,I12534,g33098,g34512,g20711,g15064,I19799,g26125,g7069,g18202,g29634,g29280,I24396,g24061,g31290,g25962,g11016,g16958,I31202,g8737,g25713,g17478,g29479,g1514,g27775,g29692,g28610,g12860,g19555,g33631,g18622,g28232,g14208,g33187,g23488,g26732,g10533,g27114,g20667,I12263,g31817,g10378,g28198,g27154,g18717,g27129,g11135,g33034,g34152,g13497,g5791,g19684,g33922,g34126,g6239,g24930,g21853,g6,g25757,g13909,g33428,g25957,g31248,g34402,g546,g12749,g12628,g26285,g15124,I32231,g33708,g25987,g22547,g18819,g9751,I32203,g17287,g23348,g6307,g29791,g10381,g2795,g6772,g15714,g28251,g23917,I31322,g15053,g2955,g18382,g232,g25901,g7891,g23716,g24561,g7461,g20093,g6573,I14579,g25423,I29236,g22117,I24364,g20448,g29970,g33926,g25865,I18543,g10475,g32607,g4899,g28629,g32976,g5591,g14018,g29886,g29262,g29905,I18168,g19517,g24803,g31616,g12819,g21977,g24152,g12252,g6513,g17200,g10074,g22170,g34636,g20535,g4843,g7558,I21100,g16844,g28121,g23421,g27450,g475,g28238,g11382,I32591,g10109,g20738,g28133,g25321,g30475,I20529,g33050,I13139,g30068,g30934,g10368,g32186,g32851,I28588,g6868,g28934,g21334,I21480,I26705,g15722,g7781,g18209,g12357,g7543,g33354,g18190,I32109,g25241,g8847,g32860,g33296,g15161,g34208,g6817,g33312,I25366,I32678,I22929,I31463,g20277,g16661,g34050,g11431,I12279,g31000,I20647,g5925,g34643,g22639,g27615,g32972,g16597,g21979,g31134,g20130,g27724,g25504,g28115,g22987,g28315,I24384,I32440,g24081,I31087,g31837,g17872,g27205,g8522,g18267,g34158,g31017,g22875,g31476,g31986,g33573,g17155,g17492,g24318,g26483,g29897,g18662,g34849,g12341,g18301,g34707,g18534,g26486,I12076,g24999,g10537,I26004,g18760,g31307,g28497,g34738,g29713,g30412,g32151,g24622,I11635,g7212,g452,g365,I14684,g11223,g10290,I16181,g13939,g23431,g11251,g25192,g19777,g24642,g18164,g1821,g17191,g16842,g32813,g20046,I18165,g16066,I22944,g1333,g8743,g5092,g32950,g20442,g30112,I31337,g28478,I18476,g12052,g5673,g6247,g4512,g33480,g12343,g29490,I12241,I32806,g16705,g19441,g7175,g23399,g22061,g27185,g18120,g30118,g33971,g13820,g23450,I22143,I17166,g29511,g30487,g30140,I12344,g16926,g10851,g6998,g21842,I22966,g19388,g613,g28569,g26055,g3546,g34873,g9012,g22851,I24461,g34787,g11674,g21271,g19906,g15090,g25923,g32174,g15739,g21290,g21742,g34045,g19471,g25929,g32471,g25944,g33468,g28081,g31187,g22220,g29944,g23260,g21888,g30181,g7907,I23360,g32235,g16621,g19386,g28298,g32465,I23979,g23720,g17121,g347,g7431,g19481,g24044,g32421,g31809,g19636,g31791,g15155,g5603,I14204,I22031,g5424,g18571,g26818,g29751,g28317,I23327,g33127,g283,g13143,g32685,g18194,I21810,g26229,g25770,g33849,I18276,g33576,g4669,g25611,g27646,g1283,g2606,g28546,g15726,g10133,g21761,g24349,g28765,g31850,g333,g12898,I26522,g6756,g18977,g7396,g16618,g25060,g32648,g18568,g33513,g24155,g2518,g21188,g27588,g20591,g19604,g11025,g18514,I13287,g33314,g19200,g13793,g19767,g34271,g14179,g25525,g15907,I17494,g33988,g12073,g20571,g25649,g16716,g24159,g25741,g20668,g11207,g20446,I14817,g20443,g14048,I23950,g21269,g27138,g4534,g29926,g24719,g30424,g21815,g22035,g18379,g34439,g28555,g20006,g18731,g11320,g10197,g25222,g14393,g24820,g6271,g20596,g21930,g20602,g34455,g11937,g17592,g30530,I27713,g19565,g9976,g16839,g34391,g34965,g15959,g11190,I12345,g4771,I22974,g9103,g32940,g9985,g12038,g20085,g25079,g20445,g34115,g16646,g24076,g25217,g21917,g30128,g29630,g9154,g24708,g9180,g19964,g20050,g2803,g29846,g18832,g25521,g25041,g34017,g13808,g13314,I22280,g29616,g26272,g10153,g28924,g7439,g32937,g2844,g27394,I27555,g34845,g16759,g25172,g12525,g5244,g32833,g23493,I18125,I31027,g18487,g34802,g26187,g30371,g29314,g24045,g31846,I12884,g18406,I17679,g21346,g12367,g28605,g21997,g33980,g25182,g21609,g8456,g12059,g16815,I13539,g10373,g21839,I22583,g33130,g5863,g18167,g13094,g28619,g13661,g19750,g25450,g18210,g16598,g27732,g32013,I31469,g23182,g26871,I27970,g33257,I31246,g9977,g22698,g29510,g1129,g29737,g33490,I27570,I13872,g12857,g13959,I23949,g3151,g14234,g31926,g26025,g1728,g5555,I18214,g26606,g28097,g16639,g15935,g21419,g4727,g17759,g34564,g32621,g26019,g8712,g25012,g32837,g12940,g29547,I22470,g25709,I33167,g3863,g29312,g12705,g16524,g29806,g15036,g13940,g9575,I16663,I27495,I17834,g27150,g19592,g6946,g30477,g34894,g19869,g34467,I31192,I19671,g13298,g27178,g29760,g29676,g34644,g34477,g17511,g14101,g30404,g29942,g7918,g8676,g34335,g18220,I18891,g27559,g13026,g18994,I13202,g12227,g18634,g3632,g23515,g26546,g7933,g31876,g30046,g21363,g18377,g21881,g28837,g26714,g24772,g19930,g26850,g10082,I15697,g16232,g9374,g14438,g28400,g18414,g12593,I29303,g24067,g27451,I18829,g7086,g24046,g26082,g34406,g32268,I17094,g9721,g13621,g21774,g22050,g33661,g19957,g14258,g27085,g18271,I33182,g128,g23825,g24761,g22624,g5937,I12240,g28456,g34591,I12289,g30729,g29244,g27589,g28576,g34269,g8088,g32492,g31189,g6828,g22844,g25157,g4826,g32548,g9728,g33927,g32630,g31184,g32904,g12143,g12779,g23262,g34375,g29953,g18894,g15708,g33387,g25801,g33820,g25003,g34133,g24913,g11779,g24287,g34871,g30461,I16541,g19740,g32988,g20178,I24552,g20567,g34486,g9226,g12198,g31813,g7469,g32592,g33461,g34123,g20916,g15091,g22670,g27998,g26087,g33978,g32176,g32637,g33883,g27991,g30375,g34350,g26836,g33083,g33322,I22571,g34870,g11128,g28161,g27779,g33470,g18474,g7880,g21402,I15382,I22921,g18703,g15799,g11741,I18086,g25925,g27537,g31224,I26785,g1239,g7841,g15849,g23782,g18987,g28358,g18793,g27229,I18778,g24564,g22003,g21802,g20239,g30419,g28701,g32336,g10610,g18570,g9640,I31177,g20188,g967,g5390,g9898,g2710,g23214,g23284,g34583,g26745,g30091,g25369,I32067,g33772,g30191,g13107,I18262,g23879,g7074,g23613,g34229,g22151,I31131,g14122,g385,g3901,g13972,g20034,g1840,g4019,g2856,g31133,g25000,g5543,g14297,I12950,I22923,g17625,g21729,g22065,g12256,g32820,g10801,g10604,g9629,g32978,g16670,g11811,g24105,g34303,g28616,g11114,g32141,g33133,g19981,g30347,I14830,I13606,g2193,g11139,g11609,g19931,I22316,g32203,g26789,g27140,I16498,g20600,g8553,g32333,g32687,g14133,g27474,g24028,g19719,g24158,g31843,g1459,g5436,g32901,g18175,I14668,g32441,g34306,g12862,g8678,g28462,g15116,g18704,g23815,g10159,g20648,g18768,g336,g12592,g23835,g29374,g25063,I22525,g25555,g34560,g26241,g34555,I31803,g20614,g34036,g2638,g34095,g5381,g7660,I22684,g8623,g34026,g4549,g28536,I31001,I14893,g18363,g18141,g34487,I27927,g27010,I12103,g16233,g6854,g14820,g23217,g8904,g12181,I19384,g28761,I20913,g2403,I31247,g29237,g10658,g24429,g33816,g2912,g19674,I12242,g13249,g23767,g20613,g26834,g24839,g11810,g16877,g32498,g23004,g6711,g10224,g31841,g31994,g6985,g21306,g25664,g22883,g33734,g19371,g12821,g7285,I31347,g18454,g31708,g8070,g17533,g28039,g25275,g34296,g20530,g10040,I14602,g7943,g24647,g14378,I11908,g32943,g32916,g17154,g34458,I32388,g17391,g34434,g5873,g29317,g32917,g18801,g13035,g7404,g23605,I13518,g22528,I14530,g34065,g28118,g28962,g31123,g11003,g28236,g29301,g30486,g30289,g29735,g26273,g16193,g11663,g23227,g30249,I33249,g29269,g25960,I17901,g27594,g6821,g25928,g28112,g29866,g32296,g16185,g10971,g28188,g27578,g933,g29927,g29765,g15830,I31807,g29316,g15094,g9184,g32125,g19487,g763,g34419,g18232,g24079,g29762,g12226,I22539,g27255,I18537,g19980,g16700,g29588,I12826,g25538,g12920,g18211,g29885,g30039,g24552,g18607,g23883,I13520,g29644,g17718,g33305,g29843,g17609,g29891,I16345,g29104,g391,g18408,g22137,I14766,g12852,g1532,g34380,g29651,g18744,g8956,I20747,g28889,g26094,g26260,g14825,g27243,g25930,g10611,g17810,g18165,g21249,I31535,g25653,g11933,g22100,g24420,g29624,g20547,g5615,g16280,g26860,I31336,g18215,g16508,g25246,g20103,g30243,I11865,g18308,g30471,g29043,g4349,g6830,g22649,g30505,g24939,I11877,g11191,g23995,g11907,g28745,I20233,g17216,g28980,g16474,I27579,g25056,g19690,g25113,g10077,g23553,g13139,g13715,g18214,g16773,g26256,g20696,g21427,g28773,g31996,g2259,g23353,g33529,g11324,g29526,g14681,g23732,g10675,g6814,g28572,I12608,g21946,g24924,I17808,g7304,g23271,g27312,g31800,g16289,g25624,g10190,g20510,I24585,g24201,g28470,g11110,g9715,g23904,g34256,g25006,g21852,g20231,g25866,g8913,g32895,g20574,g16724,g22753,g32461,I22467,g30417,g31746,g18255,g27026,g24997,g16215,g4815,g34411,g18773,I22619,g18543,I15821,I11980,g23397,g32877,g16746,g22633,g1221,g20701,g29040,g23434,g18422,g12996,g28031,g19526,g31864,I31266,g21849,g18139,g25766,I25689,g20631,g18355,g31284,g31566,g7533,g24404,g5893,g23607,I18674,g19875,g19543,g2437,g10354,g20560,g18381,g11941,g26653,g34879,g17652,g20195,g24809,g9472,g33241,I14855,g18132,g32313,g17598,g3100,g34337,g19786,g12897,I13149,g13475,I14702,g11720,g21828,g34098,g28651,g2917,g1418,g33106,g12938,g18240,g28713,g4955,g25206,g13771,g14663,g16734,g34801,g6494,g30407,I24331,g14441,g34613,g18392,g32036,g3703,g12578,g18632,g27926,g23239,g33494,g11866,g8765,g34673,g28607,g34452,I32827,g437,I26479,g32049,g4520,g20772,g21659,g23659,g13077,g14231,g27995,I33024,g344,g33838,g30048,g21744,g30179,g1404,g11410,g20579,g14232,g34408,g16707,g33588,g34485,g27074,g20562,g17086,g27240,g21060,I15872,g20993,g20537,g4076,g19585,g34481,g2241,g34932,g18780,g27009,g19343,g28620,g27266,g12136,g27134,g9630,g18521,g14272,g25532,g18541,g24717,g7322,g27316,g34807,g23630,g9753,g433,g26178,g15115,g20769,g9429,g34290,g34603,g14291,g28102,g3147,g18158,g11412,g16516,I32766,g27645,g34823,g25071,g27279,g33540,I22788,g32936,I24060,g4933,g30224,g7828,g28628,g34265,g8673,I17462,g28272,g12692,g7680,g30296,g27282,I32809,g34268,g16954,g32300,g30825,I14727,g29992,g9669,g29618,g8426,g31296,g29173,I23345,g32963,g32615,g18711,g28297,g13583,I18855,g12017,g26360,g27983,g23088,g23132,g18951,g6637,g6434,g27955,g7133,g26289,g7261,g19393,I13498,g30377,g34748,I19704,I31486,g15088,g32246,g21981,g33476,g5134,g19520,g21275,g25789,I21766,g29730,g20325,g13676,g34883,g18620,g31238,g31868,g25245,g32588,g32501,g16713,g30403,g33888,g24377,I26948,g18354,I22893,g34799,g33310,g5831,g24015,g10776,g24009,g32724,I27509,g28441,g25264,g33899,g29315,g24032,g19886,g22097,g9187,g19947,g401,g28692,g7472,g33275,g1413,g5853,g27582,g22340,g19265,g23127,g32308,g15123,g11346,g29799,g18282,g15139,g18153,g34941,g12301,g28147,g12337,g29508,g24537,g27122,I31206,g24709,g24641,g26702,g21879,g30027,I15341,g34920,g13888,g28403,I22824,g30223,g29968,g21887,g13066,I12199,g34975,g32491,g27961,I12252,g32834,g12381,I12644,g34210,g13796,g22165,g14335,g12043,g28543,g11472,g27131,g15067,g28020,g26843,g33954,I13454,g32477,g6754,g21284,I14119,g25884,g16316,g23742,g28342,g10896,g22139,g28688,g21746,g30038,g21353,g10624,I12167,g29610,g18133,g32323,g31798,g25726,g28709,I28548,g11396,g30236,g16238,I23324,g30606,g19680,g23616,g10376,g11862,g34028,g32910,g24034,g34319,g16896,g30433,g24491,g28296,g17582,g20150,g9913,g23889,g33012,g24262,g29272,g14454,g29371,g17599,g32012,g31130,g17150,g2173,g18188,g16206,g14051,g33592,g18575,g27684,g9708,g15979,g15754,g33358,g28230,g25992,g9056,g34615,I14225,I31504,g13517,I30537,I31021,g26345,g12798,g32209,g18405,g28229,g27388,g25242,g17197,g34558,g28570,g16427,I32079,g23780,g15147,I24781,g32795,g3111,g1554,g34002,g28780,I12808,g19580,g5782,g21308,I18421,g19890,g30184,g22209,g16737,g28537,g34309,g16638,g12190,g13955,g15095,g23021,g26955,g17768,g27275,g28684,g6329,g22860,g23516,g27046,g23273,g8102,g16929,g32551,g21970,g23279,g27057,g15144,I17380,g691,g18456,g21745,g28269,g1361,g13850,g26680,I19778,g27762,g19,g33887,I20116,g24921,g23563,g28288,g28622,g27525,g29983,g32403,g3518,g26667,g32111,g20230,g18283,g23167,g27931,g16655,g10420,g29657,g14927,g15723,g19502,g14851,g8310,g5523,g34472,g23961,g17410,g18497,g12002,g26276,g2756,I25907,g25596,g34469,g34509,g5084,g24444,g3905,I12064,I31072,g19442,g1500,g16866,g11559,g33537,g7166,g26294,g26511,g29787,g23229,g8565,g33405,g24757,g34847,g11467,I31121,g10037,g27145,g25144,I24597,g4204,g31124,g33686,g21010,g27535,g12778,g14953,g24378,g23435,g21835,g10369,g24208,g6098,g29147,g5965,g3195,g14543,g31785,g10266,g27572,I11626,g30922,g31144,g21377,I26643,g23258,g9326,g3602,g28137,g14665,g4489,g21421,g14679,g22526,g11845,g28116,g20663,g25040,I27749,g28687,g29940,g23629,g33051,g18432,g29881,g6977,g18692,g30247,g28715,g11915,g34642,g19505,g14252,g26547,g29895,I18581,g25492,g23549,g20977,g25160,g10160,g14520,g14750,g30506,g14216,g32256,I16618,g15589,g25399,g262,g19144,g24250,g34197,g20900,g23533,g34659,g32225,g30288,g19770,g27550,g30154,g34055,g6832,g28463,g8356,g8763,g12436,I23120,g17584,g20920,g16612,g19542,I15002,I32921,I23381,g20128,I15647,g33696,g33062,g31233,g4688,g25086,I17733,g32217,g32661,g14588,g22135,g18665,g32354,g10417,g20207,I13564,g16485,g5224,g29311,g21961,g33462,g9636,g14197,g19772,g20273,g25069,g10561,g11031,g11363,g9984,g34285,I14247,g20638,I15915,I17857,g35000,g23476,I32935,g21871,g24418,g11900,g34096,g18806,g23921,g16540,g29863,g14781,g17088,g18621,g32267,g26518,g26924,g29906,I18587,g22907,g22153,g10552,g15699,g4537,g31376,g24465,I31625,g21423,g11048,g15717,g13271,g24671,g25466,g5827,g27303,g25779,g4932,g12450,g25769,g19793,g23898,g18260,g34398,g30200,g30572,g4765,g8105,g33862,g9536,I13779,g12908,I24015,g8914,g18195,g24212,g29145,g16690,g150,g34495,I22343,I21238,g1720,g23623,g24558,g13834,g18362,g34063,g23599,g10219,g14996,g20388,g27771,g8696,g14002,g28435,g18747,g10319,g33879,g8396,g8821,g2342,g16123,g17464,g22357,g16660,g18531,g28927,g15083,g23298,g3550,g17726,g24887,I18872,g18816,g20507,g22068,I12811,g18420,g14295,I16117,g7490,g30439,g30937,g16801,g18184,g7258,g14751,g23084,g22307,g8068,g31760,g13977,g24663,g32802,g33545,g31139,g34557,g23967,g28203,g29207,g34059,g31242,g33026,g29718,g31218,g7352,g26977,g25165,g18980,g25905,I13995,g18343,g13463,g33423,g15752,g22039,g26081,g6811,I16898,g32388,g29790,g25969,g33831,g24132,g18400,g24363,g25546,g117,g8766,g27877,g32357,g25185,g9061,g30394,g10705,g12739,I16486,g26825,g21713,g31826,g29709,g22472,g28642,g34676,g24525,g12428,I14970,g31879,g12289,g21724,g22001,g25571,g28209,g32569,g921,g2999,I31162,g18891,I18900,g21330,g8854,g22006,g28307,I13317,I29977,g23307,g34051,g25051,g21067,g16031,g33087,g29060,I24078,g32483,g23188,g24415,g16128,I14229,g24346,g33517,g14359,g28153,g30926,I32158,g34172,g26887,g32144,g25368,g24141,g24915,I18301,g17475,g25715,g31988,g5120,I18482,I15620,I14518,I23387,g26880,g25023,g32039,g9960,g15903,g34496,I17121,g11773,g32809,g15798,g3408,g15721,I11750,g32088,I25586,g23226,g22493,g31126,g24402,g23201,g28510,g19779,g9911,g32305,g8180,g15068,g18517,g22308,g25640,g8663,g32159,g21415,g17325,g11715,g33228,I14633,g1714,g33350,g32530,g33700,I17585,g18385,I24128,g29491,g33527,g14164,g16625,g30444,g26967,g25135,g14655,g32593,g23541,g20532,g25733,g32493,g13267,g32869,g25765,g26252,g11380,g26391,g13412,g24849,g30297,I15284,g10356,g27324,I23163,I26051,g3639,g3103,g27103,g19873,g28867,g26204,I26394,I22461,g32850,g32693,g22835,I15587,g25738,g24307,g23221,g31166,g12522,I15869,I18671,g34833,g29231,I31622,g26972,g24118,g23358,g28135,g11512,g29166,g25084,g21416,g25548,g25138,g29092,g24063,g28172,I12954,g22920,g20056,g30045,g3661,g29766,I22400,I24448,g33616,g30507,g25670,g21181,g24203,g6259,g7873,g26902,g30612,g34860,g21861,g33507,I11816,g31858,g23223,I14213,g3586,I12994,g11193,g33544,g23896,g33328,I14885,g1612,g24407,I17750,g9821,g160,I32601,g21834,g12340,g7752,g18340,g19453,g23128,g8086,g12423,g14212,g29853,g28349,g19503,g12430,g2181,g1227,g28370,g17741,g18171,g28674,g6423,g34212,g31894,g18725,g26776,g20565,g18584,g10014,g23863,g25125,I25677,g14879,g14163,I22464,g33689,g21061,I13726,g33514,g26313,g22867,g24000,g29599,I12333,g28991,g26908,I24920,I15316,g34732,g23317,g33281,g29763,g32459,g11238,g13045,g23684,g30095,I18782,g19537,g28082,g12892,I29720,I33282,g23786,g28385,g22046,g26952,I22816,g7161,g34293,g20161,g34451,g29093,I32228,I18580,g4284,g25194,g12449,g18353,I31052,I16590,g11819,I23985,g12847,g20449,g32187,g15109,g26710,g34534,g34188,g23304,g5719,g13043,g29582,g23170,g27127,g26656,g32658,g34146,g32414,I31776,g33857,g18763,I31848,g25255,g32642,g33219,I18297,g18653,g33288,g34630,g32801,g23685,g18513,g21459,g14875,g9051,g15863,g18219,g30064,I22762,g15071,g30282,g32659,g18576,g12122,g10413,g7991,I13483,g22650,g17596,g26050,g32195,g3676,g32249,g18327,I17148,I31642,g34550,g29835,g9933,g33575,I24022,g24467,g12999,g4776,g27769,g12201,g34227,g24818,g9649,g21701,g11963,g13923,I22131,g33369,g21652,g27380,I13906,g29550,g14512,g9155,g7184,g19482,g27711,g22539,g32767,g29675,I21477,g30126,g26244,g26679,I13067,g28591,g26884,g33784,g19670,g9816,g25226,g15816,g34456,g27959,g20214,g34021,g26247,g32302,g27112,g22025,I13875,g29370,g24466,g23085,g22081,g29489,g11965,I24281,g9567,g19855,g32450,g19443,g8224,g17317,I18667,g15119,g12476,I18492,g18491,g18641,I33261,g32684,I23149,g26792,g33025,g5677,g7096,g16158,g9906,g15018,g28475,g24207,g26323,I17612,g18388,g17297,g14581,g23955,I21058,g11744,g19887,I20840,g2523,g2407,g13469,g19147,g33023,g11956,g33045,g20781,g31847,g32395,g3215,g16231,g22210,I24041,g23189,g19745,g22329,g33521,g23504,g3231,g27817,g25579,I30192,I11685,g32156,g27259,g32510,I33027,g12911,g16885,g12126,g10627,g20539,g930,g26862,g28171,g7456,g16323,g32537,g34230,g21780,g32472,g34989,g33362,g4269,g34107,g23014,g9924,I13152,g26928,g31821,g31808,I15550,g16806,g33528,g5949,g24231,g6219,g31744,g28311,g13095,g24205,g17486,g28661,g34971,g30158,g10695,g13121,I12049,g5567,g8594,g20175,g21903,g17709,g29551,g21247,I24694,g13042,g12687,g8593,g34584,g27323,g26815,g8164,g1632,g6151,g27675,g15932,g11826,I30331,g1677,g25382,g28352,g24198,I31122,g19367,I18835,g19799,g18126,g32984,I31569,g27686,g34600,g33972,I31152,g25851,g32149,g27203,g33258,g1862,g30252,g24275,g34241,g7892,g34946,g25646,g27158,g21775,g11261,g26905,g24294,I18135,g10335,g12185,g28243,g25043,g26155,g24836,g26542,g2165,g30555,g33282,g26253,I17207,g18772,g25632,g14772,g16528,g23250,g21068,g4519,g31288,g31914,g27027,I12987,g18783,g3267,I12469,g24960,g16599,g26512,g20712,g24356,g11903,I31796,I31779,g23321,g32725,g13144,g13779,g21877,g28582,g17670,g3610,g10708,g21912,I31071,g27647,g29523,g26101,g30370,I15878,g11973,g18418,g18590,g25816,g18879,g33860,g30216,g22197,g27830,g34964,g8005,g27216,g31486,g25559,g10819,g21880,g34517,g26755,g7097,g18672,g11997,g19433,g2122,g8714,g29261,g24233,g3990,g10079,g1008,g33882,g32882,g34131,g24387,g32204,g32790,I15906,g9968,g22717,I31157,g15051,g24623,g26281,g14391,g32051,g23774,g18600,g14110,g29845,g27455,g22762,g16000,g26129,g30381,g30011,g27773,g34103,g17648,g14181,g28047,g16510,g24793,g24355,g30503,g14676,g20146,g23480,I13054,g26752,g32647,g30123,g28410,g18364,g32560,g20705,g12695,I32960,g24419,g21867,g7809,g34782,g12146,g534,I15623,g24024,g18378,g25916,g12292,I26100,I15335,g26097,g22845,g24267,g33143,I31459,I31257,g25098,g17526,g10275,g33559,g26883,g30596,g758,g14090,g29552,g23542,g33951,g33247,g29882,g34213,g24499,g15650,g12944,g32193,g32070,g21762,g28513,g34248,g7992,g29732,g16075,g25771,g9888,g8639,I18694,g10542,g26650,g32273,g17296,g31788,g16695,I12776,g13999,g31475,g21786,g26180,I25594,g26929,I14790,g901,g27903,I15102,I17876,g18484,g25667,g33760,g32585,I31858,g23751,g33502,I20488,g24188,g33497,g21928,g27858,g22720,I19759,g6782,g25704,g16310,g21177,g23007,g14361,g10874,g34093,g32649,g7142,g19566,g27256,g26515,g7537,g9903,g25745,g32307,g33438,g1526,I12033,g15882,g21808,g10142,g33403,g7618,g34231,I18443,g30172,g23511,g33562,g34700,g28416,g27119,I12451,g27012,g1256,g21425,g34409,I19857,g28212,I17447,g24401,I15041,g6455,g18208,g27663,g13021,g7749,g26091,g9372,g34796,g22858,g32713,g28581,g26649,g22538,I33273,g20067,g9809,g23522,g28157,g18238,g11984,g24475,g12952,g11373,g18812,g18761,g8616,g18746,g29652,I31672,g21666,g17248,I17956,g13473,I26741,g28099,g20077,g28899,g10395,g27244,g23259,g14228,g30427,g34549,g9011,g26342,g23301,g22309,g11163,g15867,g24280,g27469,g29952,g24373,g14001,g20572,g29070,g27723,g26341,I30740,g27204,g34433,g4098,g21677,g33802,g10550,g26352,g23793,g14720,g12700,g17708,I18177,g19277,g24278,g1024,I16163,g27108,g22109,g27361,g18152,g32782,g31965,g18656,g5236,g3061,g5335,g31008,I31523,g33726,g28920,g26826,I17406,g27973,g34798,g4164,g34388,g16472,g22926,g14790,I12907,g25759,g24766,g20197,g15674,g30389,g30522,g10878,I24440,g16308,I12842,g24271,g8863,g16529,g25229,g30044,g34709,g33455,g9442,g30073,g19744,g15844,I26742,g20589,I17395,g30492,g18603,g21673,g12107,g25636,g14029,g25261,I15609,g29304,g5511,g9003,g20841,g34679,g8267,g29589,I31984,g23756,I15144,g29368,g27186,g14548,g34260,g66,g18008,g23914,g25284,g12235,g14256,g18765,I30983,g21180,g31596,g4414,g20669,g31772,I18028,g8686,g17766,g7598,g30353,g24106,I17704,g34765,g22651,g9576,g29803,g33237,g20545,g26301,g2047,g26743,g14194,g23208,g32183,g21279,g18357,g24400,g20764,g21883,g23620,g27731,g14011,g24504,g31482,g24724,g20094,g8400,g33658,g23308,g20136,g23376,g15680,g12047,g18573,g31326,g15146,g23746,I26503,g24221,g23479,g12477,g10261,I16709,g7887,I22729,g34611,g7963,g23309,g30493,g30156,g21690,g18145,g18296,g22227,g12120,g13960,g31373,g13007,g7548,g25684,g33482,g22632,g3361,g4401,g15097,g15086,g33563,g25717,g7831,g25523,g29784,g23042,g24078,g14399,g27565,g25623,g7753,g10320,g13084,I14712,g31167,g30025,I22561,g26048,g26816,g10401,g11892,g24126,g1205,g8390,g31305,g30384,g16802,g16203,g32521,g31505,g1056,I31102,g12137,g21343,g20058,I20318,I23342,g23686,g34851,g19672,I22458,g18375,g21969,g20716,g26325,g23726,g25578,g27358,g28567,g26613,g25366,g9239,g22192,g33095,I14241,g31149,g18451,g12998,g26872,I30989,g15656,g10002,g9818,g16178,g25263,g20194,g32668,g28556,g19932,g31866,g25240,g25448,g22048,I25743,g30165,g23412,g18368,g9541,g28612,g13022,I15617,g30208,g32433,g23030,I15577,g12417,g28257,g5022,g9234,g13868,g31241,g30397,g21452,g25696,g23877,g25773,g17518,g17732,g34852,g5421,g32653,g28134,g18246,g19466,g32242,g15118,g17474,g25976,g34464,g16782,g19510,g24069,g34674,g9451,g28521,g4836,g17737,g7536,g9889,g30137,I29295,g11971,g33255,g17691,g1046,g8300,I29352,g23836,g16735,g22041,g30497,g18724,g33231,g13919,g19856,g19389,g11290,g18396,g10419,g14575,g30931,g34609,I12523,I17552,g34955,g10671,g29300,g25740,g32142,g32739,g23406,g27395,g28119,g9700,g14713,g12822,g32991,g24135,g11214,I21860,g2681,g2711,I31176,g31480,g31935,g15059,g32330,g25932,g8363,g24545,g34608,I29270,g30410,g17399,g10617,g33367,g15137,g28057,g29608,g22106,g14855,g14611,g22155,g30147,g10733,g30936,g18565,g21253,g20570,g11446,g30498,g25580,I17188,g29597,g11270,g29635,g10117,g30166,g7619,g30916,I24215,g34573,g32764,g9967,g11626,g9284,g15713,g26308,g24241,g15017,I21199,g11979,g31273,g32927,g31246,I32106,I15800,g25550,I18270,g24989,g20514,g34820,I17379,g32646,g25198,g25049,g30157,g17149,g2177,g13297,g23930,g23319,I11777,g24776,g34121,g27412,I31261,I32516,g6923,g28614,g32609,g25103,g16585,g34602,g15967,g2735,g34442,g26770,g10084,g1521,g19412,I14609,g32923,g32555,g13521,I18810,g28533,g9992,g32237,g24819,g34364,g14688,g32929,g21383,g20874,g34723,I15814,g20632,I16721,g12831,g27332,g2393,g23013,I29973,g29260,g11184,g13092,g19337,I31017,g30087,g32168,g24589,g34520,g28777,g23218,I24784,g21272,g25730,g10262,g2250,g27583,g29313,I31112,g19410,g9733,g23991,I32846,g15113,g30178,g21806,g18539,g21355,I23951,g33607,g23576,g18528,g18480,g25564,g10929,g21608,g10050,g34302,g27826,g29694,g14669,g26759,g9626,g29889,g33084,I24415,g3412,g28499,g9581,g18105,g19552,g10394,g13665,g23303,g27034,g24854,g25784,g15736,g24683,g11820,g14642,g19523,g34988,g15157,g11823,g33985,g33587,g26926,g32822,g15874,g14600,g26941,g24785,I11825,I26952,g21062,g18795,g341,g10970,g32930,g34061,g7751,g34308,g18550,g34869,g34310,g32262,g24217,g33682,g26909,g27968,g12804,g25420,g33272,I13020,g30489,g16509,g34270,g29358,I22864,g18163,g33832,g19498,g25802,g31875,I32621,g25600,g25116,g28549,g26823,g33236,g24667,g14097,g17601,g28375,g30221,g20190,g31901,g27735,g18516,g25917,g27217,g7858,g21718,g29684,g19605,g13260,g10621,g21184,g1886,g22761,g29812,g28649,g29029,g18507,g33628,g8217,I23671,g29840,I32963,I17842,g34181,g21011,g33053,g18395,g11006,g28640,g5057,g30133,I14735,g25641,g16279,g32786,g12079,g13005,g5475,g10815,g27135,g15797,g33280,g34861,g10336,g20171,g18601,g30077,g30175,g32765,I22989,g33110,g32138,g31188,g11002,g10205,g21186,g19854,g24549,g17428,I20846,g34677,g24777,g5802,g18930,I12896,g25940,g32505,g13288,g18212,g23151,g33519,I22800,g27924,g34003,g33992,g24505,g19570,g25370,g29688,g32277,g30395,g24253,g31485,g10724,g23966,g24110,g6287,g26608,g9099,g26709,g22027,g19718,g24219,g12490,g22834,I22685,g16220,g1936,g15101,g4646,g28744,g20004,g34811,I20223,g27290,g32688,g28127,I13519,g29239,g32324,I25591,g11497,g33898,g26379,g34038,g14829,g30733,g34939,g7424,g27703,g19476,g12893,I25095,g13307,g26088,I32770,g24431,g7527,I20864,g34688,g23537,g33806,g31311,g32189,g20069,g28609,g24261,g20502,g17133,g12020,g24804,g27549,g9516,g34322,g13918,g13117,I25683,g23082,g33463,g12486,g4540,g32146,g34298,g9369,g27239,g4888,g11492,g34068,g15904,g11842,g16663,g33227,g10589,I32439,g15758,I23306,g34882,I33267,g9386,g8093,g32188,g12880,g12604,g20451,g32199,g20127,g32815,I12910,g18333,g25946,g25286,g14637,g19572,g14645,g33591,g7804,I21297,g27152,I28199,g31909,g6077,g34222,g26749,g22495,g30254,g10831,g2811,g24646,g18262,g23443,g24891,g1772,g34407,g16750,g25707,g2138,g3654,g11129,g18216,g13003,g31013,I15107,g29482,g17312,g22161,g21743,g604,g15027,g32897,g30116,g26598,g34504,I11655,I17507,g24482,g1816,g29536,g26869,I29371,I25847,I24603,g7134,g21945,g26026,g8255,g7517,I15262,g33100,g28322,I18376,g30551,g34970,I29218,g11786,g859,g34751,I14623,g11047,g22647,I12712,g21950,g33916,g11306,g22304,I13968,g31169,g10873,I14956,g25400,g21752,g9291,I26195,I22785,g14659,g16127,g11930,g5343,g19345,g34288,g18401,g18348,g28677,g7777,g10960,g18356,g31941,g8146,g14387,g31782,g13031,I16917,g9761,g10760,g22127,g32291,g3380,g28266,g13634,g32628,g18631,g31919,g16285,g28680,g30445,g20382,g31256,I12468,g18542,g31372,g28035,g26629,g15050,g24322,g18160,g26969,g15130,g16586,I12902,g32475,g26936,g538,I16847,g16813,g32951,g33338,g29567,g22145,g8449,g18222,g15167,g25435,g9044,g13461,g23865,g11020,g31849,g28089,g14780,g14275,g9912,g20033,g18230,g25716,I29717,g499,g14394,g21185,g20499,g17594,g31753,I24117,g16668,g26819,g23795,I16193,g12563,g4793,I16698,g20500,I29313,g18728,g31992,g23261,g11961,g24714,g17761,g5599,I17008,g13764,g32021,g24729,g22198,g9247,I28062,g27391,g6918,I13851,g24762,g31125,g18623,I20867,g12180,g9915,g27490,g22026,g9461,g32722,g12051,I32222,g23762,g19264,g34420,I24558,g18213,g13908,g28986,g31903,g23665,g19535,g4082,g23642,g22146,I17474,g33138,g21784,g28347,g33699,g33859,g20241,I23986,g30438,g27463,g24866,g10497,g32460,g33140,g17812,g15075,g6661,g26122,g32346,g28419,g31194,I29211,g27163,g13301,g24216,g28214,g18774,g32482,g21605,g26758,g26715,g15096,I14899,g14342,g3329,g13565,g6983,g22002,g25981,I12819,g18831,g12414,g12902,g7503,g33496,g12413,g31525,g8355,g6527,g9713,g5917,g34866,g33113,g32396,g17651,g34216,I17754,g32638,g7785,g30393,g15842,I22298,g30201,g17514,g25142,g15048,g18884,g19666,g33586,g5456,g20158,g26628,g9381,g25621,g21562,g10150,g27614,g121,g26090,I18104,I25005,g22218,g18579,g9456,g16588,g9574,g18439,g1542,g24001,g513,I26670,I12483,g7202,g32723,g21386,g23645,I22899,g14376,g18719,g21140,g32776,g21974,g34457,g29656,g24576,g3798,g21737,g21329,g21962,g30984,g25010,g9413,I12538,g956,g28593,g31795,g18433,g18475,g34049,g6841,g12497,g32523,I18653,g16761,I13390,g27421,g33500,g29288,g31667,g1274,g32401,g30546,g28468,g34180,g34250,g25133,g18890,g28452,g18435,I13509,g13823,g26882,g29603,g24127,g17576,I16077,I24546,g19634,g14732,g17844,g7733,g24243,g14569,g29611,g15937,g31747,g30214,g27231,g27036,g27483,g22208,I28566,I12887,g34974,g21429,g15812,g18244,g28268,g28226,g18288,I25567,g30399,g32037,g27132,g12981,I21744,g27379,g12039,g34511,g23715,g1982,g11533,I30904,I19707,g10613,g25495,g18673,g30001,g11034,g18119,I21992,g18137,g18182,g27224,g28697,g33505,g7952,g10607,g27340,g33626,g34116,g9509,g18088,g29107,g16208,g34087,g24875,g18824,g28663,g3857,g30583,g16884,g12641,g30292,g16300,g33421,g9535,g24357,g34777,g29292,g24750,g34109,g33252,g20715,g20524,I13443,g33688,g16964,g24062,g23019,g17480,g13914,g5101,g2265,g18947,g5248,g13929,g29848,g28055,g34043,g13584,g20623,g32339,g15142,g23211,g25327,g19695,g25540,g18274,g18586,g33007,g28083,g24566,g12087,g3476,g28551,g6088,g28686,g24920,g10154,g24782,g6855,g11546,g27613,g21760,g32251,g31773,g16173,g7201,g23153,g33407,g33590,g24299,g1199,g24195,I22946,g7356,g12511,g10312,g11967,g27411,g25787,g496,g33913,g22449,g29639,g14509,g34314,g33414,g23810,g6800,g21758,g13120,g32561,g17014,g26549,g18482,g28655,g19533,g17470,g21657,I19863,g7049,g16620,g17424,g25635,I14508,g33930,g27094,g32582,I14733,g24376,g24770,g16721,g1495,g18635,g21465,g34943,g34479,g10360,g33819,g34844,g27553,g32996,g30326,g29515,g22066,g25091,g22713,g21985,g29178,g13326,g19949,g34553,g27264,I25511,g18787,g26572,g1950,I19674,g31121,g7532,g28561,g7041,g13938,g28388,g28685,g11136,g34257,I31096,g14379,g25936,I32970,g9449,I26581,g32343,I18078,g29007,g18180,g33486,g14408,g10532,g12818,g18241,g7659,g7239,g27542,g13479,g33878,g28246,g22125,g28535,g22491,g19356,g30383,g22927,g20854,g29194,g23318,g21734,g26349,g10966,g28589,g34745,g23919,I14679,g13679,g25750,g32549,g15885,g33000,g28155,g34713,g21870,g27299,g5366,g28,g16770,g33960,I13740,g18574,g28584,g4405,g12054,g27427,g31971,g22872,I24839,g20732,I13206,g32768,g21960,g19866,g8136,g24990,g34454,g25274,g10551,g20702,g34800,g20699,g17671,I18832,g4917,g8186,I15918,g10141,g28034,g15042,g31301,g12021,g24584,g17733,g13873,g28406,g27667,g33335,g24965,g4045,g26232,g29094,g25117,g20542,g15978,g26346,I23587,g14032,g25151,g29612,g20186,g13313,g18545,I33079,g1624,g9657,I24619,g6065,g17469,I30755,g291,g24973,g3731,g23203,g34574,g22874,I19818,g24123,g34650,g19952,g27310,g27966,g7791,g34581,I17557,g25988,g5961,g24093,g14540,g26945,g34857,g25565,g3929,g11755,g22330,I12205,g7633,g20373,I25115,g13069,g23858,g28314,g34334,g24070,g1687,g1710,I18662,I30760,g34378,g33974,g13142,g28329,g1792,g25299,g24368,g16030,g6589,g29291,g9739,g10905,g32390,g33024,I27529,g26976,I33140,g2827,g13020,g10828,g7040,g19784,g23519,g23903,I14289,g3759,g4999,g23296,g9492,g27250,g4864,g25892,g23165,I12123,g31803,g26337,g7436,g23856,g27101,I20385,g10216,g23945,g34184,g10755,I15717,g13852,g11294,g21404,I24067,g31578,g20129,I15212,g22644,g24607,g8399,g33250,g23402,g26683,g18264,I30998,g32954,g18113,g31472,I27524,g21777,g31820,g26304,g17595,g34342,g34413,g26389,I29245,g4922,g6275,g32598,g19354,g33965,I18460,g4621,g33343,g12076,g28604,g26279,g7802,g13951,g25753,g11444,g19474,g20909,I25028,g19660,g27837,g33695,g16305,g11969,g12794,I17276,g1748,g33701,g16076,g28451,g32981,g28428,g34207,g4572,I33279,g28682,g31237,g7308,g9732,I14671,g4486,g18311,I25612,g21127,g18689,g32272,g11182,g18259,g29754,g17506,g32351,g33931,g30212,g4287,g26700,g4430,I27381,g23489,g31966,g33290,g23355,g8477,g27121,I24482,g21931,g17122,g18742,g28617,g30613,g7470,g11658,g30018,g26400,g23339,g13675,g749,I26578,g12082,g3391,g34621,g11426,g32570,g6625,g13281,g20321,g26226,I25530,g23987,g30431,I27514,I20462,I28576,g5276,g2994,g22457,g33766,g24704,g24489,g732,g24147,g23606,g18756,g6975,g24653,g27033,g33251,g16769,g26347,g17635,g30380,g24813,g16513,I22149,g13867,I24463,g23509,g34489,g25522,g20387,g21739,g8703,g33253,g23972,g542,g18934,g14313,g29834,g22527,g4197,g24408,g25997,g24723,I26356,I20584,g15080,g25634,g20672,I22892,g24518,g30160,g22129,g10821,g33555,g9670,g29672,g21958,g34183,g33390,g34744,g9620,g13217,g13795,I21941,g10676,g20135,g18917,g14187,I15702,g18360,g11169,g24436,g24411,g32137,g13102,g26424,g24372,g10078,g15508,g33542,g13637,g33549,g18916,g28779,g24059,g32966,g17721,g13295,g14365,g24720,g32845,g9683,g31186,g23965,g13932,g22138,g34638,g29540,I12790,g17611,g18181,I29441,g24725,g33365,g9498,g22635,g8417,g20166,g27556,g23124,g27223,g15005,g27527,g13745,g32974,g31816,g30213,g8296,g19712,g27180,g34810,g11962,g25718,g6195,g33694,g15824,g2571,g28601,g28871,I22124,g30553,I31361,g101,g34267,g14091,g8880,I14271,g9880,g26804,g8181,g32889,g32171,g30566,g21287,g12946,g34024,g33161,g19788,g7927,g20087,g23352,g32392,g3325,g28631,g32680,g14385,g18121,g32826,g31970,g9,g21514,g18186,g26788,g43,g13155,g8443,g11044,g12941,g16758,g16643,g24100,g31830,I24675,g7497,g6315,g25887,I24228,I18765,g34252,g29842,g15847,g31654,g21971,g34736,g13626,g18821,g31802,g20609,g33049,I22900,g21607,g14396,g32987,g21869,g22124,g13075,I12271,g11330,g1146,g18371,I17938,g30028,g7395,g29193,g8389,g17220,g18931,I12109,g3502,g32982,g34034,g25645,g794,g5969,g28046,g12785,g24056,g33429,g21897,g12364,I25576,g17367,g28647,g24443,I21042,g7823,g29167,g8905,I24704,g21387,g12812,I15533,g24674,g23969,g2204,g32719,g6904,g25149,g19717,g12954,g32103,g25900,g29959,g8219,g34057,g28955,g28316,g29533,I15494,g28575,g24608,g27218,g31314,g26654,g7834,g20580,g27569,g16535,I23162,I12089,g34672,g30614,g25081,g32821,g33311,I16747,g9974,I18224,g25491,g27404,g13946,I14305,g25179,g9092,g2024,g32855,g24850,g26329,g979,g25385,g34759,g17680,g34515,g31279,g31226,g13493,g22546,g6995,g32867,g16532,g34508,g1592,g33492,I18882,I15052,g28108,g28418,g33437,g29073,g16667,g4443,g15089,I14069,g18303,g11280,I13548,g32226,g29890,g34187,g31483,g25118,g18785,g26939,g11235,g32252,g21352,g25906,g10185,g14571,g27634,g27503,g20076,g29118,g33589,g15711,g16684,g528,g8135,g14821,g14038,I12783,g12871,g23539,g18979,I26687,g19881,I17916,I17569,g17529,g18344,g26166,g13495,g10129,g16209,g1668,I30193,I17111,g26340,g20505,g21512,g34727,g5747,g7625,g18976,g24282,g8864,g30098,g28043,g3050,g20436,g14546,g10715,g28220,g9364,g30502,g24779,g32681,g26891,g18263,g30362,g14930,g14872,I18635,g17569,I18509,g27697,g9699,g27278,g32084,g33043,g10107,I22046,g7495,g18185,g19954,g319,g25348,g21864,g5339,g21400,g24665,g13064,g19062,g26350,g33068,g12085,g31910,I18681,g28054,g33799,g21968,I16679,I31091,g7174,g29168,g30295,g21458,g12065,g33031,g34979,g13529,g16530,g28174,g16882,g24672,g29513,g7063,g23356,g33064,I21784,g26422,g20035,g18888,g29988,g2697,g12179,g20549,g31294,I18538,g34497,g13459,g6181,g30055,g10515,g18876,g29134,g22131,g32829,g2126,g20283,g2724,g2527,I24385,g32485,g9835,g24812,g2848,I14531,g31833,g8347,g25068,g26514,g32220,g26121,g34127,I22488,g21741,g24202,g13283,g29549,g7498,g11309,g13294,g34728,g10217,I26693,g23061,g25016,g32449,g20779,g22494,g30248,g26541,I20460,g29647,I27573,g2799,g28264,g24223,g23236,g29662,g9397,g3223,g25659,g22906,g146,g24080,g19518,g11666,g22626,g12431,g25875,g29041,g34161,g23843,g29697,g4717,g33413,I18120,g29036,g18061,g29351,g24636,g14740,g13028,g18782,g33729,g31491,g26095,g7411,g1094,g9862,g28156,g28429,g16026,g27540,g18953,I31597,g1216,I15636,g18802,g23942,g18093,g23651,g8340,g29303,g30388,g32240,g31151,g26517,g13100,g23895,g33665,g32128,g14773,g2227,g23016,g8804,g18827,g14307,g34841,g25266,g15426,g16960,g29142,g28087,g8844,g19468,g14867,g33244,g23978,g16211,g16757,g21712,I17885,g28323,g22974,g11355,g4125,g30519,g34501,g9283,g24957,g34173,g21399,g23086,g25744,g34147,g33909,g24574,g24853,g27575,g8097,g34149,I28597,g26921,g31936,g15753,g27377,I16417,g14035,g34370,g28120,g3933,g11846,g34518,g32915,g23692,g27331,I23969,g31672,g1548,I12106,g29995,g3558,g12521,g34682,g26903,g23949,g23254,g34664,g17785,g13080,g27378,g7670,g9174,g14366,g17786,g18473,g24644,g23770,g23456,I12227,g27141,g17585,g34041,g20639,g9220,g19569,g18799,I28147,g23906,g9060,g32554,g32415,I29939,g20213,g14683,g13299,g28874,g34607,g28540,g34708,g25061,g27232,g24300,g27669,g27017,g25129,g14210,g7515,g17713,g19948,I13473,g18537,g15158,g22010,g8948,g714,g19528,g28553,I29363,g25849,g11894,g8119,g32041,g21927,g429,g32876,g7095,g24230,g1339,g13657,g30608,g28294,g3498,g28778,g24745,g28488,g23323,g34446,g34223,g32364,I21291,g34696,g4601,g27320,I18486,I27735,g31925,g20592,g30161,g33921,g23918,g24066,g33440,g33020,I32665,g22870,g24702,g27295,g25790,I17892,g19344,I12403,g16640,I25221,I15765,I12719,g34931,g33126,g18413,g2098,g1105,I12144,g24964,g9434,g21344,g26719,g11178,g3614,g14041,g6490,g106,g28224,g15117,g14517,g29524,g11043,g16311,g22514,I18009,g27333,g25518,g34396,g15585,I31271,g7227,g27704,g25658,g19556,g18471,g595,I12877,g29287,g5352,g12013,g22172,g32785,g29565,I31232,I25908,g25948,g29836,I26438,g13133,g31540,g6005,g11893,g28895,g9962,g26392,I12611,g24039,g1422,g582,I22918,g20204,g30998,g28180,I17609,g34589,g12125,I23919,I13401,g12284,I18600,g8643,g33056,g28917,g23682,g27999,g13063,g27595,I22331,g14678,I32797,g31297,g34542,I18233,g27616,g32369,g33037,g28132,g22300,g26898,g9467,g17602,I22872,g34911,g20494,g27678,g23031,g7553,g22339,g33266,g22904,I15782,g7697,g1252,g28390,g24510,g29326,g28109,I12728,g21902,g12358,g24136,g3827,g16180,g10612,g10603,g24394,I26049,g20698,I31186,g25723,g34605,g12244,g22342,g25296,g21810,g24397,g19366,I29263,g20575,g19575,g23754,I32994,g26853,g29141,g14092,I27718,I31061,g26544,g5623,g34505,g3538,g21825,g14014,g32558,g32087,I31853,g21050,g14169,g15066,g311,g17587,g28371,g34842,g34044,g21179,g20924,I30751,g34106,I22889,g24090,g7863,g15594,g12835,g10980,g22901,g21838,I14079,g31274,I12204,g23585,g12906,g11691,g7275,I15298,I31081,g28427,g32334,g30303,g12850,g27770,g11610,I22485,g24896,I16875,g24906,g15479,g31473,g2587,g7441,g27519,I19734,g28476,g23026,g25024,I18089,g33822,g23943,I16593,g30396,I14230,g3706,g34586,g15169,g27314,g33118,g15755,g9973,g32327,I19843,g33842,g23272,g12979,I25161,g10367,g4340,g12761,g21509,g14278,g15580,g29183,I13037,g29750,g13499,g8285,g2667,g29505,g13807,I31062,g1783,g5212,g32172,g15136,g31865,I12563,I12805,g32581,g15578,I17159,g16448,g18690,g10820,g31789,g23521,g10754,g5499,g24585,g28632,g32266,g25714,g29266,g31757,g21926,g32781,g16717,I17699,g19997,g4961,g15076,g31523,g21965,I12288,g55,g33294,g30053,g33641,g15590,g13240,g26235,g34012,g33937,g21175,g17532,g17489,g11855,g17645,g30189,g27543,I15053,g6905,g18291,g13058,g16804,g10113,g28067,g12738,g18488,g32096,g34046,g33164,g24200,g9621,g27823,g20218,g8677,g14098,g26682,g3321,g9407,g30306,g25090,g23801,g30104,g5385,g28600,g20923,g33093,g27351,g25123,g20068,g29327,g7636,g13101,g27384,g15785,g10038,g24256,g33028,g31289,I31082,g9162,I31217,g1178,g17605,g32784,g23566,g33807,g22686,g22319,g14792,g27580,g12249,g28154,g18833,g7516,g18493,g1657,g14209,g15615,g7824,g3423,g27117,g6856,g17574,g16201,g32853,g6519,g32807,g25719,g17059,g23130,g19402,g26307,I33210,g14506,I31497,g34082,g6675,g21843,g23461,I18191,g17527,g30494,g14364,I13384,I17919,g18771,g33306,g33426,g27268,g30989,g28064,I11737,g9334,g18552,g34071,g20617,g10352,g14668,g34119,g27600,g18489,g18818,g1894,I33155,g34016,g29347,g24687,g19751,g30317,g21225,g8125,g14203,g11562,g21920,g9036,g29663,g3133,g6133,I20690,I30745,g6895,I21911,g15151,g5481,g16692,g24273,g16635,g27042,g11985,g34606,I12067,g25776,I18479,g18530,g17818,g10403,g30539,g31937,g27207,g16970,g13943,g20508,g28892,I32684,g32779,I33176,I15147,g33123,g33197,g21661,g32527,g22545,g30599,g9978,g9875,g2389,g29352,g23417,g32704,g17955,g30508,I11843,g32707,g20780,I17932,g24122,g2429,I14853,I14570,g27142,g8833,g17308,g30482,g24014,g25598,g28334,g19579,g21347,g18428,g23410,g8748,g23924,g28726,g8026,g19603,g20853,g18125,g11366,g17466,g20267,g15506,g12160,g8234,g19360,I22761,g3606,g30734,g32576,g8922,g8974,g14062,g25877,g18286,g20561,g31844,g31506,g14598,g26326,I12003,I32441,g24148,g753,g9599,g8715,g15848,g4358,g34658,g32381,g4944,g14253,I14258,g4653,g34011,g27408,g1319,g7897,g14573,g16119,g11761,g23439,g6505,g9185,g28953,g24968,g25109,g33579,g29177,I15073,g20374,g4417,I18495,g14065,g4035,g18322,I20861,I29261,g20526,g12453,g23453,g14800,g31915,g29930,g30022,g19902,g34151,g28751,I32274,g27489,g26751,I20929,I15572,I24689,g26690,g9853,I13010,g26312,g33522,g28527,g12910,g31921,g34200,g25341,g28286,g30554,I31561,I31292,g14968,g8123,g30130,g16616,g20184,I25399,g27821,g32478,g8431,g10556,g22447,I25845,g34684,I31272,g1878,g10808,I13730,g5495,g4119,I21162,I22502,I32871,g2878,g34758,g20629,g18252,g21277,g12875,g8059,I20035,g19372,g9433,g25517,g8666,g25758,g8898,g15749,g26901,g12432,g26077,g33357,g29331,g22763,g10351,g17498,g19862,g32419,g33433,g21332,I22725,g12951,g34384,g13009,g1233,g12844,g28262,I17495,g21820,g24799,g20852,g33232,I20744,I16762,g34524,I14427,g18229,g23172,g31755,g28548,g31479,g19761,g30611,g14205,g17062,g28819,g24025,g12437,I17228,g20710,g29282,g16291,g10862,g5228,g32627,g2152,g33798,I22973,g29369,g17643,g22400,g27431,g24528,g31287,g9688,g17366,g21669,g10353,g17707,g33052,g32289,g8818,g29179,g10288,g24157,g24186,g21830,I12855,g23009,g27730,g23248,I14749,g15572,I14789,I25146,g2070,g27238,g18415,g22756,g22123,g5176,I16371,g25680,g22919,g16224,g6978,g31323,g7514,I31201,g32828,g4812,g15732,g31138,g30069,g27977,g20452,g16200,g8287,g32787,g12041,g25158,g33038,g5905,I14517,g27263,g15701,I33258,I32116,g32385,g34689,g31223,g33379,I21246,g34604,I16526,g11479,I18709,g16197,g32743,g19470,g33902,g31468,g24680,g4633,g26987,g30374,g6163,g28143,g15106,g32287,g26021,g14418,g33516,g29306,g1277,g27492,I20221,g4616,g20624,g27692,g29298,g19905,g19637,g10890,g21049,g13125,g25507,I13403,g30458,g31960,g30310,g19691,g16745,I29582,g17175,I13708,g22054,g21296,I30686,I13452,g21283,g1266,g30443,g21430,g32468,g32484,g25676,g25783,g29176,I27777,g22005,g25908,g27544,g34376,g33457,g15911,g28977,g30467,I31126,g23257,g31509,I18323,g25031,g22166,g27183,I16468,g32699,g11149,g24369,g31961,g32278,g29365,g23578,g28405,g13638,g18811,g25453,g29377,I22967,I19345,g12730,g18753,g32961,g617,g31496,g25804,g12024,g28204,g12411,g29756,g21757,I12026,g30372,g18596,g33089,g34263,g15679,g23062,g12148,g34089,g21655,I15070,g32608,g9637,g10632,g31774,g9200,g25558,g33711,g28380,g28906,g25691,g27301,g29049,g23282,g18681,g3831,g15881,g8770,g34079,g29938,g16579,g32652,g11166,g15574,g30101,g31322,g30540,g32913,I32639,g25451,g34625,g3712,g27981,I12415,g23800,g30670,g8172,g6816,I22865,g20389,g22030,g2988,g9931,g13806,g18877,g27236,I24530,I33161,g18177,g34102,g16766,g22665,g6523,g34428,g21959,g33904,g14024,g14031,g31767,g2775,g21681,g27261,g8933,g19430,g18647,g25720,I12749,I15334,g29748,g33836,g28256,g12614,g18984,g18997,g27213,g27302,g23653,g27352,g30415,g26348,g27518,g33657,g11702,g20131,g28069,g25077,g18393,g10961,g32446,g24323,g25814,g29759,g28284,g25273,g33693,g29071,g28534,I32820,I16741,g34945,g10720,I12997,g23400,I22717,g27964,g24114,g25230,g30219,g20041,g25601,g9543,g32814,g24929,g19914,g12332,g25037,g31285,g19602,g9999,I15175,g24375,g18494,g24339,g24040,g33006,g31300,g23824,g19773,g3466,g23266,g28856,g30401,g25668,g17138,g11931,g23384,g21222,g14696,g28833,g33033,g6459,g29915,g26838,g21360,g25871,g30500,I14212,I13729,g33565,g26821,g27683,g7267,g16196,g34377,g19753,g3021,g21702,g28166,g22648,g11397,g17705,g23025,g10370,g27511,I22289,g34667,I21734,g11415,I29304,g25013,I14839,g23719,g9229,g24575,g13830,g31765,g26632,g29916,g12295,g21606,g6986,g26249,g3274,g4743,g30185,g15913,g17363,g32793,g32852,I11896,g27698,g33481,g32824,g32047,g34561,I22886,g28716,g21947,g26084,I13182,g2384,g10581,g23056,g34083,I31854,g28949,g9253,g27086,g12768,g30275,g30429,g34329,g19071,g32404,g12232,g29921,g464,g18640,I29278,g26179,g671,g16742,g23197,g16658,g25882,g27727,g33148,g25309,I24710,g18295,g29294,g2533,g32294,g31818,g32033,g1075,g8160,g3763,g28248,g29342,g24410,g10541,g20538,g1844,g23112,I18221,g1193,g20661,g24628,g27486,g27272,g16053,g13967,g30428,g11148,g33963,I32878,g25926,g12077,g32899,g26258,g32805,g23484,g157,g7586,g12955,I15929,g28217,g19449,g22757,g23195,g32261,I31302,g3025,g26930,I31236,g23028,I29182,g34545,g18599,g30143,g11867,g20240,g27597,g13594,g6390,g9598,g27177,g24726,I23300,g10384,g25050,g33717,I30735,g9965,g26604,g5983,g6263,I32950,g32908,I14647,g19210,g8497,g5320,g23382,g26365,g29722,g5216,g24073,g4216,g29996,g21054,g9690,g3813,g11935,g25665,g23524,g29514,g3247,g33884,g9015,g13901,g26694,g25168,g28727,g32095,g34716,g30561,g11832,g18629,I15932,g22492,g24139,g7591,g29149,g7693,g12460,g8284,I30995,g2819,g11429,I24549,g32545,I15088,I31838,g28579,I31197,g25700,g21909,g21715,g25941,g26096,g25993,g25380,g33569,g6819,g33373,g25136,g25224,g32946,g25619,g19519,g9551,g22859,g27552,g4232,g27128,g24324,g13573,g34794,g11413,g29772,g30490,g6322,g2495,g18875,g21999,g15740,g32683,g23840,g14977,g34316,g28245,g30299,g2837,g19355,g26130,g28199,g5112,g3065,g25027,I27391,g32928,g10377,g27592,g18112,g11441,g9316,g13324,g929,g13504,g24497,g19781,I13705,g21919,I27388,g22094,g24945,g22111,g32161,g33102,g33731,I32687,g33010,g34598,g8879,I24579,g7064,g15049,g20089,g11976,g7917,g24864,g29497,g10710,g20051,g33594,g23383,g34394,g15480,g33716,g13248,g16694,g10357,g24117,g21900,g21954,g28578,g6251,g20679,g25046,I15307,g30043,g20558,g10727,g28654,g17683,g34148,g10699,g26885,g32562,g10498,g32623,g26171,g13620,g11496,g11427,I17668,g34637,g24897,g29849,I12837,g23403,g22136,g26886,g7235,g27413,g29343,g6956,I29185,g16027,I17542,g27827,g13945,g32394,g16186,g27765,g29592,g22585,g32502,g23901,g28240,g14564,g3115,I14584,g1760,g3347,g6789,g13413,g22022,g24149,g28559,g22594,g20766,g27682,g25155,I22576,I17772,g358,g29873,g24257,g14309,g24548,g31892,g16531,g6987,g20053,g28363,g22013,g15631,g34474,g32602,g15052,g13140,g27691,g9645,g28786,I31086,g15573,g32245,g3010,g3303,I29262,g15751,I23309,I20499,g13524,g19383,I15123,g9914,g23564,I32788,g29198,g8397,g30267,I29286,g12009,g34421,I25869,g7116,g19688,g18567,g23956,g4674,g33472,g28880,I19661,g7301,g22645,g24581,g21866,g22149,g699,g24985,g25057,g31267,g17156,g19063,g10140,I31593,I32089,g19999,g26910,g1926,g15152,I13723,g25572,g28695,g13040,I17101,I13862,g490,g17644,g30000,g32664,g31518,g9104,g11590,g29485,g33261,I14576,g9694,g22105,g27690,g30309,g25199,g21994,g27234,g32358,g25169,g30035,g30927,I13374,g29385,g7601,g9820,g63,g32948,I16613,g25706,g28588,g17814,g13507,g10555,g21024,g33572,g8971,g2719,g6927,g8997,g8346,g2351,g28404,g14731,g16623,g29622,I32648,g28519,g20327,I26649,g13542,g5845,g14913,g31749,I18452,g24988,g13410,g32528,g33318,g34304,g12224,g7763,g22089,g11317,g13570,I15195,g19559,g18591,g12805,g21768,g33621,g31670,g19979,g10396,g21921,g802,g8566,g27104,g34410,g22903,g34358,g23459,g5517,g27994,g13016,I13031,g28574,g3873,g13278,g4722,g14544,I24462,g28857,g21929,g33289,g26681,g34718,g30017,g13462,g8134,g21297,g5857,g34978,g30260,g24012,g22857,g32230,g8131,g19067,g31801,g24113,I13565,g26893,g15811,g13311,g32130,g25244,g33823,g11534,g23245,g11344,g29581,g13014,g10382,g16592,g33399,g8058,g32831,g24352,g32967,g32042,g287,I15626,g33316,g7716,g31783,I20187,g29538,g19549,g22715,g16264,g32397,g222,g34480,g33430,g3787,g7293,g25211,g26293,g29598,g4931,g16322,g1768,g29569,g28184,g18652,I13937,I12799,g31292,g18277,g34166,g34639,g10738,g17570,g28938,g19539,g17589,g12108,g18683,I17460,I28567,g15060,g22358,g13048,g17307,g21899,g24124,g25708,g15741,g21721,g1087,g21273,g30242,g24209,g25938,g29337,g7315,g34862,g23695,g28281,g29001,I32119,g5283,g10379,I18885,I18740,g12883,I26070,g33109,g29157,g18500,g14730,g26386,I13852,g29788,g11450,g22142,g31706,g7162,g33944,g24272,g28557,g30132,g34924,g28987,g11216,g32132,g14406,I30400,I31817,g26914,I12401,g20644,g18440,g8479,g4165,g18470,g21349,g25470,g33892,g1736,g33094,g19546,g26131,g22217,g6191,I33300,I31166,I21918,I13236,g16652,I17154,g28458,g33287,g18667,g30573,g30434,g5156,g31653,g11978,g1582,g13436,g30365,g28402,g16307,g8721,g31213,g22305,g25699,g31750,g23812,g5689,g25764,g28391,g6755,g24664,g20611,g32827,g417,g30261,g23554,g29507,I25369,g3089,g34737,g9298,g11116,g31268,g32129,I17118,I32696,g29636,g31327,g33698,g875,g21466,g13432,g33692,g7410,g18350,g34503,I20447,g14008,g29362,g12378,g23559,g34305,I29277,g16634,g23781,g34069,g28259,g14126,g18162,g29046,g24751,g23297,g7879,I31137,g31471,g21851,I31482,g27337,g13034,g24577,I13581,g23871,g24893,I14589,g17573,g14754,g22984,g2629,g24842,g25837,g20640,g2008,g25747,g24386,g27822,g16518,g14193,g22072,g34088,g10060,g24326,g5220,g1691,g28387,g29899,g15134,g24424,g18582,g13855,g18457,g28526,g12114,g554,g25683,g24242,g15756,g34381,g18730,g25459,g30050,g5452,g20619,g30232,g30935,g21380,g29563,g23427,g8526,g30237,g33174,g2380,g28554,g10881,g24143,g27392,g3680,g6199,I21210,I16492,g21885,g19428,I21838,g23999,g33743,I18858,g19675,g10573,I33288,g25536,g23277,g34724,g32772,g23750,I32479,g24086,g34596,g11889,g28541,g31912,I31974,g31499,g16525,g17774,g19679,g7953,g25710,I31196,I25786,g21340,g26657,g25331,g12856,g34280,g19746,g30218,g9213,g7597,g18345,g25943,g14362,g14889,g12297,g33817,g34778,g10827,g11123,g32184,g30151,g22709,I11785,I18762,g7595,g12153,g24684,g18324,g29240,g58,g16720,g11325,g27574,g24682,g31477,I16217,g18250,g13968,g26052,g16739,g29187,g26855,g24765,g9050,I15837,g28748,g25615,g19267,g31118,g16306,g1724,g33917,I32309,g24987,g18397,I17098,g25566,g34533,g28699,g34903,g24211,g20655,I22128,g20052,g11276,g34977,g27541,g18231,g29925,g25603,g26083,g32939,I32681,g18403,g33981,I16438,I22819,I22096,g23550,I24685,g30590,g10402,g32578,g10415,g26950,g22169,g16282,I32062,g24659,g5933,g28100,g29267,g34136,g34259,g2504,g20662,g21422,g26857,g17508,g33515,g14761,g26849,g27570,g24095,g18269,g19596,g32669,g12211,g2028,g10358,g33119,I24474,g8906,g4521,g6311,g10371,g16956,g19553,g22592,g25465,g28671,g4122,g27461,g10033,g27984,g34369,I18868,g8938,g24797,g34992,g22530,g20215,g32024,g15120,g17504,g16617,g34465,I15238,g28516,g30996,g13103,g17650,g29981,g25021,g7685,g19557,g28721,g21813,g32740,I16610,g11543,g29334,g13394,g20546,g11115,g6867,g4291,g23514,I22792,g17495,g23931,g30093,g4239,g23953,g29975,I13510,g18615,I21013,g33805,g19681,g21764,g26299,g22591,g25832,g33048,I20321,g11371,I31604,g19739,g29188,g14177,g17057,g7451,g29922,g32106,g32657,g30468,g32880,g27927,g8163,g17135,g20112,g24249,g26971,I11697,g15817,g24290,g14497,g29537,g11356,g14453,I13731,g20054,g6941,g25749,g24425,g25821,g19564,g34663,g31281,g21819,g31015,g34153,g21411,g26145,g9014,I31041,I14818,g17015,g28453,g30531,g25937,g18688,g28573,g28219,g32557,g30217,g29775,g3072,I23918,g25439,I33041,g411,g11473,g13708,g13667,g28746,g22839,g18236,I12030,g13958,g33645,g23222,I13672,I28014,I21288,g18150,g17772,g5619,g3454,g15159,I31528,g16871,g26359,I29438,g12377,g34506,g34750,I15030,g6839,g49,I16401,g27245,g31927,g2583,g34653,g32778,g457,g25886,g31141,g14069,g31842,g26208,g12760,g13604,g26648,g27339,g28273,g14257,g34468,g18136,g24677,g33352,g12115,g16969,g20529,g24398,g17192,g26092,g10967,g3191,I32988,g28530,g17817,I20388,g32458,I18143,g33175,I12117,g32341,g8685,g15345,g26213,g22540,g12581,g19790,I12176,g19417,g18733,I13749,g3965,g32283,g32595,g19439,g15809,g33088,g17588,g9951,I26584,g8354,g24060,g8330,g20533,g26209,g4027,g26207,I14169,g17662,g25595,g3396,g29281,g7487,g28270,g33714,g18431,g24340,g33577,g2771,g22899,I29002,g1442,g33653,g25248,g34826,g25644,I30399,g5976,g19720,g9333,g22498,I22327,g32082,g7442,g19469,g27833,g29548,g30135,I14866,g405,g29268,g26020,g10916,g31219,g17479,g11952,g34262,I18385,I25613,g29871,I21002,g26176,g10158,g27664,g8774,g12099,g9864,g32474,g26358,g13087,I15121,g22838,I31161,g22905,g18469,g12293,I18313,g24266,g32512,g18558,I17374,I18571,g23324,g33388,g32522,g27359,g32200,g25909,I17416,g18935,I13094,I11623,g8297,g18975,g26287,I24527,g18625,g30062,g33443,g15820,g29152,g18174,g29650,g18524,g24764,g21350,I13360,g14448,g13997,g18664,g22112,g18122,g18157,g33485,I12850,g8584,g12967,g21978,g20114,g7738,g18320,g13887,g27538,g11036,I32352,g34717,g31867,g26257,g23842,g34085,g3139,g29607,g29679,g25131,g26089,g12900,g15121,I21294,g33125,g20608,g12116,g34382,g27313,g32514,I33134,g16596,g11949,I18304,I32284,g23848,I22512,g34864,g22228,I15732,g11875,g11910,I14991,g11652,g30558,g11374,g23687,g32796,g18358,g26270,I20895,g28477,g30915,g7611,g6848,I31056,g31067,g7361,I33152,g16613,g14861,g34935,g18808,g23416,g14664,g26160,g24144,g25163,g7998,g28586,g34300,g34047,g27237,g8806,I21930,g33876,g17790,g11394,g3969,g25371,g14415,g34139,I17461,g34973,g34140,g18974,g13239,g25216,g27586,I11716,g15810,g25616,g24197,g30342,g21910,g11292,g15706,g3470,g29271,I13718,I32470,g29153,g24320,g21326,g21923,g33625,g18144,g12053,g25140,g26292,g23335,g23015,g13083,g1036,g34572,g19352,g23337,g9340,g22318,g2255,g17392,g24846,g33416,g14918,g22019,g14034,g18779,g6850,I13857,I24051,g32756,g24944,g24792,g19540,g16424,g19874,g24279,g18272,g2831,g25101,g29032,g3401,g3554,g7219,g21700,g30117,g6917,g4742,g28903,g32169,g18330,g19489,g12239,g18898,g14321,I21300,g1811,g884,g27598,g26362,g12023,g26631,g19650,g23047,I14276,g32931,g33240,g17194,g17473,g13897,g25979,g30182,g33956,g23276,g9295,g12937,g17091,g26686,g29909,g11205,g31944,g504,g29642,g471,g12841,g4108,I14734,I18825,g13512,g34048,g17684,g22989,g33608,g16324,g11244,g15851,g32260,g11491,g27736,I26296,g11143,g4498,I23970,g28040,I31820,g25389,g102,I28185,g28544,g16313,I29225,g18234,g23027,g34363,g15745,g19500,g22856,g32728,g952,g33286,I15167,I18310,g33669,g26127,g11519,g14712,g18130,g22181,g32515,g33968,g24640,g34091,g12187,g34578,g24858,g29914,g19374,g24255,g18734,g18654,g19655,g4129,I26799,I18248,g29911,I20542,g28621,g24042,g9600,g26864,I17723,g32513,g24555,g32518,g28672,I22683,g6838,g30550,g21467,g20773,g21936,g27401,g26673,g30262,g7349,g18518,g12152,g19451,g27118,I14663,g16610,g32941,g19276,g12245,g30491,g21783,g16223,g24133,I14171,g29488,g20577,g31896,g18637,g12540,g25181,I17442,g26813,g29687,I18265,g31003,g34340,g23570,g30207,g1141,g28326,g13736,g33271,g29989,g14215,g2729,g28348,g30302,g21205,g27882,g34251,I21969,I27561,g12026,g29128,g25772,g22057,g34105,g14677,g33234,g29376,g24950,g10036,g8478,g5448,g24055,I31067,g4754,g16024,g33313,g26324,g26212,I18682,g29290,I12746,I17488,g22103,I25534,g3029,g28247,g2453,g18365,I17496,g23457,g767,g23290,g12088,g32993,g32437,g9354,g15786,I16606,g12233,g14631,g7192,g14136,g23347,g15783,g11398,g8405,I16328,g19908,g21653,g23474,I22419,g27227,g34525,g29908,I25219,g29874,I31352,g18678,g370,g8,g18618,g27717,g1902,g33321,g13108,I21067,I29337,g4297,g33715,g74,g30052,g14446,g1756,g4501,g32526,g24711,g26335,g5297,g10564,g23430,g23545,g15804,g28301,g8796,g8903,g33067,g31967,g34952,I24033,g19589,I31844,g33640,g29006,g23520,g27187,g16606,g24476,g21854,g14191,g9582,g27389,g13137,g19407,g19853,g23657,g27368,g19676,g27300,g11608,g29653,g25643,g19741,I18117,g30577,I24582,g23512,g28442,g34772,g32584,g27267,g29379,I22937,g33431,g25210,g23711,g23059,g904,g5727,g30930,g11591,g14367,g22900,g14434,g33277,g34278,g32290,g25697,g20169,g25480,g29753,g22075,g18201,g21939,g33374,g26609,g18265,g21059,g15069,g29910,g13478,g14776,g23560,g10398,g4222,g25048,I16639,I31012,g28044,g10829,g10123,I20937,g26943,g3582,g12838,g7374,g26874,g29629,g32919,g3143,g24550,g31467,I15193,g6810,g20979,I18408,g28861,g17769,g32113,g23572,g33893,I13566,g30120,g31148,g14226,g3953,I18051,g32147,I26644,g7502,g26805,g28211,g21863,g25954,g29960,g34647,g31225,g24234,g20201,I19813,g30272,g26363,g24077,g20025,g11011,g8091,g29880,g29130,g24395,I17873,g111,I31296,g33957,g6120,g34397,g45,g31260,g28073,g23776,g4188,g19685,g30041,g32425,g12345,I11892,g33159,g31007,g9891,g21468,g16512,g27179,g14767,g24579,g28205,g21138,g13091,I14687,g21913,g12207,g28931,g29242,g33982,g29503,g26519,I31356,g23954,g13025,I32364,g34004,g6972,g12287,g29600,I17626,g30544,g29539,g15833,g6682,g29322,g34430,I28419,g16584,g21433,g28071,g8057,g28542,I16629,g33761,g31315,g11170,g9506,g34797,g18547,I12935,g18337,g7812,g24807,g17725,g1620,I22000,g22216,g17292,I21006,I21769,g24602,g19713,g18314,g33568,g18581,I32476,g23878,g8165,g29121,g14183,g20060,g25995,I12841,g33796,g7026,g33680,g7581,g21300,g12872,g10177,g29710,g33065,g18887,g26625,g24244,g25005,g30343,g1964,g16732,g19493,g21303,g22448,g27555,g32622,g33811,g4375,I31555,g22332,g21604,g13974,g22116,g27393,I18252,g1430,g33691,I29279,g30081,g22711,I20355,g21841,g28287,g33371,g32691,g27445,g28724,g11028,g29984,g645,g28531,g5742,g2079,g24065,g22862,g32556,g26858,I11820,g17637,g20918,g24193,g14727,g27481,I23917,g25736,g32620,g33409,g8713,g11911,g31498,g18988,g21193,g19490,g7684,g18775,g34066,g29626,g25947,g8654,g18293,g27386,I17131,g31494,I23118,g34403,g6870,g18425,g18709,g22942,g33370,I33218,g34389,g21811,I16476,g6565,g11490,g34094,g15729,g3835,g31259,g1988,g29798,g3522,g14149,g23568,g5331,g18907,g11869,g23046,g25008,g19916,g34070,I18063,g21944,I27364,g5313,g20630,g33958,I19927,g22754,g30106,g12879,g19872,g25561,g18598,g15876,g14447,g34137,g10093,g482,g32604,g32844,g25904,g1978,g22095,g14079,g9439,g30545,g31014,g23087,g28523,g32107,g31484,I20203,I13499,g33074,g16309,g34616,g18496,I31002,g27526,g14425,g20776,I26700,g33297,g26938,I32757,g30485,g32509,I32938,g17615,g28117,I23680,g18292,g24698,g32347,g25963,g31751,g31840,g7673,g7418,g13023,g22679,g29617,g13258,g12371,I14862,g18939,I26378,g29012,I26334,g22215,g8388,g30367,g785,g8500,g18334,g22031,g9095,g4023,g13799,g32201,g16730,I12580,g29859,g15822,g21678,I22830,g23345,g33326,g20059,g13883,g24666,g11155,g33670,g23385,g25147,g8890,g1616,g18770,g13861,I15166,g30245,g21972,I29579,g14587,g34130,I17819,I32202,g24474,g976,g13273,g28812,I19487,I30766,g34768,g21833,g28611,g17820,g34331,g18561,g12483,g21767,g26865,g22406,g1061,g23963,g8462,g9662,g23698,g31814,g10203,g12318,g10204,g12081,g10430,I16129,g27825,g3457,g12837,g19755,g15149,I23963,g25528,I18627,g16052,g18169,g10112,g24399,g24011,g5180,g33541,g31526,g3317,g29660,g27028,g26824,g14639,g33620,g27426,g11959,g18143,g22450,g10178,I32074,g4372,g13044,g17418,g8056,g17657,g4434,g12865,g24409,g24716,g18281,g8928,g11200,g13882,g18248,g34671,g22200,g22055,g26297,g31775,g3976,I28336,g8075,g12443,g1798,I26667,g11469,g13527,g18680,g32223,g8728,g7437,g34215,g28471,I26439,g24421,g24111,g33581,g13062,g24384,I30055,g19734,I22866,g34022,g17119,g11134,I33137,g21785,g890,I31973,g18390,g27139,g1345,g14609,g14072,g29384,I17964,I31650,g33929,g24071,g18948,g32409,I15677,g30082,g13210,g7380,g20658,I16168,g18557,g16304,g25669,g14413,g18298,g12471,g7223,g25755,g9749,g29005,g17591,g31769,g25630,g9485,g16608,g5062,g9905,g27341,g11576,g32152,I21792,g12369,g15794,I31341,g20170,g16242,I12203,g26711,g18342,I31237,g24096,I23998,g21898,g16872,I21977,g1579,g8606,g16205,g20707,g7072,g9740,g15733,g14791,g21766,g27212,g6971,g32612,g30078,g8316,g31790,g34714,g24540,g30925,g28186,g17157,g32340,g24975,g29711,g28431,g31899,g20590,g32843,g14064,g31823,g27353,g6605,g26737,g22751,I20781,I29447,g10157,g21840,I26337,g19365,I14964,g19730,g9585,g24416,g27733,g7913,g12899,g18674,g29854,g29870,g15079,g10019,g3040,I16102,g19588,g32944,g31959,g28633,g25531,g20733,g16727,I29894,g27330,I13334,g12111,g14974,g10706,I22240,g14422,g25212,g18722,g32938,g23351,g33101,g18882,g34330,g32783,g32418,g3566,g21860,I23390,g30495,g34734,I17198,g12036,g10657,g6836,g31890,g30058,g31707,g33278,I15105,g13973,I31051,I33044,g28223,g17128,g25047,g28074,g7885,g5808,g29325,g8659,g34912,g23349,g13712,g31299,g15073,g28634,g26357,g17225,g925,I27518,g25426,g32008,g33615,g25218,g17420,g8572,I11801,g7475,g5685,g24129,I31116,g27768,g7073,I12151,g31766,g27992,g25062,g23477,g32374,g13698,g6486,I31032,I16010,g25732,g32234,g15131,g5595,g21654,g14444,g34576,g20548,g15126,I32594,g24427,g32181,g33727,I24089,g17413,I11992,I17976,g10921,g14583,g34712,g31987,g15858,g23820,g20917,g22488,g32577,g22152,g30279,g27097,g24788,g20066,g33953,g1041,g32892,g23675,g13892,g19789,g25137,g13569,g16488,g12874,g21348,g14433,g28750,g11708,g29633,g728,g31132,g30356,g17415,g26381,I25606,g34405,g28362,g14306,g1124,g29256,g29333,g5941,g29192,g32682,g21056,g9083,g34258,g29861,g25154,g30918,g18503,I32186,g4104,g21338,g32563,g13501,g8343,g22311,g25705,g28009,g31021,g15710,g20172,g22908,g4264,g32377,I26093,g19696,g28595,g29067,g30150,g30231,g34540,g16244,g20433,g13969,g22007,g32158,g18339,g11545,g18691,g29868,g17477,g27989,g32048,g32177,g28200,g14061,g11018,g20645,g2004,g30991,g12124,g29604,g33054,I11826,g22850,g32673,g10404,g32926,g24276,I31724,g34702,g32517,g18317,g32949,g26780,g28923,I16455,I19796,g29172,g7521,g17217,g19635,g34656,g10152,g34993,g12915,I24434,g25317,g33841,I14644,g28659,g27037,g7109,g10114,g30349,g30313,g18437,g33818,g22710,g29498,g17689,I23312,g27982,g34934,g15821,I33037,g34681,I31182,g28930,g13631,I12075,g11428,g25729,g27092,g21699,g26487,g29230,g28981,g14797,g23567,I24003,g29783,g25085,I26393,g8506,g10608,g29108,g23340,g11865,g29481,g17136,g32519,g34731,g3372,g21682,g34740,g17321,g12418,g26881,g26736,g32811,g19429,I16150,g23940,g9839,g32318,g19530,g16897,g34286,g16171,g9518,g31668,g33870,g29277,g10198,g16614,g11939,g31792,g14315,g22684,g17530,I31859,g33432,I14249,g11697,g28448,g18940,g12830,g12744,g9863,g29131,g22638,I11691,g25195,g3598,g14965,g18399,g16538,I28390,g34372,g24329,g10083,g31924,g34412,g23699,g32303,g11405,g25153,I23375,g34399,g28717,g19798,I12654,g33385,g20998,g27662,g10841,g27051,g15968,g33441,g28208,g16706,g22177,g32361,I23330,g33907,g13051,g21859,g27356,g5913,g15864,g9824,g33861,g3727,g33903,g23363,I23378,I14836,g5033,I19762,g843,g34030,g23935,g15114,g21037,g11621,g16699,g34053,g17430,g17302,g23496,g2823,g32348,I13464,g24137,g31609,g23875,g6831,g13662,g32363,g28935,g8407,g18804,I28162,g8561,g872,g13484,g28318,g24995,g18376,g20650,g9321,g7650,g14489,I31042,g21190,g21345,I30756,g30528,g17754,I16246,g32873,g15750,g8690,I11864,g31127,g19361,g33584,I32659,g26284,g14384,g23425,g19769,g19915,I13889,g33139,g19733,g28292,g7423,g29487,g29014,g29707,g28850,g7876,g18128,g3440,g16632,g34587,g15133,g32355,g31303,g27277,g8509,g32921,g29997,g32989,g31906,g25247,g12461,g33015,g16738,g33265,g33260,I12096,g27956,g14021,g14330,I28002,I11809,g13605,g6555,g8612,g21751,g14682,I22801,g32031,g34893,g24822,g18228,g18950,g29295,g34565,g9927,g23232,I23333,g30304,g21705,g10372,g16194,g28823,g7023,g12922,g32932,g1135,g25731,g19743,g28291,g24432,g22226,g25754,I27368,g13038,g18548,g9590,g10531,g23058,I18788,g19359,g16431,g23944,g20265,I13463,g24019,g13896,g18307,I32192,g32678,g25975,g33115,g25485,g32643,g153,g10816,I29296,g24277,g15084,g22083,g31781,g24108,g23526,g24437,g32038,g16475,g21793,g25228,I26309,g32799,g10222,g27208,g10761,I18555,I31007,g9970,g32690,g28439,g6629,g18767,g32162,g28234,g9443,g27429,I24054,I18148,g27584,g18304,g20504,g12817,g3983,I14330,g20229,g24296,g22641,g29366,g14148,g15570,g30556,g29476,g27547,g15099,g32538,g33582,g3106,g16930,g21865,g27115,g18807,g21462,g33685,g8505,g17520,g14915,I18293,g30525,g19074,g23582,g23529,g18519,g25549,g4467,g18707,g9681,g30541,g32968,g32803,g7462,g25297,g22929,g22524,g667,g4709,g32413,g10389,I29271,g13555,g10902,g19492,g25742,g33970,g25950,g9693,g32597,g34008,g17816,g10869,g24673,g20216,I17763,g2841,g5462,g32508,g32312,g10857,g21755,g14848,g2472,g34312,g24769,g6561,g30441,g13093,g4561,g23055,g661,g20102,g17571,g3618,g24351,g6958,g14539,g21922,g18796,g18790,g6657,g27649,g29864,g22456,g31321,g32635,g30452,g33924,g14739,g34220,g26917,g23289,g19499,g12308,g24254,g22148,g18140,g6845,g24289,g24627,I14428,g27962,g28973,g13046,g23678,g28918,g15856,g28426,g31754,g26102,g14320,g33723,g32127,g28283,I33050,g24588,g32344,I31770,g31286,g6049,g17488,g4975,g18257,I31317,I12372,g7857,g26693,g27820,g12976,g18129,g31881,g9916,g22884,g25678,g34366,I18909,I18449,g10939,g32520,g29757,g13994,I12262,g15077,g990,g24629,I16778,g12858,g22303,g16726,g6058,g23823,g28725,g22168,g837,g34872,g18459,g21662,g17481,I31227,g10759,g34078,g17676,g23381,g27774,g939,g32590,g19409,g27206,g21907,g27382,g18508,I15667,I16651,g34001,g21295,I31466,g7870,g8647,g33795,g24053,g10707,g6829,g26080,g6365,g3419,g24366,g7648,g25739,g32115,I18579,g20242,g24359,g34697,g24438,g22021,g28818,g25122,g28253,g18402,g33833,g32205,g3917,I33285,g32960,g33339,g34386,g26959,g32888,g26181,g20680,g31806,g8539,g18302,g29785,I12097,g25743,g11721,g21889,g33707,g27161,g4446,g13325,g21417,I19719,g25746,g10035,g16044,g11914,g11940,g28730,g26086,g29531,g32752,g17326,g27433,g20671,g27506,g25978,I16724,g10856,g16320,g6719,g4821,g22957,g7898,g34400,g8038,I17970,g6148,g20274,g12716,g26852,g8655,g11027,g4049,g3288,g23005,g6411,g32755,g29480,g32692,g22331,g20391,g28107,g23920,g15703,g13541,I13892,g703,g27666,g25258,g29855,I33264,g30454,I21993,g30032,g26195,g30436,g26267,I16538,g25534,I22880,g34559,g30255,g14832,g25178,g7443,g12889,g30246,I16660,I13383,g20603,g9685,g23941,g34531,g21036,g23768,g5611,g33744,g24041,g27148,g19951,g827,g32594,g34711,g33570,g30235,g34120,g22928,g25544,I15087,g18520,g30318,g18926,g27269,g30316,g23051,g18589,g23611,g19369,g11509,g31962,g31770,g29251,g20501,I18609,g25594,g14054,g33943,g14898,g5008,g25187,g25831,g25576,g28303,g27294,I21776,g21670,g33914,g2130,g12711,g3080,g8241,g30183,g8085,g14419,g34470,g15055,I18839,I13391,g10223,g34006,g5002,g25838,g20276,g19274,g22985,g11547,g21827,g24686,g28637,I20222,g5445,g31669,g29381,g17416,g25526,g12012,g18341,g33411,g23828,g33635,g3961,g28430,g31832,g10000,g22189,g29035,g33451,g24991,g19525,g34444,g21805,g24747,g25102,g30131,g14529,g21658,g29258,g79,g30607,I15213,I12470,g32812,g34090,g13927,g6346,g16636,g33377,I18647,g22316,g6767,g24706,g30019,g13081,g33933,g7028,g23354,g34032,g21953,g15011,I17747,g17507,g24192,g30824,g20163,I18803,g16520,g5268,g18716,g14723,g23662,g7696,g13821,g12123,g24213,g29998,g34013,g29590,g24358,g23714,g24388,g32371,g16923,g25438,g34890,g33391,g34196,g23392,g18636,g22832,g18577,I32550,g32616,g12836,g12101,g24471,g33176,I20495,g8183,g25208,g32998,g33830,I31351,g16687,I31076,g18714,I12893,g2217,g11861,g25959,I15250,g20164,g10502,g19444,g21934,I18060,g34035,I25356,g2153,g31761,I16143,I13352,I18752,g9332,g30462,I18700,g15021,g16669,g12145,I16120,g31068,I31331,g22120,g8519,g15061,g24228,g13809,g34855,I15942,g11884,I21285,g27491,g9018,g28090,I14206,g6846,I14198,I18795,g2980,g10003,g29986,g27738,I11746,g8286,g34086,g11923,g30287,g18421,g33091,g10897,I22444,I31864,g25833,g32800,g18643,g24500,g34067,g18828,g33467,g17753,g17740,g4593,g27262,g27975,g32914,g33538,g8925,g31247,g20203,g13076,g14586,g31527,g14771,I32240,g25951,g2315,g34526,g26300,g4135,I29248,g21790,g34539,g31993,g12894,g5115,g30538,g21906,g14640,g27348,g907,g24787,g34325,g8967,I32607,g32990,g28514,g34447,g29522,g22623,g27133,I26095,g24246,g23060,g34563,I13715,g9186,g33614,g10877,I17491,g31854,g34341,g34661,I13166,g14178,g18657,g34274,I23354,g20320,g18952,g27209,I30261,I24679,g19617,g18398,I28174,g32119,I14730,g18794,I13109,g28367,g23336,g15087,g12464,g10830,g18200,g24976,g1,g34735,I18138,g7251,g168,g22922,g34858,g21723,g294,g4172,g23725,I31256,g5428,g20180,g23215,g27504,g24722,g29474,g17198,g23946,g15085,g25186,g29283,I15773,g3125,g25781,g23787,g24191,g18699,g29518,g23249,g7908,g29801,g18161,g25996,g13492,g6000,g24154,g12050,g26602,g12931,g25201,g9392,g30359,g25417,g34743,I33119,g24104,I13252,g10543,g31932,g27907,g31466,g8259,g2185,g30601,g33891,g17710,g32705,g18905,g17485,g34691,g24222,g22092,I23711,g8406,g17581,g34214,g16595,g34741,g34612,g32372,g9496,g4504,g22193,g33400,I27523,g29144,g21796,g21048,g27482,I12336,g21280,g29789,g25606,g28489,g3909,g28216,g16641,g30557,I24038,g32083,I13043,g9309,g34719,g24712,g27293,g27160,g6613,g27137,g34715,g16429,g10981,g28500,g10341,g29504,g27381,g33895,g13264,g23264,g28376,g28233,g24942,g18206,I17744,g31522,g12084,g12479,I12112,g9380,g34948,g11448,g10872,g28304,g27004,g13320,g27252,g23777,g27345,g7247,g34721,g9778,g28630,g24319,g21708,g10898,I33149,I32947,g32150,g32695,g16965,g22992,g18697,g29245,g14392,g25763,I14823,g27159,I17446,I27564,g22033,g24026,I14713,g1351,g21401,g9552,g21855,g13666,g24283,g15727,I21959,g8150,g27406,g32329,g26822,g10590,g29494,g31777,I24455,I12770,g17472,g21274,g18448,g28059,g1111,g26513,I26419,g5459,g12193,g22119,g29116,g16184,g34450,g9529,g27533,g21807,g7121,I15036,g22988,g28457,g14085,g32202,g19477,g33728,g7686,g18168,g20496,I32953,g7932,g2295,g3045,g10338,g29994,g29201,g19673,I15264,g32489,g22417,g11171,I15788,g5849,g14608,g15873,g25888,g9766,g19654,g12135,g20870,g34757,g20330,g16971,I16795,g18309,g12820,g30409,g14744,g34354,g15875,g25293,g15718,g5308,g22642,I32803,g29320,g33055,g24507,g28213,g18268,I31136,g33967,g13322,I22846,g2485,g16523,g16319,g30177,g29200,g29574,g17500,g24494,g30241,g28728,g24265,g31752,I17575,g30209,g6874,g26361,g16225,g34996,g14211,g34843,g17700,I22177,g28959,g19765,g3017,g28310,g30451,g33611,g25025,g5360,g5798,g1570,g26832,g29181,g34580,g34010,g29693,g25238,g33908,g4737,g25132,g32689,g4459,I24191,g13996,g18468,g1968,g19436,g26022,g35001,g16129,g22660,g33595,g13013,g29965,I14550,g11948,g10347,g32881,g21685,g6243,g18273,g27484,g12463,g16283,g25687,g33679,g33283,g7216,g10951,g21717,g32969,g1389,g30529,g34966,g29332,g25609,I32547,g8418,g17396,g31922,g21771,g27248,g21856,g34897,g17493,g13628,g14276,g32430,I14509,g10567,g34349,g27878,g29937,g13500,g22848,g32922,g12901,g11381,g23844,g27436,g26848,g12008,g17719,g12947,g18434,g27286,g12515,g13057,g4578,g1296,g32797,g23626,g19766,g27210,g32532,g23428,g10278,g11975,g24963,g13833,g12797,g11181,g34324,g2020,g15132,g33111,g32856,g34830,g30051,g7850,g19438,g24268,I32837,g27967,g15831,g18536,g22685,g12553,g13824,g34884,g18436,g28076,I29254,g13762,g832,g32248,g19050,g25752,g5869,g28817,g23379,g11995,I31277,g24601,g24391,g21948,g7970,I33170,g4749,g34009,g2269,g11250,g27029,g23872,g24214,g22004,g33380,g20010,g33534,g3841,g34754,g31976,I20609,g6173,I27232,g16097,g29733,g11724,g14151,I31823,g19662,g8218,g33105,g11885,g29285,g7262,g30020,g28225,g23899,g28038,g16675,g12505,g30484,I17925,g30145,g26811,g28528,g32729,g23057,g22593,g14142,g26635,g13655,I31307,I22748,g19682,g28639,g11449,g20653,g34217,g32890,g20453,g20503,g23913,g24068,g17776,g16195,g32391,g32794,g34475,g22542,g14332,I13111,g32771,I28883,g14036,g29175,g23448,g13252,I20468,g7534,g7191,g10028,g9959,g34695,g7328,g13597,g20014,g7640,g29708,g26817,g33578,g16202,g22134,g30562,g31515,g12491,g26607,g13866,g29877,I18680,I28866,g19785,g28052,g28455,g16642,g22721,g15793,g22999,g13971,g13835,g28436,g20666,g24569,g7846,g19968,I11743,g29770,I15289,g24953,g34628,g9746,g8302,g30456,g30435,g33531,g4878,g18412,g33869,g19127,g18173,I31843,g23320,g9920,g33465,g30152,g15654,g16590,g27737,g33548,g27344,I31127,g9963,g8404,g18525,g31873,g25562,g6825,I12251,g28666,g30129,g25265,g15591,g9595,g21053,I26461,g19379,I12840,I15242,g14123,g32632,I32431,g21461,g9969,g4423,I15194,g27162,I27314,g1644,g24580,g14423,I12287,g34416,g29667,g11233,g27233,g8137,g34880,g7473,g24638,g7027,g22076,g32676,g23721,g28335,g34348,g15839,g24501,g215,g19574,g14585,g16728,g27088,g2197,I14400,g1608,g24759,g22707,I26459,g14570,g18193,g5485,g31835,g31009,g34649,g33393,g33424,g28173,g25695,g9197,g10361,g5260,g28496,g31318,g29205,g34812,g30405,g2767,g21209,g968,g23121,g10385,g12845,g13312,g10605,g26846,g23196,g30523,g14348,I21722,g10678,g28106,g4300,g21966,g30333,I15727,g4809,g25030,I12135,g17668,g22661,g24661,I24438,I22912,g21862,I33070,g17578,g23460,g3774,g23809,g33905,g12869,g34881,g27214,g13284,I31301,g19524,g25054,g29614,g32264,g29289,g33986,g174,g24974,g4894,g32480,g22171,g14905,g31019,g28193,g34084,g28752,g31306,g3945,g25625,g8451,g32362,g29706,g25915,g10194,g31794,g32239,g26124,g25815,g28333,g34669,g13415,g21457,g19350,g24187,I22922,g21288,g33233,g18666,g11248,g28884,g10572,g21797,g33366,g2421,g30206,g7232,g24656,g11514,g3794,I31026,g17412,g70,g8009,g24994,g33267,g12221,g7565,g32866,g16966,g16517,g24150,g22059,g12044,g27257,g25094,g29747,g16762,g24993,g34345,g10909,g10626,g25112,g29894,g29375,g31514,I13280,g24128,g34537,I24008,g14411,I26367,g32641,g30222,g34027,I31226,g24138,g25985,I17136,g32207,I16201,I15288,g13515,g31487,g24570,g19467,g12322,g32971,g31829,g13342,g5097,I15342,g16605,g13530,g16325,g25942,g4477,g25597,I15243,g30307,I22712,g17124,g28522,g31319,g33145,I32881,g8055,g20911,g25701,I18101,g24452,g2882,g34275,I32237,I29368,g25786,g21267,g32956,g32858,g14331,g24668,g10406,I14205,g29556,g28870,g31934,I12497,g27517,I12041,g18197,g5196,g10032,g34942,g6093,g4141,g22020,g22666,g33002,g8278,g26356,g21248,g27202,g11117,g29596,I14368,g15614,g9745,g31872,g460,g34760,g9402,g20706,g12629,g29844,g17734,g32754,g31639,g29170,g24794,g32552,g12539,g5921,g23819,g34432,g18553,g25850,g25432,g34195,g29496,g34132,g6668,g17249,I31287,g6633,g25931,g24477,g2551,g13483,g10935,g27925,I14259,g14416,g22534,g30290,I30728,g20432,g19396,g32219,g20181,g9910,g17433,g110,g27629,g18226,g2941,g26311,g4831,g34725,g20657,g34359,g32056,g4474,g15705,g11283,g34554,g8481,I18154,g32617,g7362,g21389,g25989,g12078,g25835,g32663,g29275,g2965,I32525,g6082,g32427,g6820,g11164,g26904,g37,g19494,g20209,g17663,g30029,g10588,g10823,g19658,I32654,g28597,g16709,g32382,g27696,g7314,g25104,g28529,g33925,g28368,g3155,g9614,g32122,g33386,g29186,g30442,g33962,g28691,g23426,g9807,g14803,g9800,g21559,g27679,g24321,I22794,g34594,I30861,g18178,g21837,g13954,I12016,g28481,g28976,g26119,g21357,g1858,g23362,g23018,g29761,g22588,g28401,g25462,g34875,g25631,g19506,g1589,g996,g29286,g32164,g18389,g7150,g12025,g13907,g10169,g9663,g22658,g15730,g28480,g30565,g33096,g28696,I14797,g34692,g30228,g9252,g32099,g29858,g32769,g31917,g562,I18588,g31481,g16920,g18638,g20751,g20622,g22044,g30233,g2279,g20234,g11201,g7957,g10359,g807,g34623,g4180,I12098,g23577,g20982,g20599,g31020,g11401,g28662,g32760,g4040,g32044,g30084,g25902,g8450,g25592,g14338,g14360,g13505,g28723,I12141,g32586,g30070,g3684,g18117,g25679,I18785,g28280,g10796,g25922,I31011,I16515,g34171,I21036,g13995,g27083,g6826,g24130,g25663,g15277,g8387,g12194,g32285,g32832,g18505,g23432,g11868,g32734,g34299,g21428,g29628,g11302,g11202,g18509,g29576,g28846,g31657,g13017,g20444,g12930,g2898,g14999,g25878,g25456,g26961,g10683,g13624,g25377,g25617,g16708,g16816,g34443,g11954,g16654,I32812,g20173,g24490,g32744,g32903,g19413,g30124,g34631,g27674,g31316,g9762,g28068,g19538,g21932,I12793,g16657,g14094,g18465,g13765,g590,g1099,g10899,I12761,I22009,g33919,g27673,g14726,g29034,g30273,g12492,g32887,g13566,g30119,g30517,g33619,g6869,g23411,g18903,g30153,I18531,I12568,g34640,g29950,g30390,g30402,g18187,g18791,I17324,g30509,g11424,g25042,g18477,g30366,g15702,I17181,g26274,g33345,g11989,g6031,g32879,g12591,I14498,I16460,g18755,g31929,g30549,g8697,g12323,g34627,g34284,g10568,I12541,I18238,g637,g10616,g32911,I13184,I24445,g13109,g9462,g23029,g26970,g28346,g32241,g23332,g24199,g13998,g30515,g32163,g8954,g23796,g24551,g5563,g33245,I23357,g16883,g23555,g31221,g7002,g29223,g7544,g7231,g32533,g30281,g24206,g26918,g16122,g29814,g23135,g24502,g26251,g9971,g24229,g24879,g29506,g26779,g15128,g11045,I31211,g650,I15663,g10350,g18313,g33941,g7118,g25408,I18180,g31497,g14160,g34827,g26190,g22017,g19458,I20951,g19771,g33639,I18379,g14113,g822,g5579,g2599,g16691,g28606,g28070,g17614,g17494,g11313,g24196,g6044,g32842,g6641,g26785,g13496,g25072,g29367,I31985,I16544,I27528,g9825,g34373,g31232,g28515,g34588,g25524,I29214,g20111,g23270,g22093,g34529,g33794,g20329,g12307,g22846,g85,g10058,g32957,g32231,g20097,I31839,g25839,g25805,g20912,g12346,I22153,g5240,g29776,g29222,g29686,g21735,g18289,g26837,g11154,g25282,g27665,g23952,g34962,g30597,g14549,g14700,g32848,g11944,g17793,g21914,g14674,g9310,g18822,g31304,g33847,g31796,g13567,g27182,g21464,g4570,g1183,g33117,I15590,g22167,g30344,g32735,g27059,g26291,I14248,g13110,g26958,g13730,g12885,g32980,g14104,g20270,g27880,g34143,I18414,g18383,I15253,g10374,g25232,g26671,g34092,g15562,g29575,g20038,g29571,g22590,g32208,g3542,I24237,g13633,g9754,g22683,g33022,g23501,g869,g25014,g25414,g11083,g27364,g16521,g27284,g34916,g24966,g12680,g24912,g3625,g34769,g21370,g21364,g12842,g23888,g20714,g17788,g887,g4304,g22455,g19435,I17999,g8571,g23023,g23733,g25017,g9000,g9007,g31920,g34185,g31786,g27879,I14050,g23647,g15936,g24621,I13326,g25642,I17671,I27238,I31267,g24483,I25351,g12370,g22760,g18670,g9390,g27710,g18646,g28739,I32868,g8292,g14984,g16856,g30578,g20081,g31517,I11617,g25173,g8742,g23964,g12197,g32438,I21757,g18612,I24018,g16666,g30449,g27721,g34273,g3243,I18728,I29239,g14687,g34326,g19913,I18160,g27184,g18460,g28231,g33800,I21242,g29475,g25872,g33057,g20232,g8130,g13877,g3092,I16555,g34776,g5256,g31748,I22564,g12918,g24790,g23771,g25927,g8237,g21354,g27126,g34367,g2763,g33418,g22029,g11675,g34108,g27568,g18993,g29967,g16615,g19631,g7661,g16511,g31591,g11913,g32116,I31701,g25881,g20210,g34990,g25409,g16582,g16228,g10609,g32053,g32726,g26399,I12269,g11367,g33329,g29204,g20005,g33993,g23886,g24605,g30107,g28360,g31122,g9823,g28558,g22147,g23191,g33292,g27219,g19128,I29297,g28830,g30351,I25598,g21268,I18822,g23666,I14993,g25092,g29619,g16243,I31282,g28816,g34502,g27554,g12487,g9908,g7995,g16893,I17420,g1437,g28644,g16479,I20487,g24052,g33525,g21384,g2834,I31117,g26783,g32924,g32194,I28591,g25610,g16278,g19737,g4191,g9826,g8534,g33070,g27700,g27014,g9037,g14522,g20105,g18896,g34294,g3004,g34244,g32191,g28539,g16736,g25513,g13763,g19483,g24755,g22034,g33532,g12780,g8990,I24684,I13750,g23420,g21991,g4531,g16725,g29745,g24884,g225,g25159,g21697,g9064,I26094,g18351,g10509,g14745,g18743,g30196,g13928,g26296,g799,g19586,g23148,g34168,g22550,g18203,g23508,g25035,g7922,g29767,g33848,g20919,g30928,g18464,g23755,g15168,g16767,g11206,g21055,g1834,I31312,g28958,g9546,g28202,g24003,g23219,g19629,g32550,g31542,g17815,I27349,g10674,g20770,g10232,g24315,g32777,g8822,g52,g3767,g32457,g18321,g32959,g18535,g24578,g9671,g31870,g17714,g31764,I23961,g7197,I12070,g8211,g31500,g26684,g10802,g28072,g34610,g11796,g33598,g29974,g18564,I24064,g13191,g28843,g19370,g33317,g23897,g22986,g13086,g5712,g28299,g2567,g19610,g8733,I25190,g29296,g31231,g24796,I16040,g12196,g20511,g22855,g28206,g11033,g18276,g23947,g28192,g19860,I22871,g30005,g25686,g20615,I14409,g25800,g21278,g20573,g12721,g27772,g30049,g7450,g26100,g24204,g32603,g19709,I12546,g18198,g13707,g10622,g13296,g25785,g31312,g1259,g27581,g32380,g3281,g24288,g31470,g29380,g22712,g26935,g13506,g7479,I12382,g10499,g23927,g24756,g18759,g29810,g10473,g21305,I22755,g10034,g34327,g18091,g25626,I16521,g13202,g34313,g12854,g16959,I22557,g13096,I23351,g17640,g25250,I33197,g18829,g30999,g7643,g32104,g27043,g8650,g10175,g34414,g3447,g28504,g32731,g18462,g2307,g10026,g28896,g26923,g9257,g10409,g316,g29057,g12929,g34170,g25612,g12796,g5441,g5011,g16072,g22064,g9030,g7616,g25111,g26236,g13041,g26098,g9842,g15781,g2657,g25298,g24037,g21844,g23617,g16176,g24335,g32817,g26394,g32496,g17141,g32196,I12253,g27523,g32197,g28712,g24775,g30406,g33797,g26259,g23608,g31277,g23267,I32234,g17771,g24291,g24450,g15728,g32610,g2563,g17221,g6541,g30109,I24439,g24089,g10375,g17782,g30286,g20576,g26397,g16296,g13522,g29501,g32717,g34344,I18852,g18227,g718,g2461,I14653,g5188,g33788,g28720,g5417,g19432,I32976,g28900,g30671,g881,g7577,g27220,g25476,g22663,g25323,g14602,g4145,g9654,g24190,g34804,g12977,I16803,g31208,g33246,g24922,g14277,g30229,g32389,I15564,g34809,g32591,g30340,g24498,I28301,g5080,g29339,g31836,g736,g28852,I22028,g12686,I25552,g28508,g21726,g10308,g32589,g22996,g18149,g24931,g15148,g31269,g30398,g12028,g24365,g9607,g26812,g32424,g23154,g9901,g14363,g9759,g32258,g31465,I29221,g17789,g8829,I31829,g18766,I18337,I26929,g26655,g13012,g28345,g28564,g12166,g30524,g28772,g7280,g29185,g14514,g28714,g30195,g24119,g34774,I31142,g12342,g34951,g29764,I15162,g33384,g14845,g33523,g20637,I16579,g20148,g4213,g15700,g17431,g29648,g31493,g10397,g32580,g5897,g19638,g19268,g26781,I27677,g12000,g25134,g21689,g21905,g21070,I18107,g18720,g24362,g13596,g7148,g17146,g34189,g29329,g25767,g21293,g1079,g20080,g15719,g27453,g30480,g25128,g34706,g33618,I26130,g14124,g31374,g20272,g14764,g31655,g6827,g16807,g26223,g34791,g18538,g9917,g28103,I22793,g9500,g8883,g15709,g28636,g16719,g10151,g8740,g13756,g25690,g32236,g30547,g25762,I11682,g27705,g33886,g19626,g27024,g17692,g21836,g14066,g27593,I22894,g33596,g25982,g30521,g23968,g26611,g6140,g30481,g23992,g29719,g29013,g24327,g27759,g28646,g15348,g18485,g33404,g27099,g31762,g18154,g15938,g10803,g27687,g32233,g4093,g27579,g22529,g13603,g32900,g3845,g23274,g8438,I18888,g20039,g10428,g27485,g27007,I27409,g23491,g27274,g18463,g30285,g26603,I32432,g22722,g18442,g24344,g27971,g13319,g13942,g34805,I16391,g28325,I33164,g28131,g32428,I33179,g28789,g17123,g2236,g29850,I27519,g550,g12982,I32967,g26159,g15800,g30453,g33704,g34575,g20584,g21814,g30548,g25554,g14107,g33681,g33511,g10606,g30099,g24354,g24676,g24140,g19351,g11858,g23256,g23971,g19776,I14480,g9073,g25482,g28754,g21299,I14301,g27273,g31891,g29875,g34629,I22302,g31257,g32660,g27548,g30376,g32375,g17847,g15093,g34577,g30420,g26712,g24075,g10598,I18713,g22521,g22408,g1696,g32884,g21333,g22681,g34111,g22042,g16428,g33624,g17687,g34033,g9510,g17603,g29620,g15693,g27648,g23108,g3574,g12945,g27325,g14173,g8841,g21426,g25287,g14536,g28237,I29269,g10179,g16886,g34156,g32398,g9975,g25780,g19795,g13514,I20569,g22036,g10619,g20101,g18651,g5489,g12285,g11432,g298,I24027,I31972,g10059,g26231,g14005,g34282,g15669,g10511,I18879,g34494,g29378,g16214,g28577,g1263,I16676,g21719,g16096,g34803,g6451,I33030,g28249,g4643,g12296,g33439,g30197,I18845,g9631,g22096,g32566,I30718,g10719,g15840,g13920,g18738,g19358,I33109,g7327,g30155,g27929,g34680,I33064,g22190,g30504,I17650,I12487,g21858,g27035,g32874,g32875,g8672,g22840,g14899,g32525,g13476,g19661,g15569,g27452,g23915,g33108,g31212,g6989,g26854,g17134,g10393,I14745,g28274,g34318,g8720,g26630,g9417,g9961,g23532,I27449,g7369,g33268,g22043,g24914,g18908,g26200,g18616,g29182,g10147,g7909,g13056,g29879,g25220,g7400,g30455,g32741,g27414,g16986,g11631,g33508,g22214,g9557,g28864,g32139,g16245,g10183,g23024,I31564,g33425,g2311,g441,I11632,g17568,g21337,g22837,g19536,g29105,g17471,g18312,g4169,g33489,g18443,g27405,g11291,g16482,g8461,g23928,g30114,g7440,g23407,g112,g21753,g31262,g17669,g13300,g32596,I15208,g22831,g16160,g19692,g6723,g18278,g25966,g34392,g12402,g24091,g20390,g6961,g18294,I24048,g31227,g25967,g28599,g27824,g32727,I17884,g18315,g29645,g24264,I22542,g22517,g14357,g24328,g16349,g29324,g18764,g16299,g25,g33609,g26949,g28124,g12936,g28138,g4012,I14395,g12067,g23527,g31001,g20082,g13067,g34243,g911,g26990,g33964,g30473,g27016,I17448,g13738,g22981,g19473,g13349,g30225,g13944,g20071,g33473,g15965,g4005,g14616,g34368,g9775,g25239,g24109,g27567,g18300,g10800,g28062,g25899,g7788,g10287,g9983,g17655,g11888,g878,g24481,g20635,I12758,I24416,g5170,g20434,g34532,g32792,g24225,g21366,g3889,I14611,g30294,g34957,g22990,g27155,g24284,g32857,g26689,g30188,g32953,g25671,g7438,g10053,I32103,g33147,g21955,g12001,g26288,g34746,g24905,g15092,g32243,g27494,g14854,g16288,I14742,g31120,g16021,I32482,g11927,I23962,g32089,g5666,I11903,g18655,g11236,g28665,I33297,g24336,I27538,g3129,g15818,g14279,g3747,g29224,g30385,g21998,g24881,g21418,g14876,g29969,g17405,I12782,g18628,g218,I30986,g23001,g24553,g12405,I20369,g30067,g15716,g22012,g29962,g13543,g26203,g18445,g8607,g21703,g9020,g25711,g16846,g12969,g30576,g24033,g29199,g16281,g13222,g33998,g19450,g24463,g1236,g19711,g28783,g24341,g13854,g32819,g20100,I23600,g21704,g22941,g23775,g29265,g2748,g31016,g14139,g19567,g33032,g24703,I14902,g10928,g23932,g24565,g18945,I30123,g33880,g29809,g13383,g28689,I32855,g30423,I22422,g20091,I22275,g18671,g12646,g32210,g23312,I26960,g24524,g28627,g23837,g26861,g26964,g10180,g10474,g11754,g29580,g9299,I31515,g34449,g28608,I28579,g8345,g12622,g31819,g14643,g14874,g34483,g28235,g20704,g20564,g12659,g34142,g31170,g23253,g28939,g33851,g13477,g32716,I26366,g23838,g32479,g20765,g31298,g29566,I15128,I17404,g15224,I21047,I14211,g27369,g14962,I32997,g34997,g29794,g26889,g27546,g5575,I26989,g2102,g23912,g27226,g19069,g16507,g8114,I15149,g25694,g25004,g22755,g19732,g33009,I14228,g27288,g16931,g30141,g23390,g2040,g17954,g11812,g24971,g12932,g10584,g25115,g25096,g23481,g14420,g12762,g8171,g20208,g12170,g30086,I12503,g17775,I22753,g17309,g29165,I19789,g27287,g10601,I15954,I12086,g21660,g18253,g6727,g32310,g12150,g10108,g24121,g21799,I31586,g20660,g24573,g32671,g9556,g22719,g10597,I31231,g9724,g9661,g6023,I22719,g27933,g3298,g33613,g32962,g10334,g9907,g24700,g31991,g7343,g13593,g9274,g21901,g22489,I18003,g27560,g34556,g11999,g26827,g21891,I26409,g20497,g32862,g31756,g21561,g16677,g29253,g29081,I32884,g6802,g10476,g6993,g19558,g27573,g25542,g22,g3096,g33085,g11714,I28458,g30121,g10518,g20516,g8227,g15792,g947,I12092,g16809,g6808,I28897,I20985,g25692,g21943,g12851,g27965,g24977,g17745,g2715,g32701,g32165,g8871,g25095,g27500,g199,g15837,g32945,g5794,g8514,I30727,g31129,g25141,g27993,g9686,g13889,g12208,g22056,g24247,g32212,g30358,g25869,g29044,g22921,I26523,g24232,g34792,g17465,g744,g32745,I18259,g29274,g20084,g12048,I15593,g23747,g5841,g31825,g29328,I15682,g1448,I30980,g18668,g34056,I12787,g3694,g26839,g34039,g20978,g25818,g12870,g11747,g9086,g2413,g20110,g28373,g22067,g21952,g16645,g23602,g28587,g17401,g11544,g24227,g24590,g20219,g32906,g34346,g34648,g32112,g14584,g6940,g28265,g27954,g23994,g11252,g24535,g10281,I33252,g14344,g27354,g28698,g26799,g23220,g30278,g20375,g10412,g18757,g18627,g24002,I12605,g26966,g32255,g34291,g6926,I19851,g10207,g29078,g22399,g20768,I24400,g23500,g17579,g26856,g20643,I31326,g33501,g376,g20566,g17525,g21896,I17695,g26922,g31812,g23357,g18661,g34601,g8848,g33814,g1959,g25868,g33122,g32011,g24390,g9491,g14417,g24298,g15628,g8033,g29689,g11042,g25171,g29196,g26310,g34417,g7649,g21456,g26994,g23761,g32178,I31610,g23821,g25650,g2370,g17174,g30291,g12755,g26831,g30113,g33509,g2907,g2946,g32546,g27064,g29235,g33867,g31142,g2595,g12524,g18332,g24389,g10041,g4698,g23648,g33134,g18708,g33375,g32935,g11881,I31172,g31871,g14237,g32270,g13037,g27958,g33504,g12983,g13480,g7046,g8182,g13247,g33813,g16653,g22087,g33697,g26610,g33539,g3782,g19529,g28735,I32904,g20656,g24620,g32553,g32583,I31251,g21750,g22199,g5630,g29255,g27668,g16763,g25547,g7690,g23926,g14636,g28820,g12046,g8945,g20233,g21829,g8205,I13442,g19594,g21558,g33580,g24325,g10029,g29702,g34813,g21412,g1848,g26963,g27100,g20235,g25498,g31709,g15160,g24652,g4555,I12666,g30513,g10721,g6419,g32279,I16535,g2112,g24094,g32773,I18417,g12286,g26053,g23859,g8107,g13990,g24926,g18614,g28603,I12730,g33333,g11960,I29314,I32170,g32028,g34918,g24814,g16526,g33702,g24546,g28668,g32328,g19387,g24911,g24557,I22873,I25555,I14398,g29773,g30352,g22032,g19495,g4194,I20467,g32140,g14567,g22156,g28467,g34005,I31849,g33627,g12037,g33016,g2319,g18374,I18031,g15712,g32979,g32749,g20651,g33885,g16673,I20891,g15694,I12767,g33137,g9716,g23228,g19385,g18792,g9259,g14207,g16,g24699,g34620,g17522,g33652,g23471,g16022,I13424,I29253,g6973,I22938,g27828,g8993,I12300,g18176,g26666,g4281,g18815,g30271,g21394,g24840,g28341,g27854,g1489,g18946,g29114,g21824,g21980,g12336,g25082,I15122,g23012,g24503,I20189,g32069,g65,g14003,g14563,g18306,g3227,g30100,I27758,g18107,g15582,g31278,g17177,g24426,g27479,g33593,g12924,g30034,I12899,g7195,g4138,g33447,g34191,g31243,g14599,g23286,g23581,g12767,g8756,I22111,g10540,g27317,g1559,I26516,g32907,I17436,g21331,g26024,g27370,g1246,g32500,g3881,g10364,g32473,g30042,g14882,g30488,g18702,g25761,g13385,g16607,g914,g10181,I11708,g29323,g29991,g30929,g23387,g34272,g6959,g24451,I12876,g24360,g9194,g17013,g14924,g25652,g9538,g27093,g27659,g10229,g26720,g24986,g21335,g28454,g17613,g21555,g15814,g16246,g22110,I14788,I29284,g34626,g6533,g7980,g24651,g27375,g10230,g34218,g19336,g23868,g14831,g7778,g17636,I29913,g25367,I31346,g25666,g32511,I25790,g16210,g34699,g13188,I31550,g30012,g22664,g34332,I25779,g20512,I33034,g17794,I12773,g18889,g34519,g24932,g7701,g12638,g18609,g18106,g34976,g12015,g14719,I12120,g22405,g28381,g14858,g8052,g10115,g26841,g18954,g28776,g71,g28969,g12225,g23000,g16703,g30595,g31989,g6609,I32909,g32244,I31619,g16589,I22366,g29913,g34473,g24334,g12997,g26488,g30526,g19606,g34668,g30426,g28160,g22662,g9444,g1802,g4462,g17744,g7634,I14800,g28736,g33353,g28425,g31838,g34347,g31182,g9547,g8530,g32854,g12083,g20905,g34868,g18449,g24348,g21291,g28520,g33936,g30170,g27800,g14202,g32780,g5805,g4157,g27415,g31889,g26153,g8064,g12222,g28774,g14308,g15672,g9748,g23104,g15100,g26965,g17738,g9264,g32192,g24984,g28210,g19601,g14641,g22040,g14449,g13464,g6954,g22668,g26387,I17392,g8249,g13886,g22000,g11833;
//# 38 inputs
//# 304 outputs
//# 1426 D-type flipflops
//# 7805 inverters
//# 11448 gates (5516 ANDs + 2126 NANDs + 2621 ORs + 1185 NORs)
//
//
//
  MSFF DFF_0(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5057),.DATA(g33046));
  MSFF DFF_1(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2771),.DATA(g34441));
  MSFF DFF_2(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1882),.DATA(g33982));
  MSFF DFF_3(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6462),.DATA(g25751));
  MSFF DFF_4(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2299),.DATA(g34007));
  MSFF DFF_5(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4040),.DATA(g24276));
  MSFF DFF_6(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2547),.DATA(g30381));
  MSFF DFF_7(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g559),.DATA(g640));
  MSFF DFF_8(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3017),.DATA(g31877));
  MSFF DFF_9(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3243),.DATA(g30405));
  MSFF DFF_10(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g452),.DATA(g25604));
  MSFF DFF_11(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g464),.DATA(g25607));
  MSFF DFF_12(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3542),.DATA(g30416));
  MSFF DFF_13(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5232),.DATA(g30466));
  MSFF DFF_14(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5813),.DATA(g25736));
  MSFF DFF_15(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2907),.DATA(g34617));
  MSFF DFF_16(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1744),.DATA(g33974));
  MSFF DFF_17(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5909),.DATA(g30505));
  MSFF DFF_18(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1802),.DATA(g33554));
  MSFF DFF_19(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3554),.DATA(g30432));
  MSFF DFF_20(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6219),.DATA(g33064));
  MSFF DFF_21(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g807),.DATA(g34881));
  MSFF DFF_22(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6031),.DATA(g6027));
  MSFF DFF_23(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g847),.DATA(g24216));
  MSFF DFF_24(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g976),.DATA(g24232));
  MSFF DFF_25(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4172),.DATA(g34733));
  MSFF DFF_26(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4372),.DATA(g34882));
  MSFF DFF_27(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3512),.DATA(g33026));
  MSFF DFF_28(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g749),.DATA(g31867));
  MSFF DFF_29(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3490),.DATA(g25668));
  MSFF DFF_30(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6005),.DATA(g24344));
  MSFF DFF_31(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4235),.DATA(g4232));
  MSFF DFF_32(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1600),.DATA(g33966));
  MSFF DFF_33(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1714),.DATA(g33550));
  MSFF DFF_34(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3649),.DATA(g3625));
  MSFF DFF_35(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3155),.DATA(g30393));
  MSFF DFF_36(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3355),.DATA(g31880));
  MSFF DFF_37(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2236),.DATA(g29248));
  MSFF DFF_38(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4555),.DATA(g4571));
  MSFF DFF_39(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3698),.DATA(g24274));
  MSFF DFF_40(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6073),.DATA(g31920));
  MSFF DFF_41(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1736),.DATA(g33973));
  MSFF DFF_42(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1968),.DATA(g30360));
  MSFF DFF_43(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4621),.DATA(g34460));
  MSFF DFF_44(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5607),.DATA(g30494));
  MSFF DFF_45(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2657),.DATA(g30384));
  MSFF DFF_46(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5659),.DATA(g24340));
  MSFF DFF_47(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g490),.DATA(g29223));
  MSFF DFF_48(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g311),.DATA(g26881));
  MSFF DFF_49(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6069),.DATA(g31925));
  MSFF DFF_50(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g772),.DATA(g34252));
  MSFF DFF_51(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5587),.DATA(g30489));
  MSFF DFF_52(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6177),.DATA(g29301));
  MSFF DFF_53(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6377),.DATA(g6373));
  MSFF DFF_54(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3167),.DATA(g33022));
  MSFF DFF_55(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5615),.DATA(g30496));
  MSFF DFF_56(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4567),.DATA(g33043));
  MSFF DFF_57(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3057),.DATA(g28062));
  MSFF DFF_58(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3457),.DATA(g29263));
  MSFF DFF_59(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6287),.DATA(g30533));
  MSFF DFF_60(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1500),.DATA(g24256));
  MSFF DFF_61(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2563),.DATA(g34015));
  MSFF DFF_62(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4776),.DATA(g34031));
  MSFF DFF_63(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4593),.DATA(g34452));
  MSFF DFF_64(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6199),.DATA(g34646));
  MSFF DFF_65(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2295),.DATA(g34001));
  MSFF DFF_66(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1384),.DATA(g25633));
  MSFF DFF_67(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1339),.DATA(g24259));
  MSFF DFF_68(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5180),.DATA(g33049));
  MSFF DFF_69(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2844),.DATA(g34609));
  MSFF DFF_70(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1024),.DATA(g31869));
  MSFF DFF_71(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5591),.DATA(g30490));
  MSFF DFF_72(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3598),.DATA(g30427));
  MSFF DFF_73(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4264),.DATA(g21894));
  MSFF DFF_74(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g767),.DATA(g33965));
  MSFF DFF_75(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5853),.DATA(g34645));
  MSFF DFF_76(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3321),.DATA(g3317));
  MSFF DFF_77(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2089),.DATA(g33571));
  MSFF DFF_78(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4933),.DATA(g34267));
  MSFF DFF_79(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4521),.DATA(g26971));
  MSFF DFF_80(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5507),.DATA(g34644));
  MSFF DFF_81(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3625),.DATA(g3618));
  MSFF DFF_82(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6291),.DATA(g30534));
  MSFF DFF_83(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g294),.DATA(g33535));
  MSFF DFF_84(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5559),.DATA(g30498));
  MSFF DFF_85(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5794),.DATA(g25728));
  MSFF DFF_86(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6144),.DATA(g25743));
  MSFF DFF_87(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3813),.DATA(g25684));
  MSFF DFF_88(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g562),.DATA(g25613));
  MSFF DFF_89(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g608),.DATA(g34438));
  MSFF DFF_90(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1205),.DATA(g24244));
  MSFF DFF_91(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3909),.DATA(g30439));
  MSFF DFF_92(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6259),.DATA(g30541));
  MSFF DFF_93(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5905),.DATA(g30519));
  MSFF DFF_94(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g921),.DATA(g25621));
  MSFF DFF_95(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2955),.DATA(g34807));
  MSFF DFF_96(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g203),.DATA(g25599));
  MSFF DFF_97(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6088),.DATA(g31924));
  MSFF DFF_98(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1099),.DATA(g24235));
  MSFF DFF_99(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4878),.DATA(g34036));
  MSFF DFF_100(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5204),.DATA(g30476));
  MSFF DFF_101(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5630),.DATA(g5623));
  MSFF DFF_102(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3606),.DATA(g30429));
  MSFF DFF_103(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1926),.DATA(g32997));
  MSFF DFF_104(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6215),.DATA(g33063));
  MSFF DFF_105(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3586),.DATA(g30424));
  MSFF DFF_106(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g291),.DATA(g32977));
  MSFF DFF_107(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4674),.DATA(g34026));
  MSFF DFF_108(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3570),.DATA(g30420));
  MSFF DFF_109(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g640),.DATA(g637));
  MSFF DFF_110(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5969),.DATA(g6012));
  MSFF DFF_111(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1862),.DATA(g33560));
  MSFF DFF_112(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g676),.DATA(g29226));
  MSFF DFF_113(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g843),.DATA(g25619));
  MSFF DFF_114(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4132),.DATA(g28076));
  MSFF DFF_115(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4332),.DATA(g34455));
  MSFF DFF_116(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4153),.DATA(g30457));
  MSFF DFF_117(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5666),.DATA(g5637));
  MSFF DFF_118(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6336),.DATA(g33625));
  MSFF DFF_119(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g622),.DATA(g34790));
  MSFF DFF_120(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3506),.DATA(g30414));
  MSFF DFF_121(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4558),.DATA(g26966));
  MSFF DFF_122(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6065),.DATA(g31923));
  MSFF DFF_123(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6322),.DATA(g6315));
  MSFF DFF_124(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3111),.DATA(g25656));
  MSFF DFF_125(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g117),.DATA(g30390));
  MSFF DFF_126(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2837),.DATA(g26935));
  MSFF DFF_127(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g939),.DATA(g34727));
  MSFF DFF_128(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g278),.DATA(g25594));
  MSFF DFF_129(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4492),.DATA(g26963));
  MSFF DFF_130(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4864),.DATA(g34034));
  MSFF DFF_131(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1036),.DATA(g33541));
  MSFF DFF_132(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g128),.DATA(g28093));
  MSFF DFF_133(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1178),.DATA(g24236));
  MSFF DFF_134(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3239),.DATA(g30404));
  MSFF DFF_135(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g718),.DATA(g28051));
  MSFF DFF_136(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6195),.DATA(g29303));
  MSFF DFF_137(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1135),.DATA(g26917));
  MSFF DFF_138(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6137),.DATA(g25741));
  MSFF DFF_139(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6395),.DATA(g33624));
  MSFF DFF_140(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3380),.DATA(g31882));
  MSFF DFF_141(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5343),.DATA(g24337));
  MSFF DFF_142(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g554),.DATA(g34911));
  MSFF DFF_143(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g496),.DATA(g33963));
  MSFF DFF_144(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3853),.DATA(g34627));
  MSFF DFF_145(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5134),.DATA(g29282));
  MSFF DFF_146(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1422),.DATA(g1418));
  MSFF DFF_147(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3794),.DATA(g25676));
  MSFF DFF_148(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2485),.DATA(g33013));
  MSFF DFF_149(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g925),.DATA(g32981));
  MSFF DFF_150(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g48),.DATA(g34993));
  MSFF DFF_151(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5555),.DATA(g30483));
  MSFF DFF_152(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g878),.DATA(g875));
  MSFF DFF_153(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1798),.DATA(g32994));
  MSFF DFF_154(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4076),.DATA(g28070));
  MSFF DFF_155(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2941),.DATA(g34806));
  MSFF DFF_156(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3905),.DATA(g30453));
  MSFF DFF_157(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g763),.DATA(g33539));
  MSFF DFF_158(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6255),.DATA(g30526));
  MSFF DFF_159(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4375),.DATA(g26951));
  MSFF DFF_160(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4871),.DATA(g34035));
  MSFF DFF_161(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4722),.DATA(g34636));
  MSFF DFF_162(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g590),.DATA(g32978));
  MSFF DFF_163(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6692),.DATA(g6668));
  MSFF DFF_164(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1632),.DATA(g30348));
  MSFF DFF_165(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5313),.DATA(g24336));
  MSFF DFF_166(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3100),.DATA(g3092));
  MSFF DFF_167(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1495),.DATA(g24250));
  MSFF DFF_168(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6497),.DATA(g6490));
  MSFF DFF_169(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1437),.DATA(g29236));
  MSFF DFF_170(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6154),.DATA(g29298));
  MSFF DFF_171(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1579),.DATA(g1576));
  MSFF DFF_172(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5567),.DATA(g30499));
  MSFF DFF_173(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1752),.DATA(g33976));
  MSFF DFF_174(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1917),.DATA(g32996));
  MSFF DFF_175(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g744),.DATA(g30335));
  MSFF DFF_176(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3040),.DATA(g31878));
  MSFF DFF_177(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4737),.DATA(g34637));
  MSFF DFF_178(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4809),.DATA(g25693));
  MSFF DFF_179(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6267),.DATA(g30528));
  MSFF DFF_180(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3440),.DATA(g25661));
  MSFF DFF_181(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3969),.DATA(g4012));
  MSFF DFF_182(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1442),.DATA(g24251));
  MSFF DFF_183(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5965),.DATA(g30521));
  MSFF DFF_184(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4477),.DATA(g26960));
  MSFF DFF_185(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1233),.DATA(g24239));
  MSFF DFF_186(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4643),.DATA(g34259));
  MSFF DFF_187(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5264),.DATA(g30474));
  MSFF DFF_188(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6329),.DATA(g6351));
  MSFF DFF_189(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2610),.DATA(g33016));
  MSFF DFF_190(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5160),.DATA(g34643));
  MSFF DFF_191(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5360),.DATA(g31905));
  MSFF DFF_192(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5933),.DATA(g30510));
  MSFF DFF_193(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1454),.DATA(g29239));
  MSFF DFF_194(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g753),.DATA(g26897));
  MSFF DFF_195(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1296),.DATA(g34729));
  MSFF DFF_196(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3151),.DATA(g34625));
  MSFF DFF_197(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2980),.DATA(g34800));
  MSFF DFF_198(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6727),.DATA(g24353));
  MSFF DFF_199(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3530),.DATA(g33029));
  MSFF DFF_200(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4742),.DATA(g21903));
  MSFF DFF_201(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4104),.DATA(g33615));
  MSFF DFF_202(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1532),.DATA(g24253));
  MSFF DFF_203(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4304),.DATA(g24281));
  MSFF DFF_204(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2177),.DATA(g33997));
  MSFF DFF_205(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3010),.DATA(g25651));
  MSFF DFF_206(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g52),.DATA(g34997));
  MSFF DFF_207(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4754),.DATA(g34263));
  MSFF DFF_208(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1189),.DATA(g24237));
  MSFF DFF_209(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2287),.DATA(g33584));
  MSFF DFF_210(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4273),.DATA(g24280));
  MSFF DFF_211(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1389),.DATA(g26920));
  MSFF DFF_212(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1706),.DATA(g33548));
  MSFF DFF_213(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5835),.DATA(g29296));
  MSFF DFF_214(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1171),.DATA(g30338));
  MSFF DFF_215(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4269),.DATA(g21895));
  MSFF DFF_216(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2399),.DATA(g33588));
  MSFF DFF_217(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3372),.DATA(g31886));
  MSFF DFF_218(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4983),.DATA(g34041));
  MSFF DFF_219(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5611),.DATA(g30495));
  MSFF DFF_220(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3618),.DATA(g3661));
  MSFF DFF_221(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4572),.DATA(g29279));
  MSFF DFF_222(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3143),.DATA(g25655));
  MSFF DFF_223(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2898),.DATA(g34795));
  MSFF DFF_224(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3343),.DATA(g24269));
  MSFF DFF_225(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3235),.DATA(g30403));
  MSFF DFF_226(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4543),.DATA(g33042));
  MSFF DFF_227(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3566),.DATA(g30419));
  MSFF DFF_228(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4534),.DATA(g34023));
  MSFF DFF_229(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4961),.DATA(g28090));
  MSFF DFF_230(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6398),.DATA(g31926));
  MSFF DFF_231(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4927),.DATA(g34642));
  MSFF DFF_232(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2259),.DATA(g30370));
  MSFF DFF_233(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2819),.DATA(g34448));
  MSFF DFF_234(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4414),.DATA(g26946));
  MSFF DFF_235(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5802),.DATA(g5794));
  MSFF DFF_236(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2852),.DATA(g34610));
  MSFF DFF_237(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g417),.DATA(g24209));
  MSFF DFF_238(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g681),.DATA(g28047));
  MSFF DFF_239(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g437),.DATA(g24206));
  MSFF DFF_240(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g351),.DATA(g26891));
  MSFF DFF_241(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5901),.DATA(g30504));
  MSFF DFF_242(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2886),.DATA(g34798));
  MSFF DFF_243(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3494),.DATA(g25669));
  MSFF DFF_244(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5511),.DATA(g30480));
  MSFF DFF_245(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3518),.DATA(g33027));
  MSFF DFF_246(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1604),.DATA(g33972));
  MSFF DFF_247(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4135),.DATA(g28077));
  MSFF DFF_248(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5092),.DATA(g25697));
  MSFF DFF_249(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4831),.DATA(g28099));
  MSFF DFF_250(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4382),.DATA(g26947));
  MSFF DFF_251(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6386),.DATA(g24350));
  MSFF DFF_252(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g479),.DATA(g24210));
  MSFF DFF_253(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3965),.DATA(g30455));
  MSFF DFF_254(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4749),.DATA(g28084));
  MSFF DFF_255(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2008),.DATA(g33993));
  MSFF DFF_256(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g736),.DATA(g802));
  MSFF DFF_257(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3933),.DATA(g30444));
  MSFF DFF_258(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g222),.DATA(g33537));
  MSFF DFF_259(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3050),.DATA(g25650));
  MSFF DFF_260(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5736),.DATA(g31915));
  MSFF DFF_261(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1052),.DATA(g25625));
  MSFF DFF_262(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g58),.DATA(g30328));
  MSFF DFF_263(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5623),.DATA(g5666));
  MSFF DFF_264(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2122),.DATA(g30366));
  MSFF DFF_265(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2465),.DATA(g33593));
  MSFF DFF_266(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6483),.DATA(g25755));
  MSFF DFF_267(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5889),.DATA(g30502));
  MSFF DFF_268(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4495),.DATA(g33036));
  MSFF DFF_269(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g365),.DATA(g25595));
  MSFF DFF_270(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4653),.DATA(g34462));
  MSFF DFF_271(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3179),.DATA(g33024));
  MSFF DFF_272(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1728),.DATA(g33552));
  MSFF DFF_273(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2433),.DATA(g34014));
  MSFF DFF_274(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3835),.DATA(g29273));
  MSFF DFF_275(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6187),.DATA(g25748));
  MSFF DFF_276(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4917),.DATA(g34638));
  MSFF DFF_277(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1070),.DATA(g30341));
  MSFF DFF_278(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g822),.DATA(g26899));
  MSFF DFF_279(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6027),.DATA(g6023));
  MSFF DFF_280(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g914),.DATA(g30336));
  MSFF DFF_281(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5339),.DATA(g5335));
  MSFF DFF_282(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4164),.DATA(g26940));
  MSFF DFF_283(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g969),.DATA(g25622));
  MSFF DFF_284(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2807),.DATA(g34447));
  MSFF DFF_285(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5424),.DATA(g25709));
  MSFF DFF_286(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4054),.DATA(g33613));
  MSFF DFF_287(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6191),.DATA(g25749));
  MSFF DFF_288(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5077),.DATA(g25704));
  MSFF DFF_289(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5523),.DATA(g33053));
  MSFF DFF_290(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3680),.DATA(g3676));
  MSFF DFF_291(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6637),.DATA(g30555));
  MSFF DFF_292(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g174),.DATA(g25601));
  MSFF DFF_293(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1682),.DATA(g33971));
  MSFF DFF_294(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g355),.DATA(g26892));
  MSFF DFF_295(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1087),.DATA(g1083));
  MSFF DFF_296(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1105),.DATA(g26915));
  MSFF DFF_297(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2342),.DATA(g33008));
  MSFF DFF_298(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6307),.DATA(g30538));
  MSFF DFF_299(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3802),.DATA(g3794));
  MSFF DFF_300(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6159),.DATA(g25750));
  MSFF DFF_301(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2255),.DATA(g30369));
  MSFF DFF_302(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2815),.DATA(g34446));
  MSFF DFF_303(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g911),.DATA(g29230));
  MSFF DFF_304(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g43),.DATA(g34789));
  MSFF DFF_305(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4012),.DATA(g3983));
  MSFF DFF_306(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1748),.DATA(g33975));
  MSFF DFF_307(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5551),.DATA(g30497));
  MSFF DFF_308(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5742),.DATA(g31917));
  MSFF DFF_309(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3558),.DATA(g30418));
  MSFF DFF_310(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5499),.DATA(g25721));
  MSFF DFF_311(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2960),.DATA(g34622));
  MSFF DFF_312(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3901),.DATA(g30438));
  MSFF DFF_313(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4888),.DATA(g34266));
  MSFF DFF_314(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6251),.DATA(g30540));
  MSFF DFF_315(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6315),.DATA(g6358));
  MSFF DFF_316(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1373),.DATA(g32986));
  MSFF DFF_317(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3092),.DATA(g25648));
  MSFF DFF_318(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g157),.DATA(g33960));
  MSFF DFF_319(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2783),.DATA(g34442));
  MSFF DFF_320(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4281),.DATA(g4277));
  MSFF DFF_321(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3574),.DATA(g30421));
  MSFF DFF_322(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2112),.DATA(g33573));
  MSFF DFF_323(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1283),.DATA(g34730));
  MSFF DFF_324(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g433),.DATA(g24205));
  MSFF DFF_325(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4297),.DATA(g4294));
  MSFF DFF_326(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5983),.DATA(g6005));
  MSFF DFF_327(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1459),.DATA(g1399));
  MSFF DFF_328(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g758),.DATA(g32979));
  MSFF DFF_329(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5712),.DATA(g25731));
  MSFF DFF_330(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4138),.DATA(g28078));
  MSFF DFF_331(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4639),.DATA(g34025));
  MSFF DFF_332(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6537),.DATA(g25763));
  MSFF DFF_333(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5543),.DATA(g30481));
  MSFF DFF_334(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1582),.DATA(g1500));
  MSFF DFF_335(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3736),.DATA(g31890));
  MSFF DFF_336(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5961),.DATA(g30517));
  MSFF DFF_337(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6243),.DATA(g30539));
  MSFF DFF_338(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g632),.DATA(g34880));
  MSFF DFF_339(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1227),.DATA(g24242));
  MSFF DFF_340(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3889),.DATA(g30436));
  MSFF DFF_341(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3476),.DATA(g29265));
  MSFF DFF_342(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1664),.DATA(g32990));
  MSFF DFF_343(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1246),.DATA(g24245));
  MSFF DFF_344(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6128),.DATA(g25739));
  MSFF DFF_345(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6629),.DATA(g30553));
  MSFF DFF_346(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g246),.DATA(g26907));
  MSFF DFF_347(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4049),.DATA(g24278));
  MSFF DFF_348(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4449),.DATA(g26955));
  MSFF DFF_349(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2932),.DATA(g24282));
  MSFF DFF_350(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4575),.DATA(g29276));
  MSFF DFF_351(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4098),.DATA(g31894));
  MSFF DFF_352(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4498),.DATA(g33037));
  MSFF DFF_353(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g528),.DATA(g26894));
  MSFF DFF_354(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5436),.DATA(g25711));
  MSFF DFF_355(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g16),.DATA(g34593));
  MSFF DFF_356(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3139),.DATA(g25654));
  MSFF DFF_357(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g102),.DATA(g33962));
  MSFF DFF_358(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4584),.DATA(g34451));
  MSFF DFF_359(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g142),.DATA(g34250));
  MSFF DFF_360(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5335),.DATA(g5331));
  MSFF DFF_361(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5831),.DATA(g29295));
  MSFF DFF_362(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g239),.DATA(g26905));
  MSFF DFF_363(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1216),.DATA(g25629));
  MSFF DFF_364(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2848),.DATA(g34792));
  MSFF DFF_365(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5805),.DATA(g5798));
  MSFF DFF_366(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5022),.DATA(g25703));
  MSFF DFF_367(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4019),.DATA(g4000));
  MSFF DFF_368(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1030),.DATA(g32983));
  MSFF DFF_369(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3672),.DATA(g3668));
  MSFF DFF_370(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3231),.DATA(g30402));
  MSFF DFF_371(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6490),.DATA(g25757));
  MSFF DFF_372(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1430),.DATA(g1426));
  MSFF DFF_373(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4452),.DATA(g4446));
  MSFF DFF_374(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2241),.DATA(g33999));
  MSFF DFF_375(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1564),.DATA(g24262));
  MSFF DFF_376(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5798),.DATA(g25729));
  MSFF DFF_377(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6148),.DATA(g6140));
  MSFF DFF_378(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6649),.DATA(g30558));
  MSFF DFF_379(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g110),.DATA(g34848));
  MSFF DFF_380(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g884),.DATA(g881));
  MSFF DFF_381(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3742),.DATA(g31892));
  MSFF DFF_382(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g225),.DATA(g26901));
  MSFF DFF_383(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4486),.DATA(g26961));
  MSFF DFF_384(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4504),.DATA(g33039));
  MSFF DFF_385(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5873),.DATA(g33059));
  MSFF DFF_386(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5037),.DATA(g31899));
  MSFF DFF_387(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2319),.DATA(g33007));
  MSFF DFF_388(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5495),.DATA(g25720));
  MSFF DFF_389(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4185),.DATA(g21891));
  MSFF DFF_390(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5208),.DATA(g30462));
  MSFF DFF_391(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2152),.DATA(g18422));
  MSFF DFF_392(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5579),.DATA(g30487));
  MSFF DFF_393(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5869),.DATA(g33058));
  MSFF DFF_394(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5719),.DATA(g31916));
  MSFF DFF_395(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1589),.DATA(g24261));
  MSFF DFF_396(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5752),.DATA(g25730));
  MSFF DFF_397(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6279),.DATA(g30531));
  MSFF DFF_398(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5917),.DATA(g30506));
  MSFF DFF_399(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2975),.DATA(g34804));
  MSFF DFF_400(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6167),.DATA(g25747));
  MSFF DFF_401(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3983),.DATA(g4005));
  MSFF DFF_402(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2599),.DATA(g33601));
  MSFF DFF_403(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1448),.DATA(g26922));
  MSFF DFF_404(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g881),.DATA(g878));
  MSFF DFF_405(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3712),.DATA(g25679));
  MSFF DFF_406(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2370),.DATA(g29250));
  MSFF DFF_407(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5164),.DATA(g30459));
  MSFF DFF_408(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1333),.DATA(g1582));
  MSFF DFF_409(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g153),.DATA(g33534));
  MSFF DFF_410(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6549),.DATA(g30543));
  MSFF DFF_411(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4087),.DATA(g29275));
  MSFF DFF_412(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4801),.DATA(g34030));
  MSFF DFF_413(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2984),.DATA(g34980));
  MSFF DFF_414(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3961),.DATA(g30451));
  MSFF DFF_415(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5770),.DATA(g25723));
  MSFF DFF_416(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g962),.DATA(g25627));
  MSFF DFF_417(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g101),.DATA(g34787));
  MSFF DFF_418(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4226),.DATA(g4222));
  MSFF DFF_419(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6625),.DATA(g30552));
  MSFF DFF_420(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g51),.DATA(g34996));
  MSFF DFF_421(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1018),.DATA(g30337));
  MSFF DFF_422(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1418),.DATA(g24254));
  MSFF DFF_423(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4045),.DATA(g24277));
  MSFF DFF_424(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1467),.DATA(g29237));
  MSFF DFF_425(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2461),.DATA(g30378));
  MSFF DFF_426(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5706),.DATA(g31912));
  MSFF DFF_427(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g457),.DATA(g25603));
  MSFF DFF_428(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2756),.DATA(g33019));
  MSFF DFF_429(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5990),.DATA(g33623));
  MSFF DFF_430(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g471),.DATA(g25608));
  MSFF DFF_431(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1256),.DATA(g29235));
  MSFF DFF_432(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5029),.DATA(g31902));
  MSFF DFF_433(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6519),.DATA(g29306));
  MSFF DFF_434(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4169),.DATA(g28080));
  MSFF DFF_435(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1816),.DATA(g33978));
  MSFF DFF_436(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4369),.DATA(g26970));
  MSFF DFF_437(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3436),.DATA(g25660));
  MSFF DFF_438(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5787),.DATA(g25726));
  MSFF DFF_439(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4578),.DATA(g29278));
  MSFF DFF_440(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4459),.DATA(g34253));
  MSFF DFF_441(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3831),.DATA(g29272));
  MSFF DFF_442(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2514),.DATA(g33595));
  MSFF DFF_443(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3288),.DATA(g33610));
  MSFF DFF_444(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2403),.DATA(g33589));
  MSFF DFF_445(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2145),.DATA(g34605));
  MSFF DFF_446(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1700),.DATA(g30350));
  MSFF DFF_447(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g513),.DATA(g25611));
  MSFF DFF_448(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2841),.DATA(g26936));
  MSFF DFF_449(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5297),.DATA(g33619));
  MSFF DFF_450(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3805),.DATA(g3798));
  MSFF DFF_451(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2763),.DATA(g34022));
  MSFF DFF_452(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4793),.DATA(g34033));
  MSFF DFF_453(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g952),.DATA(g34726));
  MSFF DFF_454(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1263),.DATA(g31870));
  MSFF DFF_455(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1950),.DATA(g33985));
  MSFF DFF_456(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5138),.DATA(g29283));
  MSFF DFF_457(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2307),.DATA(g34003));
  MSFF DFF_458(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5109),.DATA(g5101));
  MSFF DFF_459(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5791),.DATA(g25727));
  MSFF DFF_460(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3798),.DATA(g25677));
  MSFF DFF_461(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4664),.DATA(g34463));
  MSFF DFF_462(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2223),.DATA(g33006));
  MSFF DFF_463(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5808),.DATA(g29292));
  MSFF DFF_464(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6645),.DATA(g30557));
  MSFF DFF_465(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2016),.DATA(g33989));
  MSFF DFF_466(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5759),.DATA(g28098));
  MSFF DFF_467(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3873),.DATA(g33033));
  MSFF DFF_468(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3632),.DATA(g3654));
  MSFF DFF_469(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2315),.DATA(g34005));
  MSFF DFF_470(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2811),.DATA(g26932));
  MSFF DFF_471(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5957),.DATA(g30516));
  MSFF DFF_472(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2047),.DATA(g33575));
  MSFF DFF_473(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3869),.DATA(g33032));
  MSFF DFF_474(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6358),.DATA(g6329));
  MSFF DFF_475(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3719),.DATA(g31891));
  MSFF DFF_476(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5575),.DATA(g30486));
  MSFF DFF_477(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g46),.DATA(g34991));
  MSFF DFF_478(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3752),.DATA(g25678));
  MSFF DFF_479(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3917),.DATA(g30440));
  MSFF DFF_480(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4188),.DATA(g4191));
  MSFF DFF_481(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1585),.DATA(g1570));
  MSFF DFF_482(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4388),.DATA(g26949));
  MSFF DFF_483(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6275),.DATA(g30530));
  MSFF DFF_484(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6311),.DATA(g30542));
  MSFF DFF_485(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4216),.DATA(g4213));
  MSFF DFF_486(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1041),.DATA(g25624));
  MSFF DFF_487(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2595),.DATA(g30383));
  MSFF DFF_488(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2537),.DATA(g33597));
  MSFF DFF_489(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g136),.DATA(g34598));
  MSFF DFF_490(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4430),.DATA(g26957));
  MSFF DFF_491(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4564),.DATA(g26967));
  MSFF DFF_492(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3454),.DATA(g3447));
  MSFF DFF_493(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4826),.DATA(g28102));
  MSFF DFF_494(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6239),.DATA(g30524));
  MSFF DFF_495(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3770),.DATA(g25671));
  MSFF DFF_496(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g232),.DATA(g26903));
  MSFF DFF_497(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5268),.DATA(g30475));
  MSFF DFF_498(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6545),.DATA(g34647));
  MSFF DFF_499(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2417),.DATA(g30377));
  MSFF DFF_500(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1772),.DATA(g33553));
  MSFF DFF_501(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4741),.DATA(g21902));
  MSFF DFF_502(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5052),.DATA(g31903));
  MSFF DFF_503(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5452),.DATA(g25715));
  MSFF DFF_504(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1890),.DATA(g33984));
  MSFF DFF_505(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2629),.DATA(g33602));
  MSFF DFF_506(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g572),.DATA(g28045));
  MSFF DFF_507(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2130),.DATA(g34603));
  MSFF DFF_508(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4108),.DATA(g33035));
  MSFF DFF_509(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4308),.DATA(g4304));
  MSFF DFF_510(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g475),.DATA(g24208));
  MSFF DFF_511(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g990),.DATA(g1239));
  MSFF DFF_512(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g31),.DATA(g34596));
  MSFF DFF_513(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3412),.DATA(g28064));
  MSFF DFF_514(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g45),.DATA(g34990));
  MSFF DFF_515(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g799),.DATA(g24213));
  MSFF DFF_516(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3706),.DATA(g31887));
  MSFF DFF_517(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3990),.DATA(g33614));
  MSFF DFF_518(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5385),.DATA(g31907));
  MSFF DFF_519(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5881),.DATA(g33060));
  MSFF DFF_520(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1992),.DATA(g30362));
  MSFF DFF_521(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3029),.DATA(g31875));
  MSFF DFF_522(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3171),.DATA(g33023));
  MSFF DFF_523(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3787),.DATA(g25674));
  MSFF DFF_524(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g812),.DATA(g26898));
  MSFF DFF_525(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g832),.DATA(g25618));
  MSFF DFF_526(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5897),.DATA(g30518));
  MSFF DFF_527(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4165),.DATA(g28079));
  MSFF DFF_528(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4571),.DATA(g6974));
  MSFF DFF_529(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3281),.DATA(g3303));
  MSFF DFF_530(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4455),.DATA(g26959));
  MSFF DFF_531(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2902),.DATA(g34801));
  MSFF DFF_532(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g333),.DATA(g26884));
  MSFF DFF_533(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g168),.DATA(g25600));
  MSFF DFF_534(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2823),.DATA(g26933));
  MSFF DFF_535(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3684),.DATA(g28066));
  MSFF DFF_536(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3639),.DATA(g33612));
  MSFF DFF_537(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5331),.DATA(g5327));
  MSFF DFF_538(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3338),.DATA(g24268));
  MSFF DFF_539(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5406),.DATA(g25716));
  MSFF DFF_540(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3791),.DATA(g25675));
  MSFF DFF_541(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g269),.DATA(g26906));
  MSFF DFF_542(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g401),.DATA(g24203));
  MSFF DFF_543(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6040),.DATA(g24346));
  MSFF DFF_544(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g441),.DATA(g24207));
  MSFF DFF_545(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5105),.DATA(g25701));
  MSFF DFF_546(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3808),.DATA(g29269));
  MSFF DFF_547(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g9),.DATA(g34592));
  MSFF DFF_548(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3759),.DATA(g28068));
  MSFF DFF_549(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4467),.DATA(g34255));
  MSFF DFF_550(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3957),.DATA(g30450));
  MSFF DFF_551(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4093),.DATA(g30456));
  MSFF DFF_552(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1760),.DATA(g32991));
  MSFF DFF_553(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6151),.DATA(g6144));
  MSFF DFF_554(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6351),.DATA(g24348));
  MSFF DFF_555(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g160),.DATA(g34249));
  MSFF DFF_556(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5445),.DATA(g25713));
  MSFF DFF_557(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5373),.DATA(g31909));
  MSFF DFF_558(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2279),.DATA(g30371));
  MSFF DFF_559(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3498),.DATA(g29268));
  MSFF DFF_560(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g586),.DATA(g29224));
  MSFF DFF_561(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g869),.DATA(g859));
  MSFF DFF_562(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2619),.DATA(g33017));
  MSFF DFF_563(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1183),.DATA(g30339));
  MSFF DFF_564(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1608),.DATA(g33967));
  MSFF DFF_565(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4197),.DATA(g4194));
  MSFF DFF_566(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5283),.DATA(g5276));
  MSFF DFF_567(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1779),.DATA(g33559));
  MSFF DFF_568(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2652),.DATA(g29255));
  MSFF DFF_569(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5459),.DATA(g5452));
  MSFF DFF_570(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2193),.DATA(g30368));
  MSFF DFF_571(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2393),.DATA(g30375));
  MSFF DFF_572(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5767),.DATA(g25732));
  MSFF DFF_573(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g661),.DATA(g28052));
  MSFF DFF_574(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4950),.DATA(g28089));
  MSFF DFF_575(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5535),.DATA(g33055));
  MSFF DFF_576(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2834),.DATA(g30392));
  MSFF DFF_577(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1361),.DATA(g30343));
  MSFF DFF_578(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3419),.DATA(g25657));
  MSFF DFF_579(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6235),.DATA(g30523));
  MSFF DFF_580(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1146),.DATA(g24233));
  MSFF DFF_581(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2625),.DATA(g33018));
  MSFF DFF_582(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g150),.DATA(g32976));
  MSFF DFF_583(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1696),.DATA(g30349));
  MSFF DFF_584(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6555),.DATA(g33067));
  MSFF DFF_585(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g859),.DATA(g26900));
  MSFF DFF_586(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3385),.DATA(g31883));
  MSFF DFF_587(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3881),.DATA(g33034));
  MSFF DFF_588(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6621),.DATA(g30551));
  MSFF DFF_589(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3470),.DATA(g25667));
  MSFF DFF_590(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3897),.DATA(g30452));
  MSFF DFF_591(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g518),.DATA(g25612));
  MSFF DFF_592(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3025),.DATA(g31874));
  MSFF DFF_593(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g538),.DATA(g34719));
  MSFF DFF_594(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2606),.DATA(g33607));
  MSFF DFF_595(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1472),.DATA(g26923));
  MSFF DFF_596(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6113),.DATA(g25746));
  MSFF DFF_597(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g542),.DATA(g24211));
  MSFF DFF_598(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5188),.DATA(g33050));
  MSFF DFF_599(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5689),.DATA(g24341));
  MSFF DFF_600(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1116),.DATA(g1056));
  MSFF DFF_601(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g405),.DATA(g24201));
  MSFF DFF_602(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5216),.DATA(g30463));
  MSFF DFF_603(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6494),.DATA(g6486));
  MSFF DFF_604(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4669),.DATA(g34464));
  MSFF DFF_605(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5428),.DATA(g25710));
  MSFF DFF_606(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g996),.DATA(g24243));
  MSFF DFF_607(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4531),.DATA(g24335));
  MSFF DFF_608(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2860),.DATA(g34611));
  MSFF DFF_609(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4743),.DATA(g34262));
  MSFF DFF_610(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6593),.DATA(g30546));
  MSFF DFF_611(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2710),.DATA(g18527));
  MSFF DFF_612(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g215),.DATA(g25591));
  MSFF DFF_613(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4411),.DATA(g4414));
  MSFF DFF_614(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1413),.DATA(g30347));
  MSFF DFF_615(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4474),.DATA(g10384));
  MSFF DFF_616(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5308),.DATA(g5283));
  MSFF DFF_617(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6641),.DATA(g30556));
  MSFF DFF_618(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3045),.DATA(g33020));
  MSFF DFF_619(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6),.DATA(g34589));
  MSFF DFF_620(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1936),.DATA(g33562));
  MSFF DFF_621(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g55),.DATA(g35002));
  MSFF DFF_622(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g504),.DATA(g25610));
  MSFF DFF_623(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2587),.DATA(g33015));
  MSFF DFF_624(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4480),.DATA(g31896));
  MSFF DFF_625(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2311),.DATA(g34004));
  MSFF DFF_626(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3602),.DATA(g30428));
  MSFF DFF_627(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5571),.DATA(g30485));
  MSFF DFF_628(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3578),.DATA(g30422));
  MSFF DFF_629(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g468),.DATA(g25606));
  MSFF DFF_630(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5448),.DATA(g25714));
  MSFF DFF_631(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3767),.DATA(g25680));
  MSFF DFF_632(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5827),.DATA(g29294));
  MSFF DFF_633(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3582),.DATA(g30423));
  MSFF DFF_634(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6271),.DATA(g30529));
  MSFF DFF_635(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4688),.DATA(g34028));
  MSFF DFF_636(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5774),.DATA(g25724));
  MSFF DFF_637(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2380),.DATA(g33587));
  MSFF DFF_638(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5196),.DATA(g30460));
  MSFF DFF_639(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5396),.DATA(g31910));
  MSFF DFF_640(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3227),.DATA(g30401));
  MSFF DFF_641(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2020),.DATA(g33990));
  MSFF DFF_642(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4000),.DATA(g3976));
  MSFF DFF_643(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1079),.DATA(g1075));
  MSFF DFF_644(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6541),.DATA(g29309));
  MSFF DFF_645(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3203),.DATA(g30411));
  MSFF DFF_646(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1668),.DATA(g33546));
  MSFF DFF_647(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4760),.DATA(g28085));
  MSFF DFF_648(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g262),.DATA(g26904));
  MSFF DFF_649(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1840),.DATA(g33556));
  MSFF DFF_650(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g70),.DATA(g18093));
  MSFF DFF_651(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5467),.DATA(g25722));
  MSFF DFF_652(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g460),.DATA(g25605));
  MSFF DFF_653(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6209),.DATA(g33062));
  MSFF DFF_654(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g74),.DATA(g26893));
  MSFF DFF_655(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5290),.DATA(g5313));
  MSFF DFF_656(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g655),.DATA(g28050));
  MSFF DFF_657(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3502),.DATA(g34626));
  MSFF DFF_658(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2204),.DATA(g33583));
  MSFF DFF_659(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5256),.DATA(g30472));
  MSFF DFF_660(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4608),.DATA(g34454));
  MSFF DFF_661(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g794),.DATA(g34850));
  MSFF DFF_662(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4023),.DATA(g4019));
  MSFF DFF_663(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4423),.DATA(g4537));
  MSFF DFF_664(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3689),.DATA(g24272));
  MSFF DFF_665(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5381),.DATA(g31906));
  MSFF DFF_666(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5685),.DATA(g5681));
  MSFF DFF_667(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g703),.DATA(g24214));
  MSFF DFF_668(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5421),.DATA(g25718));
  MSFF DFF_669(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g862),.DATA(g26909));
  MSFF DFF_670(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3247),.DATA(g30406));
  MSFF DFF_671(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2040),.DATA(g33569));
  MSFF DFF_672(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4999),.DATA(g25694));
  MSFF DFF_673(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4146),.DATA(g34628));
  MSFF DFF_674(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4633),.DATA(g34458));
  MSFF DFF_675(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1157),.DATA(g24240));
  MSFF DFF_676(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5723),.DATA(g31918));
  MSFF DFF_677(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4732),.DATA(g34634));
  MSFF DFF_678(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5101),.DATA(g25700));
  MSFF DFF_679(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5817),.DATA(g29293));
  MSFF DFF_680(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2151),.DATA(g18421));
  MSFF DFF_681(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2351),.DATA(g33009));
  MSFF DFF_682(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2648),.DATA(g33603));
  MSFF DFF_683(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6736),.DATA(g24355));
  MSFF DFF_684(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4944),.DATA(g34268));
  MSFF DFF_685(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4072),.DATA(g25691));
  MSFF DFF_686(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g344),.DATA(g26890));
  MSFF DFF_687(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4443),.DATA(g4449));
  MSFF DFF_688(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3466),.DATA(g29264));
  MSFF DFF_689(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4116),.DATA(g28072));
  MSFF DFF_690(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5041),.DATA(g31900));
  MSFF DFF_691(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5441),.DATA(g25712));
  MSFF DFF_692(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4434),.DATA(g26956));
  MSFF DFF_693(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3827),.DATA(g29271));
  MSFF DFF_694(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6500),.DATA(g29304));
  MSFF DFF_695(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5673),.DATA(g5654));
  MSFF DFF_696(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3133),.DATA(g29261));
  MSFF DFF_697(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3333),.DATA(g28063));
  MSFF DFF_698(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g979),.DATA(g1116));
  MSFF DFF_699(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4681),.DATA(g34027));
  MSFF DFF_700(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g298),.DATA(g33961));
  MSFF DFF_701(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3774),.DATA(g25672));
  MSFF DFF_702(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2667),.DATA(g33604));
  MSFF DFF_703(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3396),.DATA(g33025));
  MSFF DFF_704(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4210),.DATA(g4207));
  MSFF DFF_705(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1894),.DATA(g32995));
  MSFF DFF_706(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2988),.DATA(g34624));
  MSFF DFF_707(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3538),.DATA(g30415));
  MSFF DFF_708(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g301),.DATA(g33536));
  MSFF DFF_709(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g341),.DATA(g26888));
  MSFF DFF_710(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g827),.DATA(g28055));
  MSFF DFF_711(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1075),.DATA(g24238));
  MSFF DFF_712(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6077),.DATA(g31921));
  MSFF DFF_713(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2555),.DATA(g33600));
  MSFF DFF_714(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5011),.DATA(g28105));
  MSFF DFF_715(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g199),.DATA(g34721));
  MSFF DFF_716(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6523),.DATA(g29307));
  MSFF DFF_717(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1526),.DATA(g30345));
  MSFF DFF_718(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4601),.DATA(g34453));
  MSFF DFF_719(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g854),.DATA(g32980));
  MSFF DFF_720(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1484),.DATA(g29238));
  MSFF DFF_721(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4922),.DATA(g34639));
  MSFF DFF_722(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5080),.DATA(g25695));
  MSFF DFF_723(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5863),.DATA(g33057));
  MSFF DFF_724(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4581),.DATA(g26969));
  MSFF DFF_725(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3021),.DATA(g31879));
  MSFF DFF_726(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2518),.DATA(g29253));
  MSFF DFF_727(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2567),.DATA(g34021));
  MSFF DFF_728(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g568),.DATA(g26895));
  MSFF DFF_729(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3263),.DATA(g30413));
  MSFF DFF_730(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6613),.DATA(g30549));
  MSFF DFF_731(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6044),.DATA(g24347));
  MSFF DFF_732(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6444),.DATA(g25758));
  MSFF DFF_733(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2965),.DATA(g34808));
  MSFF DFF_734(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5857),.DATA(g30501));
  MSFF DFF_735(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1616),.DATA(g33969));
  MSFF DFF_736(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g890),.DATA(g34440));
  MSFF DFF_737(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5976),.DATA(g5969));
  MSFF DFF_738(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3562),.DATA(g30433));
  MSFF DFF_739(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4294),.DATA(g21900));
  MSFF DFF_740(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1404),.DATA(g26921));
  MSFF DFF_741(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3723),.DATA(g31893));
  MSFF DFF_742(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3817),.DATA(g29270));
  MSFF DFF_743(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g93),.DATA(g34878));
  MSFF DFF_744(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4501),.DATA(g33038));
  MSFF DFF_745(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g287),.DATA(g31865));
  MSFF DFF_746(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2724),.DATA(g26926));
  MSFF DFF_747(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4704),.DATA(g28083));
  MSFF DFF_748(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g22),.DATA(g29209));
  MSFF DFF_749(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2878),.DATA(g34797));
  MSFF DFF_750(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5220),.DATA(g30478));
  MSFF DFF_751(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g617),.DATA(g34724));
  MSFF DFF_752(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g637),.DATA(g24212));
  MSFF DFF_753(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g316),.DATA(g26883));
  MSFF DFF_754(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1277),.DATA(g32985));
  MSFF DFF_755(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6513),.DATA(g25761));
  MSFF DFF_756(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g336),.DATA(g26886));
  MSFF DFF_757(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2882),.DATA(g34796));
  MSFF DFF_758(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g933),.DATA(g32982));
  MSFF DFF_759(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1906),.DATA(g33561));
  MSFF DFF_760(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g305),.DATA(g26880));
  MSFF DFF_761(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g8),.DATA(g34591));
  MSFF DFF_762(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3368),.DATA(g31884));
  MSFF DFF_763(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2799),.DATA(g26931));
  MSFF DFF_764(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g887),.DATA(g884));
  MSFF DFF_765(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5327),.DATA(g5308));
  MSFF DFF_766(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4912),.DATA(g34641));
  MSFF DFF_767(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4157),.DATA(g34629));
  MSFF DFF_768(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2541),.DATA(g33598));
  MSFF DFF_769(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2153),.DATA(g33576));
  MSFF DFF_770(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g550),.DATA(g34720));
  MSFF DFF_771(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g255),.DATA(g26902));
  MSFF DFF_772(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1945),.DATA(g29244));
  MSFF DFF_773(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5240),.DATA(g30468));
  MSFF DFF_774(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1478),.DATA(g26924));
  MSFF DFF_775(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3080),.DATA(g25645));
  MSFF DFF_776(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3863),.DATA(g33031));
  MSFF DFF_777(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1959),.DATA(g29245));
  MSFF DFF_778(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3480),.DATA(g29266));
  MSFF DFF_779(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6653),.DATA(g30559));
  MSFF DFF_780(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6719),.DATA(g6715));
  MSFF DFF_781(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2864),.DATA(g34794));
  MSFF DFF_782(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4894),.DATA(g28087));
  MSFF DFF_783(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5681),.DATA(g5677));
  MSFF DFF_784(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3857),.DATA(g30435));
  MSFF DFF_785(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3976),.DATA(g3969));
  MSFF DFF_786(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g499),.DATA(g25609));
  MSFF DFF_787(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5413),.DATA(g28095));
  MSFF DFF_788(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1002),.DATA(g28057));
  MSFF DFF_789(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g776),.DATA(g34439));
  MSFF DFF_790(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g28),.DATA(g34595));
  MSFF DFF_791(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1236),.DATA(g1233));
  MSFF DFF_792(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4646),.DATA(g34260));
  MSFF DFF_793(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2476),.DATA(g33012));
  MSFF DFF_794(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1657),.DATA(g32989));
  MSFF DFF_795(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2375),.DATA(g34006));
  MSFF DFF_796(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g63),.DATA(g34847));
  MSFF DFF_797(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6012),.DATA(g5983));
  MSFF DFF_798(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g358),.DATA(g365));
  MSFF DFF_799(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g896),.DATA(g26910));
  MSFF DFF_800(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g967),.DATA(g21722));
  MSFF DFF_801(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3423),.DATA(g25658));
  MSFF DFF_802(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g283),.DATA(g28043));
  MSFF DFF_803(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3161),.DATA(g33021));
  MSFF DFF_804(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2384),.DATA(g29251));
  MSFF DFF_805(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3361),.DATA(g25665));
  MSFF DFF_806(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6675),.DATA(g6697));
  MSFF DFF_807(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4616),.DATA(g34456));
  MSFF DFF_808(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4561),.DATA(g26968));
  MSFF DFF_809(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2024),.DATA(g33991));
  MSFF DFF_810(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3451),.DATA(g3443));
  MSFF DFF_811(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2795),.DATA(g26930));
  MSFF DFF_812(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g613),.DATA(g34599));
  MSFF DFF_813(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4527),.DATA(g28082));
  MSFF DFF_814(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1844),.DATA(g33557));
  MSFF DFF_815(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5937),.DATA(g30511));
  MSFF DFF_816(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4546),.DATA(g33045));
  MSFF DFF_817(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3103),.DATA(g3096));
  MSFF DFF_818(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2523),.DATA(g30379));
  MSFF DFF_819(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3303),.DATA(g24267));
  MSFF DFF_820(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2643),.DATA(g34020));
  MSFF DFF_821(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6109),.DATA(g28100));
  MSFF DFF_822(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1489),.DATA(g24249));
  MSFF DFF_823(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5390),.DATA(g31908));
  MSFF DFF_824(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g194),.DATA(g25592));
  MSFF DFF_825(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2551),.DATA(g30382));
  MSFF DFF_826(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5156),.DATA(g29285));
  MSFF DFF_827(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3072),.DATA(g25644));
  MSFF DFF_828(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1242),.DATA(g1227));
  MSFF DFF_829(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g47),.DATA(g34992));
  MSFF DFF_830(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3443),.DATA(g25662));
  MSFF DFF_831(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4277),.DATA(g21896));
  MSFF DFF_832(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1955),.DATA(g33563));
  MSFF DFF_833(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6049),.DATA(g33622));
  MSFF DFF_834(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3034),.DATA(g31876));
  MSFF DFF_835(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2273),.DATA(g33582));
  MSFF DFF_836(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6715),.DATA(g6711));
  MSFF DFF_837(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4771),.DATA(g28086));
  MSFF DFF_838(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6098),.DATA(g25744));
  MSFF DFF_839(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3147),.DATA(g29262));
  MSFF DFF_840(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3347),.DATA(g24270));
  MSFF DFF_841(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2269),.DATA(g33581));
  MSFF DFF_842(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g191),.DATA(g194));
  MSFF DFF_843(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2712),.DATA(g26937));
  MSFF DFF_844(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g626),.DATA(g34849));
  MSFF DFF_845(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2729),.DATA(g28060));
  MSFF DFF_846(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5357),.DATA(g33618));
  MSFF DFF_847(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4991),.DATA(g34038));
  MSFF DFF_848(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6019),.DATA(g6000));
  MSFF DFF_849(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4709),.DATA(g34032));
  MSFF DFF_850(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6419),.DATA(g31927));
  MSFF DFF_851(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6052),.DATA(g31919));
  MSFF DFF_852(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2927),.DATA(g34803));
  MSFF DFF_853(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4340),.DATA(g34459));
  MSFF DFF_854(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5929),.DATA(g30509));
  MSFF DFF_855(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4907),.DATA(g34640));
  MSFF DFF_856(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3317),.DATA(g3298));
  MSFF DFF_857(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4035),.DATA(g28069));
  MSFF DFF_858(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2946),.DATA(g21899));
  MSFF DFF_859(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g918),.DATA(g31868));
  MSFF DFF_860(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4082),.DATA(g26938));
  MSFF DFF_861(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6486),.DATA(g25756));
  MSFF DFF_862(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2036),.DATA(g30363));
  MSFF DFF_863(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g577),.DATA(g30334));
  MSFF DFF_864(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1620),.DATA(g33970));
  MSFF DFF_865(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2831),.DATA(g30391));
  MSFF DFF_866(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g667),.DATA(g25615));
  MSFF DFF_867(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g930),.DATA(g33540));
  MSFF DFF_868(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3937),.DATA(g30445));
  MSFF DFF_869(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5782),.DATA(g25725));
  MSFF DFF_870(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g817),.DATA(g25617));
  MSFF DFF_871(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1249),.DATA(g24247));
  MSFF DFF_872(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g837),.DATA(g24215));
  MSFF DFF_873(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3668),.DATA(g3649));
  MSFF DFF_874(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g599),.DATA(g33964));
  MSFF DFF_875(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5475),.DATA(g25719));
  MSFF DFF_876(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g739),.DATA(g29228));
  MSFF DFF_877(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5949),.DATA(g30514));
  MSFF DFF_878(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6682),.DATA(g33627));
  MSFF DFF_879(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6105),.DATA(g28101));
  MSFF DFF_880(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g904),.DATA(g24231));
  MSFF DFF_881(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2873),.DATA(g34615));
  MSFF DFF_882(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1854),.DATA(g30356));
  MSFF DFF_883(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5084),.DATA(g25696));
  MSFF DFF_884(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5603),.DATA(g30493));
  MSFF DFF_885(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4222),.DATA(g4219));
  MSFF DFF_886(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2495),.DATA(g33594));
  MSFF DFF_887(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2437),.DATA(g34009));
  MSFF DFF_888(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2102),.DATA(g30365));
  MSFF DFF_889(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2208),.DATA(g33004));
  MSFF DFF_890(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2579),.DATA(g34018));
  MSFF DFF_891(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4064),.DATA(g25685));
  MSFF DFF_892(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4899),.DATA(g34040));
  MSFF DFF_893(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2719),.DATA(g25639));
  MSFF DFF_894(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4785),.DATA(g34029));
  MSFF DFF_895(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5583),.DATA(g30488));
  MSFF DFF_896(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g781),.DATA(g34600));
  MSFF DFF_897(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6173),.DATA(g29300));
  MSFF DFF_898(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6373),.DATA(g6369));
  MSFF DFF_899(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2917),.DATA(g34802));
  MSFF DFF_900(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g686),.DATA(g25614));
  MSFF DFF_901(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1252),.DATA(g28058));
  MSFF DFF_902(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g671),.DATA(g29225));
  MSFF DFF_903(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2265),.DATA(g33580));
  MSFF DFF_904(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6283),.DATA(g30532));
  MSFF DFF_905(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6369),.DATA(g6365));
  MSFF DFF_906(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5276),.DATA(g5320));
  MSFF DFF_907(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6459),.DATA(g25760));
  MSFF DFF_908(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g901),.DATA(g25620));
  MSFF DFF_909(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4194),.DATA(g4188));
  MSFF DFF_910(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5527),.DATA(g33054));
  MSFF DFF_911(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4489),.DATA(g26962));
  MSFF DFF_912(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1974),.DATA(g33564));
  MSFF DFF_913(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1270),.DATA(g32984));
  MSFF DFF_914(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4966),.DATA(g34039));
  MSFF DFF_915(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6415),.DATA(g31932));
  MSFF DFF_916(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6227),.DATA(g33065));
  MSFF DFF_917(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3929),.DATA(g30443));
  MSFF DFF_918(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5503),.DATA(g29291));
  MSFF DFF_919(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4242),.DATA(g24279));
  MSFF DFF_920(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5925),.DATA(g30508));
  MSFF DFF_921(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1124),.DATA(g29232));
  MSFF DFF_922(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4955),.DATA(g34269));
  MSFF DFF_923(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5224),.DATA(g30464));
  MSFF DFF_924(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2012),.DATA(g33988));
  MSFF DFF_925(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6203),.DATA(g30522));
  MSFF DFF_926(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5120),.DATA(g25708));
  MSFF DFF_927(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5320),.DATA(g5290));
  MSFF DFF_928(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2389),.DATA(g30374));
  MSFF DFF_929(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4438),.DATA(g26953));
  MSFF DFF_930(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2429),.DATA(g34008));
  MSFF DFF_931(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2787),.DATA(g34444));
  MSFF DFF_932(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1287),.DATA(g34731));
  MSFF DFF_933(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2675),.DATA(g33606));
  MSFF DFF_934(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g66),.DATA(g24334));
  MSFF DFF_935(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4836),.DATA(g34265));
  MSFF DFF_936(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1199),.DATA(g30340));
  MSFF DFF_937(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1399),.DATA(g24257));
  MSFF DFF_938(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5547),.DATA(g30482));
  MSFF DFF_939(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3782),.DATA(g25673));
  MSFF DFF_940(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6428),.DATA(g31929));
  MSFF DFF_941(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2138),.DATA(g34604));
  MSFF DFF_942(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3661),.DATA(g3632));
  MSFF DFF_943(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2338),.DATA(g33591));
  MSFF DFF_944(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4229),.DATA(g4226));
  MSFF DFF_945(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6247),.DATA(g30525));
  MSFF DFF_946(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2791),.DATA(g26929));
  MSFF DFF_947(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3949),.DATA(g30448));
  MSFF DFF_948(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1291),.DATA(g34602));
  MSFF DFF_949(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5945),.DATA(g30513));
  MSFF DFF_950(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5244),.DATA(g30469));
  MSFF DFF_951(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2759),.DATA(g33608));
  MSFF DFF_952(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6741),.DATA(g33626));
  MSFF DFF_953(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g785),.DATA(g34725));
  MSFF DFF_954(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1259),.DATA(g30342));
  MSFF DFF_955(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3484),.DATA(g29267));
  MSFF DFF_956(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g209),.DATA(g25593));
  MSFF DFF_957(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6609),.DATA(g30548));
  MSFF DFF_958(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5517),.DATA(g33052));
  MSFF DFF_959(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2449),.DATA(g34012));
  MSFF DFF_960(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2575),.DATA(g34017));
  MSFF DFF_961(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g65),.DATA(g34785));
  MSFF DFF_962(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2715),.DATA(g24263));
  MSFF DFF_963(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g936),.DATA(g26912));
  MSFF DFF_964(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2098),.DATA(g30364));
  MSFF DFF_965(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4462),.DATA(g34254));
  MSFF DFF_966(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g604),.DATA(g34251));
  MSFF DFF_967(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6589),.DATA(g30560));
  MSFF DFF_968(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1886),.DATA(g33983));
  MSFF DFF_969(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6466),.DATA(g25752));
  MSFF DFF_970(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6365),.DATA(g6346));
  MSFF DFF_971(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6711),.DATA(g6692));
  MSFF DFF_972(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g429),.DATA(g24204));
  MSFF DFF_973(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1870),.DATA(g33980));
  MSFF DFF_974(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4249),.DATA(g34631));
  MSFF DFF_975(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6455),.DATA(g28103));
  MSFF DFF_976(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3004),.DATA(g31873));
  MSFF DFF_977(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1825),.DATA(g29243));
  MSFF DFF_978(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6133),.DATA(g25740));
  MSFF DFF_979(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1008),.DATA(g25623));
  MSFF DFF_980(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4392),.DATA(g26950));
  MSFF DFF_981(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5002),.DATA(g4999));
  MSFF DFF_982(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3546),.DATA(g30431));
  MSFF DFF_983(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5236),.DATA(g30467));
  MSFF DFF_984(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1768),.DATA(g30353));
  MSFF DFF_985(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4854),.DATA(g34467));
  MSFF DFF_986(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3925),.DATA(g30442));
  MSFF DFF_987(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6509),.DATA(g29305));
  MSFF DFF_988(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g732),.DATA(g25616));
  MSFF DFF_989(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2504),.DATA(g29252));
  MSFF DFF_990(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1322),.DATA(g1459));
  MSFF DFF_991(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4520),.DATA(g6972));
  MSFF DFF_992(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4219),.DATA(g4216));
  MSFF DFF_993(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2185),.DATA(g33003));
  MSFF DFF_994(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g37),.DATA(g34613));
  MSFF DFF_995(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4031),.DATA(g4027));
  MSFF DFF_996(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2070),.DATA(g33570));
  MSFF DFF_997(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4812),.DATA(g4809));
  MSFF DFF_998(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6093),.DATA(g33061));
  MSFF DFF_999(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g968),.DATA(g21723));
  MSFF DFF_1000(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4176),.DATA(g34734));
  MSFF DFF_1001(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4005),.DATA(g24275));
  MSFF DFF_1002(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4405),.DATA(g4408));
  MSFF DFF_1003(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g872),.DATA(g887));
  MSFF DFF_1004(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6181),.DATA(g29302));
  MSFF DFF_1005(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6381),.DATA(g24349));
  MSFF DFF_1006(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4765),.DATA(g34264));
  MSFF DFF_1007(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5563),.DATA(g30484));
  MSFF DFF_1008(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1395),.DATA(g25634));
  MSFF DFF_1009(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1913),.DATA(g33567));
  MSFF DFF_1010(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2331),.DATA(g33585));
  MSFF DFF_1011(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6263),.DATA(g30527));
  MSFF DFF_1012(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g50),.DATA(g34995));
  MSFF DFF_1013(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3945),.DATA(g30447));
  MSFF DFF_1014(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g347),.DATA(g344));
  MSFF DFF_1015(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5731),.DATA(g31914));
  MSFF DFF_1016(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4473),.DATA(g34256));
  MSFF DFF_1017(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1266),.DATA(g25630));
  MSFF DFF_1018(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5489),.DATA(g29290));
  MSFF DFF_1019(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g714),.DATA(g29227));
  MSFF DFF_1020(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2748),.DATA(g31872));
  MSFF DFF_1021(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5471),.DATA(g29287));
  MSFF DFF_1022(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4540),.DATA(g31897));
  MSFF DFF_1023(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6723),.DATA(g6719));
  MSFF DFF_1024(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6605),.DATA(g30562));
  MSFF DFF_1025(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2445),.DATA(g34011));
  MSFF DFF_1026(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2173),.DATA(g33996));
  MSFF DFF_1027(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4287),.DATA(g21898));
  MSFF DFF_1028(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2491),.DATA(g33014));
  MSFF DFF_1029(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4849),.DATA(g34465));
  MSFF DFF_1030(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2169),.DATA(g33995));
  MSFF DFF_1031(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2283),.DATA(g30372));
  MSFF DFF_1032(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6585),.DATA(g30545));
  MSFF DFF_1033(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g121),.DATA(g30389));
  MSFF DFF_1034(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2407),.DATA(g33590));
  MSFF DFF_1035(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2868),.DATA(g34616));
  MSFF DFF_1036(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2767),.DATA(g26927));
  MSFF DFF_1037(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1783),.DATA(g32992));
  MSFF DFF_1038(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3310),.DATA(g3281));
  MSFF DFF_1039(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1312),.DATA(g25631));
  MSFF DFF_1040(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5212),.DATA(g30477));
  MSFF DFF_1041(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4245),.DATA(g34632));
  MSFF DFF_1042(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g645),.DATA(g28046));
  MSFF DFF_1043(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4291),.DATA(g4287));
  MSFF DFF_1044(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g79),.DATA(g26896));
  MSFF DFF_1045(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g182),.DATA(g25602));
  MSFF DFF_1046(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1129),.DATA(g26916));
  MSFF DFF_1047(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2227),.DATA(g33578));
  MSFF DFF_1048(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6058),.DATA(g25745));
  MSFF DFF_1049(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4207),.DATA(g4204));
  MSFF DFF_1050(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2246),.DATA(g33579));
  MSFF DFF_1051(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1830),.DATA(g30354));
  MSFF DFF_1052(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3590),.DATA(g30425));
  MSFF DFF_1053(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g392),.DATA(g24200));
  MSFF DFF_1054(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1592),.DATA(g33544));
  MSFF DFF_1055(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6505),.DATA(g25764));
  MSFF DFF_1056(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6411),.DATA(g31930));
  MSFF DFF_1057(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1221),.DATA(g24246));
  MSFF DFF_1058(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5921),.DATA(g30507));
  MSFF DFF_1059(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g106),.DATA(g26889));
  MSFF DFF_1060(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g146),.DATA(g30333));
  MSFF DFF_1061(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g218),.DATA(g215));
  MSFF DFF_1062(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6474),.DATA(g25753));
  MSFF DFF_1063(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1932),.DATA(g32998));
  MSFF DFF_1064(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1624),.DATA(g32987));
  MSFF DFF_1065(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5062),.DATA(g25702));
  MSFF DFF_1066(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5462),.DATA(g29286));
  MSFF DFF_1067(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2689),.DATA(g34606));
  MSFF DFF_1068(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6573),.DATA(g33070));
  MSFF DFF_1069(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1677),.DATA(g29240));
  MSFF DFF_1070(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2028),.DATA(g32999));
  MSFF DFF_1071(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2671),.DATA(g33605));
  MSFF DFF_1072(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1576),.DATA(g24255));
  MSFF DFF_1073(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4408),.DATA(g26945));
  MSFF DFF_1074(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g34),.DATA(g34877));
  MSFF DFF_1075(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1848),.DATA(g33558));
  MSFF DFF_1076(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3089),.DATA(g25647));
  MSFF DFF_1077(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3731),.DATA(g31889));
  MSFF DFF_1078(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g86),.DATA(g25699));
  MSFF DFF_1079(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5485),.DATA(g29289));
  MSFF DFF_1080(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2741),.DATA(g30388));
  MSFF DFF_1081(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g802),.DATA(g799));
  MSFF DFF_1082(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2638),.DATA(g29254));
  MSFF DFF_1083(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4122),.DATA(g28074));
  MSFF DFF_1084(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4322),.DATA(g34450));
  MSFF DFF_1085(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5941),.DATA(g30512));
  MSFF DFF_1086(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2108),.DATA(g33572));
  MSFF DFF_1087(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6000),.DATA(g5976));
  MSFF DFF_1088(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g25),.DATA(g15048));
  MSFF DFF_1089(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1644),.DATA(g33551));
  MSFF DFF_1090(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g595),.DATA(g33538));
  MSFF DFF_1091(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2217),.DATA(g33005));
  MSFF DFF_1092(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1319),.DATA(g24248));
  MSFF DFF_1093(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2066),.DATA(g33002));
  MSFF DFF_1094(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1152),.DATA(g24234));
  MSFF DFF_1095(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5252),.DATA(g30471));
  MSFF DFF_1096(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2165),.DATA(g34000));
  MSFF DFF_1097(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2571),.DATA(g34016));
  MSFF DFF_1098(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5176),.DATA(g33048));
  MSFF DFF_1099(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g391),.DATA(g26911));
  MSFF DFF_1100(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5005),.DATA(g5002));
  MSFF DFF_1101(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2711),.DATA(g18528));
  MSFF DFF_1102(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6023),.DATA(g6019));
  MSFF DFF_1103(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1211),.DATA(g25628));
  MSFF DFF_1104(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2827),.DATA(g26934));
  MSFF DFF_1105(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6423),.DATA(g31928));
  MSFF DFF_1106(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g875),.DATA(g869));
  MSFF DFF_1107(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4859),.DATA(g34468));
  MSFF DFF_1108(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g424),.DATA(g24202));
  MSFF DFF_1109(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1274),.DATA(g33542));
  MSFF DFF_1110(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1426),.DATA(g1422));
  MSFF DFF_1111(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g85),.DATA(g34717));
  MSFF DFF_1112(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2803),.DATA(g34445));
  MSFF DFF_1113(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6451),.DATA(g28104));
  MSFF DFF_1114(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1821),.DATA(g33555));
  MSFF DFF_1115(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2509),.DATA(g34013));
  MSFF DFF_1116(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5073),.DATA(g28091));
  MSFF DFF_1117(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1280),.DATA(g26919));
  MSFF DFF_1118(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4815),.DATA(g4812));
  MSFF DFF_1119(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6346),.DATA(g6322));
  MSFF DFF_1120(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6633),.DATA(g30554));
  MSFF DFF_1121(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5124),.DATA(g29281));
  MSFF DFF_1122(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1083),.DATA(g1079));
  MSFF DFF_1123(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6303),.DATA(g30537));
  MSFF DFF_1124(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5069),.DATA(g28092));
  MSFF DFF_1125(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2994),.DATA(g34732));
  MSFF DFF_1126(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g650),.DATA(g28049));
  MSFF DFF_1127(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1636),.DATA(g33545));
  MSFF DFF_1128(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3921),.DATA(g30441));
  MSFF DFF_1129(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2093),.DATA(g29247));
  MSFF DFF_1130(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6732),.DATA(g24354));
  MSFF DFF_1131(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1306),.DATA(g25636));
  MSFF DFF_1132(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5377),.DATA(g31911));
  MSFF DFF_1133(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1061),.DATA(g26914));
  MSFF DFF_1134(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3462),.DATA(g25670));
  MSFF DFF_1135(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2181),.DATA(g33998));
  MSFF DFF_1136(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g956),.DATA(g25626));
  MSFF DFF_1137(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1756),.DATA(g33977));
  MSFF DFF_1138(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5849),.DATA(g29297));
  MSFF DFF_1139(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4112),.DATA(g28071));
  MSFF DFF_1140(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2685),.DATA(g30387));
  MSFF DFF_1141(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2197),.DATA(g33577));
  MSFF DFF_1142(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6116),.DATA(g25737));
  MSFF DFF_1143(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2421),.DATA(g33592));
  MSFF DFF_1144(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1046),.DATA(g26913));
  MSFF DFF_1145(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g482),.DATA(g28044));
  MSFF DFF_1146(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4401),.DATA(g26948));
  MSFF DFF_1147(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6434),.DATA(g31931));
  MSFF DFF_1148(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1514),.DATA(g30344));
  MSFF DFF_1149(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g329),.DATA(g26885));
  MSFF DFF_1150(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6565),.DATA(g33069));
  MSFF DFF_1151(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2950),.DATA(g34621));
  MSFF DFF_1152(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4129),.DATA(g28075));
  MSFF DFF_1153(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1345),.DATA(g28059));
  MSFF DFF_1154(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6533),.DATA(g25762));
  MSFF DFF_1155(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3298),.DATA(g3274));
  MSFF DFF_1156(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3085),.DATA(g25646));
  MSFF DFF_1157(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4727),.DATA(g34633));
  MSFF DFF_1158(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6697),.DATA(g24352));
  MSFF DFF_1159(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1536),.DATA(g26925));
  MSFF DFF_1160(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3941),.DATA(g30446));
  MSFF DFF_1161(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g370),.DATA(g25597));
  MSFF DFF_1162(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5694),.DATA(g24342));
  MSFF DFF_1163(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1858),.DATA(g30357));
  MSFF DFF_1164(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g446),.DATA(g26908));
  MSFF DFF_1165(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4932),.DATA(g21905));
  MSFF DFF_1166(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3219),.DATA(g30399));
  MSFF DFF_1167(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1811),.DATA(g29242));
  MSFF DFF_1168(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3431),.DATA(g25659));
  MSFF DFF_1169(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6601),.DATA(g30547));
  MSFF DFF_1170(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3376),.DATA(g31881));
  MSFF DFF_1171(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2441),.DATA(g34010));
  MSFF DFF_1172(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1874),.DATA(g33986));
  MSFF DFF_1173(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4349),.DATA(g34257));
  MSFF DFF_1174(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6581),.DATA(g30544));
  MSFF DFF_1175(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6597),.DATA(g30561));
  MSFF DFF_1176(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5008),.DATA(g5005));
  MSFF DFF_1177(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3610),.DATA(g30430));
  MSFF DFF_1178(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2890),.DATA(g34799));
  MSFF DFF_1179(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1978),.DATA(g33565));
  MSFF DFF_1180(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1612),.DATA(g33968));
  MSFF DFF_1181(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g112),.DATA(g34879));
  MSFF DFF_1182(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2856),.DATA(g34793));
  MSFF DFF_1183(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6479),.DATA(g25754));
  MSFF DFF_1184(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1982),.DATA(g33566));
  MSFF DFF_1185(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6668),.DATA(g6661));
  MSFF DFF_1186(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5228),.DATA(g30465));
  MSFF DFF_1187(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4119),.DATA(g28073));
  MSFF DFF_1188(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6390),.DATA(g24351));
  MSFF DFF_1189(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1542),.DATA(g30346));
  MSFF DFF_1190(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4258),.DATA(g21893));
  MSFF DFF_1191(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4818),.DATA(g4815));
  MSFF DFF_1192(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5033),.DATA(g31904));
  MSFF DFF_1193(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4717),.DATA(g34635));
  MSFF DFF_1194(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1554),.DATA(g25637));
  MSFF DFF_1195(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3849),.DATA(g29274));
  MSFF DFF_1196(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6704),.DATA(g6675));
  MSFF DFF_1197(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3199),.DATA(g30396));
  MSFF DFF_1198(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5845),.DATA(g25735));
  MSFF DFF_1199(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4975),.DATA(g34037));
  MSFF DFF_1200(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g790),.DATA(g34791));
  MSFF DFF_1201(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5913),.DATA(g30520));
  MSFF DFF_1202(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1902),.DATA(g30358));
  MSFF DFF_1203(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6163),.DATA(g29299));
  MSFF DFF_1204(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4125),.DATA(g28081));
  MSFF DFF_1205(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4821),.DATA(g28096));
  MSFF DFF_1206(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4939),.DATA(g28088));
  MSFF DFF_1207(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1056),.DATA(g24241));
  MSFF DFF_1208(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3207),.DATA(g30397));
  MSFF DFF_1209(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4483),.DATA(g4520));
  MSFF DFF_1210(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3259),.DATA(g30409));
  MSFF DFF_1211(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5142),.DATA(g29284));
  MSFF DFF_1212(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5248),.DATA(g30470));
  MSFF DFF_1213(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2126),.DATA(g30367));
  MSFF DFF_1214(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3694),.DATA(g24273));
  MSFF DFF_1215(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5481),.DATA(g29288));
  MSFF DFF_1216(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1964),.DATA(g30359));
  MSFF DFF_1217(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5097),.DATA(g25698));
  MSFF DFF_1218(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3215),.DATA(g30398));
  MSFF DFF_1219(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4027),.DATA(g4023));
  MSFF DFF_1220(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g111),.DATA(g34718));
  MSFF DFF_1221(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4427),.DATA(g26952));
  MSFF DFF_1222(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g7),.DATA(g34590));
  MSFF DFF_1223(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2779),.DATA(g26928));
  MSFF DFF_1224(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4200),.DATA(g4197));
  MSFF DFF_1225(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4446),.DATA(g26954));
  MSFF DFF_1226(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1720),.DATA(g30351));
  MSFF DFF_1227(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1367),.DATA(g31871));
  MSFF DFF_1228(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5112),.DATA(g5105));
  MSFF DFF_1229(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g19),.DATA(g34594));
  MSFF DFF_1230(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4145),.DATA(g26939));
  MSFF DFF_1231(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2161),.DATA(g33994));
  MSFF DFF_1232(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g376),.DATA(g25596));
  MSFF DFF_1233(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2361),.DATA(g33586));
  MSFF DFF_1234(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4191),.DATA(g21901));
  MSFF DFF_1235(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g582),.DATA(g31866));
  MSFF DFF_1236(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2051),.DATA(g33000));
  MSFF DFF_1237(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1193),.DATA(g26918));
  MSFF DFF_1238(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5401),.DATA(g33051));
  MSFF DFF_1239(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3408),.DATA(g28065));
  MSFF DFF_1240(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2327),.DATA(g30373));
  MSFF DFF_1241(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g907),.DATA(g28056));
  MSFF DFF_1242(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g947),.DATA(g34601));
  MSFF DFF_1243(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1834),.DATA(g30355));
  MSFF DFF_1244(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3594),.DATA(g30426));
  MSFF DFF_1245(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2999),.DATA(g34805));
  MSFF DFF_1246(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5727),.DATA(g31913));
  MSFF DFF_1247(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2303),.DATA(g34002));
  MSFF DFF_1248(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6661),.DATA(g6704));
  MSFF DFF_1249(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3065),.DATA(g25652));
  MSFF DFF_1250(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g699),.DATA(g28053));
  MSFF DFF_1251(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g723),.DATA(g29229));
  MSFF DFF_1252(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5703),.DATA(g33620));
  MSFF DFF_1253(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g546),.DATA(g34722));
  MSFF DFF_1254(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2472),.DATA(g33599));
  MSFF DFF_1255(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5953),.DATA(g30515));
  MSFF DFF_1256(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3096),.DATA(g25649));
  MSFF DFF_1257(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6439),.DATA(g33066));
  MSFF DFF_1258(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1740),.DATA(g33979));
  MSFF DFF_1259(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3550),.DATA(g30417));
  MSFF DFF_1260(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3845),.DATA(g25683));
  MSFF DFF_1261(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2116),.DATA(g33574));
  MSFF DFF_1262(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5677),.DATA(g5673));
  MSFF DFF_1263(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3195),.DATA(g30410));
  MSFF DFF_1264(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3913),.DATA(g30454));
  MSFF DFF_1265(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4537),.DATA(g34024));
  MSFF DFF_1266(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1687),.DATA(g33547));
  MSFF DFF_1267(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2681),.DATA(g30386));
  MSFF DFF_1268(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2533),.DATA(g33596));
  MSFF DFF_1269(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g324),.DATA(g26887));
  MSFF DFF_1270(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2697),.DATA(g34607));
  MSFF DFF_1271(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5747),.DATA(g33056));
  MSFF DFF_1272(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4417),.DATA(g31895));
  MSFF DFF_1273(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6561),.DATA(g33068));
  MSFF DFF_1274(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1141),.DATA(g29233));
  MSFF DFF_1275(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1570),.DATA(g24258));
  MSFF DFF_1276(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2413),.DATA(g30376));
  MSFF DFF_1277(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1710),.DATA(g33549));
  MSFF DFF_1278(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6527),.DATA(g29308));
  MSFF DFF_1279(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6404),.DATA(g25759));
  MSFF DFF_1280(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3255),.DATA(g30408));
  MSFF DFF_1281(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1691),.DATA(g29241));
  MSFF DFF_1282(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2936),.DATA(g34620));
  MSFF DFF_1283(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5644),.DATA(g33621));
  MSFF DFF_1284(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5152),.DATA(g25707));
  MSFF DFF_1285(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5352),.DATA(g24339));
  MSFF DFF_1286(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4213),.DATA(g4185));
  MSFF DFF_1287(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6120),.DATA(g25738));
  MSFF DFF_1288(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2775),.DATA(g34443));
  MSFF DFF_1289(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2922),.DATA(g34619));
  MSFF DFF_1290(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1111),.DATA(g29234));
  MSFF DFF_1291(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5893),.DATA(g30503));
  MSFF DFF_1292(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1311),.DATA(g21724));
  MSFF DFF_1293(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3267),.DATA(g3310));
  MSFF DFF_1294(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6617),.DATA(g30550));
  MSFF DFF_1295(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2060),.DATA(g33001));
  MSFF DFF_1296(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4512),.DATA(g33040));
  MSFF DFF_1297(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5599),.DATA(g30492));
  MSFF DFF_1298(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3401),.DATA(g25664));
  MSFF DFF_1299(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4366),.DATA(g26944));
  MSFF DFF_1300(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3676),.DATA(g3672));
  MSFF DFF_1301(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g94),.DATA(g34614));
  MSFF DFF_1302(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3129),.DATA(g29260));
  MSFF DFF_1303(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3329),.DATA(g3325));
  MSFF DFF_1304(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5170),.DATA(g33047));
  MSFF DFF_1305(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4456),.DATA(g25692));
  MSFF DFF_1306(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5821),.DATA(g25733));
  MSFF DFF_1307(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6299),.DATA(g30536));
  MSFF DFF_1308(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1239),.DATA(g1157));
  MSFF DFF_1309(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3727),.DATA(g31888));
  MSFF DFF_1310(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2079),.DATA(g29246));
  MSFF DFF_1311(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4698),.DATA(g34261));
  MSFF DFF_1312(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3703),.DATA(g33611));
  MSFF DFF_1313(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1559),.DATA(g25638));
  MSFF DFF_1314(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g943),.DATA(g34728));
  MSFF DFF_1315(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g411),.DATA(g29222));
  MSFF DFF_1316(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6140),.DATA(g25742));
  MSFF DFF_1317(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3953),.DATA(g30449));
  MSFF DFF_1318(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3068),.DATA(g25643));
  MSFF DFF_1319(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2704),.DATA(g34608));
  MSFF DFF_1320(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6035),.DATA(g24345));
  MSFF DFF_1321(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6082),.DATA(g31922));
  MSFF DFF_1322(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g49),.DATA(g34994));
  MSFF DFF_1323(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1300),.DATA(g25635));
  MSFF DFF_1324(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4057),.DATA(g25686));
  MSFF DFF_1325(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5200),.DATA(g30461));
  MSFF DFF_1326(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4843),.DATA(g34466));
  MSFF DFF_1327(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5046),.DATA(g31901));
  MSFF DFF_1328(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2250),.DATA(g29249));
  MSFF DFF_1329(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g319),.DATA(g26882));
  MSFF DFF_1330(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4549),.DATA(g33041));
  MSFF DFF_1331(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2453),.DATA(g33011));
  MSFF DFF_1332(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5841),.DATA(g25734));
  MSFF DFF_1333(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5763),.DATA(g28097));
  MSFF DFF_1334(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3747),.DATA(g33030));
  MSFF DFF_1335(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5637),.DATA(g5659));
  MSFF DFF_1336(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2912),.DATA(g34618));
  MSFF DFF_1337(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2357),.DATA(g33010));
  MSFF DFF_1338(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4232),.DATA(g4229));
  MSFF DFF_1339(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g164),.DATA(g31864));
  MSFF DFF_1340(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4253),.DATA(g34630));
  MSFF DFF_1341(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5016),.DATA(g31898));
  MSFF DFF_1342(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3119),.DATA(g25653));
  MSFF DFF_1343(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1351),.DATA(g25632));
  MSFF DFF_1344(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1648),.DATA(g32988));
  MSFF DFF_1345(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4519),.DATA(g33616));
  MSFF DFF_1346(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5115),.DATA(g29280));
  MSFF DFF_1347(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3352),.DATA(g33609));
  MSFF DFF_1348(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6657),.DATA(g30563));
  MSFF DFF_1349(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4552),.DATA(g33044));
  MSFF DFF_1350(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3893),.DATA(g30437));
  MSFF DFF_1351(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3211),.DATA(g30412));
  MSFF DFF_1352(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5654),.DATA(g5630));
  MSFF DFF_1353(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g929),.DATA(g21725));
  MSFF DFF_1354(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3274),.DATA(g3267));
  MSFF DFF_1355(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5595),.DATA(g30491));
  MSFF DFF_1356(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3614),.DATA(g30434));
  MSFF DFF_1357(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2894),.DATA(g34612));
  MSFF DFF_1358(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3125),.DATA(g29259));
  MSFF DFF_1359(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3325),.DATA(g3321));
  MSFF DFF_1360(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3821),.DATA(g25681));
  MSFF DFF_1361(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4141),.DATA(g25687));
  MSFF DFF_1362(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4570),.DATA(g33617));
  MSFF DFF_1363(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5272),.DATA(g30479));
  MSFF DFF_1364(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2735),.DATA(g29256));
  MSFF DFF_1365(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g728),.DATA(g28054));
  MSFF DFF_1366(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6295),.DATA(g30535));
  MSFF DFF_1367(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5417),.DATA(g28094));
  MSFF DFF_1368(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2661),.DATA(g30385));
  MSFF DFF_1369(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1988),.DATA(g30361));
  MSFF DFF_1370(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5128),.DATA(g25705));
  MSFF DFF_1371(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1548),.DATA(g24260));
  MSFF DFF_1372(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3106),.DATA(g29257));
  MSFF DFF_1373(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4659),.DATA(g34461));
  MSFF DFF_1374(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4358),.DATA(g34258));
  MSFF DFF_1375(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1792),.DATA(g32993));
  MSFF DFF_1376(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2084),.DATA(g33992));
  MSFF DFF_1377(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3061),.DATA(g28061));
  MSFF DFF_1378(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3187),.DATA(g30394));
  MSFF DFF_1379(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4311),.DATA(g34449));
  MSFF DFF_1380(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2583),.DATA(g34019));
  MSFF DFF_1381(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3003),.DATA(g21726));
  MSFF DFF_1382(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1094),.DATA(g29231));
  MSFF DFF_1383(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3841),.DATA(g25682));
  MSFF DFF_1384(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4284),.DATA(g21897));
  MSFF DFF_1385(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3763),.DATA(g28067));
  MSFF DFF_1386(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3191),.DATA(g30395));
  MSFF DFF_1387(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4239),.DATA(g21892));
  MSFF DFF_1388(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3391),.DATA(g31885));
  MSFF DFF_1389(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4180),.DATA(g4210));
  MSFF DFF_1390(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g691),.DATA(g28048));
  MSFF DFF_1391(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g534),.DATA(g34723));
  MSFF DFF_1392(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5366),.DATA(g25717));
  MSFF DFF_1393(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g385),.DATA(g25598));
  MSFF DFF_1394(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2004),.DATA(g33987));
  MSFF DFF_1395(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2527),.DATA(g30380));
  MSFF DFF_1396(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5456),.DATA(g5448));
  MSFF DFF_1397(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4420),.DATA(g26965));
  MSFF DFF_1398(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5148),.DATA(g25706));
  MSFF DFF_1399(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4507),.DATA(g30458));
  MSFF DFF_1400(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5348),.DATA(g24338));
  MSFF DFF_1401(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3223),.DATA(g30400));
  MSFF DFF_1402(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4931),.DATA(g21904));
  MSFF DFF_1403(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2970),.DATA(g34623));
  MSFF DFF_1404(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5698),.DATA(g24343));
  MSFF DFF_1405(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3416),.DATA(g25666));
  MSFF DFF_1406(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5260),.DATA(g30473));
  MSFF DFF_1407(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1521),.DATA(g24252));
  MSFF DFF_1408(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3522),.DATA(g33028));
  MSFF DFF_1409(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3115),.DATA(g29258));
  MSFF DFF_1410(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3251),.DATA(g30407));
  MSFF DFF_1411(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1),.DATA(g26958));
  MSFF DFF_1412(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4628),.DATA(g34457));
  MSFF DFF_1413(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1996),.DATA(g33568));
  MSFF DFF_1414(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3447),.DATA(g25663));
  MSFF DFF_1415(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4515),.DATA(g26964));
  MSFF DFF_1416(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4204),.DATA(g4200));
  MSFF DFF_1417(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4300),.DATA(g34735));
  MSFF DFF_1418(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1724),.DATA(g30352));
  MSFF DFF_1419(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1379),.DATA(g33543));
  MSFF DFF_1420(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3654),.DATA(g24271));
  MSFF DFF_1421(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g12),.DATA(g30326));
  MSFF DFF_1422(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1878),.DATA(g33981));
  MSFF DFF_1423(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5619),.DATA(g30500));
  MSFF DFF_1424(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g71),.DATA(g34786));
  MSFF DFF_1425(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g59),.DATA(g29277));
//
  NOT NOT1_0(.VSS(VSS),.VDD(VDD),.Y(I28349),.A(g28367));
  NOT NOT1_1(.VSS(VSS),.VDD(VDD),.Y(g19408),.A(g16066));
  NOT NOT1_2(.VSS(VSS),.VDD(VDD),.Y(I21294),.A(g18274));
  NOT NOT1_3(.VSS(VSS),.VDD(VDD),.Y(g13297),.A(g10831));
  NOT NOT1_4(.VSS(VSS),.VDD(VDD),.Y(g19635),.A(g16349));
  NOT NOT1_5(.VSS(VSS),.VDD(VDD),.Y(g32394),.A(g30601));
  NOT NOT1_6(.VSS(VSS),.VDD(VDD),.Y(I19778),.A(g17781));
  NOT NOT1_7(.VSS(VSS),.VDD(VDD),.Y(g9900),.A(g6));
  NOT NOT1_8(.VSS(VSS),.VDD(VDD),.Y(g11889),.A(g9954));
  NOT NOT1_9(.VSS(VSS),.VDD(VDD),.Y(g13103),.A(g10905));
  NOT NOT1_10(.VSS(VSS),.VDD(VDD),.Y(g17470),.A(g14454));
  NOT NOT1_11(.VSS(VSS),.VDD(VDD),.Y(g23499),.A(g20785));
  NOT NOT1_12(.VSS(VSS),.VDD(VDD),.Y(g6895),.A(g3288));
  NOT NOT1_13(.VSS(VSS),.VDD(VDD),.Y(g9797),.A(g5441));
  NOT NOT1_14(.VSS(VSS),.VDD(VDD),.Y(g31804),.A(g29385));
  NOT NOT1_15(.VSS(VSS),.VDD(VDD),.Y(g6837),.A(g968));
  NOT NOT1_16(.VSS(VSS),.VDD(VDD),.Y(I15824),.A(g1116));
  NOT NOT1_17(.VSS(VSS),.VDD(VDD),.Y(g20066),.A(g17433));
  NOT NOT1_18(.VSS(VSS),.VDD(VDD),.Y(g33804),.A(g33250));
  NOT NOT1_19(.VSS(VSS),.VDD(VDD),.Y(g20231),.A(g17821));
  NOT NOT1_20(.VSS(VSS),.VDD(VDD),.Y(I19786),.A(g17844));
  NOT NOT1_21(.VSS(VSS),.VDD(VDD),.Y(g24066),.A(g21127));
  NOT NOT1_22(.VSS(VSS),.VDD(VDD),.Y(g11888),.A(g10160));
  NOT NOT1_23(.VSS(VSS),.VDD(VDD),.Y(g9510),.A(g5835));
  NOT NOT1_24(.VSS(VSS),.VDD(VDD),.Y(I22692),.A(g21308));
  NOT NOT1_25(.VSS(VSS),.VDD(VDD),.Y(g12884),.A(g10392));
  NOT NOT1_26(.VSS(VSS),.VDD(VDD),.Y(g22494),.A(g19801));
  NOT NOT1_27(.VSS(VSS),.VDD(VDD),.Y(g9245),.A(I13031));
  NOT NOT1_28(.VSS(VSS),.VDD(VDD),.Y(g8925),.A(I12910));
  NOT NOT1_29(.VSS(VSS),.VDD(VDD),.Y(g34248),.A(I32243));
  NOT NOT1_30(.VSS(VSS),.VDD(VDD),.Y(g10289),.A(g1319));
  NOT NOT1_31(.VSS(VSS),.VDD(VDD),.Y(g11181),.A(g8134));
  NOT NOT1_32(.VSS(VSS),.VDD(VDD),.Y(I20116),.A(g15737));
  NOT NOT1_33(.VSS(VSS),.VDD(VDD),.Y(g7888),.A(g1536));
  NOT NOT1_34(.VSS(VSS),.VDD(VDD),.Y(g9291),.A(g3021));
  NOT NOT1_35(.VSS(VSS),.VDD(VDD),.Y(g28559),.A(g27700));
  NOT NOT1_36(.VSS(VSS),.VDD(VDD),.Y(g21056),.A(g15426));
  NOT NOT1_37(.VSS(VSS),.VDD(VDD),.Y(I33246),.A(g34970));
  NOT NOT1_38(.VSS(VSS),.VDD(VDD),.Y(g10288),.A(I13718));
  NOT NOT1_39(.VSS(VSS),.VDD(VDD),.Y(g8224),.A(g3774));
  NOT NOT1_40(.VSS(VSS),.VDD(VDD),.Y(g21611),.A(I21210));
  NOT NOT1_41(.VSS(VSS),.VDD(VDD),.Y(g16718),.A(I17932));
  NOT NOT1_42(.VSS(VSS),.VDD(VDD),.Y(g21722),.A(I21285));
  NOT NOT1_43(.VSS(VSS),.VDD(VDD),.Y(I12530),.A(g4815));
  NOT NOT1_44(.VSS(VSS),.VDD(VDD),.Y(g16521),.A(g13543));
  NOT NOT1_45(.VSS(VSS),.VDD(VDD),.Y(I22400),.A(g19620));
  NOT NOT1_46(.VSS(VSS),.VDD(VDD),.Y(g23611),.A(g18833));
  NOT NOT1_47(.VSS(VSS),.VDD(VDD),.Y(g10571),.A(g10233));
  NOT NOT1_48(.VSS(VSS),.VDD(VDD),.Y(g17467),.A(g14339));
  NOT NOT1_49(.VSS(VSS),.VDD(VDD),.Y(g17494),.A(g14339));
  NOT NOT1_50(.VSS(VSS),.VDD(VDD),.Y(g10308),.A(g4459));
  NOT NOT1_51(.VSS(VSS),.VDD(VDD),.Y(g27015),.A(g26869));
  NOT NOT1_52(.VSS(VSS),.VDD(VDD),.Y(g23988),.A(g19277));
  NOT NOT1_53(.VSS(VSS),.VDD(VDD),.Y(g23924),.A(g18997));
  NOT NOT1_54(.VSS(VSS),.VDD(VDD),.Y(g12217),.A(I15070));
  NOT NOT1_55(.VSS(VSS),.VDD(VDD),.Y(g14571),.A(I16688));
  NOT NOT1_56(.VSS(VSS),.VDD(VDD),.Y(g32318),.A(g31596));
  NOT NOT1_57(.VSS(VSS),.VDD(VDD),.Y(g32446),.A(g31596));
  NOT NOT1_58(.VSS(VSS),.VDD(VDD),.Y(g14308),.A(I16471));
  NOT NOT1_59(.VSS(VSS),.VDD(VDD),.Y(I24041),.A(g22182));
  NOT NOT1_60(.VSS(VSS),.VDD(VDD),.Y(I14935),.A(g9902));
  NOT NOT1_61(.VSS(VSS),.VDD(VDD),.Y(g34778),.A(I32976));
  NOT NOT1_62(.VSS(VSS),.VDD(VDD),.Y(g20511),.A(g17929));
  NOT NOT1_63(.VSS(VSS),.VDD(VDD),.Y(g26672),.A(g25275));
  NOT NOT1_64(.VSS(VSS),.VDD(VDD),.Y(g11931),.A(I14749));
  NOT NOT1_65(.VSS(VSS),.VDD(VDD),.Y(g20763),.A(I20816));
  NOT NOT1_66(.VSS(VSS),.VDD(VDD),.Y(g23432),.A(g21514));
  NOT NOT1_67(.VSS(VSS),.VDD(VDD),.Y(I18165),.A(g13177));
  NOT NOT1_68(.VSS(VSS),.VDD(VDD),.Y(I18523),.A(g14443));
  NOT NOT1_69(.VSS(VSS),.VDD(VDD),.Y(g21271),.A(I21002));
  NOT NOT1_70(.VSS(VSS),.VDD(VDD),.Y(I31776),.A(g33204));
  NOT NOT1_71(.VSS(VSS),.VDD(VDD),.Y(g23271),.A(g20785));
  NOT NOT1_72(.VSS(VSS),.VDD(VDD),.Y(g22155),.A(g19074));
  NOT NOT1_73(.VSS(VSS),.VDD(VDD),.Y(I22539),.A(g19606));
  NOT NOT1_74(.VSS(VSS),.VDD(VDD),.Y(I32231),.A(g34123));
  NOT NOT1_75(.VSS(VSS),.VDD(VDD),.Y(g34786),.A(I32988));
  NOT NOT1_76(.VSS(VSS),.VDD(VDD),.Y(g9259),.A(g5176));
  NOT NOT1_77(.VSS(VSS),.VDD(VDD),.Y(I15190),.A(g6005));
  NOT NOT1_78(.VSS(VSS),.VDD(VDD),.Y(g17782),.A(I18788));
  NOT NOT1_79(.VSS(VSS),.VDD(VDD),.Y(g8277),.A(I12483));
  NOT NOT1_80(.VSS(VSS),.VDD(VDD),.Y(g9819),.A(g92));
  NOT NOT1_81(.VSS(VSS),.VDD(VDD),.Y(I16969),.A(g13943));
  NOT NOT1_82(.VSS(VSS),.VDD(VDD),.Y(g32540),.A(g30614));
  NOT NOT1_83(.VSS(VSS),.VDD(VDD),.Y(g25027),.A(I24191));
  NOT NOT1_84(.VSS(VSS),.VDD(VDD),.Y(g19711),.A(g17062));
  NOT NOT1_85(.VSS(VSS),.VDD(VDD),.Y(g22170),.A(g19210));
  NOT NOT1_86(.VSS(VSS),.VDD(VDD),.Y(g13190),.A(g10939));
  NOT NOT1_87(.VSS(VSS),.VDD(VDD),.Y(g7297),.A(g6069));
  NOT NOT1_88(.VSS(VSS),.VDD(VDD),.Y(g17419),.A(g14965));
  NOT NOT1_89(.VSS(VSS),.VDD(VDD),.Y(g20660),.A(g17873));
  NOT NOT1_90(.VSS(VSS),.VDD(VDD),.Y(g16861),.A(I18051));
  NOT NOT1_91(.VSS(VSS),.VDD(VDD),.Y(g21461),.A(g15348));
  NOT NOT1_92(.VSS(VSS),.VDD(VDD),.Y(g10816),.A(I14054));
  NOT NOT1_93(.VSS(VSS),.VDD(VDD),.Y(g28713),.A(g27907));
  NOT NOT1_94(.VSS(VSS),.VDD(VDD),.Y(g15755),.A(g13134));
  NOT NOT1_95(.VSS(VSS),.VDD(VDD),.Y(g23461),.A(g18833));
  NOT NOT1_96(.VSS(VSS),.VDD(VDD),.Y(I24237),.A(g23823));
  NOT NOT1_97(.VSS(VSS),.VDD(VDD),.Y(g34945),.A(g34933));
  NOT NOT1_98(.VSS(VSS),.VDD(VDD),.Y(g8789),.A(I12779));
  NOT NOT1_99(.VSS(VSS),.VDD(VDD),.Y(g31833),.A(g29385));
  NOT NOT1_100(.VSS(VSS),.VDD(VDD),.Y(I18006),.A(g13638));
  NOT NOT1_101(.VSS(VSS),.VDD(VDD),.Y(I20035),.A(g15706));
  NOT NOT1_102(.VSS(VSS),.VDD(VDD),.Y(I17207),.A(g13835));
  NOT NOT1_103(.VSS(VSS),.VDD(VDD),.Y(g30999),.A(g29722));
  NOT NOT1_104(.VSS(VSS),.VDD(VDD),.Y(g25249),.A(g22228));
  NOT NOT1_105(.VSS(VSS),.VDD(VDD),.Y(g9488),.A(g1878));
  NOT NOT1_106(.VSS(VSS),.VDD(VDD),.Y(g19537),.A(g15938));
  NOT NOT1_107(.VSS(VSS),.VDD(VDD),.Y(g17155),.A(I18205));
  NOT NOT1_108(.VSS(VSS),.VDD(VDD),.Y(I16855),.A(g10473));
  NOT NOT1_109(.VSS(VSS),.VDD(VDD),.Y(g15563),.A(I17140));
  NOT NOT1_110(.VSS(VSS),.VDD(VDD),.Y(g23031),.A(g19801));
  NOT NOT1_111(.VSS(VSS),.VDD(VDD),.Y(g30090),.A(g29134));
  NOT NOT1_112(.VSS(VSS),.VDD(VDD),.Y(g30998),.A(g29719));
  NOT NOT1_113(.VSS(VSS),.VDD(VDD),.Y(g25248),.A(g22228));
  NOT NOT1_114(.VSS(VSS),.VDD(VDD),.Y(g23650),.A(g20653));
  NOT NOT1_115(.VSS(VSS),.VDD(VDD),.Y(g7138),.A(g5360));
  NOT NOT1_116(.VSS(VSS),.VDD(VDD),.Y(g16099),.A(g13437));
  NOT NOT1_117(.VSS(VSS),.VDD(VDD),.Y(g34998),.A(g34981));
  NOT NOT1_118(.VSS(VSS),.VDD(VDD),.Y(g23887),.A(g18997));
  NOT NOT1_119(.VSS(VSS),.VDD(VDD),.Y(g25552),.A(g22594));
  NOT NOT1_120(.VSS(VSS),.VDD(VDD),.Y(g20916),.A(g18008));
  NOT NOT1_121(.VSS(VSS),.VDD(VDD),.Y(g27084),.A(g26673));
  NOT NOT1_122(.VSS(VSS),.VDD(VDD),.Y(g30182),.A(I28419));
  NOT NOT1_123(.VSS(VSS),.VDD(VDD),.Y(g7963),.A(g4146));
  NOT NOT1_124(.VSS(VSS),.VDD(VDD),.Y(g10374),.A(g6903));
  NOT NOT1_125(.VSS(VSS),.VDD(VDD),.Y(I32763),.A(g34511));
  NOT NOT1_126(.VSS(VSS),.VDD(VDD),.Y(g19606),.A(g17614));
  NOT NOT1_127(.VSS(VSS),.VDD(VDD),.Y(g19492),.A(g16349));
  NOT NOT1_128(.VSS(VSS),.VDD(VDD),.Y(g22167),.A(g19074));
  NOT NOT1_129(.VSS(VSS),.VDD(VDD),.Y(g22194),.A(I21776));
  NOT NOT1_130(.VSS(VSS),.VDD(VDD),.Y(g7109),.A(g5011));
  NOT NOT1_131(.VSS(VSS),.VDD(VDD),.Y(g7791),.A(I12199));
  NOT NOT1_132(.VSS(VSS),.VDD(VDD),.Y(g34672),.A(I32800));
  NOT NOT1_133(.VSS(VSS),.VDD(VDD),.Y(g16777),.A(I18003));
  NOT NOT1_134(.VSS(VSS),.VDD(VDD),.Y(g20550),.A(g15864));
  NOT NOT1_135(.VSS(VSS),.VDD(VDD),.Y(g23529),.A(g20558));
  NOT NOT1_136(.VSS(VSS),.VDD(VDD),.Y(g6854),.A(g2685));
  NOT NOT1_137(.VSS(VSS),.VDD(VDD),.Y(g18930),.A(g15789));
  NOT NOT1_138(.VSS(VSS),.VDD(VDD),.Y(g13024),.A(g11900));
  NOT NOT1_139(.VSS(VSS),.VDD(VDD),.Y(g32902),.A(g30673));
  NOT NOT1_140(.VSS(VSS),.VDD(VDD),.Y(g6941),.A(g3990));
  NOT NOT1_141(.VSS(VSS),.VDD(VDD),.Y(g12110),.A(I14970));
  NOT NOT1_142(.VSS(VSS),.VDD(VDD),.Y(g32957),.A(g31672));
  NOT NOT1_143(.VSS(VSS),.VDD(VDD),.Y(g9951),.A(g6133));
  NOT NOT1_144(.VSS(VSS),.VDD(VDD),.Y(g32377),.A(g30984));
  NOT NOT1_145(.VSS(VSS),.VDD(VDD),.Y(g12922),.A(g12297));
  NOT NOT1_146(.VSS(VSS),.VDD(VDD),.Y(g23528),.A(g18833));
  NOT NOT1_147(.VSS(VSS),.VDD(VDD),.Y(g12321),.A(g9637));
  NOT NOT1_148(.VSS(VSS),.VDD(VDD),.Y(g28678),.A(g27800));
  NOT NOT1_149(.VSS(VSS),.VDD(VDD),.Y(g32739),.A(g30735));
  NOT NOT1_150(.VSS(VSS),.VDD(VDD),.Y(g21393),.A(g17264));
  NOT NOT1_151(.VSS(VSS),.VDD(VDD),.Y(g23843),.A(g19147));
  NOT NOT1_152(.VSS(VSS),.VDD(VDD),.Y(g26026),.A(I25105));
  NOT NOT1_153(.VSS(VSS),.VDD(VDD),.Y(g25081),.A(g22342));
  NOT NOT1_154(.VSS(VSS),.VDD(VDD),.Y(g20085),.A(g16187));
  NOT NOT1_155(.VSS(VSS),.VDD(VDD),.Y(g23393),.A(g20739));
  NOT NOT1_156(.VSS(VSS),.VDD(VDD),.Y(g19750),.A(g16326));
  NOT NOT1_157(.VSS(VSS),.VDD(VDD),.Y(g30331),.A(I28594));
  NOT NOT1_158(.VSS(VSS),.VDD(VDD),.Y(g24076),.A(g19984));
  NOT NOT1_159(.VSS(VSS),.VDD(VDD),.Y(g24085),.A(g20857));
  NOT NOT1_160(.VSS(VSS),.VDD(VDD),.Y(g17589),.A(g14981));
  NOT NOT1_161(.VSS(VSS),.VDD(VDD),.Y(g20596),.A(I20690));
  NOT NOT1_162(.VSS(VSS),.VDD(VDD),.Y(g34932),.A(g34914));
  NOT NOT1_163(.VSS(VSS),.VDD(VDD),.Y(g23764),.A(g21308));
  NOT NOT1_164(.VSS(VSS),.VDD(VDD),.Y(g25786),.A(g24518));
  NOT NOT1_165(.VSS(VSS),.VDD(VDD),.Y(I25869),.A(g25851));
  NOT NOT1_166(.VSS(VSS),.VDD(VDD),.Y(g32738),.A(g31376));
  NOT NOT1_167(.VSS(VSS),.VDD(VDD),.Y(g32562),.A(g30673));
  NOT NOT1_168(.VSS(VSS),.VDD(VDD),.Y(g32645),.A(g30825));
  NOT NOT1_169(.VSS(VSS),.VDD(VDD),.Y(g14669),.A(g12301));
  NOT NOT1_170(.VSS(VSS),.VDD(VDD),.Y(g20054),.A(g17328));
  NOT NOT1_171(.VSS(VSS),.VDD(VDD),.Y(I26337),.A(g26835));
  NOT NOT1_172(.VSS(VSS),.VDD(VDD),.Y(g24054),.A(g19919));
  NOT NOT1_173(.VSS(VSS),.VDD(VDD),.Y(I20130),.A(g15748));
  NOT NOT1_174(.VSS(VSS),.VDD(VDD),.Y(g17588),.A(g14782));
  NOT NOT1_175(.VSS(VSS),.VDD(VDD),.Y(g17524),.A(g14933));
  NOT NOT1_176(.VSS(VSS),.VDD(VDD),.Y(I18600),.A(g5335));
  NOT NOT1_177(.VSS(VSS),.VDD(VDD),.Y(g23869),.A(g19277));
  NOT NOT1_178(.VSS(VSS),.VDD(VDD),.Y(g32699),.A(g31528));
  NOT NOT1_179(.VSS(VSS),.VDD(VDD),.Y(g10392),.A(g6989));
  NOT NOT1_180(.VSS(VSS),.VDD(VDD),.Y(I28576),.A(g28431));
  NOT NOT1_181(.VSS(VSS),.VDD(VDD),.Y(I28585),.A(g30217));
  NOT NOT1_182(.VSS(VSS),.VDD(VDD),.Y(I15987),.A(g12381));
  NOT NOT1_183(.VSS(VSS),.VDD(VDD),.Y(g14668),.A(g12450));
  NOT NOT1_184(.VSS(VSS),.VDD(VDD),.Y(g25356),.A(g22763));
  NOT NOT1_185(.VSS(VSS),.VDD(VDD),.Y(g24431),.A(g22722));
  NOT NOT1_186(.VSS(VSS),.VDD(VDD),.Y(g29725),.A(g28349));
  NOT NOT1_187(.VSS(VSS),.VDD(VDD),.Y(I15250),.A(g9152));
  NOT NOT1_188(.VSS(VSS),.VDD(VDD),.Y(g28294),.A(g27295));
  NOT NOT1_189(.VSS(VSS),.VDD(VDD),.Y(g8945),.A(g608));
  NOT NOT1_190(.VSS(VSS),.VDD(VDD),.Y(g10489),.A(g9259));
  NOT NOT1_191(.VSS(VSS),.VDD(VDD),.Y(g11987),.A(I14833));
  NOT NOT1_192(.VSS(VSS),.VDD(VDD),.Y(g13625),.A(g10971));
  NOT NOT1_193(.VSS(VSS),.VDD(VDD),.Y(I25161),.A(g24920));
  NOT NOT1_194(.VSS(VSS),.VDD(VDD),.Y(g17477),.A(g14848));
  NOT NOT1_195(.VSS(VSS),.VDD(VDD),.Y(g23868),.A(g19277));
  NOT NOT1_196(.VSS(VSS),.VDD(VDD),.Y(g32698),.A(g30614));
  NOT NOT1_197(.VSS(VSS),.VDD(VDD),.Y(g31812),.A(g29385));
  NOT NOT1_198(.VSS(VSS),.VDD(VDD),.Y(g11250),.A(g7502));
  NOT NOT1_199(.VSS(VSS),.VDD(VDD),.Y(g25380),.A(g23776));
  NOT NOT1_200(.VSS(VSS),.VDD(VDD),.Y(I32550),.A(g34398));
  NOT NOT1_201(.VSS(VSS),.VDD(VDD),.Y(g7957),.A(g1252));
  NOT NOT1_202(.VSS(VSS),.VDD(VDD),.Y(g13250),.A(I15811));
  NOT NOT1_203(.VSS(VSS),.VDD(VDD),.Y(g20269),.A(g15844));
  NOT NOT1_204(.VSS(VSS),.VDD(VDD),.Y(g34505),.A(g34409));
  NOT NOT1_205(.VSS(VSS),.VDD(VDD),.Y(g7049),.A(g5853));
  NOT NOT1_206(.VSS(VSS),.VDD(VDD),.Y(g20773),.A(I20830));
  NOT NOT1_207(.VSS(VSS),.VDD(VDD),.Y(g25090),.A(g23630));
  NOT NOT1_208(.VSS(VSS),.VDD(VDD),.Y(g6958),.A(g4372));
  NOT NOT1_209(.VSS(VSS),.VDD(VDD),.Y(g20268),.A(g18008));
  NOT NOT1_210(.VSS(VSS),.VDD(VDD),.Y(g14424),.A(g11136));
  NOT NOT1_211(.VSS(VSS),.VDD(VDD),.Y(g34717),.A(I32881));
  NOT NOT1_212(.VSS(VSS),.VDD(VDD),.Y(g12417),.A(g7175));
  NOT NOT1_213(.VSS(VSS),.VDD(VDD),.Y(g25182),.A(g22763));
  NOT NOT1_214(.VSS(VSS),.VDD(VDD),.Y(g12936),.A(g12601));
  NOT NOT1_215(.VSS(VSS),.VDD(VDD),.Y(g20655),.A(I20753));
  NOT NOT1_216(.VSS(VSS),.VDD(VDD),.Y(g8340),.A(g3050));
  NOT NOT1_217(.VSS(VSS),.VDD(VDD),.Y(g13943),.A(I16231));
  NOT NOT1_218(.VSS(VSS),.VDD(VDD),.Y(g21225),.A(g17428));
  NOT NOT1_219(.VSS(VSS),.VDD(VDD),.Y(g24156),.A(I23312));
  NOT NOT1_220(.VSS(VSS),.VDD(VDD),.Y(g23259),.A(g21070));
  NOT NOT1_221(.VSS(VSS),.VDD(VDD),.Y(g24655),.A(g23067));
  NOT NOT1_222(.VSS(VSS),.VDD(VDD),.Y(I12109),.A(g749));
  NOT NOT1_223(.VSS(VSS),.VDD(VDD),.Y(I18063),.A(g14357));
  NOT NOT1_224(.VSS(VSS),.VDD(VDD),.Y(g7715),.A(g1178));
  NOT NOT1_225(.VSS(VSS),.VDD(VDD),.Y(g29744),.A(g28431));
  NOT NOT1_226(.VSS(VSS),.VDD(VDD),.Y(g8478),.A(g3103));
  NOT NOT1_227(.VSS(VSS),.VDD(VDD),.Y(g20180),.A(g17533));
  NOT NOT1_228(.VSS(VSS),.VDD(VDD),.Y(g17616),.A(g14309));
  NOT NOT1_229(.VSS(VSS),.VDD(VDD),.Y(g20670),.A(g15426));
  NOT NOT1_230(.VSS(VSS),.VDD(VDD),.Y(I29447),.A(g30729));
  NOT NOT1_231(.VSS(VSS),.VDD(VDD),.Y(g10830),.A(g10087));
  NOT NOT1_232(.VSS(VSS),.VDD(VDD),.Y(I32243),.A(g34134));
  NOT NOT1_233(.VSS(VSS),.VDD(VDD),.Y(g22305),.A(g19801));
  NOT NOT1_234(.VSS(VSS),.VDD(VDD),.Y(g24180),.A(I23384));
  NOT NOT1_235(.VSS(VSS),.VDD(VDD),.Y(g32632),.A(g31070));
  NOT NOT1_236(.VSS(VSS),.VDD(VDD),.Y(g31795),.A(I29371));
  NOT NOT1_237(.VSS(VSS),.VDD(VDD),.Y(g9594),.A(g2307));
  NOT NOT1_238(.VSS(VSS),.VDD(VDD),.Y(g6829),.A(g1319));
  NOT NOT1_239(.VSS(VSS),.VDD(VDD),.Y(g7498),.A(g6675));
  NOT NOT1_240(.VSS(VSS),.VDD(VDD),.Y(g23258),.A(g20924));
  NOT NOT1_241(.VSS(VSS),.VDD(VDD),.Y(g26811),.A(g25206));
  NOT NOT1_242(.VSS(VSS),.VDD(VDD),.Y(I16590),.A(g11966));
  NOT NOT1_243(.VSS(VSS),.VDD(VDD),.Y(g10544),.A(I13906));
  NOT NOT1_244(.VSS(VSS),.VDD(VDD),.Y(g15573),.A(I17154));
  NOT NOT1_245(.VSS(VSS),.VDD(VDD),.Y(I27492),.A(g27511));
  NOT NOT1_246(.VSS(VSS),.VDD(VDD),.Y(g9806),.A(g5782));
  NOT NOT1_247(.VSS(VSS),.VDD(VDD),.Y(g14544),.A(I16663));
  NOT NOT1_248(.VSS(VSS),.VDD(VDD),.Y(I14653),.A(g9417));
  NOT NOT1_249(.VSS(VSS),.VDD(VDD),.Y(I33044),.A(g34775));
  NOT NOT1_250(.VSS(VSS),.VDD(VDD),.Y(I16741),.A(g5677));
  NOT NOT1_251(.VSS(VSS),.VDD(VDD),.Y(g25513),.A(g23870));
  NOT NOT1_252(.VSS(VSS),.VDD(VDD),.Y(g32661),.A(g31070));
  NOT NOT1_253(.VSS(VSS),.VDD(VDD),.Y(g20993),.A(g15615));
  NOT NOT1_254(.VSS(VSS),.VDD(VDD),.Y(g32547),.A(g30614));
  NOT NOT1_255(.VSS(VSS),.VDD(VDD),.Y(g32895),.A(g30673));
  NOT NOT1_256(.VSS(VSS),.VDD(VDD),.Y(g8876),.A(I12855));
  NOT NOT1_257(.VSS(VSS),.VDD(VDD),.Y(g24839),.A(g23436));
  NOT NOT1_258(.VSS(VSS),.VDD(VDD),.Y(g23244),.A(I22343));
  NOT NOT1_259(.VSS(VSS),.VDD(VDD),.Y(g24993),.A(g22384));
  NOT NOT1_260(.VSS(VSS),.VDD(VDD),.Y(g22177),.A(g19074));
  NOT NOT1_261(.VSS(VSS),.VDD(VDD),.Y(g16162),.A(g13437));
  NOT NOT1_262(.VSS(VSS),.VDD(VDD),.Y(g11855),.A(I14671));
  NOT NOT1_263(.VSS(VSS),.VDD(VDD),.Y(g20667),.A(g15224));
  NOT NOT1_264(.VSS(VSS),.VDD(VDD),.Y(g17466),.A(g12983));
  NOT NOT1_265(.VSS(VSS),.VDD(VDD),.Y(g9887),.A(g5802));
  NOT NOT1_266(.VSS(VSS),.VDD(VDD),.Y(g6974),.A(I11746));
  NOT NOT1_267(.VSS(VSS),.VDD(VDD),.Y(g24667),.A(g23112));
  NOT NOT1_268(.VSS(VSS),.VDD(VDD),.Y(g9934),.A(g5849));
  NOT NOT1_269(.VSS(VSS),.VDD(VDD),.Y(g21069),.A(g15277));
  NOT NOT1_270(.VSS(VSS),.VDD(VDD),.Y(g25505),.A(g22228));
  NOT NOT1_271(.VSS(VSS),.VDD(VDD),.Y(g34433),.A(I32470));
  NOT NOT1_272(.VSS(VSS),.VDD(VDD),.Y(g34387),.A(g34188));
  NOT NOT1_273(.VSS(VSS),.VDD(VDD),.Y(g10042),.A(g2671));
  NOT NOT1_274(.VSS(VSS),.VDD(VDD),.Y(g24131),.A(g21209));
  NOT NOT1_275(.VSS(VSS),.VDD(VDD),.Y(g32481),.A(g31194));
  NOT NOT1_276(.VSS(VSS),.VDD(VDD),.Y(g14705),.A(I16803));
  NOT NOT1_277(.VSS(VSS),.VDD(VDD),.Y(I13321),.A(g6486));
  NOT NOT1_278(.VSS(VSS),.VDD(VDD),.Y(g18975),.A(g15938));
  NOT NOT1_279(.VSS(VSS),.VDD(VDD),.Y(g19553),.A(g16782));
  NOT NOT1_280(.VSS(VSS),.VDD(VDD),.Y(g19862),.A(I20233));
  NOT NOT1_281(.VSS(VSS),.VDD(VDD),.Y(g30097),.A(g29118));
  NOT NOT1_282(.VSS(VSS),.VDD(VDD),.Y(g8915),.A(I12884));
  NOT NOT1_283(.VSS(VSS),.VDD(VDD),.Y(g16629),.A(g13990));
  NOT NOT1_284(.VSS(VSS),.VDD(VDD),.Y(I16150),.A(g10430));
  NOT NOT1_285(.VSS(VSS),.VDD(VDD),.Y(g21657),.A(g17657));
  NOT NOT1_286(.VSS(VSS),.VDD(VDD),.Y(g16472),.A(g14098));
  NOT NOT1_287(.VSS(VSS),.VDD(VDD),.Y(I20781),.A(g17155));
  NOT NOT1_288(.VSS(VSS),.VDD(VDD),.Y(g21068),.A(g15277));
  NOT NOT1_289(.VSS(VSS),.VDD(VDD),.Y(g14255),.A(g12381));
  NOT NOT1_290(.VSS(VSS),.VDD(VDD),.Y(I21477),.A(g18695));
  NOT NOT1_291(.VSS(VSS),.VDD(VDD),.Y(g14189),.A(I16391));
  NOT NOT1_292(.VSS(VSS),.VDD(VDD),.Y(g32551),.A(g30735));
  NOT NOT1_293(.VSS(VSS),.VDD(VDD),.Y(g32572),.A(g30735));
  NOT NOT1_294(.VSS(VSS),.VDD(VDD),.Y(g23375),.A(g20924));
  NOT NOT1_295(.VSS(VSS),.VDD(VDD),.Y(I24781),.A(g24264));
  NOT NOT1_296(.VSS(VSS),.VDD(VDD),.Y(I33146),.A(g34903));
  NOT NOT1_297(.VSS(VSS),.VDD(VDD),.Y(g7162),.A(g4521));
  NOT NOT1_298(.VSS(VSS),.VDD(VDD),.Y(g25212),.A(g22763));
  NOT NOT1_299(.VSS(VSS),.VDD(VDD),.Y(g7268),.A(g1636));
  NOT NOT1_300(.VSS(VSS),.VDD(VDD),.Y(I11740),.A(g4519));
  NOT NOT1_301(.VSS(VSS),.VDD(VDD),.Y(g7362),.A(g1906));
  NOT NOT1_302(.VSS(VSS),.VDD(VDD),.Y(g12909),.A(g10412));
  NOT NOT1_303(.VSS(VSS),.VDD(VDD),.Y(g9433),.A(g5148));
  NOT NOT1_304(.VSS(VSS),.VDD(VDD),.Y(g26850),.A(I25576));
  NOT NOT1_305(.VSS(VSS),.VDD(VDD),.Y(g12543),.A(g9417));
  NOT NOT1_306(.VSS(VSS),.VDD(VDD),.Y(g17642),.A(g14691));
  NOT NOT1_307(.VSS(VSS),.VDD(VDD),.Y(g20502),.A(g15373));
  NOT NOT1_308(.VSS(VSS),.VDD(VDD),.Y(g10678),.A(I13990));
  NOT NOT1_309(.VSS(VSS),.VDD(VDD),.Y(I22725),.A(g21250));
  NOT NOT1_310(.VSS(VSS),.VDD(VDD),.Y(I13740),.A(g85));
  NOT NOT1_311(.VSS(VSS),.VDD(VDD),.Y(g23879),.A(g19210));
  NOT NOT1_312(.VSS(VSS),.VDD(VDD),.Y(g20557),.A(I20647));
  NOT NOT1_313(.VSS(VSS),.VDD(VDD),.Y(g23970),.A(g19277));
  NOT NOT1_314(.VSS(VSS),.VDD(VDD),.Y(g34343),.A(g34089));
  NOT NOT1_315(.VSS(VSS),.VDD(VDD),.Y(g20210),.A(g16897));
  NOT NOT1_316(.VSS(VSS),.VDD(VDD),.Y(I22114),.A(g19935));
  NOT NOT1_317(.VSS(VSS),.VDD(VDD),.Y(g12908),.A(g10414));
  NOT NOT1_318(.VSS(VSS),.VDD(VDD),.Y(g20618),.A(g15277));
  NOT NOT1_319(.VSS(VSS),.VDD(VDD),.Y(g11867),.A(I14679));
  NOT NOT1_320(.VSS(VSS),.VDD(VDD),.Y(g11894),.A(I14702));
  NOT NOT1_321(.VSS(VSS),.VDD(VDD),.Y(I11685),.A(g117));
  NOT NOT1_322(.VSS(VSS),.VDD(VDD),.Y(g8310),.A(g2051));
  NOT NOT1_323(.VSS(VSS),.VDD(VDD),.Y(g23878),.A(g19147));
  NOT NOT1_324(.VSS(VSS),.VDD(VDD),.Y(g21337),.A(g15758));
  NOT NOT1_325(.VSS(VSS),.VDD(VDD),.Y(g20443),.A(g15171));
  NOT NOT1_326(.VSS(VSS),.VDD(VDD),.Y(g10383),.A(g6978));
  NOT NOT1_327(.VSS(VSS),.VDD(VDD),.Y(g23337),.A(g20924));
  NOT NOT1_328(.VSS(VSS),.VDD(VDD),.Y(g19757),.A(g17224));
  NOT NOT1_329(.VSS(VSS),.VDD(VDD),.Y(g9496),.A(g3303));
  NOT NOT1_330(.VSS(VSS),.VDD(VDD),.Y(g14383),.A(I16535));
  NOT NOT1_331(.VSS(VSS),.VDD(VDD),.Y(g17733),.A(g14238));
  NOT NOT1_332(.VSS(VSS),.VDD(VDD),.Y(I16526),.A(g10430));
  NOT NOT1_333(.VSS(VSS),.VDD(VDD),.Y(g8663),.A(g3343));
  NOT NOT1_334(.VSS(VSS),.VDD(VDD),.Y(g10030),.A(g116));
  NOT NOT1_335(.VSS(VSS),.VDD(VDD),.Y(g23886),.A(g21468));
  NOT NOT1_336(.VSS(VSS),.VDD(VDD),.Y(I18614),.A(g6315));
  NOT NOT1_337(.VSS(VSS),.VDD(VDD),.Y(g32490),.A(g30673));
  NOT NOT1_338(.VSS(VSS),.VDD(VDD),.Y(g10093),.A(g5703));
  NOT NOT1_339(.VSS(VSS),.VDD(VDD),.Y(g18884),.A(g15938));
  NOT NOT1_340(.VSS(VSS),.VDD(VDD),.Y(g27242),.A(g26183));
  NOT NOT1_341(.VSS(VSS),.VDD(VDD),.Y(I14576),.A(g8791));
  NOT NOT1_342(.VSS(VSS),.VDD(VDD),.Y(g11714),.A(g8107));
  NOT NOT1_343(.VSS(VSS),.VDD(VDD),.Y(g22166),.A(g18997));
  NOT NOT1_344(.VSS(VSS),.VDD(VDD),.Y(g11450),.A(I14455));
  NOT NOT1_345(.VSS(VSS),.VDD(VDD),.Y(I17114),.A(g14358));
  NOT NOT1_346(.VSS(VSS),.VDD(VDD),.Y(I27192),.A(g27662));
  NOT NOT1_347(.VSS(VSS),.VDD(VDD),.Y(g23792),.A(g19074));
  NOT NOT1_348(.VSS(VSS),.VDD(VDD),.Y(g23967),.A(g19210));
  NOT NOT1_349(.VSS(VSS),.VDD(VDD),.Y(g23994),.A(g19277));
  NOT NOT1_350(.VSS(VSS),.VDD(VDD),.Y(g32784),.A(g31672));
  NOT NOT1_351(.VSS(VSS),.VDD(VDD),.Y(g9891),.A(g6173));
  NOT NOT1_352(.VSS(VSS),.VDD(VDD),.Y(I18320),.A(g13605));
  NOT NOT1_353(.VSS(VSS),.VDD(VDD),.Y(g28037),.A(g26365));
  NOT NOT1_354(.VSS(VSS),.VDD(VDD),.Y(g8002),.A(g1389));
  NOT NOT1_355(.VSS(VSS),.VDD(VDD),.Y(g9337),.A(g1608));
  NOT NOT1_356(.VSS(VSS),.VDD(VDD),.Y(g9913),.A(g2403));
  NOT NOT1_357(.VSS(VSS),.VDD(VDD),.Y(g32956),.A(g30825));
  NOT NOT1_358(.VSS(VSS),.VDD(VDD),.Y(I21285),.A(g18215));
  NOT NOT1_359(.VSS(VSS),.VDD(VDD),.Y(g11819),.A(g7717));
  NOT NOT1_360(.VSS(VSS),.VDD(VDD),.Y(g11910),.A(g10185));
  NOT NOT1_361(.VSS(VSS),.VDD(VDD),.Y(g14065),.A(g11048));
  NOT NOT1_362(.VSS(VSS),.VDD(VDD),.Y(g7086),.A(g4826));
  NOT NOT1_363(.VSS(VSS),.VDD(VDD),.Y(g13707),.A(g11360));
  NOT NOT1_364(.VSS(VSS),.VDD(VDD),.Y(g31829),.A(g29385));
  NOT NOT1_365(.VSS(VSS),.VDD(VDD),.Y(g32889),.A(g31376));
  NOT NOT1_366(.VSS(VSS),.VDD(VDD),.Y(g11202),.A(I14267));
  NOT NOT1_367(.VSS(VSS),.VDD(VDD),.Y(g8236),.A(g4812));
  NOT NOT1_368(.VSS(VSS),.VDD(VDD),.Y(g33920),.A(I31786));
  NOT NOT1_369(.VSS(VSS),.VDD(VDD),.Y(I21254),.A(g16540));
  NOT NOT1_370(.VSS(VSS),.VDD(VDD),.Y(g24039),.A(g21256));
  NOT NOT1_371(.VSS(VSS),.VDD(VDD),.Y(g25620),.A(I24759));
  NOT NOT1_372(.VSS(VSS),.VDD(VDD),.Y(g21425),.A(g15509));
  NOT NOT1_373(.VSS(VSS),.VDD(VDD),.Y(g29221),.A(I27579));
  NOT NOT1_374(.VSS(VSS),.VDD(VDD),.Y(I17744),.A(g14912));
  NOT NOT1_375(.VSS(VSS),.VDD(VDD),.Y(g23459),.A(g21611));
  NOT NOT1_376(.VSS(VSS),.VDD(VDD),.Y(I16917),.A(g10582));
  NOT NOT1_377(.VSS(VSS),.VDD(VDD),.Y(g20038),.A(g17328));
  NOT NOT1_378(.VSS(VSS),.VDD(VDD),.Y(g23425),.A(g20751));
  NOT NOT1_379(.VSS(VSS),.VDD(VDD),.Y(g31828),.A(g29385));
  NOT NOT1_380(.VSS(VSS),.VDD(VDD),.Y(g32888),.A(g30673));
  NOT NOT1_381(.VSS(VSS),.VDD(VDD),.Y(I15070),.A(g10108));
  NOT NOT1_382(.VSS(VSS),.VDD(VDD),.Y(g25097),.A(g22342));
  NOT NOT1_383(.VSS(VSS),.VDD(VDD),.Y(g32824),.A(g31376));
  NOT NOT1_384(.VSS(VSS),.VDD(VDD),.Y(g10219),.A(g2697));
  NOT NOT1_385(.VSS(VSS),.VDD(VDD),.Y(g13055),.A(I15682));
  NOT NOT1_386(.VSS(VSS),.VDD(VDD),.Y(g9807),.A(g5712));
  NOT NOT1_387(.VSS(VSS),.VDD(VDD),.Y(I30901),.A(g32407));
  NOT NOT1_388(.VSS(VSS),.VDD(VDD),.Y(g19673),.A(g16931));
  NOT NOT1_389(.VSS(VSS),.VDD(VDD),.Y(g24038),.A(g21193));
  NOT NOT1_390(.VSS(VSS),.VDD(VDD),.Y(g14219),.A(g12381));
  NOT NOT1_391(.VSS(VSS),.VDD(VDD),.Y(g19397),.A(g16449));
  NOT NOT1_392(.VSS(VSS),.VDD(VDD),.Y(g21458),.A(g15758));
  NOT NOT1_393(.VSS(VSS),.VDD(VDD),.Y(g6849),.A(g2551));
  NOT NOT1_394(.VSS(VSS),.VDD(VDD),.Y(I15590),.A(g11988));
  NOT NOT1_395(.VSS(VSS),.VDD(VDD),.Y(g28155),.A(I26664));
  NOT NOT1_396(.VSS(VSS),.VDD(VDD),.Y(I13762),.A(g6755));
  NOT NOT1_397(.VSS(VSS),.VDD(VDD),.Y(g13070),.A(g11984));
  NOT NOT1_398(.VSS(VSS),.VDD(VDD),.Y(g23458),.A(I22583));
  NOT NOT1_399(.VSS(VSS),.VDD(VDD),.Y(g32671),.A(g31528));
  NOT NOT1_400(.VSS(VSS),.VDD(VDD),.Y(I21036),.A(g17221));
  NOT NOT1_401(.VSS(VSS),.VDD(VDD),.Y(g34229),.A(g33936));
  NOT NOT1_402(.VSS(VSS),.VDD(VDD),.Y(g10218),.A(g2527));
  NOT NOT1_403(.VSS(VSS),.VDD(VDD),.Y(I18034),.A(g13680));
  NOT NOT1_404(.VSS(VSS),.VDD(VDD),.Y(g16172),.A(g13584));
  NOT NOT1_405(.VSS(VSS),.VDD(VDD),.Y(g20601),.A(g17433));
  NOT NOT1_406(.VSS(VSS),.VDD(VDD),.Y(g21010),.A(g15634));
  NOT NOT1_407(.VSS(VSS),.VDD(VDD),.Y(g11986),.A(I14830));
  NOT NOT1_408(.VSS(VSS),.VDD(VDD),.Y(g7470),.A(g5623));
  NOT NOT1_409(.VSS(VSS),.VDD(VDD),.Y(I12483),.A(g3096));
  NOT NOT1_410(.VSS(VSS),.VDD(VDD),.Y(g17476),.A(g14665));
  NOT NOT1_411(.VSS(VSS),.VDD(VDD),.Y(g17485),.A(I18408));
  NOT NOT1_412(.VSS(VSS),.VDD(VDD),.Y(I16077),.A(g10430));
  NOT NOT1_413(.VSS(VSS),.VDD(VDD),.Y(I14745),.A(g10029));
  NOT NOT1_414(.VSS(VSS),.VDD(VDD),.Y(g11741),.A(g10033));
  NOT NOT1_415(.VSS(VSS),.VDD(VDD),.Y(g22907),.A(g20453));
  NOT NOT1_416(.VSS(VSS),.VDD(VDD),.Y(g23545),.A(g21562));
  NOT NOT1_417(.VSS(VSS),.VDD(VDD),.Y(g23444),.A(I22561));
  NOT NOT1_418(.VSS(VSS),.VDD(VDD),.Y(g25369),.A(g22228));
  NOT NOT1_419(.VSS(VSS),.VDD(VDD),.Y(g32931),.A(g30937));
  NOT NOT1_420(.VSS(VSS),.VDD(VDD),.Y(g33682),.A(I31515));
  NOT NOT1_421(.VSS(VSS),.VDD(VDD),.Y(g6900),.A(g3440));
  NOT NOT1_422(.VSS(VSS),.VDD(VDD),.Y(g19634),.A(g16349));
  NOT NOT1_423(.VSS(VSS),.VDD(VDD),.Y(g19872),.A(g17015));
  NOT NOT1_424(.VSS(VSS),.VDD(VDD),.Y(g34716),.A(I32878));
  NOT NOT1_425(.VSS(VSS),.VDD(VDD),.Y(I20542),.A(g16508));
  NOT NOT1_426(.VSS(VSS),.VDD(VDD),.Y(I25598),.A(g25424));
  NOT NOT1_427(.VSS(VSS),.VDD(VDD),.Y(g8928),.A(g4340));
  NOT NOT1_428(.VSS(VSS),.VDD(VDD),.Y(g29812),.A(g28381));
  NOT NOT1_429(.VSS(VSS),.VDD(VDD),.Y(I28241),.A(g28709));
  NOT NOT1_430(.VSS(VSS),.VDD(VDD),.Y(g12841),.A(g10357));
  NOT NOT1_431(.VSS(VSS),.VDD(VDD),.Y(g22594),.A(I21934));
  NOT NOT1_432(.VSS(VSS),.VDD(VDD),.Y(I16688),.A(g10981));
  NOT NOT1_433(.VSS(VSS),.VDD(VDD),.Y(g9815),.A(g6098));
  NOT NOT1_434(.VSS(VSS),.VDD(VDD),.Y(g8064),.A(g3376));
  NOT NOT1_435(.VSS(VSS),.VDD(VDD),.Y(I18408),.A(g13017));
  NOT NOT1_436(.VSS(VSS),.VDD(VDD),.Y(I20913),.A(g16964));
  NOT NOT1_437(.VSS(VSS),.VDD(VDD),.Y(g23086),.A(g20283));
  NOT NOT1_438(.VSS(VSS),.VDD(VDD),.Y(I32815),.A(g34470));
  NOT NOT1_439(.VSS(VSS),.VDD(VDD),.Y(g30310),.A(g28830));
  NOT NOT1_440(.VSS(VSS),.VDD(VDD),.Y(g8899),.A(g807));
  NOT NOT1_441(.VSS(VSS),.VDD(VDD),.Y(g11735),.A(g8534));
  NOT NOT1_442(.VSS(VSS),.VDD(VDD),.Y(g29371),.A(I27735));
  NOT NOT1_443(.VSS(VSS),.VDD(VDD),.Y(I11908),.A(g4449));
  NOT NOT1_444(.VSS(VSS),.VDD(VDD),.Y(g9692),.A(g1756));
  NOT NOT1_445(.VSS(VSS),.VDD(VDD),.Y(g13877),.A(g11350));
  NOT NOT1_446(.VSS(VSS),.VDD(VDD),.Y(I32601),.A(g34319));
  NOT NOT1_447(.VSS(VSS),.VDD(VDD),.Y(g8785),.A(I12767));
  NOT NOT1_448(.VSS(VSS),.VDD(VDD),.Y(g24169),.A(I23351));
  NOT NOT1_449(.VSS(VSS),.VDD(VDD),.Y(g24791),.A(g23850));
  NOT NOT1_450(.VSS(VSS),.VDD(VDD),.Y(g9497),.A(I13166));
  NOT NOT1_451(.VSS(VSS),.VDD(VDD),.Y(I16102),.A(g10430));
  NOT NOT1_452(.VSS(VSS),.VDD(VDD),.Y(g26681),.A(g25396));
  NOT NOT1_453(.VSS(VSS),.VDD(VDD),.Y(g20168),.A(g17533));
  NOT NOT1_454(.VSS(VSS),.VDD(VDD),.Y(g9154),.A(I12994));
  NOT NOT1_455(.VSS(VSS),.VDD(VDD),.Y(g25133),.A(g23733));
  NOT NOT1_456(.VSS(VSS),.VDD(VDD),.Y(g34925),.A(I33167));
  NOT NOT1_457(.VSS(VSS),.VDD(VDD),.Y(I26309),.A(g26825));
  NOT NOT1_458(.VSS(VSS),.VDD(VDD),.Y(g9354),.A(g2719));
  NOT NOT1_459(.VSS(VSS),.VDD(VDD),.Y(g27014),.A(g25888));
  NOT NOT1_460(.VSS(VSS),.VDD(VDD),.Y(I27564),.A(g28166));
  NOT NOT1_461(.VSS(VSS),.VDD(VDD),.Y(g24168),.A(I23348));
  NOT NOT1_462(.VSS(VSS),.VDD(VDD),.Y(g23322),.A(I22425));
  NOT NOT1_463(.VSS(VSS),.VDD(VDD),.Y(g32546),.A(g31170));
  NOT NOT1_464(.VSS(VSS),.VDD(VDD),.Y(g9960),.A(g6474));
  NOT NOT1_465(.VSS(VSS),.VDD(VDD),.Y(g22519),.A(g19801));
  NOT NOT1_466(.VSS(VSS),.VDD(VDD),.Y(g22176),.A(g18997));
  NOT NOT1_467(.VSS(VSS),.VDD(VDD),.Y(g14201),.A(I16401));
  NOT NOT1_468(.VSS(VSS),.VDD(VDD),.Y(g26802),.A(I25514));
  NOT NOT1_469(.VSS(VSS),.VDD(VDD),.Y(g28119),.A(g27008));
  NOT NOT1_470(.VSS(VSS),.VDD(VDD),.Y(g12835),.A(g10352));
  NOT NOT1_471(.VSS(VSS),.VDD(VDD),.Y(g7635),.A(g1002));
  NOT NOT1_472(.VSS(VSS),.VDD(VDD),.Y(g14277),.A(I16455));
  NOT NOT1_473(.VSS(VSS),.VDD(VDD),.Y(g20666),.A(g15224));
  NOT NOT1_474(.VSS(VSS),.VDD(VDD),.Y(g13018),.A(I15636));
  NOT NOT1_475(.VSS(VSS),.VDD(VDD),.Y(I16231),.A(g10520));
  NOT NOT1_476(.VSS(VSS),.VDD(VDD),.Y(g32024),.A(I29582));
  NOT NOT1_477(.VSS(VSS),.VDD(VDD),.Y(g25228),.A(g23828));
  NOT NOT1_478(.VSS(VSS),.VDD(VDD),.Y(I19802),.A(g15727));
  NOT NOT1_479(.VSS(VSS),.VDD(VDD),.Y(g19574),.A(g16826));
  NOT NOT1_480(.VSS(VSS),.VDD(VDD),.Y(g7766),.A(I12189));
  NOT NOT1_481(.VSS(VSS),.VDD(VDD),.Y(g19452),.A(g16326));
  NOT NOT1_482(.VSS(VSS),.VDD(VDD),.Y(g6819),.A(g1046));
  NOT NOT1_483(.VSS(VSS),.VDD(VDD),.Y(g16540),.A(I17744));
  NOT NOT1_484(.VSS(VSS),.VDD(VDD),.Y(I19857),.A(g16640));
  NOT NOT1_485(.VSS(VSS),.VDD(VDD),.Y(g22154),.A(g19074));
  NOT NOT1_486(.VSS(VSS),.VDD(VDD),.Y(g7087),.A(g6336));
  NOT NOT1_487(.VSS(VSS),.VDD(VDD),.Y(I33297),.A(g35000));
  NOT NOT1_488(.VSS(VSS),.VDD(VDD),.Y(g25011),.A(g22763));
  NOT NOT1_489(.VSS(VSS),.VDD(VDD),.Y(g32860),.A(g30673));
  NOT NOT1_490(.VSS(VSS),.VDD(VDD),.Y(I18891),.A(g16676));
  NOT NOT1_491(.VSS(VSS),.VDD(VDD),.Y(g7487),.A(g1259));
  NOT NOT1_492(.VSS(VSS),.VDD(VDD),.Y(I33103),.A(g34846));
  NOT NOT1_493(.VSS(VSS),.VDD(VDD),.Y(g8237),.A(g255));
  NOT NOT1_494(.VSS(VSS),.VDD(VDD),.Y(g18953),.A(g16077));
  NOT NOT1_495(.VSS(VSS),.VDD(VDD),.Y(I14761),.A(g7753));
  NOT NOT1_496(.VSS(VSS),.VDD(VDD),.Y(g19912),.A(g17328));
  NOT NOT1_497(.VSS(VSS),.VDD(VDD),.Y(g17519),.A(I18460));
  NOT NOT1_498(.VSS(VSS),.VDD(VDD),.Y(g21561),.A(g15595));
  NOT NOT1_499(.VSS(VSS),.VDD(VDD),.Y(I12183),.A(g2719));
  NOT NOT1_500(.VSS(VSS),.VDD(VDD),.Y(g21656),.A(g17700));
  NOT NOT1_501(.VSS(VSS),.VDD(VDD),.Y(g6923),.A(g3791));
  NOT NOT1_502(.VSS(VSS),.VDD(VDD),.Y(g26765),.A(g25309));
  NOT NOT1_503(.VSS(VSS),.VDD(VDD),.Y(I25680),.A(g25641));
  NOT NOT1_504(.VSS(VSS),.VDD(VDD),.Y(g22935),.A(g20283));
  NOT NOT1_505(.VSS(VSS),.VDD(VDD),.Y(g17092),.A(g14011));
  NOT NOT1_506(.VSS(VSS),.VDD(VDD),.Y(g34944),.A(g34932));
  NOT NOT1_507(.VSS(VSS),.VDD(VDD),.Y(g10037),.A(g1848));
  NOT NOT1_508(.VSS(VSS),.VDD(VDD),.Y(I32791),.A(g34578));
  NOT NOT1_509(.VSS(VSS),.VDD(VDD),.Y(g32497),.A(g30673));
  NOT NOT1_510(.VSS(VSS),.VDD(VDD),.Y(g21295),.A(g17533));
  NOT NOT1_511(.VSS(VSS),.VDD(VDD),.Y(g23353),.A(g20924));
  NOT NOT1_512(.VSS(VSS),.VDD(VDD),.Y(g29507),.A(g28353));
  NOT NOT1_513(.VSS(VSS),.VDD(VDD),.Y(I32884),.A(g34690));
  NOT NOT1_514(.VSS(VSS),.VDD(VDD),.Y(g8844),.A(I12826));
  NOT NOT1_515(.VSS(VSS),.VDD(VDD),.Y(g11402),.A(g7594));
  NOT NOT1_516(.VSS(VSS),.VDD(VDD),.Y(g17518),.A(g14918));
  NOT NOT1_517(.VSS(VSS),.VDD(VDD),.Y(g26549),.A(I25391));
  NOT NOT1_518(.VSS(VSS),.VDD(VDD),.Y(g17154),.A(g14348));
  NOT NOT1_519(.VSS(VSS),.VDD(VDD),.Y(g22883),.A(g20391));
  NOT NOT1_520(.VSS(VSS),.VDD(VDD),.Y(g20556),.A(g15483));
  NOT NOT1_521(.VSS(VSS),.VDD(VDD),.Y(g23823),.A(I22989));
  NOT NOT1_522(.VSS(VSS),.VDD(VDD),.Y(g17637),.A(g12933));
  NOT NOT1_523(.VSS(VSS),.VDD(VDD),.Y(g20580),.A(g17328));
  NOT NOT1_524(.VSS(VSS),.VDD(VDD),.Y(g26548),.A(g25255));
  NOT NOT1_525(.VSS(VSS),.VDD(VDD),.Y(g10419),.A(g8821));
  NOT NOT1_526(.VSS(VSS),.VDD(VDD),.Y(g11866),.A(g9883));
  NOT NOT1_527(.VSS(VSS),.VDD(VDD),.Y(g11917),.A(I14727));
  NOT NOT1_528(.VSS(VSS),.VDD(VDD),.Y(g32700),.A(g31579));
  NOT NOT1_529(.VSS(VSS),.VDD(VDD),.Y(I26687),.A(g27880));
  NOT NOT1_530(.VSS(VSS),.VDD(VDD),.Y(g32659),.A(g30735));
  NOT NOT1_531(.VSS(VSS),.VDD(VDD),.Y(g21336),.A(g17367));
  NOT NOT1_532(.VSS(VSS),.VDD(VDD),.Y(g32625),.A(g31070));
  NOT NOT1_533(.VSS(VSS),.VDD(VDD),.Y(g10352),.A(g6804));
  NOT NOT1_534(.VSS(VSS),.VDD(VDD),.Y(g23336),.A(g20924));
  NOT NOT1_535(.VSS(VSS),.VDD(VDD),.Y(I32479),.A(g34302));
  NOT NOT1_536(.VSS(VSS),.VDD(VDD),.Y(g19592),.A(I20035));
  NOT NOT1_537(.VSS(VSS),.VDD(VDD),.Y(g34429),.A(I32458));
  NOT NOT1_538(.VSS(VSS),.VDD(VDD),.Y(g10155),.A(g2643));
  NOT NOT1_539(.VSS(VSS),.VDD(VDD),.Y(g10418),.A(g8818));
  NOT NOT1_540(.VSS(VSS),.VDD(VDD),.Y(g12041),.A(I14905));
  NOT NOT1_541(.VSS(VSS),.VDD(VDD),.Y(g32658),.A(g31579));
  NOT NOT1_542(.VSS(VSS),.VDD(VDD),.Y(g19780),.A(g16449));
  NOT NOT1_543(.VSS(VSS),.VDD(VDD),.Y(g16739),.A(g13223));
  NOT NOT1_544(.VSS(VSS),.VDD(VDD),.Y(g12430),.A(I15250));
  NOT NOT1_545(.VSS(VSS),.VDD(VDD),.Y(I16660),.A(g10981));
  NOT NOT1_546(.VSS(VSS),.VDD(VDD),.Y(g34428),.A(I32455));
  NOT NOT1_547(.VSS(VSS),.VDD(VDD),.Y(I21074),.A(g17766));
  NOT NOT1_548(.VSS(VSS),.VDD(VDD),.Y(g23966),.A(g19210));
  NOT NOT1_549(.VSS(VSS),.VDD(VDD),.Y(g22215),.A(g19277));
  NOT NOT1_550(.VSS(VSS),.VDD(VDD),.Y(g28036),.A(g26365));
  NOT NOT1_551(.VSS(VSS),.VDD(VDD),.Y(g27237),.A(g26162));
  NOT NOT1_552(.VSS(VSS),.VDD(VDD),.Y(g32943),.A(g31710));
  NOT NOT1_553(.VSS(VSS),.VDD(VDD),.Y(g20110),.A(g16897));
  NOT NOT1_554(.VSS(VSS),.VDD(VDD),.Y(g11706),.A(I14579));
  NOT NOT1_555(.VSS(VSS),.VDD(VDD),.Y(g24084),.A(g20720));
  NOT NOT1_556(.VSS(VSS),.VDD(VDD),.Y(g16738),.A(I17956));
  NOT NOT1_557(.VSS(VSS),.VDD(VDD),.Y(g9761),.A(g2445));
  NOT NOT1_558(.VSS(VSS),.VDD(VDD),.Y(g13706),.A(g11280));
  NOT NOT1_559(.VSS(VSS),.VDD(VDD),.Y(g16645),.A(g13756));
  NOT NOT1_560(.VSS(VSS),.VDD(VDD),.Y(g12465),.A(g7192));
  NOT NOT1_561(.VSS(VSS),.VDD(VDD),.Y(I11992),.A(g763));
  NOT NOT1_562(.VSS(VSS),.VDD(VDD),.Y(g24110),.A(g21209));
  NOT NOT1_563(.VSS(VSS),.VDD(VDD),.Y(g20922),.A(I20891));
  NOT NOT1_564(.VSS(VSS),.VDD(VDD),.Y(g27983),.A(g26725));
  NOT NOT1_565(.VSS(VSS),.VDD(VDD),.Y(g20321),.A(g17821));
  NOT NOT1_566(.VSS(VSS),.VDD(VDD),.Y(g23017),.A(g20453));
  NOT NOT1_567(.VSS(VSS),.VDD(VDD),.Y(g32644),.A(g30735));
  NOT NOT1_568(.VSS(VSS),.VDD(VDD),.Y(g33648),.A(I31482));
  NOT NOT1_569(.VSS(VSS),.VDD(VDD),.Y(I21238),.A(g16540));
  NOT NOT1_570(.VSS(VSS),.VDD(VDD),.Y(g34690),.A(I32840));
  NOT NOT1_571(.VSS(VSS),.VDD(VDD),.Y(g6870),.A(g3089));
  NOT NOT1_572(.VSS(VSS),.VDD(VDD),.Y(g9828),.A(g2024));
  NOT NOT1_573(.VSS(VSS),.VDD(VDD),.Y(g20179),.A(g17249));
  NOT NOT1_574(.VSS(VSS),.VDD(VDD),.Y(g34549),.A(I32617));
  NOT NOT1_575(.VSS(VSS),.VDD(VDD),.Y(g8948),.A(g785));
  NOT NOT1_576(.VSS(VSS),.VDD(VDD),.Y(g20531),.A(g15907));
  NOT NOT1_577(.VSS(VSS),.VDD(VDD),.Y(g12983),.A(I15600));
  NOT NOT1_578(.VSS(VSS),.VDD(VDD),.Y(g24179),.A(I23381));
  NOT NOT1_579(.VSS(VSS),.VDD(VDD),.Y(g16290),.A(g13260));
  NOT NOT1_580(.VSS(VSS),.VDD(VDD),.Y(g32969),.A(g30735));
  NOT NOT1_581(.VSS(VSS),.VDD(VDD),.Y(g13280),.A(I15846));
  NOT NOT1_582(.VSS(VSS),.VDD(VDD),.Y(g6825),.A(g979));
  NOT NOT1_583(.VSS(VSS),.VDD(VDD),.Y(g33755),.A(I31610));
  NOT NOT1_584(.VSS(VSS),.VDD(VDD),.Y(g17501),.A(I18434));
  NOT NOT1_585(.VSS(VSS),.VDD(VDD),.Y(g7369),.A(g1996));
  NOT NOT1_586(.VSS(VSS),.VDD(VDD),.Y(g27142),.A(g26105));
  NOT NOT1_587(.VSS(VSS),.VDD(VDD),.Y(g8955),.A(g1418));
  NOT NOT1_588(.VSS(VSS),.VDD(VDD),.Y(g20178),.A(g16971));
  NOT NOT1_589(.VSS(VSS),.VDD(VDD),.Y(g10194),.A(g6741));
  NOT NOT1_590(.VSS(VSS),.VDD(VDD),.Y(g19396),.A(g16431));
  NOT NOT1_591(.VSS(VSS),.VDD(VDD),.Y(g17577),.A(I18504));
  NOT NOT1_592(.VSS(VSS),.VDD(VDD),.Y(g13624),.A(g10951));
  NOT NOT1_593(.VSS(VSS),.VDD(VDD),.Y(I14241),.A(g8356));
  NOT NOT1_594(.VSS(VSS),.VDD(VDD),.Y(I21941),.A(g18918));
  NOT NOT1_595(.VSS(VSS),.VDD(VDD),.Y(g24178),.A(I23378));
  NOT NOT1_596(.VSS(VSS),.VDD(VDD),.Y(g14167),.A(I16371));
  NOT NOT1_597(.VSS(VSS),.VDD(VDD),.Y(g32968),.A(g31376));
  NOT NOT1_598(.VSS(VSS),.VDD(VDD),.Y(g19731),.A(g17093));
  NOT NOT1_599(.VSS(VSS),.VDD(VDD),.Y(g29920),.A(g28824));
  NOT NOT1_600(.VSS(VSS),.VDD(VDD),.Y(g34504),.A(g34408));
  NOT NOT1_601(.VSS(VSS),.VDD(VDD),.Y(g29358),.A(I27718));
  NOT NOT1_602(.VSS(VSS),.VDD(VDD),.Y(g7868),.A(g1099));
  NOT NOT1_603(.VSS(VSS),.VDD(VDD),.Y(I15102),.A(g5313));
  NOT NOT1_604(.VSS(VSS),.VDD(VDD),.Y(I26195),.A(g26260));
  NOT NOT1_605(.VSS(VSS),.VDD(VDD),.Y(I11835),.A(g101));
  NOT NOT1_606(.VSS(VSS),.VDD(VDD),.Y(I20891),.A(g17700));
  NOT NOT1_607(.VSS(VSS),.VDD(VDD),.Y(g9746),.A(I13326));
  NOT NOT1_608(.VSS(VSS),.VDD(VDD),.Y(g20373),.A(g17929));
  NOT NOT1_609(.VSS(VSS),.VDD(VDD),.Y(g32855),.A(g30825));
  NOT NOT1_610(.VSS(VSS),.VDD(VDD),.Y(g23289),.A(g20924));
  NOT NOT1_611(.VSS(VSS),.VDD(VDD),.Y(g24685),.A(g23139));
  NOT NOT1_612(.VSS(VSS),.VDD(VDD),.Y(g24373),.A(g22908));
  NOT NOT1_613(.VSS(VSS),.VDD(VDD),.Y(I33024),.A(g34783));
  NOT NOT1_614(.VSS(VSS),.VDD(VDD),.Y(g8150),.A(g2185));
  NOT NOT1_615(.VSS(VSS),.VDD(VDD),.Y(g10401),.A(g7041));
  NOT NOT1_616(.VSS(VSS),.VDD(VDD),.Y(g22906),.A(g20453));
  NOT NOT1_617(.VSS(VSS),.VDD(VDD),.Y(g20654),.A(I20750));
  NOT NOT1_618(.VSS(VSS),.VDD(VDD),.Y(I16596),.A(g12640));
  NOT NOT1_619(.VSS(VSS),.VDD(VDD),.Y(g34317),.A(g34115));
  NOT NOT1_620(.VSS(VSS),.VDD(VDD),.Y(g8350),.A(g4646));
  NOT NOT1_621(.VSS(VSS),.VDD(VDD),.Y(g18908),.A(g16100));
  NOT NOT1_622(.VSS(VSS),.VDD(VDD),.Y(g32870),.A(g31021));
  NOT NOT1_623(.VSS(VSS),.VDD(VDD),.Y(g7535),.A(g1500));
  NOT NOT1_624(.VSS(VSS),.VDD(VDD),.Y(g32527),.A(g30673));
  NOT NOT1_625(.VSS(VSS),.VDD(VDD),.Y(I13007),.A(g65));
  NOT NOT1_626(.VSS(VSS),.VDD(VDD),.Y(g8038),.A(I12360));
  NOT NOT1_627(.VSS(VSS),.VDD(VDD),.Y(g10119),.A(g2841));
  NOT NOT1_628(.VSS(VSS),.VDD(VDD),.Y(I24474),.A(g22546));
  NOT NOT1_629(.VSS(VSS),.VDD(VDD),.Y(g16632),.A(g14454));
  NOT NOT1_630(.VSS(VSS),.VDD(VDD),.Y(g21308),.A(g17485));
  NOT NOT1_631(.VSS(VSS),.VDD(VDD),.Y(g8438),.A(g3100));
  NOT NOT1_632(.VSS(VSS),.VDD(VDD),.Y(g23571),.A(g18833));
  NOT NOT1_633(.VSS(VSS),.VDD(VDD),.Y(g28693),.A(g27837));
  NOT NOT1_634(.VSS(VSS),.VDD(VDD),.Y(g23308),.A(g21024));
  NOT NOT1_635(.VSS(VSS),.VDD(VDD),.Y(g31794),.A(I29368));
  NOT NOT1_636(.VSS(VSS),.VDD(VDD),.Y(g6972),.A(I11740));
  NOT NOT1_637(.VSS(VSS),.VDD(VDD),.Y(g31845),.A(g29385));
  NOT NOT1_638(.VSS(VSS),.VDD(VDD),.Y(g8009),.A(g3106));
  NOT NOT1_639(.VSS(VSS),.VDD(VDD),.Y(I31497),.A(g33187));
  NOT NOT1_640(.VSS(VSS),.VDD(VDD),.Y(g7261),.A(g4449));
  NOT NOT1_641(.VSS(VSS),.VDD(VDD),.Y(g24417),.A(g22171));
  NOT NOT1_642(.VSS(VSS),.VDD(VDD),.Y(g33845),.A(I31694));
  NOT NOT1_643(.VSS(VSS),.VDD(VDD),.Y(g10118),.A(g2541));
  NOT NOT1_644(.VSS(VSS),.VDD(VDD),.Y(I19775),.A(g17780));
  NOT NOT1_645(.VSS(VSS),.VDD(VDD),.Y(g9932),.A(g5805));
  NOT NOT1_646(.VSS(VSS),.VDD(VDD),.Y(g28166),.A(I26687));
  NOT NOT1_647(.VSS(VSS),.VDD(VDD),.Y(g28009),.A(I26516));
  NOT NOT1_648(.VSS(VSS),.VDD(VDD),.Y(g16661),.A(g14454));
  NOT NOT1_649(.VSS(VSS),.VDD(VDD),.Y(I17507),.A(g13416));
  NOT NOT1_650(.VSS(VSS),.VDD(VDD),.Y(g25549),.A(g22763));
  NOT NOT1_651(.VSS(VSS),.VDD(VDD),.Y(g13876),.A(g11432));
  NOT NOT1_652(.VSS(VSS),.VDD(VDD),.Y(g13885),.A(g10862));
  NOT NOT1_653(.VSS(VSS),.VDD(VDD),.Y(g32503),.A(g31194));
  NOT NOT1_654(.VSS(VSS),.VDD(VDD),.Y(g23495),.A(I22622));
  NOT NOT1_655(.VSS(VSS),.VDD(VDD),.Y(I31659),.A(g33219));
  NOT NOT1_656(.VSS(VSS),.VDD(VDD),.Y(g14749),.A(I16829));
  NOT NOT1_657(.VSS(VSS),.VDD(VDD),.Y(g32867),.A(g30673));
  NOT NOT1_658(.VSS(VSS),.VDD(VDD),.Y(g32894),.A(g30614));
  NOT NOT1_659(.VSS(VSS),.VDD(VDD),.Y(I31625),.A(g33197));
  NOT NOT1_660(.VSS(VSS),.VDD(VDD),.Y(g14616),.A(I16733));
  NOT NOT1_661(.VSS(VSS),.VDD(VDD),.Y(g34245),.A(I32234));
  NOT NOT1_662(.VSS(VSS),.VDD(VDD),.Y(I32953),.A(g34656));
  NOT NOT1_663(.VSS(VSS),.VDD(VDD),.Y(g8836),.A(g736));
  NOT NOT1_664(.VSS(VSS),.VDD(VDD),.Y(g30299),.A(g28765));
  NOT NOT1_665(.VSS(VSS),.VDD(VDD),.Y(g6887),.A(g3333));
  NOT NOT1_666(.VSS(VSS),.VDD(VDD),.Y(g23816),.A(g21308));
  NOT NOT1_667(.VSS(VSS),.VDD(VDD),.Y(g25548),.A(g22550));
  NOT NOT1_668(.VSS(VSS),.VDD(VDD),.Y(g34323),.A(g34105));
  NOT NOT1_669(.VSS(VSS),.VDD(VDD),.Y(g34299),.A(g34080));
  NOT NOT1_670(.VSS(VSS),.VDD(VDD),.Y(I32654),.A(g34378));
  NOT NOT1_671(.VSS(VSS),.VDD(VDD),.Y(g22139),.A(I21722));
  NOT NOT1_672(.VSS(VSS),.VDD(VDD),.Y(g8918),.A(I12893));
  NOT NOT1_673(.VSS(VSS),.VDD(VDD),.Y(g24964),.A(I24128));
  NOT NOT1_674(.VSS(VSS),.VDD(VDD),.Y(g7246),.A(g4446));
  NOT NOT1_675(.VSS(VSS),.VDD(VDD),.Y(I11746),.A(g4570));
  NOT NOT1_676(.VSS(VSS),.VDD(VDD),.Y(g26856),.A(I25586));
  NOT NOT1_677(.VSS(VSS),.VDD(VDD),.Y(g13763),.A(g10971));
  NOT NOT1_678(.VSS(VSS),.VDD(VDD),.Y(g14276),.A(I16452));
  NOT NOT1_679(.VSS(VSS),.VDD(VDD),.Y(g31521),.A(I29182));
  NOT NOT1_680(.VSS(VSS),.VDD(VDD),.Y(I32800),.A(g34582));
  NOT NOT1_681(.VSS(VSS),.VDD(VDD),.Y(g32581),.A(g31070));
  NOT NOT1_682(.VSS(VSS),.VDD(VDD),.Y(g32714),.A(g31528));
  NOT NOT1_683(.VSS(VSS),.VDD(VDD),.Y(g32450),.A(g31591));
  NOT NOT1_684(.VSS(VSS),.VDD(VDD),.Y(g10053),.A(g6381));
  NOT NOT1_685(.VSS(VSS),.VDD(VDD),.Y(g23985),.A(g19210));
  NOT NOT1_686(.VSS(VSS),.VDD(VDD),.Y(g22138),.A(g21370));
  NOT NOT1_687(.VSS(VSS),.VDD(VDD),.Y(g15739),.A(g13284));
  NOT NOT1_688(.VSS(VSS),.VDD(VDD),.Y(I26705),.A(g27967));
  NOT NOT1_689(.VSS(VSS),.VDD(VDD),.Y(g34775),.A(I32967));
  NOT NOT1_690(.VSS(VSS),.VDD(VDD),.Y(I20750),.A(g16677));
  NOT NOT1_691(.VSS(VSS),.VDD(VDD),.Y(g20587),.A(g15373));
  NOT NOT1_692(.VSS(VSS),.VDD(VDD),.Y(g32707),.A(g31579));
  NOT NOT1_693(.VSS(VSS),.VDD(VDD),.Y(g32819),.A(g30825));
  NOT NOT1_694(.VSS(VSS),.VDD(VDD),.Y(g9576),.A(g6565));
  NOT NOT1_695(.VSS(VSS),.VDD(VDD),.Y(g31832),.A(g29385));
  NOT NOT1_696(.VSS(VSS),.VDD(VDD),.Y(I20982),.A(g16300));
  NOT NOT1_697(.VSS(VSS),.VDD(VDD),.Y(g23954),.A(I23099));
  NOT NOT1_698(.VSS(VSS),.VDD(VDD),.Y(g24587),.A(g23112));
  NOT NOT1_699(.VSS(VSS),.VDD(VDD),.Y(g8229),.A(g3881));
  NOT NOT1_700(.VSS(VSS),.VDD(VDD),.Y(g9716),.A(g5057));
  NOT NOT1_701(.VSS(VSS),.VDD(VDD),.Y(I22788),.A(g18940));
  NOT NOT1_702(.VSS(VSS),.VDD(VDD),.Y(I26679),.A(g27773));
  NOT NOT1_703(.VSS(VSS),.VDD(VDD),.Y(g12863),.A(g10371));
  NOT NOT1_704(.VSS(VSS),.VDD(VDD),.Y(g8993),.A(g385));
  NOT NOT1_705(.VSS(VSS),.VDD(VDD),.Y(g15562),.A(g14943));
  NOT NOT1_706(.VSS(VSS),.VDD(VDD),.Y(g32818),.A(g30735));
  NOT NOT1_707(.VSS(VSS),.VDD(VDD),.Y(g10036),.A(g1816));
  NOT NOT1_708(.VSS(VSS),.VDD(VDD),.Y(g32496),.A(g30614));
  NOT NOT1_709(.VSS(VSS),.VDD(VDD),.Y(g19787),.A(g17096));
  NOT NOT1_710(.VSS(VSS),.VDD(VDD),.Y(g16127),.A(g13437));
  NOT NOT1_711(.VSS(VSS),.VDD(VDD),.Y(g8822),.A(g4975));
  NOT NOT1_712(.VSS(VSS),.VDD(VDD),.Y(g10177),.A(g1834));
  NOT NOT1_713(.VSS(VSS),.VDD(VDD),.Y(g20909),.A(g17955));
  NOT NOT1_714(.VSS(VSS),.VDD(VDD),.Y(g20543),.A(g17955));
  NOT NOT1_715(.VSS(VSS),.VDD(VDD),.Y(I13684),.A(g128));
  NOT NOT1_716(.VSS(VSS),.VDD(VDD),.Y(g31861),.A(I29441));
  NOT NOT1_717(.VSS(VSS),.VDD(VDD),.Y(g9848),.A(g4462));
  NOT NOT1_718(.VSS(VSS),.VDD(VDD),.Y(g21669),.A(I21230));
  NOT NOT1_719(.VSS(VSS),.VDD(VDD),.Y(g19357),.A(I19837));
  NOT NOT1_720(.VSS(VSS),.VDD(VDD),.Y(g17415),.A(g14797));
  NOT NOT1_721(.VSS(VSS),.VDD(VDD),.Y(g6845),.A(g2126));
  NOT NOT1_722(.VSS(VSS),.VDD(VDD),.Y(g7502),.A(I11992));
  NOT NOT1_723(.VSS(VSS),.VDD(VDD),.Y(I15550),.A(g10430));
  NOT NOT1_724(.VSS(VSS),.VDD(VDD),.Y(g32590),.A(g31154));
  NOT NOT1_725(.VSS(VSS),.VDD(VDD),.Y(g9699),.A(g2311));
  NOT NOT1_726(.VSS(VSS),.VDD(VDD),.Y(g9747),.A(I13329));
  NOT NOT1_727(.VSS(VSS),.VDD(VDD),.Y(g24117),.A(g21209));
  NOT NOT1_728(.VSS(VSS),.VDD(VDD),.Y(g24000),.A(g19277));
  NOT NOT1_729(.VSS(VSS),.VDD(VDD),.Y(I33197),.A(g34930));
  NOT NOT1_730(.VSS(VSS),.VDD(VDD),.Y(g23260),.A(g21070));
  NOT NOT1_731(.VSS(VSS),.VDD(VDD),.Y(g19743),.A(g17125));
  NOT NOT1_732(.VSS(VSS),.VDD(VDD),.Y(I14584),.A(g9766));
  NOT NOT1_733(.VSS(VSS),.VDD(VDD),.Y(g33926),.A(I31796));
  NOT NOT1_734(.VSS(VSS),.VDD(VDD),.Y(g25245),.A(g22763));
  NOT NOT1_735(.VSS(VSS),.VDD(VDD),.Y(g34697),.A(g34545));
  NOT NOT1_736(.VSS(VSS),.VDD(VDD),.Y(g26831),.A(g24836));
  NOT NOT1_737(.VSS(VSS),.VDD(VDD),.Y(g20569),.A(g15277));
  NOT NOT1_738(.VSS(VSS),.VDD(VDD),.Y(I20840),.A(g17727));
  NOT NOT1_739(.VSS(VSS),.VDD(VDD),.Y(g34995),.A(I33285));
  NOT NOT1_740(.VSS(VSS),.VDD(VDD),.Y(g23842),.A(g19147));
  NOT NOT1_741(.VSS(VSS),.VDD(VDD),.Y(g32741),.A(g31710));
  NOT NOT1_742(.VSS(VSS),.VDD(VDD),.Y(g13314),.A(g10893));
  NOT NOT1_743(.VSS(VSS),.VDD(VDD),.Y(I23348),.A(g23384));
  NOT NOT1_744(.VSS(VSS),.VDD(VDD),.Y(g25299),.A(g22763));
  NOT NOT1_745(.VSS(VSS),.VDD(VDD),.Y(g32384),.A(g31666));
  NOT NOT1_746(.VSS(VSS),.VDD(VDD),.Y(I19831),.A(g16533));
  NOT NOT1_747(.VSS(VSS),.VDD(VDD),.Y(g33388),.A(g32382));
  NOT NOT1_748(.VSS(VSS),.VDD(VDD),.Y(I18252),.A(g13177));
  NOT NOT1_749(.VSS(VSS),.VDD(VDD),.Y(I16502),.A(g10430));
  NOT NOT1_750(.VSS(VSS),.VDD(VDD),.Y(g20568),.A(g15509));
  NOT NOT1_751(.VSS(VSS),.VDD(VDD),.Y(g23489),.A(g21468));
  NOT NOT1_752(.VSS(VSS),.VDD(VDD),.Y(g25533),.A(g22550));
  NOT NOT1_753(.VSS(VSS),.VDD(VDD),.Y(g13085),.A(I15717));
  NOT NOT1_754(.VSS(VSS),.VDD(VDD),.Y(g19769),.A(g16987));
  NOT NOT1_755(.VSS(VSS),.VDD(VDD),.Y(g24568),.A(g22942));
  NOT NOT1_756(.VSS(VSS),.VDD(VDD),.Y(g20242),.A(g16308));
  NOT NOT1_757(.VSS(VSS),.VDD(VDD),.Y(g25298),.A(g23760));
  NOT NOT1_758(.VSS(VSS),.VDD(VDD),.Y(g11721),.A(g10074));
  NOT NOT1_759(.VSS(VSS),.VDD(VDD),.Y(g7689),.A(I12159));
  NOT NOT1_760(.VSS(VSS),.VDD(VDD),.Y(g29927),.A(g28861));
  NOT NOT1_761(.VSS(VSS),.VDD(VDD),.Y(I17121),.A(g14366));
  NOT NOT1_762(.VSS(VSS),.VDD(VDD),.Y(g34512),.A(g34420));
  NOT NOT1_763(.VSS(VSS),.VDD(VDD),.Y(g21424),.A(g15426));
  NOT NOT1_764(.VSS(VSS),.VDD(VDD),.Y(g23559),.A(g21070));
  NOT NOT1_765(.VSS(VSS),.VDD(VDD),.Y(g13596),.A(g10971));
  NOT NOT1_766(.VSS(VSS),.VDD(VDD),.Y(g23525),.A(g21562));
  NOT NOT1_767(.VSS(VSS),.VDD(VDD),.Y(g23488),.A(g21468));
  NOT NOT1_768(.VSS(VSS),.VDD(VDD),.Y(g28675),.A(g27779));
  NOT NOT1_769(.VSS(VSS),.VDD(VDD),.Y(g23016),.A(g20453));
  NOT NOT1_770(.VSS(VSS),.VDD(VDD),.Y(I32909),.A(g34712));
  NOT NOT1_771(.VSS(VSS),.VDD(VDD),.Y(g7216),.A(g822));
  NOT NOT1_772(.VSS(VSS),.VDD(VDD),.Y(g11431),.A(g7618));
  NOT NOT1_773(.VSS(VSS),.VDD(VDD),.Y(g12952),.A(I15572));
  NOT NOT1_774(.VSS(VSS),.VDD(VDD),.Y(g23558),.A(g20924));
  NOT NOT1_775(.VSS(VSS),.VDD(VDD),.Y(g13431),.A(I15932));
  NOT NOT1_776(.VSS(VSS),.VDD(VDD),.Y(g32801),.A(g30937));
  NOT NOT1_777(.VSS(VSS),.VDD(VDD),.Y(g14630),.A(g12402));
  NOT NOT1_778(.VSS(VSS),.VDD(VDD),.Y(g32735),.A(g31021));
  NOT NOT1_779(.VSS(VSS),.VDD(VDD),.Y(g24123),.A(g21143));
  NOT NOT1_780(.VSS(VSS),.VDD(VDD),.Y(g32877),.A(g30825));
  NOT NOT1_781(.VSS(VSS),.VDD(VDD),.Y(g7028),.A(I11785));
  NOT NOT1_782(.VSS(VSS),.VDD(VDD),.Y(I30686),.A(g32381));
  NOT NOT1_783(.VSS(VSS),.VDD(VDD),.Y(g8895),.A(g599));
  NOT NOT1_784(.VSS(VSS),.VDD(VDD),.Y(g10166),.A(g6040));
  NOT NOT1_785(.VSS(VSS),.VDD(VDD),.Y(g17576),.A(g14953));
  NOT NOT1_786(.VSS(VSS),.VDD(VDD),.Y(g17585),.A(g14974));
  NOT NOT1_787(.VSS(VSS),.VDD(VDD),.Y(g20772),.A(g15171));
  NOT NOT1_788(.VSS(VSS),.VDD(VDD),.Y(g9644),.A(g2016));
  NOT NOT1_789(.VSS(VSS),.VDD(VDD),.Y(g22200),.A(g19277));
  NOT NOT1_790(.VSS(VSS),.VDD(VDD),.Y(g23893),.A(g19074));
  NOT NOT1_791(.VSS(VSS),.VDD(VDD),.Y(I15773),.A(g10430));
  NOT NOT1_792(.VSS(VSS),.VDD(VDD),.Y(g11269),.A(g7516));
  NOT NOT1_793(.VSS(VSS),.VDD(VDD),.Y(I15942),.A(g12381));
  NOT NOT1_794(.VSS(VSS),.VDD(VDD),.Y(g14166),.A(g11048));
  NOT NOT1_795(.VSS(VSS),.VDD(VDD),.Y(g8620),.A(g3065));
  NOT NOT1_796(.VSS(VSS),.VDD(VDD),.Y(g19881),.A(g15915));
  NOT NOT1_797(.VSS(VSS),.VDD(VDD),.Y(g8462),.A(g1183));
  NOT NOT1_798(.VSS(VSS),.VDD(VDD),.Y(g25232),.A(g22228));
  NOT NOT1_799(.VSS(VSS),.VDD(VDD),.Y(g29491),.A(I27777));
  NOT NOT1_800(.VSS(VSS),.VDD(VDD),.Y(g7247),.A(g5377));
  NOT NOT1_801(.VSS(VSS),.VDD(VDD),.Y(g20639),.A(g15224));
  NOT NOT1_802(.VSS(VSS),.VDD(VDD),.Y(I17173),.A(g13716));
  NOT NOT1_803(.VSS(VSS),.VDD(VDD),.Y(g16931),.A(I18101));
  NOT NOT1_804(.VSS(VSS),.VDD(VDD),.Y(I16468),.A(g12760));
  NOT NOT1_805(.VSS(VSS),.VDD(VDD),.Y(g23544),.A(g21562));
  NOT NOT1_806(.VSS(VSS),.VDD(VDD),.Y(g23865),.A(g21308));
  NOT NOT1_807(.VSS(VSS),.VDD(VDD),.Y(I12046),.A(g613));
  NOT NOT1_808(.VSS(VSS),.VDD(VDD),.Y(g32695),.A(g30735));
  NOT NOT1_809(.VSS(VSS),.VDD(VDD),.Y(I31581),.A(g33164));
  NOT NOT1_810(.VSS(VSS),.VDD(VDD),.Y(g11268),.A(g7515));
  NOT NOT1_811(.VSS(VSS),.VDD(VDD),.Y(g20230),.A(I20499));
  NOT NOT1_812(.VSS(VSS),.VDD(VDD),.Y(g12790),.A(g7097));
  NOT NOT1_813(.VSS(VSS),.VDD(VDD),.Y(g17609),.A(g14817));
  NOT NOT1_814(.VSS(VSS),.VDD(VDD),.Y(g29755),.A(I28002));
  NOT NOT1_815(.VSS(VSS),.VDD(VDD),.Y(g7564),.A(g336));
  NOT NOT1_816(.VSS(VSS),.VDD(VDD),.Y(g9152),.A(g2834));
  NOT NOT1_817(.VSS(VSS),.VDD(VDD),.Y(g20638),.A(g15224));
  NOT NOT1_818(.VSS(VSS),.VDD(VDD),.Y(I18509),.A(g5623));
  NOT NOT1_819(.VSS(VSS),.VDD(VDD),.Y(g9818),.A(g6490));
  NOT NOT1_820(.VSS(VSS),.VDD(VDD),.Y(g13655),.A(g10573));
  NOT NOT1_821(.VSS(VSS),.VDD(VDD),.Y(g34316),.A(g34093));
  NOT NOT1_822(.VSS(VSS),.VDD(VDD),.Y(g17200),.A(I18238));
  NOT NOT1_823(.VSS(VSS),.VDD(VDD),.Y(g32526),.A(g30614));
  NOT NOT1_824(.VSS(VSS),.VDD(VDD),.Y(g20265),.A(g17821));
  NOT NOT1_825(.VSS(VSS),.VDD(VDD),.Y(g29981),.A(g28942));
  NOT NOT1_826(.VSS(VSS),.VDD(VDD),.Y(g6815),.A(g929));
  NOT NOT1_827(.VSS(VSS),.VDD(VDD),.Y(I12787),.A(g4311));
  NOT NOT1_828(.VSS(VSS),.VDD(VDD),.Y(g12873),.A(g10380));
  NOT NOT1_829(.VSS(VSS),.VDD(VDD),.Y(I22028),.A(g20204));
  NOT NOT1_830(.VSS(VSS),.VDD(VDD),.Y(I29211),.A(g30298));
  NOT NOT1_831(.VSS(VSS),.VDD(VDD),.Y(g8788),.A(I12776));
  NOT NOT1_832(.VSS(VSS),.VDD(VDD),.Y(I18872),.A(g13745));
  NOT NOT1_833(.VSS(VSS),.VDD(VDD),.Y(I23333),.A(g22683));
  NOT NOT1_834(.VSS(VSS),.VDD(VDD),.Y(g30989),.A(g29672));
  NOT NOT1_835(.VSS(VSS),.VDD(VDD),.Y(g33766),.A(I31619));
  NOT NOT1_836(.VSS(VSS),.VDD(VDD),.Y(g19662),.A(g17432));
  NOT NOT1_837(.VSS(VSS),.VDD(VDD),.Y(g21610),.A(g15615));
  NOT NOT1_838(.VSS(VSS),.VDD(VDD),.Y(g14454),.A(I16613));
  NOT NOT1_839(.VSS(VSS),.VDD(VDD),.Y(g23610),.A(g18833));
  NOT NOT1_840(.VSS(VSS),.VDD(VDD),.Y(g10570),.A(g9021));
  NOT NOT1_841(.VSS(VSS),.VDD(VDD),.Y(g34989),.A(I33267));
  NOT NOT1_842(.VSS(VSS),.VDD(VDD),.Y(g8249),.A(g1917));
  NOT NOT1_843(.VSS(VSS),.VDD(VDD),.Y(g20391),.A(I20562));
  NOT NOT1_844(.VSS(VSS),.VDD(VDD),.Y(g32457),.A(g30735));
  NOT NOT1_845(.VSS(VSS),.VDD(VDD),.Y(g21189),.A(g15634));
  NOT NOT1_846(.VSS(VSS),.VDD(VDD),.Y(g24992),.A(g22417));
  NOT NOT1_847(.VSS(VSS),.VDD(VDD),.Y(I33070),.A(g34810));
  NOT NOT1_848(.VSS(VSS),.VDD(VDD),.Y(g20510),.A(g17226));
  NOT NOT1_849(.VSS(VSS),.VDD(VDD),.Y(g23189),.A(g20060));
  NOT NOT1_850(.VSS(VSS),.VDD(VDD),.Y(g11930),.A(g9281));
  NOT NOT1_851(.VSS(VSS),.VDD(VDD),.Y(g12422),.A(I15238));
  NOT NOT1_852(.VSS(VSS),.VDD(VDD),.Y(g26736),.A(g25349));
  NOT NOT1_853(.VSS(VSS),.VDD(VDD),.Y(g9186),.A(I13010));
  NOT NOT1_854(.VSS(VSS),.VDD(VDD),.Y(g17745),.A(g14978));
  NOT NOT1_855(.VSS(VSS),.VDD(VDD),.Y(g34988),.A(I33264));
  NOT NOT1_856(.VSS(VSS),.VDD(VDD),.Y(g22973),.A(g20330));
  NOT NOT1_857(.VSS(VSS),.VDD(VDD),.Y(g34924),.A(I33164));
  NOT NOT1_858(.VSS(VSS),.VDD(VDD),.Y(g6960),.A(g1));
  NOT NOT1_859(.VSS(VSS),.VDD(VDD),.Y(g9386),.A(g5727));
  NOT NOT1_860(.VSS(VSS),.VDD(VDD),.Y(I15667),.A(g12143));
  NOT NOT1_861(.VSS(VSS),.VDD(VDD),.Y(I32639),.A(g34345));
  NOT NOT1_862(.VSS(VSS),.VDD(VDD),.Y(g21270),.A(I20999));
  NOT NOT1_863(.VSS(VSS),.VDD(VDD),.Y(g32866),.A(g30614));
  NOT NOT1_864(.VSS(VSS),.VDD(VDD),.Y(g32917),.A(g30937));
  NOT NOT1_865(.VSS(VSS),.VDD(VDD),.Y(g23270),.A(g20785));
  NOT NOT1_866(.VSS(VSS),.VDD(VDD),.Y(g19482),.A(g16349));
  NOT NOT1_867(.VSS(VSS),.VDD(VDD),.Y(g21678),.A(g16540));
  NOT NOT1_868(.VSS(VSS),.VDD(VDD),.Y(g17813),.A(I18813));
  NOT NOT1_869(.VSS(VSS),.VDD(VDD),.Y(g12834),.A(g10349));
  NOT NOT1_870(.VSS(VSS),.VDD(VDD),.Y(g20579),.A(g17249));
  NOT NOT1_871(.VSS(VSS),.VDD(VDD),.Y(g34432),.A(I32467));
  NOT NOT1_872(.VSS(VSS),.VDD(VDD),.Y(g7308),.A(g1668));
  NOT NOT1_873(.VSS(VSS),.VDD(VDD),.Y(g11965),.A(I14797));
  NOT NOT1_874(.VSS(VSS),.VDD(VDD),.Y(g8085),.A(I12382));
  NOT NOT1_875(.VSS(VSS),.VDD(VDD),.Y(g9599),.A(g3310));
  NOT NOT1_876(.VSS(VSS),.VDD(VDD),.Y(g10074),.A(g718));
  NOT NOT1_877(.VSS(VSS),.VDD(VDD),.Y(g19710),.A(g17059));
  NOT NOT1_878(.VSS(VSS),.VDD(VDD),.Y(g18983),.A(g16077));
  NOT NOT1_879(.VSS(VSS),.VDD(VDD),.Y(g24579),.A(g23067));
  NOT NOT1_880(.VSS(VSS),.VDD(VDD),.Y(g34271),.A(g34160));
  NOT NOT1_881(.VSS(VSS),.VDD(VDD),.Y(g19552),.A(g16856));
  NOT NOT1_882(.VSS(VSS),.VDD(VDD),.Y(g21460),.A(g15628));
  NOT NOT1_883(.VSS(VSS),.VDD(VDD),.Y(g21686),.A(g16540));
  NOT NOT1_884(.VSS(VSS),.VDD(VDD),.Y(g9274),.A(g5857));
  NOT NOT1_885(.VSS(VSS),.VDD(VDD),.Y(g20578),.A(g15563));
  NOT NOT1_886(.VSS(VSS),.VDD(VDD),.Y(g26843),.A(I25567));
  NOT NOT1_887(.VSS(VSS),.VDD(VDD),.Y(g23460),.A(g21611));
  NOT NOT1_888(.VSS(VSS),.VDD(VDD),.Y(g23939),.A(g19074));
  NOT NOT1_889(.VSS(VSS),.VDD(VDD),.Y(g21383),.A(g17367));
  NOT NOT1_890(.VSS(VSS),.VDD(VDD),.Y(g19779),.A(g16431));
  NOT NOT1_891(.VSS(VSS),.VDD(VDD),.Y(I19843),.A(g16594));
  NOT NOT1_892(.VSS(VSS),.VDD(VDD),.Y(g9614),.A(g5128));
  NOT NOT1_893(.VSS(VSS),.VDD(VDD),.Y(I33067),.A(g34812));
  NOT NOT1_894(.VSS(VSS),.VDD(VDD),.Y(g17674),.A(I18647));
  NOT NOT1_895(.VSS(VSS),.VDD(VDD),.Y(g12021),.A(g9543));
  NOT NOT1_896(.VSS(VSS),.VDD(VDD),.Y(g14238),.A(g10823));
  NOT NOT1_897(.VSS(VSS),.VDD(VDD),.Y(g20586),.A(g15171));
  NOT NOT1_898(.VSS(VSS),.VDD(VDD),.Y(g23030),.A(g20453));
  NOT NOT1_899(.VSS(VSS),.VDD(VDD),.Y(g32706),.A(g30673));
  NOT NOT1_900(.VSS(VSS),.VDD(VDD),.Y(g23938),.A(g18997));
  NOT NOT1_901(.VSS(VSS),.VDD(VDD),.Y(g32597),.A(g31154));
  NOT NOT1_902(.VSS(VSS),.VDD(VDD),.Y(I18574),.A(g13075));
  NOT NOT1_903(.VSS(VSS),.VDD(VDD),.Y(g25316),.A(g22763));
  NOT NOT1_904(.VSS(VSS),.VDD(VDD),.Y(g8854),.A(g613));
  NOT NOT1_905(.VSS(VSS),.VDD(VDD),.Y(g21267),.A(g15680));
  NOT NOT1_906(.VSS(VSS),.VDD(VDD),.Y(g24586),.A(g23067));
  NOT NOT1_907(.VSS(VSS),.VDD(VDD),.Y(I32391),.A(g34153));
  NOT NOT1_908(.VSS(VSS),.VDD(VDD),.Y(g23267),.A(g20097));
  NOT NOT1_909(.VSS(VSS),.VDD(VDD),.Y(g9821),.A(g115));
  NOT NOT1_910(.VSS(VSS),.VDD(VDD),.Y(I13236),.A(g5452));
  NOT NOT1_911(.VSS(VSS),.VDD(VDD),.Y(I18205),.A(g14563));
  NOT NOT1_912(.VSS(VSS),.VDD(VDD),.Y(g34145),.A(I32096));
  NOT NOT1_913(.VSS(VSS),.VDD(VDD),.Y(I16168),.A(g3321));
  NOT NOT1_914(.VSS(VSS),.VDD(VDD),.Y(g26869),.A(g24842));
  NOT NOT1_915(.VSS(VSS),.VDD(VDD),.Y(g32689),.A(g30825));
  NOT NOT1_916(.VSS(VSS),.VDD(VDD),.Y(g15824),.A(I17324));
  NOT NOT1_917(.VSS(VSS),.VDD(VDD),.Y(g20442),.A(g15171));
  NOT NOT1_918(.VSS(VSS),.VDD(VDD),.Y(g10382),.A(g6958));
  NOT NOT1_919(.VSS(VSS),.VDD(VDD),.Y(I18912),.A(g15050));
  NOT NOT1_920(.VSS(VSS),.VDD(VDD),.Y(I22240),.A(g20086));
  NOT NOT1_921(.VSS(VSS),.VDD(VDD),.Y(g32923),.A(g31021));
  NOT NOT1_922(.VSS(VSS),.VDD(VDD),.Y(g33451),.A(g32132));
  NOT NOT1_923(.VSS(VSS),.VDD(VDD),.Y(g19786),.A(g17062));
  NOT NOT1_924(.VSS(VSS),.VDD(VDD),.Y(I14833),.A(g10142));
  NOT NOT1_925(.VSS(VSS),.VDD(VDD),.Y(g16659),.A(I17857));
  NOT NOT1_926(.VSS(VSS),.VDD(VDD),.Y(g12614),.A(g9935));
  NOT NOT1_927(.VSS(VSS),.VDD(VDD),.Y(g22761),.A(g21024));
  NOT NOT1_928(.VSS(VSS),.VDD(VDD),.Y(g9280),.A(I13054));
  NOT NOT1_929(.VSS(VSS),.VDD(VDD),.Y(g10519),.A(g9326));
  NOT NOT1_930(.VSS(VSS),.VDD(VDD),.Y(g34736),.A(I32904));
  NOT NOT1_931(.VSS(VSS),.VDD(VDD),.Y(g10176),.A(g44));
  NOT NOT1_932(.VSS(VSS),.VDD(VDD),.Y(I16479),.A(g10430));
  NOT NOT1_933(.VSS(VSS),.VDD(VDD),.Y(g27320),.A(I26004));
  NOT NOT1_934(.VSS(VSS),.VDD(VDD),.Y(g16987),.A(I18135));
  NOT NOT1_935(.VSS(VSS),.VDD(VDD),.Y(g32688),.A(g30735));
  NOT NOT1_936(.VSS(VSS),.VDD(VDD),.Y(g32624),.A(g30825));
  NOT NOT1_937(.VSS(VSS),.VDD(VDD),.Y(I23312),.A(g21681));
  NOT NOT1_938(.VSS(VSS),.VDD(VDD),.Y(g13279),.A(I15843));
  NOT NOT1_939(.VSS(VSS),.VDD(VDD),.Y(I16217),.A(g3632));
  NOT NOT1_940(.VSS(VSS),.VDD(VDD),.Y(I21115),.A(g15714));
  NOT NOT1_941(.VSS(VSS),.VDD(VDD),.Y(g16658),.A(g14157));
  NOT NOT1_942(.VSS(VSS),.VDD(VDD),.Y(I22604),.A(g21143));
  NOT NOT1_943(.VSS(VSS),.VDD(VDD),.Y(g10518),.A(g9311));
  NOT NOT1_944(.VSS(VSS),.VDD(VDD),.Y(g10154),.A(g2547));
  NOT NOT1_945(.VSS(VSS),.VDD(VDD),.Y(g12905),.A(g10408));
  NOT NOT1_946(.VSS(VSS),.VDD(VDD),.Y(g20615),.A(g15509));
  NOT NOT1_947(.VSS(VSS),.VDD(VDD),.Y(g33246),.A(g32212));
  NOT NOT1_948(.VSS(VSS),.VDD(VDD),.Y(g9083),.A(g626));
  NOT NOT1_949(.VSS(VSS),.VDD(VDD),.Y(g23875),.A(g18997));
  NOT NOT1_950(.VSS(VSS),.VDD(VDD),.Y(g25080),.A(g23742));
  NOT NOT1_951(.VSS(VSS),.VDD(VDD),.Y(g24116),.A(g21143));
  NOT NOT1_952(.VSS(VSS),.VDD(VDD),.Y(g14518),.A(I16639));
  NOT NOT1_953(.VSS(VSS),.VDD(VDD),.Y(g23219),.A(I22316));
  NOT NOT1_954(.VSS(VSS),.VDD(VDD),.Y(I18051),.A(g13680));
  NOT NOT1_955(.VSS(VSS),.VDD(VDD),.Y(g30330),.A(I28591));
  NOT NOT1_956(.VSS(VSS),.VDD(VDD),.Y(g13278),.A(g10738));
  NOT NOT1_957(.VSS(VSS),.VDD(VDD),.Y(g26709),.A(g25435));
  NOT NOT1_958(.VSS(VSS),.VDD(VDD),.Y(I29969),.A(g30991));
  NOT NOT1_959(.VSS(VSS),.VDD(VDD),.Y(g8219),.A(g3731));
  NOT NOT1_960(.VSS(VSS),.VDD(VDD),.Y(g27565),.A(g26645));
  NOT NOT1_961(.VSS(VSS),.VDD(VDD),.Y(I17491),.A(g13416));
  NOT NOT1_962(.VSS(VSS),.VDD(VDD),.Y(I16486),.A(g11204));
  NOT NOT1_963(.VSS(VSS),.VDD(VDD),.Y(g20041),.A(g15569));
  NOT NOT1_964(.VSS(VSS),.VDD(VDD),.Y(g9636),.A(g72));
  NOT NOT1_965(.VSS(VSS),.VDD(VDD),.Y(g22214),.A(g19210));
  NOT NOT1_966(.VSS(VSS),.VDD(VDD),.Y(g7827),.A(g4688));
  NOT NOT1_967(.VSS(VSS),.VDD(VDD),.Y(g12122),.A(g9705));
  NOT NOT1_968(.VSS(VSS),.VDD(VDD),.Y(g20275),.A(g17929));
  NOT NOT1_969(.VSS(VSS),.VDD(VDD),.Y(g24041),.A(g19968));
  NOT NOT1_970(.VSS(VSS),.VDD(VDD),.Y(g19998),.A(g15915));
  NOT NOT1_971(.VSS(VSS),.VDD(VDD),.Y(g8431),.A(g3085));
  NOT NOT1_972(.VSS(VSS),.VDD(VDD),.Y(g11468),.A(g7624));
  NOT NOT1_973(.VSS(VSS),.VDD(VDD),.Y(g16644),.A(I17842));
  NOT NOT1_974(.VSS(VSS),.VDD(VDD),.Y(g13039),.A(I15663));
  NOT NOT1_975(.VSS(VSS),.VDD(VDD),.Y(g8812),.A(I12805));
  NOT NOT1_976(.VSS(VSS),.VDD(VDD),.Y(g15426),.A(I17121));
  NOT NOT1_977(.VSS(VSS),.VDD(VDD),.Y(g22207),.A(I21787));
  NOT NOT1_978(.VSS(VSS),.VDD(VDD),.Y(g6828),.A(g1300));
  NOT NOT1_979(.VSS(VSS),.VDD(VDD),.Y(g19672),.A(g16931));
  NOT NOT1_980(.VSS(VSS),.VDD(VDD),.Y(g34132),.A(g33831));
  NOT NOT1_981(.VSS(VSS),.VDD(VDD),.Y(g17400),.A(I18333));
  NOT NOT1_982(.VSS(VSS),.VDD(VDD),.Y(I12890),.A(g4219));
  NOT NOT1_983(.VSS(VSS),.VDD(VDD),.Y(g29045),.A(g27779));
  NOT NOT1_984(.VSS(VSS),.VDD(VDD),.Y(g34960),.A(I33218));
  NOT NOT1_985(.VSS(VSS),.VDD(VDD),.Y(g11038),.A(g8632));
  NOT NOT1_986(.VSS(VSS),.VDD(VDD),.Y(g16969),.A(g14262));
  NOT NOT1_987(.VSS(VSS),.VDD(VDD),.Y(g6830),.A(g1389));
  NOT NOT1_988(.VSS(VSS),.VDD(VDD),.Y(g17013),.A(g14262));
  NOT NOT1_989(.VSS(VSS),.VDD(VDD),.Y(I18350),.A(g13716));
  NOT NOT1_990(.VSS(VSS),.VDD(VDD),.Y(g8005),.A(g3025));
  NOT NOT1_991(.VSS(VSS),.VDD(VDD),.Y(g20237),.A(g17213));
  NOT NOT1_992(.VSS(VSS),.VDD(VDD),.Y(g21160),.A(g17508));
  NOT NOT1_993(.VSS(VSS),.VDD(VDD),.Y(g7196),.A(I11860));
  NOT NOT1_994(.VSS(VSS),.VDD(VDD),.Y(g11815),.A(g7582));
  NOT NOT1_995(.VSS(VSS),.VDD(VDD),.Y(g8405),.A(I12572));
  NOT NOT1_996(.VSS(VSS),.VDD(VDD),.Y(g9187),.A(g518));
  NOT NOT1_997(.VSS(VSS),.VDD(VDD),.Y(g16968),.A(g14238));
  NOT NOT1_998(.VSS(VSS),.VDD(VDD),.Y(I27552),.A(g28162));
  NOT NOT1_999(.VSS(VSS),.VDD(VDD),.Y(I15677),.A(g5654));
  NOT NOT1_1000(.VSS(VSS),.VDD(VDD),.Y(g31859),.A(g29385));
  NOT NOT1_1001(.VSS(VSS),.VDD(VDD),.Y(I32116),.A(g33937));
  NOT NOT1_1002(.VSS(VSS),.VDD(VDD),.Y(g20035),.A(g16430));
  NOT NOT1_1003(.VSS(VSS),.VDD(VDD),.Y(g31825),.A(g29385));
  NOT NOT1_1004(.VSS(VSS),.VDD(VDD),.Y(g32876),.A(g30735));
  NOT NOT1_1005(.VSS(VSS),.VDD(VDD),.Y(g32885),.A(g31021));
  NOT NOT1_1006(.VSS(VSS),.VDD(VDD),.Y(g34161),.A(g33851));
  NOT NOT1_1007(.VSS(VSS),.VDD(VDD),.Y(g16197),.A(g13861));
  NOT NOT1_1008(.VSS(VSS),.VDD(VDD),.Y(g24035),.A(g20841));
  NOT NOT1_1009(.VSS(VSS),.VDD(VDD),.Y(g11677),.A(g7689));
  NOT NOT1_1010(.VSS(VSS),.VDD(VDD),.Y(g21455),.A(g15426));
  NOT NOT1_1011(.VSS(VSS),.VDD(VDD),.Y(I12003),.A(g767));
  NOT NOT1_1012(.VSS(VSS),.VDD(VDD),.Y(g8286),.A(g53));
  NOT NOT1_1013(.VSS(VSS),.VDD(VDD),.Y(g8765),.A(g3333));
  NOT NOT1_1014(.VSS(VSS),.VDD(VDD),.Y(g17328),.A(I18313));
  NOT NOT1_1015(.VSS(VSS),.VDD(VDD),.Y(g31858),.A(g29385));
  NOT NOT1_1016(.VSS(VSS),.VDD(VDD),.Y(g13975),.A(g11048));
  NOT NOT1_1017(.VSS(VSS),.VDD(VDD),.Y(g32854),.A(g30735));
  NOT NOT1_1018(.VSS(VSS),.VDD(VDD),.Y(g7780),.A(g2878));
  NOT NOT1_1019(.VSS(VSS),.VDD(VDD),.Y(I12779),.A(g4210));
  NOT NOT1_1020(.VSS(VSS),.VDD(VDD),.Y(g16527),.A(g14048));
  NOT NOT1_1021(.VSS(VSS),.VDD(VDD),.Y(g25198),.A(g22228));
  NOT NOT1_1022(.VSS(VSS),.VDD(VDD),.Y(g30259),.A(g28463));
  NOT NOT1_1023(.VSS(VSS),.VDD(VDD),.Y(g25529),.A(g22763));
  NOT NOT1_1024(.VSS(VSS),.VDD(VDD),.Y(g14215),.A(g12198));
  NOT NOT1_1025(.VSS(VSS),.VDD(VDD),.Y(g32511),.A(g30614));
  NOT NOT1_1026(.VSS(VSS),.VDD(VDD),.Y(g23915),.A(g19277));
  NOT NOT1_1027(.VSS(VSS),.VDD(VDD),.Y(g32763),.A(g31710));
  NOT NOT1_1028(.VSS(VSS),.VDD(VDD),.Y(I15937),.A(g11676));
  NOT NOT1_1029(.VSS(VSS),.VDD(VDD),.Y(I17395),.A(g12952));
  NOT NOT1_1030(.VSS(VSS),.VDD(VDD),.Y(I28434),.A(g28114));
  NOT NOT1_1031(.VSS(VSS),.VDD(VDD),.Y(g30087),.A(g29121));
  NOT NOT1_1032(.VSS(VSS),.VDD(VDD),.Y(g11143),.A(g8032));
  NOT NOT1_1033(.VSS(VSS),.VDD(VDD),.Y(g19961),.A(g17328));
  NOT NOT1_1034(.VSS(VSS),.VDD(VDD),.Y(g26810),.A(g25220));
  NOT NOT1_1035(.VSS(VSS),.VDD(VDD),.Y(I29894),.A(g31771));
  NOT NOT1_1036(.VSS(VSS),.VDD(VDD),.Y(I14033),.A(g8912));
  NOT NOT1_1037(.VSS(VSS),.VDD(VDD),.Y(g34471),.A(g34423));
  NOT NOT1_1038(.VSS(VSS),.VDD(VDD),.Y(g9200),.A(g1548));
  NOT NOT1_1039(.VSS(VSS),.VDD(VDD),.Y(g25528),.A(g22594));
  NOT NOT1_1040(.VSS(VSS),.VDD(VDD),.Y(I21934),.A(g21273));
  NOT NOT1_1041(.VSS(VSS),.VDD(VDD),.Y(g31844),.A(g29385));
  NOT NOT1_1042(.VSS(VSS),.VDD(VDD),.Y(I31597),.A(g33187));
  NOT NOT1_1043(.VSS(VSS),.VDD(VDD),.Y(g8733),.A(g3698));
  NOT NOT1_1044(.VSS(VSS),.VDD(VDD),.Y(g19505),.A(g16349));
  NOT NOT1_1045(.VSS(VSS),.VDD(VDD),.Y(g23277),.A(I22380));
  NOT NOT1_1046(.VSS(VSS),.VDD(VDD),.Y(g7018),.A(g5297));
  NOT NOT1_1047(.VSS(VSS),.VDD(VDD),.Y(g8974),.A(I12930));
  NOT NOT1_1048(.VSS(VSS),.VDD(VDD),.Y(I11726),.A(g4273));
  NOT NOT1_1049(.VSS(VSS),.VDD(VDD),.Y(I32237),.A(g34130));
  NOT NOT1_1050(.VSS(VSS),.VDD(VDD),.Y(I17633),.A(g13258));
  NOT NOT1_1051(.VSS(VSS),.VDD(VDD),.Y(g32660),.A(g30825));
  NOT NOT1_1052(.VSS(VSS),.VDD(VDD),.Y(g7418),.A(g2361));
  NOT NOT1_1053(.VSS(VSS),.VDD(VDD),.Y(I13726),.A(g4537));
  NOT NOT1_1054(.VSS(VSS),.VDD(VDD),.Y(g9003),.A(g790));
  NOT NOT1_1055(.VSS(VSS),.VDD(VDD),.Y(g6953),.A(g4157));
  NOT NOT1_1056(.VSS(VSS),.VDD(VDD),.Y(g7994),.A(I12336));
  NOT NOT1_1057(.VSS(VSS),.VDD(VDD),.Y(g29997),.A(g29060));
  NOT NOT1_1058(.VSS(VSS),.VDD(VDD),.Y(g11884),.A(g8125));
  NOT NOT1_1059(.VSS(VSS),.VDD(VDD),.Y(g21467),.A(g15758));
  NOT NOT1_1060(.VSS(VSS),.VDD(VDD),.Y(I16676),.A(g10588));
  NOT NOT1_1061(.VSS(VSS),.VDD(VDD),.Y(g25869),.A(g25250));
  NOT NOT1_1062(.VSS(VSS),.VDD(VDD),.Y(g10349),.A(g6956));
  NOT NOT1_1063(.VSS(VSS),.VDD(VDD),.Y(g23494),.A(I22619));
  NOT NOT1_1064(.VSS(VSS),.VDD(VDD),.Y(g26337),.A(g24818));
  NOT NOT1_1065(.VSS(VSS),.VDD(VDD),.Y(I32806),.A(g34585));
  NOT NOT1_1066(.VSS(VSS),.VDD(VDD),.Y(g8796),.A(g4785));
  NOT NOT1_1067(.VSS(VSS),.VDD(VDD),.Y(I32684),.A(g34430));
  NOT NOT1_1068(.VSS(VSS),.VDD(VDD),.Y(g32456),.A(g31376));
  NOT NOT1_1069(.VSS(VSS),.VDD(VDD),.Y(g34244),.A(I32231));
  NOT NOT1_1070(.VSS(VSS),.VDD(VDD),.Y(I33300),.A(g35001));
  NOT NOT1_1071(.VSS(VSS),.VDD(VDD),.Y(g20130),.A(g17328));
  NOT NOT1_1072(.VSS(VSS),.VDD(VDD),.Y(g22683),.A(I22000));
  NOT NOT1_1073(.VSS(VSS),.VDD(VDD),.Y(g13410),.A(I15921));
  NOT NOT1_1074(.VSS(VSS),.VDD(VDD),.Y(I12826),.A(g4349));
  NOT NOT1_1075(.VSS(VSS),.VDD(VDD),.Y(g21037),.A(I20913));
  NOT NOT1_1076(.VSS(VSS),.VDD(VDD),.Y(g24130),.A(g20998));
  NOT NOT1_1077(.VSS(VSS),.VDD(VDD),.Y(g32480),.A(g31070));
  NOT NOT1_1078(.VSS(VSS),.VDD(VDD),.Y(g10083),.A(g2407));
  NOT NOT1_1079(.VSS(VSS),.VDD(VDD),.Y(g10348),.A(I13762));
  NOT NOT1_1080(.VSS(VSS),.VDD(VDD),.Y(g32916),.A(g31021));
  NOT NOT1_1081(.VSS(VSS),.VDD(VDD),.Y(g14348),.A(g10887));
  NOT NOT1_1082(.VSS(VSS),.VDD(VDD),.Y(g12891),.A(g10399));
  NOT NOT1_1083(.VSS(VSS),.VDD(VDD),.Y(g8324),.A(g2476));
  NOT NOT1_1084(.VSS(VSS),.VDD(VDD),.Y(g26792),.A(g25439));
  NOT NOT1_1085(.VSS(VSS),.VDD(VDD),.Y(g20523),.A(g17821));
  NOT NOT1_1086(.VSS(VSS),.VDD(VDD),.Y(I16417),.A(g875));
  NOT NOT1_1087(.VSS(VSS),.VDD(VDD),.Y(I21013),.A(g15806));
  NOT NOT1_1088(.VSS(VSS),.VDD(VDD),.Y(g32550),.A(g31376));
  NOT NOT1_1089(.VSS(VSS),.VDD(VDD),.Y(g9637),.A(I13252));
  NOT NOT1_1090(.VSS(VSS),.VDD(VDD),.Y(g23984),.A(g19210));
  NOT NOT1_1091(.VSS(VSS),.VDD(VDD),.Y(g18952),.A(g16053));
  NOT NOT1_1092(.VSS(VSS),.VDD(VDD),.Y(g24165),.A(I23339));
  NOT NOT1_1093(.VSS(VSS),.VDD(VDD),.Y(g30068),.A(g29157));
  NOT NOT1_1094(.VSS(VSS),.VDD(VDD),.Y(g34810),.A(I33020));
  NOT NOT1_1095(.VSS(VSS),.VDD(VDD),.Y(g31227),.A(g29744));
  NOT NOT1_1096(.VSS(VSS),.VDD(VDD),.Y(g17683),.A(g15027));
  NOT NOT1_1097(.VSS(VSS),.VDD(VDD),.Y(g23419),.A(g21468));
  NOT NOT1_1098(.VSS(VSS),.VDD(VDD),.Y(g34068),.A(g33728));
  NOT NOT1_1099(.VSS(VSS),.VDD(VDD),.Y(g21352),.A(g16322));
  NOT NOT1_1100(.VSS(VSS),.VDD(VDD),.Y(g13015),.A(g11875));
  NOT NOT1_1101(.VSS(VSS),.VDD(VDD),.Y(g8540),.A(g3408));
  NOT NOT1_1102(.VSS(VSS),.VDD(VDD),.Y(g23352),.A(g20924));
  NOT NOT1_1103(.VSS(VSS),.VDD(VDD),.Y(g25259),.A(I24445));
  NOT NOT1_1104(.VSS(VSS),.VDD(VDD),.Y(g25225),.A(g23802));
  NOT NOT1_1105(.VSS(VSS),.VDD(VDD),.Y(g21155),.A(g15656));
  NOT NOT1_1106(.VSS(VSS),.VDD(VDD),.Y(g34879),.A(I33109));
  NOT NOT1_1107(.VSS(VSS),.VDD(VDD),.Y(g21418),.A(g17821));
  NOT NOT1_1108(.VSS(VSS),.VDD(VDD),.Y(g22882),.A(g20391));
  NOT NOT1_1109(.VSS(VSS),.VDD(VDD),.Y(g28608),.A(g27670));
  NOT NOT1_1110(.VSS(VSS),.VDD(VDD),.Y(g23418),.A(g21468));
  NOT NOT1_1111(.VSS(VSS),.VDD(VDD),.Y(g32721),.A(g31021));
  NOT NOT1_1112(.VSS(VSS),.VDD(VDD),.Y(g20006),.A(g17328));
  NOT NOT1_1113(.VSS(VSS),.VDD(VDD),.Y(I26466),.A(g26870));
  NOT NOT1_1114(.VSS(VSS),.VDD(VDD),.Y(I15556),.A(g11928));
  NOT NOT1_1115(.VSS(VSS),.VDD(VDD),.Y(g32596),.A(g31070));
  NOT NOT1_1116(.VSS(VSS),.VDD(VDD),.Y(g9223),.A(g1216));
  NOT NOT1_1117(.VSS(VSS),.VDD(VDD),.Y(g12109),.A(I14967));
  NOT NOT1_1118(.VSS(VSS),.VDD(VDD),.Y(g19433),.A(g15915));
  NOT NOT1_1119(.VSS(VSS),.VDD(VDD),.Y(g23170),.A(g20046));
  NOT NOT1_1120(.VSS(VSS),.VDD(VDD),.Y(g7197),.A(g812));
  NOT NOT1_1121(.VSS(VSS),.VDD(VDD),.Y(g22407),.A(g19455));
  NOT NOT1_1122(.VSS(VSS),.VDD(VDD),.Y(g34878),.A(I33106));
  NOT NOT1_1123(.VSS(VSS),.VDD(VDD),.Y(g19387),.A(g16431));
  NOT NOT1_1124(.VSS(VSS),.VDD(VDD),.Y(I16762),.A(g5290));
  NOT NOT1_1125(.VSS(VSS),.VDD(VDD),.Y(g6848),.A(g2417));
  NOT NOT1_1126(.VSS(VSS),.VDD(VDD),.Y(g7397),.A(g890));
  NOT NOT1_1127(.VSS(VSS),.VDD(VDD),.Y(I27449),.A(g27737));
  NOT NOT1_1128(.VSS(VSS),.VDD(VDD),.Y(g15969),.A(I17416));
  NOT NOT1_1129(.VSS(VSS),.VDD(VDD),.Y(I20846),.A(g16923));
  NOT NOT1_1130(.VSS(VSS),.VDD(VDD),.Y(g19620),.A(g17296));
  NOT NOT1_1131(.VSS(VSS),.VDD(VDD),.Y(g12108),.A(I14964));
  NOT NOT1_1132(.VSS(VSS),.VDD(VDD),.Y(g10139),.A(g136));
  NOT NOT1_1133(.VSS(VSS),.VDD(VDD),.Y(I15223),.A(g10119));
  NOT NOT1_1134(.VSS(VSS),.VDD(VDD),.Y(I17612),.A(g13250));
  NOT NOT1_1135(.VSS(VSS),.VDD(VDD),.Y(I24396),.A(g23453));
  NOT NOT1_1136(.VSS(VSS),.VDD(VDD),.Y(g6855),.A(g2711));
  NOT NOT1_1137(.VSS(VSS),.VDD(VDD),.Y(g17414),.A(g14627));
  NOT NOT1_1138(.VSS(VSS),.VDD(VDD),.Y(g27492),.A(g26598));
  NOT NOT1_1139(.VSS(VSS),.VDD(VDD),.Y(g8287),.A(g160));
  NOT NOT1_1140(.VSS(VSS),.VDD(VDD),.Y(I17324),.A(g14119));
  NOT NOT1_1141(.VSS(VSS),.VDD(VDD),.Y(g9416),.A(g2429));
  NOT NOT1_1142(.VSS(VSS),.VDD(VDD),.Y(g13223),.A(I15800));
  NOT NOT1_1143(.VSS(VSS),.VDD(VDD),.Y(g24437),.A(g22654));
  NOT NOT1_1144(.VSS(VSS),.VDD(VDD),.Y(g25244),.A(g23802));
  NOT NOT1_1145(.VSS(VSS),.VDD(VDD),.Y(g19343),.A(g16136));
  NOT NOT1_1146(.VSS(VSS),.VDD(VDD),.Y(g34994),.A(I33282));
  NOT NOT1_1147(.VSS(VSS),.VDD(VDD),.Y(I17098),.A(g14336));
  NOT NOT1_1148(.VSS(VSS),.VDD(VDD),.Y(g32773),.A(g31376));
  NOT NOT1_1149(.VSS(VSS),.VDD(VDD),.Y(g32942),.A(g30825));
  NOT NOT1_1150(.VSS(VSS),.VDD(VDD),.Y(g9251),.A(I13037));
  NOT NOT1_1151(.VSS(VSS),.VDD(VDD),.Y(g20703),.A(g15373));
  NOT NOT1_1152(.VSS(VSS),.VDD(VDD),.Y(g29220),.A(I27576));
  NOT NOT1_1153(.VSS(VSS),.VDD(VDD),.Y(I11635),.A(g9));
  NOT NOT1_1154(.VSS(VSS),.VDD(VDD),.Y(g23589),.A(g21468));
  NOT NOT1_1155(.VSS(VSS),.VDD(VDD),.Y(g10415),.A(g7109));
  NOT NOT1_1156(.VSS(VSS),.VDD(VDD),.Y(g18422),.A(I19238));
  NOT NOT1_1157(.VSS(VSS),.VDD(VDD),.Y(g32655),.A(g30614));
  NOT NOT1_1158(.VSS(VSS),.VDD(VDD),.Y(g8399),.A(g3798));
  NOT NOT1_1159(.VSS(VSS),.VDD(VDD),.Y(g11110),.A(g8728));
  NOT NOT1_1160(.VSS(VSS),.VDD(VDD),.Y(g29911),.A(g28780));
  NOT NOT1_1161(.VSS(VSS),.VDD(VDD),.Y(g19369),.A(g15995));
  NOT NOT1_1162(.VSS(VSS),.VDD(VDD),.Y(g33377),.A(I30901));
  NOT NOT1_1163(.VSS(VSS),.VDD(VDD),.Y(g34425),.A(I32446));
  NOT NOT1_1164(.VSS(VSS),.VDD(VDD),.Y(g12381),.A(I15223));
  NOT NOT1_1165(.VSS(VSS),.VDD(VDD),.Y(g23524),.A(g21562));
  NOT NOT1_1166(.VSS(VSS),.VDD(VDD),.Y(g27091),.A(g26725));
  NOT NOT1_1167(.VSS(VSS),.VDD(VDD),.Y(g28184),.A(I26705));
  NOT NOT1_1168(.VSS(VSS),.VDD(VDD),.Y(g32670),.A(g30673));
  NOT NOT1_1169(.VSS(VSS),.VDD(VDD),.Y(g33120),.A(I30686));
  NOT NOT1_1170(.VSS(VSS),.VDD(VDD),.Y(I12026),.A(g344));
  NOT NOT1_1171(.VSS(VSS),.VDD(VDD),.Y(I21100),.A(g16284));
  NOT NOT1_1172(.VSS(VSS),.VDD(VDD),.Y(g8898),.A(g676));
  NOT NOT1_1173(.VSS(VSS),.VDD(VDD),.Y(g20600),.A(g15348));
  NOT NOT1_1174(.VSS(VSS),.VDD(VDD),.Y(I16117),.A(g10430));
  NOT NOT1_1175(.VSS(VSS),.VDD(VDD),.Y(g34919),.A(I33149));
  NOT NOT1_1176(.VSS(VSS),.VDD(VDD),.Y(g19368),.A(g16326));
  NOT NOT1_1177(.VSS(VSS),.VDD(VDD),.Y(I32222),.A(g34118));
  NOT NOT1_1178(.VSS(VSS),.VDD(VDD),.Y(g20781),.A(I20840));
  NOT NOT1_1179(.VSS(VSS),.VDD(VDD),.Y(g16877),.A(I18071));
  NOT NOT1_1180(.VSS(VSS),.VDD(VDD),.Y(g23477),.A(g21468));
  NOT NOT1_1181(.VSS(VSS),.VDD(VDD),.Y(g32734),.A(g31710));
  NOT NOT1_1182(.VSS(VSS),.VDD(VDD),.Y(g33645),.A(I31477));
  NOT NOT1_1183(.VSS(VSS),.VDD(VDD),.Y(g22759),.A(g19857));
  NOT NOT1_1184(.VSS(VSS),.VDD(VDD),.Y(I17140),.A(g13835));
  NOT NOT1_1185(.VSS(VSS),.VDD(VDD),.Y(g26817),.A(g25242));
  NOT NOT1_1186(.VSS(VSS),.VDD(VDD),.Y(g7631),.A(g74));
  NOT NOT1_1187(.VSS(VSS),.VDD(VDD),.Y(g34918),.A(I33146));
  NOT NOT1_1188(.VSS(VSS),.VDD(VDD),.Y(g17584),.A(g14773));
  NOT NOT1_1189(.VSS(VSS),.VDD(VDD),.Y(I26693),.A(g27930));
  NOT NOT1_1190(.VSS(VSS),.VDD(VDD),.Y(g10664),.A(g8928));
  NOT NOT1_1191(.VSS(VSS),.VDD(VDD),.Y(I20929),.A(g17663));
  NOT NOT1_1192(.VSS(VSS),.VDD(VDD),.Y(g32839),.A(g30735));
  NOT NOT1_1193(.VSS(VSS),.VDD(VDD),.Y(g32930),.A(g31021));
  NOT NOT1_1194(.VSS(VSS),.VDD(VDD),.Y(g20372),.A(g17847));
  NOT NOT1_1195(.VSS(VSS),.VDD(VDD),.Y(g30079),.A(g29097));
  NOT NOT1_1196(.VSS(VSS),.VDD(VDD),.Y(g19412),.A(g16489));
  NOT NOT1_1197(.VSS(VSS),.VDD(VDD),.Y(g7257),.A(I11903));
  NOT NOT1_1198(.VSS(VSS),.VDD(VDD),.Y(g22758),.A(g20330));
  NOT NOT1_1199(.VSS(VSS),.VDD(VDD),.Y(g24372),.A(g22885));
  NOT NOT1_1200(.VSS(VSS),.VDD(VDD),.Y(g16695),.A(g14454));
  NOT NOT1_1201(.VSS(VSS),.VDD(VDD),.Y(g25171),.A(g22228));
  NOT NOT1_1202(.VSS(VSS),.VDD(VDD),.Y(g20175),.A(I20433));
  NOT NOT1_1203(.VSS(VSS),.VDD(VDD),.Y(g7301),.A(g925));
  NOT NOT1_1204(.VSS(VSS),.VDD(VDD),.Y(I16747),.A(g12729));
  NOT NOT1_1205(.VSS(VSS),.VDD(VDD),.Y(g8291),.A(I12503));
  NOT NOT1_1206(.VSS(VSS),.VDD(VDD),.Y(g11373),.A(g7566));
  NOT NOT1_1207(.VSS(VSS),.VDD(VDD),.Y(g23864),.A(g19210));
  NOT NOT1_1208(.VSS(VSS),.VDD(VDD),.Y(g25886),.A(g24537));
  NOT NOT1_1209(.VSS(VSS),.VDD(VDD),.Y(g23022),.A(g20283));
  NOT NOT1_1210(.VSS(VSS),.VDD(VDD),.Y(g32667),.A(g30825));
  NOT NOT1_1211(.VSS(VSS),.VDD(VDD),.Y(g32694),.A(g31376));
  NOT NOT1_1212(.VSS(VSS),.VDD(VDD),.Y(g32838),.A(g31376));
  NOT NOT1_1213(.VSS(VSS),.VDD(VDD),.Y(I31550),.A(g33204));
  NOT NOT1_1214(.VSS(VSS),.VDD(VDD),.Y(g33698),.A(I31539));
  NOT NOT1_1215(.VSS(VSS),.VDD(VDD),.Y(g24175),.A(I23369));
  NOT NOT1_1216(.VSS(VSS),.VDD(VDD),.Y(g29147),.A(I27449));
  NOT NOT1_1217(.VSS(VSS),.VDD(VDD),.Y(g32965),.A(g31710));
  NOT NOT1_1218(.VSS(VSS),.VDD(VDD),.Y(g12840),.A(g10356));
  NOT NOT1_1219(.VSS(VSS),.VDD(VDD),.Y(g6818),.A(g976));
  NOT NOT1_1220(.VSS(VSS),.VDD(VDD),.Y(g17759),.A(g14864));
  NOT NOT1_1221(.VSS(VSS),.VDD(VDD),.Y(g6867),.A(I11685));
  NOT NOT1_1222(.VSS(VSS),.VDD(VDD),.Y(g16526),.A(g13898));
  NOT NOT1_1223(.VSS(VSS),.VDD(VDD),.Y(g23749),.A(g18997));
  NOT NOT1_1224(.VSS(VSS),.VDD(VDD),.Y(I15800),.A(g11607));
  NOT NOT1_1225(.VSS(VSS),.VDD(VDD),.Y(g15714),.A(I17228));
  NOT NOT1_1226(.VSS(VSS),.VDD(VDD),.Y(g9880),.A(g5787));
  NOT NOT1_1227(.VSS(VSS),.VDD(VDD),.Y(g23313),.A(g21070));
  NOT NOT1_1228(.VSS(VSS),.VDD(VDD),.Y(g25994),.A(g24575));
  NOT NOT1_1229(.VSS(VSS),.VDD(VDD),.Y(g8344),.A(I12523));
  NOT NOT1_1230(.VSS(VSS),.VDD(VDD),.Y(g9537),.A(g1748));
  NOT NOT1_1231(.VSS(VSS),.VDD(VDD),.Y(g29950),.A(g28896));
  NOT NOT1_1232(.VSS(VSS),.VDD(VDD),.Y(g24063),.A(g20014));
  NOT NOT1_1233(.VSS(VSS),.VDD(VDD),.Y(g17758),.A(g14861));
  NOT NOT1_1234(.VSS(VSS),.VDD(VDD),.Y(g26656),.A(g25495));
  NOT NOT1_1235(.VSS(VSS),.VDD(VDD),.Y(g20516),.A(I20609));
  NOT NOT1_1236(.VSS(VSS),.VDD(VDD),.Y(g10554),.A(g8974));
  NOT NOT1_1237(.VSS(VSS),.VDD(VDD),.Y(g18905),.A(g16077));
  NOT NOT1_1238(.VSS(VSS),.VDD(VDD),.Y(g24137),.A(g20998));
  NOT NOT1_1239(.VSS(VSS),.VDD(VDD),.Y(g32487),.A(g30825));
  NOT NOT1_1240(.VSS(VSS),.VDD(VDD),.Y(g24516),.A(g22670));
  NOT NOT1_1241(.VSS(VSS),.VDD(VDD),.Y(g7751),.A(g1521));
  NOT NOT1_1242(.VSS(VSS),.VDD(VDD),.Y(g23285),.A(g20887));
  NOT NOT1_1243(.VSS(VSS),.VDD(VDD),.Y(g26680),.A(g25300));
  NOT NOT1_1244(.VSS(VSS),.VDD(VDD),.Y(g32619),.A(g30614));
  NOT NOT1_1245(.VSS(VSS),.VDD(VDD),.Y(g8259),.A(g2217));
  NOT NOT1_1246(.VSS(VSS),.VDD(VDD),.Y(g21305),.A(g15758));
  NOT NOT1_1247(.VSS(VSS),.VDD(VDD),.Y(g21053),.A(g15373));
  NOT NOT1_1248(.VSS(VSS),.VDD(VDD),.Y(g32502),.A(g31070));
  NOT NOT1_1249(.VSS(VSS),.VDD(VDD),.Y(g14609),.A(I16724));
  NOT NOT1_1250(.VSS(VSS),.VDD(VDD),.Y(g15979),.A(I17420));
  NOT NOT1_1251(.VSS(VSS),.VDD(VDD),.Y(g10200),.A(g2138));
  NOT NOT1_1252(.VSS(VSS),.VDD(VDD),.Y(g23305),.A(g20391));
  NOT NOT1_1253(.VSS(VSS),.VDD(VDD),.Y(g32557),.A(g31376));
  NOT NOT1_1254(.VSS(VSS),.VDD(VDD),.Y(g13334),.A(g11048));
  NOT NOT1_1255(.VSS(VSS),.VDD(VDD),.Y(g29151),.A(g27858));
  NOT NOT1_1256(.VSS(VSS),.VDD(VDD),.Y(g29172),.A(g27020));
  NOT NOT1_1257(.VSS(VSS),.VDD(VDD),.Y(I24787),.A(g24266));
  NOT NOT1_1258(.VSS(VSS),.VDD(VDD),.Y(g9978),.A(g2756));
  NOT NOT1_1259(.VSS(VSS),.VDD(VDD),.Y(g30322),.A(g28431));
  NOT NOT1_1260(.VSS(VSS),.VDD(VDD),.Y(g10608),.A(g9155));
  NOT NOT1_1261(.VSS(VSS),.VDD(VDD),.Y(g29996),.A(g28962));
  NOT NOT1_1262(.VSS(VSS),.VDD(VDD),.Y(I12811),.A(g4340));
  NOT NOT1_1263(.VSS(VSS),.VDD(VDD),.Y(g10115),.A(g2283));
  NOT NOT1_1264(.VSS(VSS),.VDD(VDD),.Y(I16639),.A(g4000));
  NOT NOT1_1265(.VSS(VSS),.VDD(VDD),.Y(g21466),.A(g15509));
  NOT NOT1_1266(.VSS(VSS),.VDD(VDD),.Y(g32618),.A(g31154));
  NOT NOT1_1267(.VSS(VSS),.VDD(VDD),.Y(I18662),.A(g6322));
  NOT NOT1_1268(.VSS(VSS),.VDD(VDD),.Y(g8088),.A(g1554));
  NOT NOT1_1269(.VSS(VSS),.VDD(VDD),.Y(g6975),.A(g4507));
  NOT NOT1_1270(.VSS(VSS),.VDD(VDD),.Y(g9417),.A(I13124));
  NOT NOT1_1271(.VSS(VSS),.VDD(VDD),.Y(g34159),.A(I32116));
  NOT NOT1_1272(.VSS(VSS),.VDD(VDD),.Y(g11762),.A(g7964));
  NOT NOT1_1273(.VSS(VSS),.VDD(VDD),.Y(g7041),.A(g5644));
  NOT NOT1_1274(.VSS(VSS),.VDD(VDD),.Y(g9935),.A(I13483));
  NOT NOT1_1275(.VSS(VSS),.VDD(VDD),.Y(I13606),.A(g74));
  NOT NOT1_1276(.VSS(VSS),.VDD(VDD),.Y(g11964),.A(g9154));
  NOT NOT1_1277(.VSS(VSS),.VDD(VDD),.Y(g21036),.A(I20910));
  NOT NOT1_1278(.VSS(VSS),.VDD(VDD),.Y(g7441),.A(g862));
  NOT NOT1_1279(.VSS(VSS),.VDD(VDD),.Y(g20209),.A(g17821));
  NOT NOT1_1280(.VSS(VSS),.VDD(VDD),.Y(g33661),.A(I31497));
  NOT NOT1_1281(.VSS(VSS),.VDD(VDD),.Y(g33895),.A(I31751));
  NOT NOT1_1282(.VSS(VSS),.VDD(VDD),.Y(g9982),.A(g3976));
  NOT NOT1_1283(.VSS(VSS),.VDD(VDD),.Y(g21177),.A(I20957));
  NOT NOT1_1284(.VSS(VSS),.VDD(VDD),.Y(g21560),.A(g17873));
  NOT NOT1_1285(.VSS(VSS),.VDD(VDD),.Y(g16077),.A(I17456));
  NOT NOT1_1286(.VSS(VSS),.VDD(VDD),.Y(g9234),.A(g5170));
  NOT NOT1_1287(.VSS(VSS),.VDD(VDD),.Y(I15587),.A(g11985));
  NOT NOT1_1288(.VSS(VSS),.VDD(VDD),.Y(g32469),.A(g30673));
  NOT NOT1_1289(.VSS(VSS),.VDD(VDD),.Y(I27368),.A(g27881));
  NOT NOT1_1290(.VSS(VSS),.VDD(VDD),.Y(I18482),.A(g13350));
  NOT NOT1_1291(.VSS(VSS),.VDD(VDD),.Y(g20208),.A(g17533));
  NOT NOT1_1292(.VSS(VSS),.VDD(VDD),.Y(g14745),.A(g12423));
  NOT NOT1_1293(.VSS(VSS),.VDD(VDD),.Y(g13216),.A(g10939));
  NOT NOT1_1294(.VSS(VSS),.VDD(VDD),.Y(g17141),.A(I18191));
  NOT NOT1_1295(.VSS(VSS),.VDD(VDD),.Y(I11750),.A(g4474));
  NOT NOT1_1296(.VSS(VSS),.VDD(VDD),.Y(I18248),.A(g12938));
  NOT NOT1_1297(.VSS(VSS),.VDD(VDD),.Y(g19379),.A(g17327));
  NOT NOT1_1298(.VSS(VSS),.VDD(VDD),.Y(g26631),.A(g25467));
  NOT NOT1_1299(.VSS(VSS),.VDD(VDD),.Y(g12862),.A(g10370));
  NOT NOT1_1300(.VSS(VSS),.VDD(VDD),.Y(g17652),.A(g15033));
  NOT NOT1_1301(.VSS(VSS),.VDD(VDD),.Y(g34656),.A(I32770));
  NOT NOT1_1302(.VSS(VSS),.VDD(VDD),.Y(g8215),.A(I12451));
  NOT NOT1_1303(.VSS(VSS),.VDD(VDD),.Y(g30295),.A(I28540));
  NOT NOT1_1304(.VSS(VSS),.VDD(VDD),.Y(g22332),.A(I21838));
  NOT NOT1_1305(.VSS(VSS),.VDD(VDD),.Y(g9542),.A(g2173));
  NOT NOT1_1306(.VSS(VSS),.VDD(VDD),.Y(I16391),.A(g859));
  NOT NOT1_1307(.VSS(VSS),.VDD(VDD),.Y(g26364),.A(I25327));
  NOT NOT1_1308(.VSS(VSS),.VDD(VDD),.Y(g32468),.A(g30614));
  NOT NOT1_1309(.VSS(VSS),.VDD(VDD),.Y(g6821),.A(I11655));
  NOT NOT1_1310(.VSS(VSS),.VDD(VDD),.Y(I18003),.A(g13638));
  NOT NOT1_1311(.VSS(VSS),.VDD(VDD),.Y(g19050),.A(I19759));
  NOT NOT1_1312(.VSS(VSS),.VDD(VDD),.Y(g34680),.A(I32820));
  NOT NOT1_1313(.VSS(VSS),.VDD(VDD),.Y(g8951),.A(g554));
  NOT NOT1_1314(.VSS(VSS),.VDD(VDD),.Y(g16689),.A(g13923));
  NOT NOT1_1315(.VSS(VSS),.VDD(VDD),.Y(g34144),.A(I32093));
  NOT NOT1_1316(.VSS(VSS),.VDD(VDD),.Y(g34823),.A(I33037));
  NOT NOT1_1317(.VSS(VSS),.VDD(VDD),.Y(g20542),.A(g17873));
  NOT NOT1_1318(.VSS(VSS),.VDD(VDD),.Y(g16923),.A(I18089));
  NOT NOT1_1319(.VSS(VSS),.VDD(VDD),.Y(g20453),.A(I20584));
  NOT NOT1_1320(.VSS(VSS),.VDD(VDD),.Y(g16280),.A(g13330));
  NOT NOT1_1321(.VSS(VSS),.VDD(VDD),.Y(g6984),.A(g4709));
  NOT NOT1_1322(.VSS(VSS),.VDD(VDD),.Y(g32038),.A(g30934));
  NOT NOT1_1323(.VSS(VSS),.VDD(VDD),.Y(g24021),.A(g20841));
  NOT NOT1_1324(.VSS(VSS),.VDD(VDD),.Y(g28241),.A(g27064));
  NOT NOT1_1325(.VSS(VSS),.VDD(VDD),.Y(g29318),.A(g29029));
  NOT NOT1_1326(.VSS(VSS),.VDD(VDD),.Y(g16688),.A(g14045));
  NOT NOT1_1327(.VSS(VSS),.VDD(VDD),.Y(g16624),.A(I17814));
  NOT NOT1_1328(.VSS(VSS),.VDD(VDD),.Y(g22406),.A(g19506));
  NOT NOT1_1329(.VSS(VSS),.VDD(VDD),.Y(g8114),.A(g3522));
  NOT NOT1_1330(.VSS(VSS),.VDD(VDD),.Y(g10184),.A(g4486));
  NOT NOT1_1331(.VSS(VSS),.VDD(VDD),.Y(g12040),.A(I14902));
  NOT NOT1_1332(.VSS(VSS),.VDD(VDD),.Y(I16579),.A(g10981));
  NOT NOT1_1333(.VSS(VSS),.VDD(VDD),.Y(g16300),.A(I17626));
  NOT NOT1_1334(.VSS(VSS),.VDD(VDD),.Y(g19386),.A(g16431));
  NOT NOT1_1335(.VSS(VSS),.VDD(VDD),.Y(g10805),.A(I14046));
  NOT NOT1_1336(.VSS(VSS),.VDD(VDD),.Y(I22785),.A(g18940));
  NOT NOT1_1337(.VSS(VSS),.VDD(VDD),.Y(g20913),.A(g15373));
  NOT NOT1_1338(.VSS(VSS),.VDD(VDD),.Y(I18778),.A(g6704));
  NOT NOT1_1339(.VSS(VSS),.VDD(VDD),.Y(g34336),.A(g34112));
  NOT NOT1_1340(.VSS(VSS),.VDD(VDD),.Y(g32815),.A(g30937));
  NOT NOT1_1341(.VSS(VSS),.VDD(VDD),.Y(g14184),.A(g12381));
  NOT NOT1_1342(.VSS(VSS),.VDD(VDD),.Y(g19603),.A(g16349));
  NOT NOT1_1343(.VSS(VSS),.VDD(VDD),.Y(g19742),.A(g17096));
  NOT NOT1_1344(.VSS(VSS),.VDD(VDD),.Y(g13117),.A(g10981));
  NOT NOT1_1345(.VSS(VSS),.VDD(VDD),.Y(g17135),.A(g14297));
  NOT NOT1_1346(.VSS(VSS),.VDD(VDD),.Y(g12904),.A(g10410));
  NOT NOT1_1347(.VSS(VSS),.VDD(VDD),.Y(g20614),.A(g15426));
  NOT NOT1_1348(.VSS(VSS),.VDD(VDD),.Y(g32601),.A(g31376));
  NOT NOT1_1349(.VSS(VSS),.VDD(VDD),.Y(I15569),.A(g11965));
  NOT NOT1_1350(.VSS(VSS),.VDD(VDD),.Y(g9554),.A(g5105));
  NOT NOT1_1351(.VSS(VSS),.VDD(VDD),.Y(g20436),.A(I20569));
  NOT NOT1_1352(.VSS(VSS),.VDD(VDD),.Y(g23874),.A(g18997));
  NOT NOT1_1353(.VSS(VSS),.VDD(VDD),.Y(g8870),.A(I12837));
  NOT NOT1_1354(.VSS(VSS),.VDD(VDD),.Y(g32677),.A(g30673));
  NOT NOT1_1355(.VSS(VSS),.VDD(VDD),.Y(g33127),.A(g31950));
  NOT NOT1_1356(.VSS(VSS),.VDD(VDD),.Y(g25322),.A(I24497));
  NOT NOT1_1357(.VSS(VSS),.VDD(VDD),.Y(I31694),.A(g33176));
  NOT NOT1_1358(.VSS(VSS),.VDD(VDD),.Y(I32834),.A(g34472));
  NOT NOT1_1359(.VSS(VSS),.VDD(VDD),.Y(g32975),.A(I30537));
  NOT NOT1_1360(.VSS(VSS),.VDD(VDD),.Y(g21693),.A(I21254));
  NOT NOT1_1361(.VSS(VSS),.VDD(VDD),.Y(g20607),.A(g17955));
  NOT NOT1_1362(.VSS(VSS),.VDD(VDD),.Y(g13569),.A(g10951));
  NOT NOT1_1363(.VSS(VSS),.VDD(VDD),.Y(g8650),.A(g4664));
  NOT NOT1_1364(.VSS(VSS),.VDD(VDD),.Y(I12896),.A(g4229));
  NOT NOT1_1365(.VSS(VSS),.VDD(VDD),.Y(g20320),.A(g17015));
  NOT NOT1_1366(.VSS(VSS),.VDD(VDD),.Y(I18647),.A(g5320));
  NOT NOT1_1367(.VSS(VSS),.VDD(VDD),.Y(g20073),.A(g16540));
  NOT NOT1_1368(.VSS(VSS),.VDD(VDD),.Y(I28832),.A(g30301));
  NOT NOT1_1369(.VSS(VSS),.VDD(VDD),.Y(I33131),.A(g34906));
  NOT NOT1_1370(.VSS(VSS),.VDD(VDD),.Y(g30017),.A(g29085));
  NOT NOT1_1371(.VSS(VSS),.VDD(VDD),.Y(g20274),.A(g17847));
  NOT NOT1_1372(.VSS(VSS),.VDD(VDD),.Y(g9213),.A(I13020));
  NOT NOT1_1373(.VSS(VSS),.VDD(VDD),.Y(g24073),.A(g21127));
  NOT NOT1_1374(.VSS(VSS),.VDD(VDD),.Y(g20530),.A(g15509));
  NOT NOT1_1375(.VSS(VSS),.VDD(VDD),.Y(g21665),.A(I21226));
  NOT NOT1_1376(.VSS(VSS),.VDD(VDD),.Y(g25158),.A(g22228));
  NOT NOT1_1377(.VSS(VSS),.VDD(VDD),.Y(I21744),.A(g19338));
  NOT NOT1_1378(.VSS(VSS),.VDD(VDD),.Y(g20593),.A(g15277));
  NOT NOT1_1379(.VSS(VSS),.VDD(VDD),.Y(I17754),.A(g13494));
  NOT NOT1_1380(.VSS(VSS),.VDD(VDD),.Y(g23665),.A(g21562));
  NOT NOT1_1381(.VSS(VSS),.VDD(VDD),.Y(g25783),.A(g25250));
  NOT NOT1_1382(.VSS(VSS),.VDD(VDD),.Y(I17355),.A(g14591));
  NOT NOT1_1383(.VSS(VSS),.VDD(VDD),.Y(g32937),.A(g31021));
  NOT NOT1_1384(.VSS(VSS),.VDD(VDD),.Y(g19429),.A(g16489));
  NOT NOT1_1385(.VSS(VSS),.VDD(VDD),.Y(I23345),.A(g23320));
  NOT NOT1_1386(.VSS(VSS),.VDD(VDD),.Y(g33385),.A(g32038));
  NOT NOT1_1387(.VSS(VSS),.VDD(VDD),.Y(I21849),.A(g19620));
  NOT NOT1_1388(.VSS(VSS),.VDD(VDD),.Y(g29044),.A(g27742));
  NOT NOT1_1389(.VSS(VSS),.VDD(VDD),.Y(g10761),.A(g8411));
  NOT NOT1_1390(.VSS(VSS),.VDD(VDD),.Y(g7411),.A(g2040));
  NOT NOT1_1391(.VSS(VSS),.VDD(VDD),.Y(g25561),.A(g22550));
  NOT NOT1_1392(.VSS(VSS),.VDD(VDD),.Y(g18891),.A(g16053));
  NOT NOT1_1393(.VSS(VSS),.VDD(VDD),.Y(g20565),.A(g18008));
  NOT NOT1_1394(.VSS(VSS),.VDD(VDD),.Y(I31619),.A(g33212));
  NOT NOT1_1395(.VSS(VSS),.VDD(VDD),.Y(I15814),.A(g11129));
  NOT NOT1_1396(.VSS(VSS),.VDD(VDD),.Y(g24122),.A(g20857));
  NOT NOT1_1397(.VSS(VSS),.VDD(VDD),.Y(I23399),.A(g23450));
  NOT NOT1_1398(.VSS(VSS),.VDD(VDD),.Y(g8136),.A(g269));
  NOT NOT1_1399(.VSS(VSS),.VDD(VDD),.Y(g19730),.A(g17062));
  NOT NOT1_1400(.VSS(VSS),.VDD(VDD),.Y(g19428),.A(g16090));
  NOT NOT1_1401(.VSS(VSS),.VDD(VDD),.Y(g12183),.A(I15033));
  NOT NOT1_1402(.VSS(VSS),.VDD(VDD),.Y(g9902),.A(g100));
  NOT NOT1_1403(.VSS(VSS),.VDD(VDD),.Y(I18233),.A(g14639));
  NOT NOT1_1404(.VSS(VSS),.VDD(VDD),.Y(g33354),.A(g32329));
  NOT NOT1_1405(.VSS(VSS),.VDD(VDD),.Y(I33210),.A(g34943));
  NOT NOT1_1406(.VSS(VSS),.VDD(VDD),.Y(g32791),.A(g31672));
  NOT NOT1_1407(.VSS(VSS),.VDD(VDD),.Y(g23476),.A(g21468));
  NOT NOT1_1408(.VSS(VSS),.VDD(VDD),.Y(g23485),.A(g20785));
  NOT NOT1_1409(.VSS(VSS),.VDD(VDD),.Y(I25555),.A(g25241));
  NOT NOT1_1410(.VSS(VSS),.VDD(VDD),.Y(g31824),.A(g29385));
  NOT NOT1_1411(.VSS(VSS),.VDD(VDD),.Y(g32884),.A(g30825));
  NOT NOT1_1412(.VSS(VSS),.VDD(VDD),.Y(g33888),.A(g33346));
  NOT NOT1_1413(.VSS(VSS),.VDD(VDD),.Y(g8594),.A(g3849));
  NOT NOT1_1414(.VSS(VSS),.VDD(VDD),.Y(g19765),.A(g16897));
  NOT NOT1_1415(.VSS(VSS),.VDD(VDD),.Y(g6756),.A(I11623));
  NOT NOT1_1416(.VSS(VSS),.VDD(VDD),.Y(g24034),.A(g19968));
  NOT NOT1_1417(.VSS(VSS),.VDD(VDD),.Y(g7074),.A(I11801));
  NOT NOT1_1418(.VSS(VSS),.VDD(VDD),.Y(g11772),.A(I14623));
  NOT NOT1_1419(.VSS(VSS),.VDD(VDD),.Y(g10400),.A(g7002));
  NOT NOT1_1420(.VSS(VSS),.VDD(VDD),.Y(g20641),.A(g15509));
  NOT NOT1_1421(.VSS(VSS),.VDD(VDD),.Y(g26816),.A(g25260));
  NOT NOT1_1422(.VSS(VSS),.VDD(VDD),.Y(g21454),.A(g15373));
  NOT NOT1_1423(.VSS(VSS),.VDD(VDD),.Y(I33279),.A(g34986));
  NOT NOT1_1424(.VSS(VSS),.VDD(VDD),.Y(g23555),.A(I22692));
  NOT NOT1_1425(.VSS(VSS),.VDD(VDD),.Y(I32607),.A(g34358));
  NOT NOT1_1426(.VSS(VSS),.VDD(VDD),.Y(g7474),.A(I11980));
  NOT NOT1_1427(.VSS(VSS),.VDD(VDD),.Y(g17221),.A(I18245));
  NOT NOT1_1428(.VSS(VSS),.VDD(VDD),.Y(g19690),.A(g16826));
  NOT NOT1_1429(.VSS(VSS),.VDD(VDD),.Y(g30309),.A(g28959));
  NOT NOT1_1430(.VSS(VSS),.VDD(VDD),.Y(g7992),.A(g5008));
  NOT NOT1_1431(.VSS(VSS),.VDD(VDD),.Y(g9490),.A(g2563));
  NOT NOT1_1432(.VSS(VSS),.VDD(VDD),.Y(I14563),.A(g802));
  NOT NOT1_1433(.VSS(VSS),.VDD(VDD),.Y(g16511),.A(g14130));
  NOT NOT1_1434(.VSS(VSS),.VDD(VDD),.Y(g9166),.A(g837));
  NOT NOT1_1435(.VSS(VSS),.VDD(VDD),.Y(g20153),.A(g16782));
  NOT NOT1_1436(.VSS(VSS),.VDD(VDD),.Y(g23570),.A(g18833));
  NOT NOT1_1437(.VSS(VSS),.VDD(VDD),.Y(I32274),.A(g34195));
  NOT NOT1_1438(.VSS(VSS),.VDD(VDD),.Y(g23914),.A(g19210));
  NOT NOT1_1439(.VSS(VSS),.VDD(VDD),.Y(g32479),.A(g30735));
  NOT NOT1_1440(.VSS(VSS),.VDD(VDD),.Y(g32666),.A(g31376));
  NOT NOT1_1441(.VSS(VSS),.VDD(VDD),.Y(I13483),.A(g6035));
  NOT NOT1_1442(.VSS(VSS),.VDD(VDD),.Y(g11293),.A(g7527));
  NOT NOT1_1443(.VSS(VSS),.VDD(VDD),.Y(g24153),.A(I23303));
  NOT NOT1_1444(.VSS(VSS),.VDD(VDD),.Y(I31469),.A(g33388));
  NOT NOT1_1445(.VSS(VSS),.VDD(VDD),.Y(g6904),.A(g3494));
  NOT NOT1_1446(.VSS(VSS),.VDD(VDD),.Y(g32363),.A(I29891));
  NOT NOT1_1447(.VSS(VSS),.VDD(VDD),.Y(I12112),.A(g794));
  NOT NOT1_1448(.VSS(VSS),.VDD(VDD),.Y(g12872),.A(g10379));
  NOT NOT1_1449(.VSS(VSS),.VDD(VDD),.Y(g13638),.A(I16057));
  NOT NOT1_1450(.VSS(VSS),.VDD(VDD),.Y(g34308),.A(g34088));
  NOT NOT1_1451(.VSS(VSS),.VDD(VDD),.Y(g9056),.A(g3017));
  NOT NOT1_1452(.VSS(VSS),.VDD(VDD),.Y(g23907),.A(g19074));
  NOT NOT1_1453(.VSS(VSS),.VDD(VDD),.Y(g32478),.A(g31376));
  NOT NOT1_1454(.VSS(VSS),.VDD(VDD),.Y(g32015),.A(I29571));
  NOT NOT1_1455(.VSS(VSS),.VDD(VDD),.Y(g19504),.A(g16349));
  NOT NOT1_1456(.VSS(VSS),.VDD(VDD),.Y(g9456),.A(g6073));
  NOT NOT1_1457(.VSS(VSS),.VDD(VDD),.Y(g33931),.A(I31807));
  NOT NOT1_1458(.VSS(VSS),.VDD(VDD),.Y(I32464),.A(g34245));
  NOT NOT1_1459(.VSS(VSS),.VDD(VDD),.Y(g8228),.A(g3835));
  NOT NOT1_1460(.VSS(VSS),.VDD(VDD),.Y(g9529),.A(g6561));
  NOT NOT1_1461(.VSS(VSS),.VDD(VDD),.Y(g7863),.A(g1249));
  NOT NOT1_1462(.VSS(VSS),.VDD(VDD),.Y(g20136),.A(I20399));
  NOT NOT1_1463(.VSS(VSS),.VDD(VDD),.Y(g20635),.A(g18008));
  NOT NOT1_1464(.VSS(VSS),.VDD(VDD),.Y(I27742),.A(g28819));
  NOT NOT1_1465(.VSS(VSS),.VDD(VDD),.Y(g13416),.A(I15929));
  NOT NOT1_1466(.VSS(VSS),.VDD(VDD),.Y(g25017),.A(g23699));
  NOT NOT1_1467(.VSS(VSS),.VDD(VDD),.Y(I25567),.A(g25272));
  NOT NOT1_1468(.VSS(VSS),.VDD(VDD),.Y(I25594),.A(g25531));
  NOT NOT1_1469(.VSS(VSS),.VDD(VDD),.Y(I18897),.A(g16738));
  NOT NOT1_1470(.VSS(VSS),.VDD(VDD),.Y(g24136),.A(g20857));
  NOT NOT1_1471(.VSS(VSS),.VDD(VDD),.Y(g32486),.A(g30735));
  NOT NOT1_1472(.VSS(VSS),.VDD(VDD),.Y(I13326),.A(g66));
  NOT NOT1_1473(.VSS(VSS),.VDD(VDD),.Y(g23239),.A(g21308));
  NOT NOT1_1474(.VSS(VSS),.VDD(VDD),.Y(g33426),.A(g32017));
  NOT NOT1_1475(.VSS(VSS),.VDD(VDD),.Y(g11841),.A(g9800));
  NOT NOT1_1476(.VSS(VSS),.VDD(VDD),.Y(g9155),.A(I12997));
  NOT NOT1_1477(.VSS(VSS),.VDD(VDD),.Y(I14395),.A(g3654));
  NOT NOT1_1478(.VSS(VSS),.VDD(VDD),.Y(g6841),.A(g2145));
  NOT NOT1_1479(.VSS(VSS),.VDD(VDD),.Y(I17420),.A(g13394));
  NOT NOT1_1480(.VSS(VSS),.VDD(VDD),.Y(g23567),.A(g21562));
  NOT NOT1_1481(.VSS(VSS),.VDD(VDD),.Y(g32556),.A(g31554));
  NOT NOT1_1482(.VSS(VSS),.VDD(VDD),.Y(I32797),.A(g34581));
  NOT NOT1_1483(.VSS(VSS),.VDD(VDD),.Y(I14899),.A(g10198));
  NOT NOT1_1484(.VSS(VSS),.VDD(VDD),.Y(g8033),.A(g157));
  NOT NOT1_1485(.VSS(VSS),.VDD(VDD),.Y(g23238),.A(g20924));
  NOT NOT1_1486(.VSS(VSS),.VDD(VDD),.Y(g11510),.A(g7633));
  NOT NOT1_1487(.VSS(VSS),.VDD(VDD),.Y(g13510),.A(I15981));
  NOT NOT1_1488(.VSS(VSS),.VDD(VDD),.Y(g17812),.A(I18810));
  NOT NOT1_1489(.VSS(VSS),.VDD(VDD),.Y(g34816),.A(I33030));
  NOT NOT1_1490(.VSS(VSS),.VDD(VDD),.Y(I20647),.A(g17010));
  NOT NOT1_1491(.VSS(VSS),.VDD(VDD),.Y(g32580),.A(g30825));
  NOT NOT1_1492(.VSS(VSS),.VDD(VDD),.Y(g9698),.A(g2181));
  NOT NOT1_1493(.VSS(VSS),.VDD(VDD),.Y(g28441),.A(g27629));
  NOT NOT1_1494(.VSS(VSS),.VDD(VDD),.Y(g26260),.A(g24759));
  NOT NOT1_1495(.VSS(VSS),.VDD(VDD),.Y(I14633),.A(g9340));
  NOT NOT1_1496(.VSS(VSS),.VDD(VDD),.Y(g9964),.A(g126));
  NOT NOT1_1497(.VSS(VSS),.VDD(VDD),.Y(I13252),.A(g6751));
  NOT NOT1_1498(.VSS(VSS),.VDD(VDD),.Y(g20164),.A(g16826));
  NOT NOT1_1499(.VSS(VSS),.VDD(VDD),.Y(g34985),.A(I33255));
  NOT NOT1_1500(.VSS(VSS),.VDD(VDD),.Y(I20999),.A(g16709));
  NOT NOT1_1501(.VSS(VSS),.VDD(VDD),.Y(g23941),.A(g19074));
  NOT NOT1_1502(.VSS(VSS),.VDD(VDD),.Y(g18091),.A(I18879));
  NOT NOT1_1503(.VSS(VSS),.VDD(VDD),.Y(g19128),.A(I19778));
  NOT NOT1_1504(.VSS(VSS),.VDD(VDD),.Y(g23382),.A(g20682));
  NOT NOT1_1505(.VSS(VSS),.VDD(VDD),.Y(g24164),.A(I23336));
  NOT NOT1_1506(.VSS(VSS),.VDD(VDD),.Y(g25289),.A(g22228));
  NOT NOT1_1507(.VSS(VSS),.VDD(VDD),.Y(g21176),.A(I20954));
  NOT NOT1_1508(.VSS(VSS),.VDD(VDD),.Y(g21185),.A(g15277));
  NOT NOT1_1509(.VSS(VSS),.VDD(VDD),.Y(g23519),.A(g21468));
  NOT NOT1_1510(.VSS(VSS),.VDD(VDD),.Y(I27730),.A(g28752));
  NOT NOT1_1511(.VSS(VSS),.VDD(VDD),.Y(g12047),.A(g9591));
  NOT NOT1_1512(.VSS(VSS),.VDD(VDD),.Y(g16307),.A(I17633));
  NOT NOT1_1513(.VSS(VSS),.VDD(VDD),.Y(g13835),.A(I16150));
  NOT NOT1_1514(.VSS(VSS),.VDD(VDD),.Y(g34954),.A(I33210));
  NOT NOT1_1515(.VSS(VSS),.VDD(VDD),.Y(g13014),.A(g11872));
  NOT NOT1_1516(.VSS(VSS),.VDD(VDD),.Y(g25023),.A(g22457));
  NOT NOT1_1517(.VSS(VSS),.VDD(VDD),.Y(g24891),.A(g23231));
  NOT NOT1_1518(.VSS(VSS),.VDD(VDD),.Y(I33143),.A(g34903));
  NOT NOT1_1519(.VSS(VSS),.VDD(VDD),.Y(g19626),.A(g17409));
  NOT NOT1_1520(.VSS(VSS),.VDD(VDD),.Y(g25288),.A(g22228));
  NOT NOT1_1521(.VSS(VSS),.VDD(VDD),.Y(g25224),.A(g22763));
  NOT NOT1_1522(.VSS(VSS),.VDD(VDD),.Y(I20233),.A(g17487));
  NOT NOT1_1523(.VSS(VSS),.VDD(VDD),.Y(g16721),.A(g14072));
  NOT NOT1_1524(.VSS(VSS),.VDD(VDD),.Y(I12793),.A(g4578));
  NOT NOT1_1525(.VSS(VSS),.VDD(VDD),.Y(g23518),.A(g21070));
  NOT NOT1_1526(.VSS(VSS),.VDD(VDD),.Y(g23154),.A(I22264));
  NOT NOT1_1527(.VSS(VSS),.VDD(VDD),.Y(g26488),.A(I25366));
  NOT NOT1_1528(.VSS(VSS),.VDD(VDD),.Y(g26424),.A(I25356));
  NOT NOT1_1529(.VSS(VSS),.VDD(VDD),.Y(g20575),.A(g17929));
  NOT NOT1_1530(.VSS(VSS),.VDD(VDD),.Y(g31860),.A(I29438));
  NOT NOT1_1531(.VSS(VSS),.VDD(VDD),.Y(g13007),.A(g11852));
  NOT NOT1_1532(.VSS(VSS),.VDD(VDD),.Y(g25308),.A(g22763));
  NOT NOT1_1533(.VSS(VSS),.VDD(VDD),.Y(g8195),.A(g1783));
  NOT NOT1_1534(.VSS(VSS),.VDD(VDD),.Y(g8137),.A(g411));
  NOT NOT1_1535(.VSS(VSS),.VDD(VDD),.Y(g32922),.A(g31710));
  NOT NOT1_1536(.VSS(VSS),.VDD(VDD),.Y(g8891),.A(g582));
  NOT NOT1_1537(.VSS(VSS),.VDD(VDD),.Y(g19533),.A(g16261));
  NOT NOT1_1538(.VSS(VSS),.VDD(VDD),.Y(g24474),.A(g23620));
  NOT NOT1_1539(.VSS(VSS),.VDD(VDD),.Y(g20711),.A(g15509));
  NOT NOT1_1540(.VSS(VSS),.VDD(VDD),.Y(I16193),.A(g3281));
  NOT NOT1_1541(.VSS(VSS),.VDD(VDD),.Y(g16431),.A(I17675));
  NOT NOT1_1542(.VSS(VSS),.VDD(VDD),.Y(I27549),.A(g28161));
  NOT NOT1_1543(.VSS(VSS),.VDD(VDD),.Y(g27051),.A(I25779));
  NOT NOT1_1544(.VSS(VSS),.VDD(VDD),.Y(g32531),.A(g31070));
  NOT NOT1_1545(.VSS(VSS),.VDD(VDD),.Y(I13847),.A(g7266));
  NOT NOT1_1546(.VSS(VSS),.VDD(VDD),.Y(I31791),.A(g33354));
  NOT NOT1_1547(.VSS(VSS),.VDD(VDD),.Y(g20327),.A(g15224));
  NOT NOT1_1548(.VSS(VSS),.VDD(VDD),.Y(g23935),.A(g19210));
  NOT NOT1_1549(.VSS(VSS),.VDD(VDD),.Y(g24711),.A(g23139));
  NOT NOT1_1550(.VSS(VSS),.VDD(VDD),.Y(g34669),.A(I32791));
  NOT NOT1_1551(.VSS(VSS),.VDD(VDD),.Y(g26830),.A(g24411));
  NOT NOT1_1552(.VSS(VSS),.VDD(VDD),.Y(g27592),.A(g26715));
  NOT NOT1_1553(.VSS(VSS),.VDD(VDD),.Y(g12051),.A(g9595));
  NOT NOT1_1554(.VSS(VSS),.VDD(VDD),.Y(g20537),.A(g15345));
  NOT NOT1_1555(.VSS(VSS),.VDD(VDD),.Y(g24109),.A(g21143));
  NOT NOT1_1556(.VSS(VSS),.VDD(VDD),.Y(g32740),.A(g31672));
  NOT NOT1_1557(.VSS(VSS),.VDD(VDD),.Y(g15885),.A(I17374));
  NOT NOT1_1558(.VSS(VSS),.VDD(VDD),.Y(g8807),.A(g79));
  NOT NOT1_1559(.VSS(VSS),.VDD(VDD),.Y(g11615),.A(g6875));
  NOT NOT1_1560(.VSS(VSS),.VDD(VDD),.Y(g9619),.A(g5845));
  NOT NOT1_1561(.VSS(VSS),.VDD(VDD),.Y(g17507),.A(g15030));
  NOT NOT1_1562(.VSS(VSS),.VDD(VDD),.Y(I24331),.A(g22976));
  NOT NOT1_1563(.VSS(VSS),.VDD(VDD),.Y(g34668),.A(I32788));
  NOT NOT1_1564(.VSS(VSS),.VDD(VDD),.Y(g13116),.A(g10935));
  NOT NOT1_1565(.VSS(VSS),.VDD(VDD),.Y(g16773),.A(g14021));
  NOT NOT1_1566(.VSS(VSS),.VDD(VDD),.Y(I18148),.A(g13526));
  NOT NOT1_1567(.VSS(VSS),.VDD(VDD),.Y(g24108),.A(g20998));
  NOT NOT1_1568(.VSS(VSS),.VDD(VDD),.Y(I28162),.A(g28803));
  NOT NOT1_1569(.VSS(VSS),.VDD(VDD),.Y(g32186),.A(I29720));
  NOT NOT1_1570(.VSS(VSS),.VDD(VDD),.Y(g34392),.A(g34202));
  NOT NOT1_1571(.VSS(VSS),.VDD(VDD),.Y(g32676),.A(g30614));
  NOT NOT1_1572(.VSS(VSS),.VDD(VDD),.Y(g32685),.A(g31528));
  NOT NOT1_1573(.VSS(VSS),.VDD(VDD),.Y(g33659),.A(I31491));
  NOT NOT1_1574(.VSS(VSS),.VDD(VDD),.Y(g28399),.A(g27074));
  NOT NOT1_1575(.VSS(VSS),.VDD(VDD),.Y(g30195),.A(I28434));
  NOT NOT1_1576(.VSS(VSS),.VDD(VDD),.Y(g7400),.A(g911));
  NOT NOT1_1577(.VSS(VSS),.VDD(VDD),.Y(g8859),.A(g772));
  NOT NOT1_1578(.VSS(VSS),.VDD(VDD),.Y(g32953),.A(g31327));
  NOT NOT1_1579(.VSS(VSS),.VDD(VDD),.Y(g19737),.A(g17015));
  NOT NOT1_1580(.VSS(VSS),.VDD(VDD),.Y(g11720),.A(I14589));
  NOT NOT1_1581(.VSS(VSS),.VDD(VDD),.Y(g20283),.A(I20529));
  NOT NOT1_1582(.VSS(VSS),.VDD(VDD),.Y(g6811),.A(g714));
  NOT NOT1_1583(.VSS(VSS),.VDD(VDD),.Y(g34195),.A(I32150));
  NOT NOT1_1584(.VSS(VSS),.VDD(VDD),.Y(g20606),.A(g17955));
  NOT NOT1_1585(.VSS(VSS),.VDD(VDD),.Y(g33250),.A(g32186));
  NOT NOT1_1586(.VSS(VSS),.VDD(VDD),.Y(g16655),.A(g14151));
  NOT NOT1_1587(.VSS(VSS),.VDD(VDD),.Y(g10882),.A(g7601));
  NOT NOT1_1588(.VSS(VSS),.VDD(VDD),.Y(I18104),.A(g13177));
  NOT NOT1_1589(.VSS(VSS),.VDD(VDD),.Y(g10414),.A(g7092));
  NOT NOT1_1590(.VSS(VSS),.VDD(VDD),.Y(I13634),.A(g79));
  NOT NOT1_1591(.VSS(VSS),.VDD(VDD),.Y(g31658),.A(I29242));
  NOT NOT1_1592(.VSS(VSS),.VDD(VDD),.Y(I13872),.A(g7474));
  NOT NOT1_1593(.VSS(VSS),.VDD(VDD),.Y(g13041),.A(I15667));
  NOT NOT1_1594(.VSS(VSS),.VDD(VDD),.Y(g32654),.A(g31070));
  NOT NOT1_1595(.VSS(VSS),.VDD(VDD),.Y(g9843),.A(g4311));
  NOT NOT1_1596(.VSS(VSS),.VDD(VDD),.Y(g33658),.A(g33080));
  NOT NOT1_1597(.VSS(VSS),.VDD(VDD),.Y(g16180),.A(g13437));
  NOT NOT1_1598(.VSS(VSS),.VDD(VDD),.Y(g30016),.A(g29049));
  NOT NOT1_1599(.VSS(VSS),.VDD(VDD),.Y(g9989),.A(g5077));
  NOT NOT1_1600(.VSS(VSS),.VDD(VDD),.Y(I24448),.A(g22923));
  NOT NOT1_1601(.VSS(VSS),.VDD(VDD),.Y(g11430),.A(g7617));
  NOT NOT1_1602(.VSS(VSS),.VDD(VDD),.Y(g22541),.A(I21911));
  NOT NOT1_1603(.VSS(VSS),.VDD(VDD),.Y(g34559),.A(g34384));
  NOT NOT1_1604(.VSS(VSS),.VDD(VDD),.Y(g12350),.A(I15190));
  NOT NOT1_1605(.VSS(VSS),.VDD(VDD),.Y(g10407),.A(g7063));
  NOT NOT1_1606(.VSS(VSS),.VDD(VDD),.Y(g32800),.A(g31021));
  NOT NOT1_1607(.VSS(VSS),.VDD(VDD),.Y(g32936),.A(g31710));
  NOT NOT1_1608(.VSS(VSS),.VDD(VDD),.Y(g19697),.A(g16886));
  NOT NOT1_1609(.VSS(VSS),.VDD(VDD),.Y(I31486),.A(g33197));
  NOT NOT1_1610(.VSS(VSS),.VDD(VDD),.Y(g23215),.A(g20785));
  NOT NOT1_1611(.VSS(VSS),.VDD(VDD),.Y(g12820),.A(g10233));
  NOT NOT1_1612(.VSS(VSS),.VDD(VDD),.Y(I17699),.A(g13416));
  NOT NOT1_1613(.VSS(VSS),.VDD(VDD),.Y(g23501),.A(g20924));
  NOT NOT1_1614(.VSS(VSS),.VDD(VDD),.Y(g6874),.A(g3143));
  NOT NOT1_1615(.VSS(VSS),.VDD(VDD),.Y(I29965),.A(g31189));
  NOT NOT1_1616(.VSS(VSS),.VDD(VDD),.Y(I32109),.A(g33631));
  NOT NOT1_1617(.VSS(VSS),.VDD(VDD),.Y(I21033),.A(g17221));
  NOT NOT1_1618(.VSS(VSS),.VDD(VDD),.Y(g20381),.A(g17955));
  NOT NOT1_1619(.VSS(VSS),.VDD(VDD),.Y(g8342),.A(I12519));
  NOT NOT1_1620(.VSS(VSS),.VDD(VDD),.Y(g11237),.A(I14305));
  NOT NOT1_1621(.VSS(VSS),.VDD(VDD),.Y(g9834),.A(g2579));
  NOT NOT1_1622(.VSS(VSS),.VDD(VDD),.Y(g9971),.A(g2093));
  NOT NOT1_1623(.VSS(VSS),.VDD(VDD),.Y(I21234),.A(g16540));
  NOT NOT1_1624(.VSS(VSS),.VDD(VDD),.Y(g24982),.A(g22763));
  NOT NOT1_1625(.VSS(VSS),.VDD(VDD),.Y(g26679),.A(g25385));
  NOT NOT1_1626(.VSS(VSS),.VDD(VDD),.Y(g34830),.A(I33044));
  NOT NOT1_1627(.VSS(VSS),.VDD(VDD),.Y(g34893),.A(I33119));
  NOT NOT1_1628(.VSS(VSS),.VDD(VDD),.Y(g9686),.A(g73));
  NOT NOT1_1629(.VSS(VSS),.VDD(VDD),.Y(g22359),.A(g19495));
  NOT NOT1_1630(.VSS(VSS),.VDD(VDD),.Y(g8255),.A(g2028));
  NOT NOT1_1631(.VSS(VSS),.VDD(VDD),.Y(g17473),.A(g14841));
  NOT NOT1_1632(.VSS(VSS),.VDD(VDD),.Y(g20091),.A(g17328));
  NOT NOT1_1633(.VSS(VSS),.VDD(VDD),.Y(I22366),.A(g19757));
  NOT NOT1_1634(.VSS(VSS),.VDD(VDD),.Y(g24091),.A(g20720));
  NOT NOT1_1635(.VSS(VSS),.VDD(VDD),.Y(g7183),.A(g4608));
  NOT NOT1_1636(.VSS(VSS),.VDD(VDD),.Y(g8481),.A(I12618));
  NOT NOT1_1637(.VSS(VSS),.VDD(VDD),.Y(I12128),.A(g4253));
  NOT NOT1_1638(.VSS(VSS),.VDD(VDD),.Y(g17789),.A(g14321));
  NOT NOT1_1639(.VSS(VSS),.VDD(VDD),.Y(g29956),.A(I28185));
  NOT NOT1_1640(.VSS(VSS),.VDD(VDD),.Y(g29385),.A(g28180));
  NOT NOT1_1641(.VSS(VSS),.VDD(VDD),.Y(g34544),.A(I32613));
  NOT NOT1_1642(.VSS(VSS),.VDD(VDD),.Y(g15480),.A(I17125));
  NOT NOT1_1643(.VSS(VSS),.VDD(VDD),.Y(I26664),.A(g27708));
  NOT NOT1_1644(.VSS(VSS),.VDD(VDD),.Y(g22358),.A(g19801));
  NOT NOT1_1645(.VSS(VSS),.VDD(VDD),.Y(g32762),.A(g31672));
  NOT NOT1_1646(.VSS(VSS),.VDD(VDD),.Y(g9598),.A(g2571));
  NOT NOT1_1647(.VSS(VSS),.VDD(VDD),.Y(g24174),.A(I23366));
  NOT NOT1_1648(.VSS(VSS),.VDD(VDD),.Y(g8097),.A(g3029));
  NOT NOT1_1649(.VSS(VSS),.VDD(VDD),.Y(g25260),.A(I24448));
  NOT NOT1_1650(.VSS(VSS),.VDD(VDD),.Y(g32964),.A(g31672));
  NOT NOT1_1651(.VSS(VSS),.VDD(VDD),.Y(g29980),.A(g28935));
  NOT NOT1_1652(.VSS(VSS),.VDD(VDD),.Y(g7779),.A(g1413));
  NOT NOT1_1653(.VSS(VSS),.VDD(VDD),.Y(g34713),.A(I32871));
  NOT NOT1_1654(.VSS(VSS),.VDD(VDD),.Y(g8497),.A(g3436));
  NOT NOT1_1655(.VSS(VSS),.VDD(VDD),.Y(g13142),.A(g10632));
  NOT NOT1_1656(.VSS(VSS),.VDD(VDD),.Y(g21349),.A(g15758));
  NOT NOT1_1657(.VSS(VSS),.VDD(VDD),.Y(g8154),.A(g3139));
  NOT NOT1_1658(.VSS(VSS),.VDD(VDD),.Y(I28591),.A(g29371));
  NOT NOT1_1659(.VSS(VSS),.VDD(VDD),.Y(g17325),.A(I18304));
  NOT NOT1_1660(.VSS(VSS),.VDD(VDD),.Y(g8354),.A(g4815));
  NOT NOT1_1661(.VSS(VSS),.VDD(VDD),.Y(g18948),.A(g15800));
  NOT NOT1_1662(.VSS(VSS),.VDD(VDD),.Y(g7023),.A(g5445));
  NOT NOT1_1663(.VSS(VSS),.VDD(VDD),.Y(g31855),.A(g29385));
  NOT NOT1_1664(.VSS(VSS),.VDD(VDD),.Y(g10206),.A(g4489));
  NOT NOT1_1665(.VSS(VSS),.VDD(VDD),.Y(g14441),.A(I16590));
  NOT NOT1_1666(.VSS(VSS),.VDD(VDD),.Y(g14584),.A(g11048));
  NOT NOT1_1667(.VSS(VSS),.VDD(VDD),.Y(g9321),.A(g5863));
  NOT NOT1_1668(.VSS(VSS),.VDD(VDD),.Y(g7423),.A(g2433));
  NOT NOT1_1669(.VSS(VSS),.VDD(VDD),.Y(g9670),.A(g5022));
  NOT NOT1_1670(.VSS(VSS),.VDD(VDD),.Y(I22547),.A(g20720));
  NOT NOT1_1671(.VSS(VSS),.VDD(VDD),.Y(g25195),.A(g22763));
  NOT NOT1_1672(.VSS(VSS),.VDD(VDD),.Y(g16487),.A(I17695));
  NOT NOT1_1673(.VSS(VSS),.VDD(VDD),.Y(g23906),.A(g19074));
  NOT NOT1_1674(.VSS(VSS),.VDD(VDD),.Y(g26093),.A(g24814));
  NOT NOT1_1675(.VSS(VSS),.VDD(VDD),.Y(g30610),.A(I28872));
  NOT NOT1_1676(.VSS(VSS),.VDD(VDD),.Y(g18904),.A(g16053));
  NOT NOT1_1677(.VSS(VSS),.VDD(VDD),.Y(g32587),.A(g30735));
  NOT NOT1_1678(.VSS(VSS),.VDD(VDD),.Y(g15085),.A(I17008));
  NOT NOT1_1679(.VSS(VSS),.VDD(VDD),.Y(I32982),.A(g34749));
  NOT NOT1_1680(.VSS(VSS),.VDD(VDD),.Y(g23284),.A(g20785));
  NOT NOT1_1681(.VSS(VSS),.VDD(VDD),.Y(g19445),.A(g15915));
  NOT NOT1_1682(.VSS(VSS),.VDD(VDD),.Y(g10725),.A(g7846));
  NOT NOT1_1683(.VSS(VSS),.VDD(VDD),.Y(g21304),.A(g17367));
  NOT NOT1_1684(.VSS(VSS),.VDD(VDD),.Y(g25525),.A(g22550));
  NOT NOT1_1685(.VSS(VSS),.VDD(VDD),.Y(g34042),.A(g33674));
  NOT NOT1_1686(.VSS(VSS),.VDD(VDD),.Y(g25424),.A(g23800));
  NOT NOT1_1687(.VSS(VSS),.VDD(VDD),.Y(I20433),.A(g16234));
  NOT NOT1_1688(.VSS(VSS),.VDD(VDD),.Y(g23304),.A(g20785));
  NOT NOT1_1689(.VSS(VSS),.VDD(VDD),.Y(g25016),.A(g23666));
  NOT NOT1_1690(.VSS(VSS),.VDD(VDD),.Y(g6978),.A(g4616));
  NOT NOT1_1691(.VSS(VSS),.VDD(VDD),.Y(I33179),.A(g34893));
  NOT NOT1_1692(.VSS(VSS),.VDD(VDD),.Y(g7161),.A(I11843));
  NOT NOT1_1693(.VSS(VSS),.VDD(VDD),.Y(g19499),.A(g16782));
  NOT NOT1_1694(.VSS(VSS),.VDD(VDD),.Y(g17121),.A(g14321));
  NOT NOT1_1695(.VSS(VSS),.VDD(VDD),.Y(g7361),.A(g1874));
  NOT NOT1_1696(.VSS(VSS),.VDD(VDD),.Y(g22682),.A(g19379));
  NOT NOT1_1697(.VSS(VSS),.VDD(VDD),.Y(g10114),.A(g2116));
  NOT NOT1_1698(.VSS(VSS),.VDD(VDD),.Y(g20192),.A(g17268));
  NOT NOT1_1699(.VSS(VSS),.VDD(VDD),.Y(g9253),.A(g5037));
  NOT NOT1_1700(.VSS(VSS),.VDD(VDD),.Y(I16821),.A(g5983));
  NOT NOT1_1701(.VSS(VSS),.VDD(VDD),.Y(I17661),.A(g13329));
  NOT NOT1_1702(.VSS(VSS),.VDD(VDD),.Y(g27929),.A(I26448));
  NOT NOT1_1703(.VSS(VSS),.VDD(VDD),.Y(g25558),.A(g22594));
  NOT NOT1_1704(.VSS(VSS),.VDD(VDD),.Y(g23566),.A(g21562));
  NOT NOT1_1705(.VSS(VSS),.VDD(VDD),.Y(g32909),.A(g30614));
  NOT NOT1_1706(.VSS(VSS),.VDD(VDD),.Y(g10082),.A(g2375));
  NOT NOT1_1707(.VSS(VSS),.VDD(VDD),.Y(g32543),.A(g31376));
  NOT NOT1_1708(.VSS(VSS),.VDD(VDD),.Y(g34270),.A(g34159));
  NOT NOT1_1709(.VSS(VSS),.VDD(VDD),.Y(I27232),.A(g27993));
  NOT NOT1_1710(.VSS(VSS),.VDD(VDD),.Y(g19498),.A(g16752));
  NOT NOT1_1711(.VSS(VSS),.VDD(VDD),.Y(g34188),.A(g33875));
  NOT NOT1_1712(.VSS(VSS),.VDD(VDD),.Y(g7051),.A(I11793));
  NOT NOT1_1713(.VSS(VSS),.VDD(VDD),.Y(g10107),.A(I13606));
  NOT NOT1_1714(.VSS(VSS),.VDD(VDD),.Y(g22173),.A(I21757));
  NOT NOT1_1715(.VSS(VSS),.VDD(VDD),.Y(g34124),.A(g33819));
  NOT NOT1_1716(.VSS(VSS),.VDD(VDD),.Y(g9909),.A(g1978));
  NOT NOT1_1717(.VSS(VSS),.VDD(VDD),.Y(g12929),.A(g12550));
  NOT NOT1_1718(.VSS(VSS),.VDD(VDD),.Y(g25830),.A(g24485));
  NOT NOT1_1719(.VSS(VSS),.VDD(VDD),.Y(g27583),.A(g26686));
  NOT NOT1_1720(.VSS(VSS),.VDD(VDD),.Y(g20663),.A(g15373));
  NOT NOT1_1721(.VSS(VSS),.VDD(VDD),.Y(g27928),.A(g26810));
  NOT NOT1_1722(.VSS(VSS),.VDD(VDD),.Y(g25893),.A(g24541));
  NOT NOT1_1723(.VSS(VSS),.VDD(VDD),.Y(g8783),.A(I12761));
  NOT NOT1_1724(.VSS(VSS),.VDD(VDD),.Y(g7451),.A(g2070));
  NOT NOT1_1725(.VSS(VSS),.VDD(VDD),.Y(g32908),.A(g31327));
  NOT NOT1_1726(.VSS(VSS),.VDD(VDD),.Y(g6982),.A(g4531));
  NOT NOT1_1727(.VSS(VSS),.VDD(VDD),.Y(g7327),.A(g2165));
  NOT NOT1_1728(.VSS(VSS),.VDD(VDD),.Y(g24522),.A(g22689));
  NOT NOT1_1729(.VSS(VSS),.VDD(VDD),.Y(g33894),.A(I31748));
  NOT NOT1_1730(.VSS(VSS),.VDD(VDD),.Y(g11165),.A(I14222));
  NOT NOT1_1731(.VSS(VSS),.VDD(VDD),.Y(g8112),.A(g3419));
  NOT NOT1_1732(.VSS(VSS),.VDD(VDD),.Y(g8218),.A(g3490));
  NOT NOT1_1733(.VSS(VSS),.VDD(VDD),.Y(g34939),.A(g34922));
  NOT NOT1_1734(.VSS(VSS),.VDD(VDD),.Y(g9740),.A(g5821));
  NOT NOT1_1735(.VSS(VSS),.VDD(VDD),.Y(g8267),.A(g2342));
  NOT NOT1_1736(.VSS(VSS),.VDD(VDD),.Y(g25544),.A(g22594));
  NOT NOT1_1737(.VSS(VSS),.VDD(VDD),.Y(g32569),.A(g30673));
  NOT NOT1_1738(.VSS(VSS),.VDD(VDD),.Y(g34383),.A(I32388));
  NOT NOT1_1739(.VSS(VSS),.VDD(VDD),.Y(g29190),.A(g27046));
  NOT NOT1_1740(.VSS(VSS),.VDD(VDD),.Y(I32840),.A(g34480));
  NOT NOT1_1741(.VSS(VSS),.VDD(VDD),.Y(g17291),.A(I18276));
  NOT NOT1_1742(.VSS(VSS),.VDD(VDD),.Y(g14744),.A(g12578));
  NOT NOT1_1743(.VSS(VSS),.VDD(VDD),.Y(g16286),.A(I17615));
  NOT NOT1_1744(.VSS(VSS),.VDD(VDD),.Y(g21139),.A(g15634));
  NOT NOT1_1745(.VSS(VSS),.VDD(VDD),.Y(g21653),.A(g17663));
  NOT NOT1_1746(.VSS(VSS),.VDD(VDD),.Y(g26837),.A(g24869));
  NOT NOT1_1747(.VSS(VSS),.VDD(VDD),.Y(g7633),.A(I12120));
  NOT NOT1_1748(.VSS(VSS),.VDD(VDD),.Y(g34938),.A(g34920));
  NOT NOT1_1749(.VSS(VSS),.VDD(VDD),.Y(g23653),.A(I22788));
  NOT NOT1_1750(.VSS(VSS),.VDD(VDD),.Y(g9552),.A(g3654));
  NOT NOT1_1751(.VSS(VSS),.VDD(VDD),.Y(g15655),.A(g13202));
  NOT NOT1_1752(.VSS(VSS),.VDD(VDD),.Y(I31800),.A(g33164));
  NOT NOT1_1753(.VSS(VSS),.VDD(VDD),.Y(g10399),.A(g7017));
  NOT NOT1_1754(.VSS(VSS),.VDD(VDD),.Y(g32568),.A(g31170));
  NOT NOT1_1755(.VSS(VSS),.VDD(VDD),.Y(g32747),.A(g30825));
  NOT NOT1_1756(.VSS(VSS),.VDD(VDD),.Y(I18310),.A(g12978));
  NOT NOT1_1757(.VSS(VSS),.VDD(VDD),.Y(I20369),.A(g17690));
  NOT NOT1_1758(.VSS(VSS),.VDD(VDD),.Y(g18062),.A(I18872));
  NOT NOT1_1759(.VSS(VSS),.VDD(VDD),.Y(g21138),.A(g15634));
  NOT NOT1_1760(.VSS(VSS),.VDD(VDD),.Y(g24483),.A(I23688));
  NOT NOT1_1761(.VSS(VSS),.VDD(VDD),.Y(g19432),.A(g15885));
  NOT NOT1_1762(.VSS(VSS),.VDD(VDD),.Y(I19837),.A(g1399));
  NOT NOT1_1763(.VSS(VSS),.VDD(VDD),.Y(g30065),.A(g29049));
  NOT NOT1_1764(.VSS(VSS),.VDD(VDD),.Y(I11820),.A(g3869));
  NOT NOT1_1765(.VSS(VSS),.VDD(VDD),.Y(g23138),.A(g20453));
  NOT NOT1_1766(.VSS(VSS),.VDD(VDD),.Y(I26799),.A(g27660));
  NOT NOT1_1767(.VSS(VSS),.VDD(VDD),.Y(g20553),.A(g17929));
  NOT NOT1_1768(.VSS(VSS),.VDD(VDD),.Y(g31819),.A(g29385));
  NOT NOT1_1769(.VSS(VSS),.VDD(VDD),.Y(g8676),.A(g4821));
  NOT NOT1_1770(.VSS(VSS),.VDD(VDD),.Y(I15727),.A(g10981));
  NOT NOT1_1771(.VSS(VSS),.VDD(VDD),.Y(I32192),.A(g33628));
  NOT NOT1_1772(.VSS(VSS),.VDD(VDD),.Y(g10398),.A(g6999));
  NOT NOT1_1773(.VSS(VSS),.VDD(VDD),.Y(I18379),.A(g13012));
  NOT NOT1_1774(.VSS(VSS),.VDD(VDD),.Y(g14398),.A(I16555));
  NOT NOT1_1775(.VSS(VSS),.VDD(VDD),.Y(g10141),.A(I13634));
  NOT NOT1_1776(.VSS(VSS),.VDD(VDD),.Y(g29211),.A(I27549));
  NOT NOT1_1777(.VSS(VSS),.VDD(VDD),.Y(g10652),.A(g7601));
  NOT NOT1_1778(.VSS(VSS),.VDD(VDD),.Y(g10804),.A(g9772));
  NOT NOT1_1779(.VSS(VSS),.VDD(VDD),.Y(g6800),.A(g203));
  NOT NOT1_1780(.VSS(VSS),.VDD(VDD),.Y(I13152),.A(g6746));
  NOT NOT1_1781(.VSS(VSS),.VDD(VDD),.Y(g9687),.A(I13287));
  NOT NOT1_1782(.VSS(VSS),.VDD(VDD),.Y(g31818),.A(g29385));
  NOT NOT1_1783(.VSS(VSS),.VDD(VDD),.Y(g32814),.A(g31021));
  NOT NOT1_1784(.VSS(VSS),.VDD(VDD),.Y(g20326),.A(g18008));
  NOT NOT1_1785(.VSS(VSS),.VDD(VDD),.Y(g23333),.A(g20785));
  NOT NOT1_1786(.VSS(VSS),.VDD(VDD),.Y(g13222),.A(g10590));
  NOT NOT1_1787(.VSS(VSS),.VDD(VDD),.Y(g19753),.A(g16987));
  NOT NOT1_1788(.VSS(VSS),.VDD(VDD),.Y(g16601),.A(I17783));
  NOT NOT1_1789(.VSS(VSS),.VDD(VDD),.Y(g17760),.A(I18752));
  NOT NOT1_1790(.VSS(VSS),.VDD(VDD),.Y(g16677),.A(I17879));
  NOT NOT1_1791(.VSS(VSS),.VDD(VDD),.Y(I22889),.A(g18926));
  NOT NOT1_1792(.VSS(VSS),.VDD(VDD),.Y(g20536),.A(g18065));
  NOT NOT1_1793(.VSS(VSS),.VDD(VDD),.Y(g20040),.A(g17271));
  NOT NOT1_1794(.VSS(VSS),.VDD(VDD),.Y(g13437),.A(I15937));
  NOT NOT1_1795(.VSS(VSS),.VDD(VDD),.Y(I20412),.A(g16213));
  NOT NOT1_1796(.VSS(VSS),.VDD(VDD),.Y(g32751),.A(g31327));
  NOT NOT1_1797(.VSS(VSS),.VDD(VDD),.Y(g32807),.A(g31021));
  NOT NOT1_1798(.VSS(VSS),.VDD(VDD),.Y(g32772),.A(g31327));
  NOT NOT1_1799(.VSS(VSS),.VDD(VDD),.Y(g28463),.A(I26952));
  NOT NOT1_1800(.VSS(VSS),.VDD(VDD),.Y(g32974),.A(g30937));
  NOT NOT1_1801(.VSS(VSS),.VDD(VDD),.Y(g8830),.A(g767));
  NOT NOT1_1802(.VSS(VSS),.VDD(VDD),.Y(g24040),.A(g19919));
  NOT NOT1_1803(.VSS(VSS),.VDD(VDD),.Y(g7753),.A(I12183));
  NOT NOT1_1804(.VSS(VSS),.VDD(VDD),.Y(g20702),.A(g17955));
  NOT NOT1_1805(.VSS(VSS),.VDD(VDD),.Y(g30218),.A(g28918));
  NOT NOT1_1806(.VSS(VSS),.VDD(VDD),.Y(g25188),.A(g23909));
  NOT NOT1_1807(.VSS(VSS),.VDD(VDD),.Y(g32639),.A(g31070));
  NOT NOT1_1808(.VSS(VSS),.VDD(VDD),.Y(g20904),.A(g17433));
  NOT NOT1_1809(.VSS(VSS),.VDD(VDD),.Y(I17956),.A(g14562));
  NOT NOT1_1810(.VSS(VSS),.VDD(VDD),.Y(g23963),.A(g19147));
  NOT NOT1_1811(.VSS(VSS),.VDD(VDD),.Y(g19650),.A(g16971));
  NOT NOT1_1812(.VSS(VSS),.VDD(VDD),.Y(g28033),.A(g26365));
  NOT NOT1_1813(.VSS(VSS),.VDD(VDD),.Y(g8592),.A(g3805));
  NOT NOT1_1814(.VSS(VSS),.VDD(VDD),.Y(g7072),.A(g6199));
  NOT NOT1_1815(.VSS(VSS),.VDD(VDD),.Y(g14332),.A(I16492));
  NOT NOT1_1816(.VSS(VSS),.VDD(VDD),.Y(I11691),.A(g36));
  NOT NOT1_1817(.VSS(VSS),.VDD(VDD),.Y(I28540),.A(g28954));
  NOT NOT1_1818(.VSS(VSS),.VDD(VDD),.Y(g32638),.A(g30825));
  NOT NOT1_1819(.VSS(VSS),.VDD(VDD),.Y(g7472),.A(g6329));
  NOT NOT1_1820(.VSS(VSS),.VDD(VDD),.Y(g19529),.A(g16349));
  NOT NOT1_1821(.VSS(VSS),.VDD(VDD),.Y(g12640),.A(I15382));
  NOT NOT1_1822(.VSS(VSS),.VDD(VDD),.Y(I15600),.A(g10430));
  NOT NOT1_1823(.VSS(VSS),.VDD(VDD),.Y(g22927),.A(I22128));
  NOT NOT1_1824(.VSS(VSS),.VDD(VDD),.Y(g9860),.A(g5417));
  NOT NOT1_1825(.VSS(VSS),.VDD(VDD),.Y(g10406),.A(g7046));
  NOT NOT1_1826(.VSS(VSS),.VDD(VDD),.Y(I24228),.A(g22409));
  NOT NOT1_1827(.VSS(VSS),.VDD(VDD),.Y(g20564),.A(g15373));
  NOT NOT1_1828(.VSS(VSS),.VDD(VDD),.Y(g10361),.A(g6841));
  NOT NOT1_1829(.VSS(VSS),.VDD(VDD),.Y(I25576),.A(g25296));
  NOT NOT1_1830(.VSS(VSS),.VDD(VDD),.Y(g7443),.A(g914));
  NOT NOT1_1831(.VSS(VSS),.VDD(VDD),.Y(g8703),.A(I12709));
  NOT NOT1_1832(.VSS(VSS),.VDD(VDD),.Y(g14406),.A(g12249));
  NOT NOT1_1833(.VSS(VSS),.VDD(VDD),.Y(g19528),.A(g16349));
  NOT NOT1_1834(.VSS(VSS),.VDD(VDD),.Y(g19696),.A(g17015));
  NOT NOT1_1835(.VSS(VSS),.VDD(VDD),.Y(g34160),.A(I32119));
  NOT NOT1_1836(.VSS(VSS),.VDD(VDD),.Y(g25267),.A(g22228));
  NOT NOT1_1837(.VSS(VSS),.VDD(VDD),.Y(g19330),.A(g17326));
  NOT NOT1_1838(.VSS(VSS),.VDD(VDD),.Y(I17181),.A(g13745));
  NOT NOT1_1839(.VSS(VSS),.VDD(VDD),.Y(I17671),.A(g13280));
  NOT NOT1_1840(.VSS(VSS),.VDD(VDD),.Y(I29363),.A(g30218));
  NOT NOT1_1841(.VSS(VSS),.VDD(VDD),.Y(g23585),.A(g21070));
  NOT NOT1_1842(.VSS(VSS),.VDD(VDD),.Y(g32841),.A(g31672));
  NOT NOT1_1843(.VSS(VSS),.VDD(VDD),.Y(g11236),.A(g8357));
  NOT NOT1_1844(.VSS(VSS),.VDD(VDD),.Y(I21291),.A(g18273));
  NOT NOT1_1845(.VSS(VSS),.VDD(VDD),.Y(g7116),.A(g22));
  NOT NOT1_1846(.VSS(VSS),.VDD(VDD),.Y(g22649),.A(g19063));
  NOT NOT1_1847(.VSS(VSS),.VDD(VDD),.Y(g10500),.A(I13875));
  NOT NOT1_1848(.VSS(VSS),.VDD(VDD),.Y(g27881),.A(I26430));
  NOT NOT1_1849(.VSS(VSS),.VDD(VDD),.Y(g19365),.A(g16249));
  NOT NOT1_1850(.VSS(VSS),.VDD(VDD),.Y(g20673),.A(g15277));
  NOT NOT1_1851(.VSS(VSS),.VDD(VDD),.Y(g32510),.A(g31194));
  NOT NOT1_1852(.VSS(VSS),.VDD(VDD),.Y(g9691),.A(g1706));
  NOT NOT1_1853(.VSS(VSS),.VDD(VDD),.Y(g31801),.A(g29385));
  NOT NOT1_1854(.VSS(VSS),.VDD(VDD),.Y(I15821),.A(g11143));
  NOT NOT1_1855(.VSS(VSS),.VDD(VDD),.Y(I12056),.A(g2748));
  NOT NOT1_1856(.VSS(VSS),.VDD(VDD),.Y(g24183),.A(I23393));
  NOT NOT1_1857(.VSS(VSS),.VDD(VDD),.Y(I32904),.A(g34708));
  NOT NOT1_1858(.VSS(VSS),.VDD(VDD),.Y(g14833),.A(g11405));
  NOT NOT1_1859(.VSS(VSS),.VDD(VDD),.Y(g19869),.A(g16540));
  NOT NOT1_1860(.VSS(VSS),.VDD(VDD),.Y(g21609),.A(g18008));
  NOT NOT1_1861(.VSS(VSS),.VDD(VDD),.Y(g19960),.A(g17433));
  NOT NOT1_1862(.VSS(VSS),.VDD(VDD),.Y(g23609),.A(g21611));
  NOT NOT1_1863(.VSS(VSS),.VDD(VDD),.Y(g24397),.A(g22908));
  NOT NOT1_1864(.VSS(VSS),.VDD(VDD),.Y(g29339),.A(g28274));
  NOT NOT1_1865(.VSS(VSS),.VDD(VDD),.Y(g12881),.A(g10388));
  NOT NOT1_1866(.VSS(VSS),.VDD(VDD),.Y(g7565),.A(I12046));
  NOT NOT1_1867(.VSS(VSS),.VDD(VDD),.Y(g22903),.A(g20330));
  NOT NOT1_1868(.VSS(VSS),.VDD(VDD),.Y(g13175),.A(g10909));
  NOT NOT1_1869(.VSS(VSS),.VDD(VDD),.Y(g34915),.A(I33137));
  NOT NOT1_1870(.VSS(VSS),.VDD(VDD),.Y(I16593),.A(g10498));
  NOT NOT1_1871(.VSS(VSS),.VDD(VDD),.Y(I25115),.A(g25322));
  NOT NOT1_1872(.VSS(VSS),.VDD(VDD),.Y(g32579),.A(g30735));
  NOT NOT1_1873(.VSS(VSS),.VDD(VDD),.Y(g8068),.A(g3457));
  NOT NOT1_1874(.VSS(VSS),.VDD(VDD),.Y(I13020),.A(g6750));
  NOT NOT1_1875(.VSS(VSS),.VDD(VDD),.Y(I32621),.A(g34335));
  NOT NOT1_1876(.VSS(VSS),.VDD(VDD),.Y(g23312),.A(g21070));
  NOT NOT1_1877(.VSS(VSS),.VDD(VDD),.Y(I31569),.A(g33197));
  NOT NOT1_1878(.VSS(VSS),.VDD(VDD),.Y(I28301),.A(g29042));
  NOT NOT1_1879(.VSS(VSS),.VDD(VDD),.Y(g25219),.A(I24393));
  NOT NOT1_1880(.VSS(VSS),.VDD(VDD),.Y(I27271),.A(g27998));
  NOT NOT1_1881(.VSS(VSS),.VDD(VDD),.Y(g21608),.A(g17955));
  NOT NOT1_1882(.VSS(VSS),.VDD(VDD),.Y(g24062),.A(g19968));
  NOT NOT1_1883(.VSS(VSS),.VDD(VDD),.Y(g17649),.A(I18614));
  NOT NOT1_1884(.VSS(VSS),.VDD(VDD),.Y(g20509),.A(g15277));
  NOT NOT1_1885(.VSS(VSS),.VDD(VDD),.Y(g23608),.A(g21611));
  NOT NOT1_1886(.VSS(VSS),.VDD(VDD),.Y(g34201),.A(I32158));
  NOT NOT1_1887(.VSS(VSS),.VDD(VDD),.Y(g9607),.A(g5046));
  NOT NOT1_1888(.VSS(VSS),.VDD(VDD),.Y(g24509),.A(g22689));
  NOT NOT1_1889(.VSS(VSS),.VDD(VDD),.Y(g32578),.A(g31376));
  NOT NOT1_1890(.VSS(VSS),.VDD(VDD),.Y(g32835),.A(g31710));
  NOT NOT1_1891(.VSS(VSS),.VDD(VDD),.Y(g33695),.A(g33187));
  NOT NOT1_1892(.VSS(VSS),.VDD(VDD),.Y(g34277),.A(I32274));
  NOT NOT1_1893(.VSS(VSS),.VDD(VDD),.Y(g25218),.A(g23949));
  NOT NOT1_1894(.VSS(VSS),.VDD(VDD),.Y(g9962),.A(g6519));
  NOT NOT1_1895(.VSS(VSS),.VDD(VDD),.Y(g11790),.A(I14630));
  NOT NOT1_1896(.VSS(VSS),.VDD(VDD),.Y(g14004),.A(g11149));
  NOT NOT1_1897(.VSS(VSS),.VDD(VDD),.Y(g17648),.A(g15024));
  NOT NOT1_1898(.VSS(VSS),.VDD(VDD),.Y(g20508),.A(g15277));
  NOT NOT1_1899(.VSS(VSS),.VDD(VDD),.Y(g9158),.A(g513));
  NOT NOT1_1900(.VSS(VSS),.VDD(VDD),.Y(g27662),.A(I26296));
  NOT NOT1_1901(.VSS(VSS),.VDD(VDD),.Y(g17491),.A(g12983));
  NOT NOT1_1902(.VSS(VSS),.VDD(VDD),.Y(g22981),.A(g20283));
  NOT NOT1_1903(.VSS(VSS),.VDD(VDD),.Y(g20634),.A(g15373));
  NOT NOT1_1904(.VSS(VSS),.VDD(VDD),.Y(I21029),.A(g15816));
  NOT NOT1_1905(.VSS(VSS),.VDD(VDD),.Y(g21052),.A(g15373));
  NOT NOT1_1906(.VSS(VSS),.VDD(VDD),.Y(g28163),.A(I26682));
  NOT NOT1_1907(.VSS(VSS),.VDD(VDD),.Y(g8677),.A(g4854));
  NOT NOT1_1908(.VSS(VSS),.VDD(VDD),.Y(g25837),.A(g25064));
  NOT NOT1_1909(.VSS(VSS),.VDD(VDD),.Y(g7533),.A(g1306));
  NOT NOT1_1910(.VSS(VSS),.VDD(VDD),.Y(g19709),.A(g16987));
  NOT NOT1_1911(.VSS(VSS),.VDD(VDD),.Y(g32586),.A(g31376));
  NOT NOT1_1912(.VSS(VSS),.VDD(VDD),.Y(I22211),.A(g21463));
  NOT NOT1_1913(.VSS(VSS),.VDD(VDD),.Y(g9506),.A(g5774));
  NOT NOT1_1914(.VSS(VSS),.VDD(VDD),.Y(g17604),.A(I18555));
  NOT NOT1_1915(.VSS(VSS),.VDD(VDD),.Y(g34595),.A(I32693));
  NOT NOT1_1916(.VSS(VSS),.VDD(VDD),.Y(g7697),.A(g4087));
  NOT NOT1_1917(.VSS(VSS),.VDD(VDD),.Y(g10613),.A(g10233));
  NOT NOT1_1918(.VSS(VSS),.VDD(VDD),.Y(g23745),.A(g20900));
  NOT NOT1_1919(.VSS(VSS),.VDD(VDD),.Y(I18504),.A(g5283));
  NOT NOT1_1920(.VSS(VSS),.VDD(VDD),.Y(I22024),.A(g19350));
  NOT NOT1_1921(.VSS(VSS),.VDD(VDD),.Y(g32442),.A(g31213));
  NOT NOT1_1922(.VSS(VSS),.VDD(VDD),.Y(I31814),.A(g33149));
  NOT NOT1_1923(.VSS(VSS),.VDD(VDD),.Y(g19471),.A(g16449));
  NOT NOT1_1924(.VSS(VSS),.VDD(VDD),.Y(g30037),.A(g29121));
  NOT NOT1_1925(.VSS(VSS),.VDD(VDD),.Y(g12890),.A(g10397));
  NOT NOT1_1926(.VSS(VSS),.VDD(VDD),.Y(g16580),.A(I17754));
  NOT NOT1_1927(.VSS(VSS),.VDD(VDD),.Y(g23813),.A(g18997));
  NOT NOT1_1928(.VSS(VSS),.VDD(VDD),.Y(g7596),.A(I12070));
  NOT NOT1_1929(.VSS(VSS),.VDD(VDD),.Y(I31751),.A(g33228));
  NOT NOT1_1930(.VSS(VSS),.VDD(VDD),.Y(I31807),.A(g33149));
  NOT NOT1_1931(.VSS(VSS),.VDD(VDD),.Y(g16223),.A(g13437));
  NOT NOT1_1932(.VSS(VSS),.VDD(VDD),.Y(g10273),.A(I13708));
  NOT NOT1_1933(.VSS(VSS),.VDD(VDD),.Y(g33457),.A(I30989));
  NOT NOT1_1934(.VSS(VSS),.VDD(VDD),.Y(I32062),.A(g33653));
  NOT NOT1_1935(.VSS(VSS),.VDD(VDD),.Y(I12199),.A(g6215));
  NOT NOT1_1936(.VSS(VSS),.VDD(VDD),.Y(g10106),.A(g16));
  NOT NOT1_1937(.VSS(VSS),.VDD(VDD),.Y(g9311),.A(g5523));
  NOT NOT1_1938(.VSS(VSS),.VDD(VDD),.Y(I11743),.A(g4564));
  NOT NOT1_1939(.VSS(VSS),.VDD(VDD),.Y(g22845),.A(g20682));
  NOT NOT1_1940(.VSS(VSS),.VDD(VDD),.Y(I12887),.A(g4216));
  NOT NOT1_1941(.VSS(VSS),.VDD(VDD),.Y(g34984),.A(I33252));
  NOT NOT1_1942(.VSS(VSS),.VDD(VDD),.Y(g32615),.A(g31376));
  NOT NOT1_1943(.VSS(VSS),.VDD(VDD),.Y(I15834),.A(g11164));
  NOT NOT1_1944(.VSS(VSS),.VDD(VDD),.Y(g13209),.A(g10632));
  NOT NOT1_1945(.VSS(VSS),.VDD(VDD),.Y(g8848),.A(g358));
  NOT NOT1_1946(.VSS(VSS),.VDD(VDD),.Y(g20213),.A(g17062));
  NOT NOT1_1947(.VSS(VSS),.VDD(VDD),.Y(I15208),.A(g637));
  NOT NOT1_1948(.VSS(VSS),.VDD(VDD),.Y(g33917),.A(I31779));
  NOT NOT1_1949(.VSS(VSS),.VDD(VDD),.Y(g21184),.A(g15509));
  NOT NOT1_1950(.VSS(VSS),.VDD(VDD),.Y(g34419),.A(g34151));
  NOT NOT1_1951(.VSS(VSS),.VDD(VDD),.Y(g9615),.A(I13236));
  NOT NOT1_1952(.VSS(VSS),.VDD(VDD),.Y(g21674),.A(g16540));
  NOT NOT1_1953(.VSS(VSS),.VDD(VDD),.Y(g10812),.A(I14050));
  NOT NOT1_1954(.VSS(VSS),.VDD(VDD),.Y(g32720),.A(g31710));
  NOT NOT1_1955(.VSS(VSS),.VDD(VDD),.Y(g30155),.A(I28390));
  NOT NOT1_1956(.VSS(VSS),.VDD(VDD),.Y(g8398),.A(I12563));
  NOT NOT1_1957(.VSS(VSS),.VDD(VDD),.Y(g28325),.A(g27463));
  NOT NOT1_1958(.VSS(VSS),.VDD(VDD),.Y(g12779),.A(g9444));
  NOT NOT1_1959(.VSS(VSS),.VDD(VDD),.Y(g22898),.A(g20283));
  NOT NOT1_1960(.VSS(VSS),.VDD(VDD),.Y(g9174),.A(g1205));
  NOT NOT1_1961(.VSS(VSS),.VDD(VDD),.Y(g34418),.A(g34150));
  NOT NOT1_1962(.VSS(VSS),.VDD(VDD),.Y(g17794),.A(g13350));
  NOT NOT1_1963(.VSS(VSS),.VDD(VDD),.Y(g26836),.A(g24866));
  NOT NOT1_1964(.VSS(VSS),.VDD(VDD),.Y(g17845),.A(I18835));
  NOT NOT1_1965(.VSS(VSS),.VDD(VDD),.Y(g9374),.A(g5188));
  NOT NOT1_1966(.VSS(VSS),.VDD(VDD),.Y(g20574),.A(g17847));
  NOT NOT1_1967(.VSS(VSS),.VDD(VDD),.Y(g20452),.A(g17200));
  NOT NOT1_1968(.VSS(VSS),.VDD(VDD),.Y(I15542),.A(g1570));
  NOT NOT1_1969(.VSS(VSS),.VDD(VDD),.Y(g32430),.A(g30984));
  NOT NOT1_1970(.VSS(VSS),.VDD(VDD),.Y(g10033),.A(g655));
  NOT NOT1_1971(.VSS(VSS),.VDD(VDD),.Y(g10371),.A(g6918));
  NOT NOT1_1972(.VSS(VSS),.VDD(VDD),.Y(g32746),.A(g30735));
  NOT NOT1_1973(.VSS(VSS),.VDD(VDD),.Y(g32493),.A(g30735));
  NOT NOT1_1974(.VSS(VSS),.VDD(VDD),.Y(g22719),.A(I22024));
  NOT NOT1_1975(.VSS(VSS),.VDD(VDD),.Y(g24452),.A(g22722));
  NOT NOT1_1976(.VSS(VSS),.VDD(VDD),.Y(I26100),.A(g26365));
  NOT NOT1_1977(.VSS(VSS),.VDD(VDD),.Y(g7936),.A(g1061));
  NOT NOT1_1978(.VSS(VSS),.VDD(VDD),.Y(g9985),.A(g4332));
  NOT NOT1_1979(.VSS(VSS),.VDD(VDD),.Y(g24047),.A(g19919));
  NOT NOT1_1980(.VSS(VSS),.VDD(VDD),.Y(g12778),.A(g9856));
  NOT NOT1_1981(.VSS(VSS),.VDD(VDD),.Y(I18245),.A(g14676));
  NOT NOT1_1982(.VSS(VSS),.VDD(VDD),.Y(I12764),.A(g4194));
  NOT NOT1_1983(.VSS(VSS),.VDD(VDD),.Y(g23732),.A(g18833));
  NOT NOT1_1984(.VSS(VSS),.VDD(VDD),.Y(g8241),.A(g1792));
  NOT NOT1_1985(.VSS(VSS),.VDD(VDD),.Y(I20793),.A(g17694));
  NOT NOT1_1986(.VSS(VSS),.VDD(VDD),.Y(g20912),.A(g15171));
  NOT NOT1_1987(.VSS(VSS),.VDD(VDD),.Y(g19602),.A(g16349));
  NOT NOT1_1988(.VSS(VSS),.VDD(VDD),.Y(g32465),.A(g30825));
  NOT NOT1_1989(.VSS(VSS),.VDD(VDD),.Y(g7117),.A(I11816));
  NOT NOT1_1990(.VSS(VSS),.VDD(VDD),.Y(I18323),.A(g13680));
  NOT NOT1_1991(.VSS(VSS),.VDD(VDD),.Y(g19657),.A(g16349));
  NOT NOT1_1992(.VSS(VSS),.VDD(VDD),.Y(g22718),.A(g20887));
  NOT NOT1_1993(.VSS(VSS),.VDD(VDD),.Y(g16740),.A(g13980));
  NOT NOT1_1994(.VSS(VSS),.VDD(VDD),.Y(I12132),.A(g577));
  NOT NOT1_1995(.VSS(VSS),.VDD(VDD),.Y(g19068),.A(g16031));
  NOT NOT1_1996(.VSS(VSS),.VDD(VDD),.Y(g15169),.A(I17094));
  NOT NOT1_1997(.VSS(VSS),.VDD(VDD),.Y(g28121),.A(g27093));
  NOT NOT1_1998(.VSS(VSS),.VDD(VDD),.Y(g9284),.A(g2161));
  NOT NOT1_1999(.VSS(VSS),.VDD(VDD),.Y(g19375),.A(I19863));
  NOT NOT1_2000(.VSS(VSS),.VDD(VDD),.Y(g10795),.A(g7202));
  NOT NOT1_2001(.VSS(VSS),.VDD(VDD),.Y(I25692),.A(g25689));
  NOT NOT1_2002(.VSS(VSS),.VDD(VDD),.Y(g9239),.A(g5511));
  NOT NOT1_2003(.VSS(VSS),.VDD(VDD),.Y(g33923),.A(I31791));
  NOT NOT1_2004(.VSS(VSS),.VDD(VDD),.Y(g9180),.A(g3719));
  NOT NOT1_2005(.VSS(VSS),.VDD(VDD),.Y(g16186),.A(g13555));
  NOT NOT1_2006(.VSS(VSS),.VDD(VDD),.Y(g16676),.A(I17876));
  NOT NOT1_2007(.VSS(VSS),.VDD(VDD),.Y(g16685),.A(g14038));
  NOT NOT1_2008(.VSS(VSS),.VDD(VDD),.Y(I20690),.A(g15733));
  NOT NOT1_2009(.VSS(VSS),.VDD(VDD),.Y(I29936),.A(g30606));
  NOT NOT1_2010(.VSS(VSS),.VDD(VDD),.Y(I17658),.A(g13394));
  NOT NOT1_2011(.VSS(VSS),.VDD(VDD),.Y(g9380),.A(g5471));
  NOT NOT1_2012(.VSS(VSS),.VDD(VDD),.Y(g12945),.A(g12467));
  NOT NOT1_2013(.VSS(VSS),.VDD(VDD),.Y(g31624),.A(I29218));
  NOT NOT1_2014(.VSS(VSS),.VDD(VDD),.Y(g32806),.A(g31710));
  NOT NOT1_2015(.VSS(VSS),.VDD(VDD),.Y(g20072),.A(g17384));
  NOT NOT1_2016(.VSS(VSS),.VDD(VDD),.Y(g32684),.A(g30673));
  NOT NOT1_2017(.VSS(VSS),.VDD(VDD),.Y(g33688),.A(I31523));
  NOT NOT1_2018(.VSS(VSS),.VDD(VDD),.Y(g29707),.A(g28504));
  NOT NOT1_2019(.VSS(VSS),.VDD(VDD),.Y(g9832),.A(g2399));
  NOT NOT1_2020(.VSS(VSS),.VDD(VDD),.Y(I15073),.A(g10109));
  NOT NOT1_2021(.VSS(VSS),.VDD(VDD),.Y(g19878),.A(g17271));
  NOT NOT1_2022(.VSS(VSS),.VDD(VDD),.Y(g24051),.A(g21127));
  NOT NOT1_2023(.VSS(VSS),.VDD(VDD),.Y(g24072),.A(g20982));
  NOT NOT1_2024(.VSS(VSS),.VDD(VDD),.Y(g34589),.A(I32675));
  NOT NOT1_2025(.VSS(VSS),.VDD(VDD),.Y(g17718),.A(g14776));
  NOT NOT1_2026(.VSS(VSS),.VDD(VDD),.Y(g17521),.A(g14727));
  NOT NOT1_2027(.VSS(VSS),.VDD(VDD),.Y(g16654),.A(g14136));
  NOT NOT1_2028(.VSS(VSS),.VDD(VDD),.Y(g20592),.A(g15277));
  NOT NOT1_2029(.VSS(VSS),.VDD(VDD),.Y(g27998),.A(I26512));
  NOT NOT1_2030(.VSS(VSS),.VDD(VDD),.Y(I16575),.A(g3298));
  NOT NOT1_2031(.VSS(VSS),.VDD(VDD),.Y(g15479),.A(g14895));
  NOT NOT1_2032(.VSS(VSS),.VDD(VDD),.Y(g9853),.A(g5297));
  NOT NOT1_2033(.VSS(VSS),.VDD(VDD),.Y(I15593),.A(g11989));
  NOT NOT1_2034(.VSS(VSS),.VDD(VDD),.Y(g8644),.A(g3352));
  NOT NOT1_2035(.VSS(VSS),.VDD(VDD),.Y(g6989),.A(g4575));
  NOT NOT1_2036(.VSS(VSS),.VDD(VDD),.Y(g9020),.A(g4287));
  NOT NOT1_2037(.VSS(VSS),.VDD(VDD),.Y(g24756),.A(g22763));
  NOT NOT1_2038(.VSS(VSS),.VDD(VDD),.Y(I32452),.A(g34241));
  NOT NOT1_2039(.VSS(VSS),.VDD(VDD),.Y(I12709),.A(g4284));
  NOT NOT1_2040(.VSS(VSS),.VDD(VDD),.Y(g21400),.A(g17847));
  NOT NOT1_2041(.VSS(VSS),.VDD(VDD),.Y(g20780),.A(g15509));
  NOT NOT1_2042(.VSS(VSS),.VDD(VDD),.Y(g7922),.A(g1312));
  NOT NOT1_2043(.VSS(VSS),.VDD(VDD),.Y(g8119),.A(g3727));
  NOT NOT1_2044(.VSS(VSS),.VDD(VDD),.Y(g13530),.A(g12641));
  NOT NOT1_2045(.VSS(VSS),.VDD(VDD),.Y(g23400),.A(g20676));
  NOT NOT1_2046(.VSS(VSS),.VDD(VDD),.Y(g12998),.A(g11829));
  NOT NOT1_2047(.VSS(VSS),.VDD(VDD),.Y(g34836),.A(I33050));
  NOT NOT1_2048(.VSS(VSS),.VDD(VDD),.Y(g13593),.A(g10556));
  NOT NOT1_2049(.VSS(VSS),.VDD(VDD),.Y(g28173),.A(I26693));
  NOT NOT1_2050(.VSS(VSS),.VDD(VDD),.Y(g18929),.A(g16100));
  NOT NOT1_2051(.VSS(VSS),.VDD(VDD),.Y(g32517),.A(g31194));
  NOT NOT1_2052(.VSS(VSS),.VDD(VDD),.Y(g23013),.A(g20330));
  NOT NOT1_2053(.VSS(VSS),.VDD(VDD),.Y(I28572),.A(g28274));
  NOT NOT1_2054(.VSS(VSS),.VDD(VDD),.Y(g12233),.A(g10338));
  NOT NOT1_2055(.VSS(VSS),.VDD(VDD),.Y(I31586),.A(g33149));
  NOT NOT1_2056(.VSS(VSS),.VDD(VDD),.Y(g23214),.A(g20785));
  NOT NOT1_2057(.VSS(VSS),.VDD(VDD),.Y(g11122),.A(g8751));
  NOT NOT1_2058(.VSS(VSS),.VDD(VDD),.Y(I14902),.A(g9821));
  NOT NOT1_2059(.VSS(VSS),.VDD(VDD),.Y(I14301),.A(g8571));
  NOT NOT1_2060(.VSS(VSS),.VDD(VDD),.Y(g12182),.A(I15030));
  NOT NOT1_2061(.VSS(VSS),.VDD(VDD),.Y(g29978),.A(g28927));
  NOT NOT1_2062(.VSS(VSS),.VDD(VDD),.Y(g12672),.A(g10003));
  NOT NOT1_2063(.VSS(VSS),.VDD(VDD),.Y(g7581),.A(g1379));
  NOT NOT1_2064(.VSS(VSS),.VDD(VDD),.Y(g21329),.A(g16577));
  NOT NOT1_2065(.VSS(VSS),.VDD(VDD),.Y(g22926),.A(g20391));
  NOT NOT1_2066(.VSS(VSS),.VDD(VDD),.Y(g25155),.A(g22472));
  NOT NOT1_2067(.VSS(VSS),.VDD(VDD),.Y(g9559),.A(g6077));
  NOT NOT1_2068(.VSS(VSS),.VDD(VDD),.Y(g13565),.A(g11006));
  NOT NOT1_2069(.VSS(VSS),.VDD(VDD),.Y(g6971),.A(I11737));
  NOT NOT1_2070(.VSS(VSS),.VDD(VDD),.Y(g8818),.A(I12808));
  NOT NOT1_2071(.VSS(VSS),.VDD(VDD),.Y(I25005),.A(g24417));
  NOT NOT1_2072(.VSS(VSS),.VDD(VDD),.Y(g14421),.A(I16575));
  NOT NOT1_2073(.VSS(VSS),.VDD(VDD),.Y(I19704),.A(g17653));
  NOT NOT1_2074(.VSS(VSS),.VDD(VDD),.Y(g25266),.A(g22228));
  NOT NOT1_2075(.VSS(VSS),.VDD(VDD),.Y(g25170),.A(g22498));
  NOT NOT1_2076(.VSS(VSS),.VDD(VDD),.Y(g9931),.A(g5763));
  NOT NOT1_2077(.VSS(VSS),.VDD(VDD),.Y(g23539),.A(g21070));
  NOT NOT1_2078(.VSS(VSS),.VDD(VDD),.Y(g17573),.A(g12911));
  NOT NOT1_2079(.VSS(VSS),.VDD(VDD),.Y(g7597),.A(g952));
  NOT NOT1_2080(.VSS(VSS),.VDD(VDD),.Y(g11034),.A(g7611));
  NOT NOT1_2081(.VSS(VSS),.VDD(VDD),.Y(g23005),.A(g20283));
  NOT NOT1_2082(.VSS(VSS),.VDD(VDD),.Y(g13034),.A(g11920));
  NOT NOT1_2083(.VSS(VSS),.VDD(VDD),.Y(g17247),.A(I18259));
  NOT NOT1_2084(.VSS(VSS),.VDD(VDD),.Y(I32051),.A(g33631));
  NOT NOT1_2085(.VSS(VSS),.VDD(VDD),.Y(g30022),.A(g29001));
  NOT NOT1_2086(.VSS(VSS),.VDD(VDD),.Y(g34118),.A(I32051));
  NOT NOT1_2087(.VSS(VSS),.VDD(VDD),.Y(I16606),.A(g3649));
  NOT NOT1_2088(.VSS(VSS),.VDD(VDD),.Y(g15580),.A(g13242));
  NOT NOT1_2089(.VSS(VSS),.VDD(VDD),.Y(g12932),.A(I15550));
  NOT NOT1_2090(.VSS(VSS),.VDD(VDD),.Y(g23538),.A(g20924));
  NOT NOT1_2091(.VSS(VSS),.VDD(VDD),.Y(g34864),.A(g34840));
  NOT NOT1_2092(.VSS(VSS),.VDD(VDD),.Y(I16492),.A(g12430));
  NOT NOT1_2093(.VSS(VSS),.VDD(VDD),.Y(g17389),.A(g14915));
  NOT NOT1_2094(.VSS(VSS),.VDD(VDD),.Y(g17926),.A(I18852));
  NOT NOT1_2095(.VSS(VSS),.VDD(VDD),.Y(g16964),.A(I18120));
  NOT NOT1_2096(.VSS(VSS),.VDD(VDD),.Y(g24152),.A(I23300));
  NOT NOT1_2097(.VSS(VSS),.VDD(VDD),.Y(g19458),.A(I19927));
  NOT NOT1_2098(.VSS(VSS),.VDD(VDD),.Y(g30313),.A(g28843));
  NOT NOT1_2099(.VSS(VSS),.VDD(VDD),.Y(g34749),.A(I32921));
  NOT NOT1_2100(.VSS(VSS),.VDD(VDD),.Y(g17612),.A(g15014));
  NOT NOT1_2101(.VSS(VSS),.VDD(VDD),.Y(g24396),.A(g22885));
  NOT NOT1_2102(.VSS(VSS),.VDD(VDD),.Y(g8211),.A(g2319));
  NOT NOT1_2103(.VSS(VSS),.VDD(VDD),.Y(g29067),.A(I27401));
  NOT NOT1_2104(.VSS(VSS),.VDD(VDD),.Y(g9905),.A(g802));
  NOT NOT1_2105(.VSS(VSS),.VDD(VDD),.Y(g10541),.A(g9407));
  NOT NOT1_2106(.VSS(VSS),.VDD(VDD),.Y(g16423),.A(g14066));
  NOT NOT1_2107(.VSS(VSS),.VDD(VDD),.Y(g27961),.A(g26816));
  NOT NOT1_2108(.VSS(VSS),.VDD(VDD),.Y(g8186),.A(g990));
  NOT NOT1_2109(.VSS(VSS),.VDD(VDD),.Y(g34313),.A(g34086));
  NOT NOT1_2110(.VSS(VSS),.VDD(VDD),.Y(I13552),.A(g121));
  NOT NOT1_2111(.VSS(VSS),.VDD(VDD),.Y(g10473),.A(I13857));
  NOT NOT1_2112(.VSS(VSS),.VDD(VDD),.Y(g17324),.A(I18301));
  NOT NOT1_2113(.VSS(VSS),.VDD(VDD),.Y(g32523),.A(g30825));
  NOT NOT1_2114(.VSS(VSS),.VDD(VDD),.Y(I24128),.A(g23009));
  NOT NOT1_2115(.VSS(VSS),.VDD(VDD),.Y(g31854),.A(g29385));
  NOT NOT1_2116(.VSS(VSS),.VDD(VDD),.Y(g14541),.A(g11405));
  NOT NOT1_2117(.VSS(VSS),.VDD(VDD),.Y(g16216),.A(I17557));
  NOT NOT1_2118(.VSS(VSS),.VDD(VDD),.Y(I29909),.A(g31791));
  NOT NOT1_2119(.VSS(VSS),.VDD(VDD),.Y(I33041),.A(g34772));
  NOT NOT1_2120(.VSS(VSS),.VDD(VDD),.Y(g12897),.A(g10400));
  NOT NOT1_2121(.VSS(VSS),.VDD(VDD),.Y(g13409),.A(I15918));
  NOT NOT1_2122(.VSS(VSS),.VDD(VDD),.Y(g16587),.A(I17763));
  NOT NOT1_2123(.VSS(VSS),.VDD(VDD),.Y(g17777),.A(g14908));
  NOT NOT1_2124(.VSS(VSS),.VDD(VDD),.Y(g25167),.A(I24331));
  NOT NOT1_2125(.VSS(VSS),.VDD(VDD),.Y(g25194),.A(g22763));
  NOT NOT1_2126(.VSS(VSS),.VDD(VDD),.Y(I13779),.A(g6868));
  NOT NOT1_2127(.VSS(VSS),.VDD(VDD),.Y(I26584),.A(g26943));
  NOT NOT1_2128(.VSS(VSS),.VDD(VDD),.Y(g9630),.A(g6527));
  NOT NOT1_2129(.VSS(VSS),.VDD(VDD),.Y(g29150),.A(g27886));
  NOT NOT1_2130(.VSS(VSS),.VDD(VDD),.Y(g34276),.A(g34058));
  NOT NOT1_2131(.VSS(VSS),.VDD(VDD),.Y(g34285),.A(I32284));
  NOT NOT1_2132(.VSS(VSS),.VDD(VDD),.Y(g7995),.A(g153));
  NOT NOT1_2133(.VSS(VSS),.VDD(VDD),.Y(g30305),.A(g28939));
  NOT NOT1_2134(.VSS(VSS),.VDD(VDD),.Y(g11136),.A(I14192));
  NOT NOT1_2135(.VSS(VSS),.VDD(VDD),.Y(g30053),.A(g29121));
  NOT NOT1_2136(.VSS(VSS),.VDD(VDD),.Y(g8026),.A(g3857));
  NOT NOT1_2137(.VSS(VSS),.VDD(VDD),.Y(g25524),.A(g22228));
  NOT NOT1_2138(.VSS(VSS),.VDD(VDD),.Y(I27970),.A(g28803));
  NOT NOT1_2139(.VSS(VSS),.VDD(VDD),.Y(g18827),.A(g16000));
  NOT NOT1_2140(.VSS(VSS),.VDD(VDD),.Y(g34053),.A(g33683));
  NOT NOT1_2141(.VSS(VSS),.VDD(VDD),.Y(g7479),.A(g1008));
  NOT NOT1_2142(.VSS(VSS),.VDD(VDD),.Y(g9300),.A(g5180));
  NOT NOT1_2143(.VSS(VSS),.VDD(VDD),.Y(g10359),.A(g6830));
  NOT NOT1_2144(.VSS(VSS),.VDD(VDD),.Y(I32820),.A(g34474));
  NOT NOT1_2145(.VSS(VSS),.VDD(VDD),.Y(g8426),.A(g3045));
  NOT NOT1_2146(.VSS(VSS),.VDD(VDD),.Y(g32475),.A(g30614));
  NOT NOT1_2147(.VSS(VSS),.VDD(VDD),.Y(g14359),.A(I16515));
  NOT NOT1_2148(.VSS(VSS),.VDD(VDD),.Y(g8170),.A(g3770));
  NOT NOT1_2149(.VSS(VSS),.VDD(VDD),.Y(g7840),.A(g4878));
  NOT NOT1_2150(.VSS(VSS),.VDD(VDD),.Y(g22997),.A(g20391));
  NOT NOT1_2151(.VSS(VSS),.VDD(VDD),.Y(g32727),.A(g31710));
  NOT NOT1_2152(.VSS(VSS),.VDD(VDD),.Y(g10358),.A(g6827));
  NOT NOT1_2153(.VSS(VSS),.VDD(VDD),.Y(g33660),.A(I31494));
  NOT NOT1_2154(.VSS(VSS),.VDD(VDD),.Y(g32863),.A(g31021));
  NOT NOT1_2155(.VSS(VSS),.VDD(VDD),.Y(g29196),.A(g27059));
  NOT NOT1_2156(.VSS(VSS),.VDD(VDD),.Y(I32846),.A(g34502));
  NOT NOT1_2157(.VSS(VSS),.VDD(VDD),.Y(g14535),.A(g12318));
  NOT NOT1_2158(.VSS(VSS),.VDD(VDD),.Y(g24405),.A(g22722));
  NOT NOT1_2159(.VSS(VSS),.VDD(VDD),.Y(g8125),.A(g3869));
  NOT NOT1_2160(.VSS(VSS),.VDD(VDD),.Y(g30036),.A(g29085));
  NOT NOT1_2161(.VSS(VSS),.VDD(VDD),.Y(g14358),.A(I16512));
  NOT NOT1_2162(.VSS(VSS),.VDD(VDD),.Y(g25119),.A(g22384));
  NOT NOT1_2163(.VSS(VSS),.VDD(VDD),.Y(I22819),.A(g19862));
  NOT NOT1_2164(.VSS(VSS),.VDD(VDD),.Y(g8821),.A(I12811));
  NOT NOT1_2165(.VSS(VSS),.VDD(VDD),.Y(g16000),.A(I17425));
  NOT NOT1_2166(.VSS(VSS),.VDD(VDD),.Y(g15740),.A(g13342));
  NOT NOT1_2167(.VSS(VSS),.VDD(VDD),.Y(I25683),.A(g25642));
  NOT NOT1_2168(.VSS(VSS),.VDD(VDD),.Y(I29242),.A(g29313));
  NOT NOT1_2169(.VSS(VSS),.VDD(VDD),.Y(g32437),.A(I29965));
  NOT NOT1_2170(.VSS(VSS),.VDD(VDD),.Y(g14828),.A(I16875));
  NOT NOT1_2171(.VSS(VSS),.VDD(VDD),.Y(g23235),.A(g20785));
  NOT NOT1_2172(.VSS(VSS),.VDD(VDD),.Y(g33456),.A(I30986));
  NOT NOT1_2173(.VSS(VSS),.VDD(VDD),.Y(g10121),.A(g2327));
  NOT NOT1_2174(.VSS(VSS),.VDD(VDD),.Y(g11164),.A(g8085));
  NOT NOT1_2175(.VSS(VSS),.VDD(VDD),.Y(g25118),.A(g22417));
  NOT NOT1_2176(.VSS(VSS),.VDD(VDD),.Y(g26693),.A(g25300));
  NOT NOT1_2177(.VSS(VSS),.VDD(VDD),.Y(g8280),.A(g3443));
  NOT NOT1_2178(.VSS(VSS),.VDD(VDD),.Y(g23683),.A(I22816));
  NOT NOT1_2179(.VSS(VSS),.VDD(VDD),.Y(g15373),.A(I17118));
  NOT NOT1_2180(.VSS(VSS),.VDD(VDD),.Y(g9973),.A(g2112));
  NOT NOT1_2181(.VSS(VSS),.VDD(VDD),.Y(g33916),.A(I31776));
  NOT NOT1_2182(.VSS(VSS),.VDD(VDD),.Y(I22111),.A(g19919));
  NOT NOT1_2183(.VSS(VSS),.VDD(VDD),.Y(g7356),.A(g1802));
  NOT NOT1_2184(.VSS(VSS),.VDD(VDD),.Y(I17819),.A(g3618));
  NOT NOT1_2185(.VSS(VSS),.VDD(VDD),.Y(g16747),.A(g14113));
  NOT NOT1_2186(.VSS(VSS),.VDD(VDD),.Y(g20583),.A(g17873));
  NOT NOT1_2187(.VSS(VSS),.VDD(VDD),.Y(g32703),.A(g30825));
  NOT NOT1_2188(.VSS(VSS),.VDD(VDD),.Y(I12994),.A(g6748));
  NOT NOT1_2189(.VSS(VSS),.VDD(VDD),.Y(I15474),.A(g10364));
  NOT NOT1_2190(.VSS(VSS),.VDD(VDD),.Y(g24020),.A(g20014));
  NOT NOT1_2191(.VSS(VSS),.VDD(VDD),.Y(g19532),.A(g16821));
  NOT NOT1_2192(.VSS(VSS),.VDD(VDD),.Y(g22360),.A(I21849));
  NOT NOT1_2193(.VSS(VSS),.VDD(VDD),.Y(g9040),.A(g499));
  NOT NOT1_2194(.VSS(VSS),.VDD(VDD),.Y(g28648),.A(g27693));
  NOT NOT1_2195(.VSS(VSS),.VDD(VDD),.Y(g18881),.A(I19671));
  NOT NOT1_2196(.VSS(VSS),.VDD(VDD),.Y(I13672),.A(g106));
  NOT NOT1_2197(.VSS(VSS),.VDD(VDD),.Y(g13474),.A(g11048));
  NOT NOT1_2198(.VSS(VSS),.VDD(VDD),.Y(I25882),.A(g25776));
  NOT NOT1_2199(.VSS(VSS),.VDD(VDD),.Y(g20046),.A(g16540));
  NOT NOT1_2200(.VSS(VSS),.VDD(VDD),.Y(g9969),.A(g1682));
  NOT NOT1_2201(.VSS(VSS),.VDD(VDD),.Y(g19783),.A(g16931));
  NOT NOT1_2202(.VSS(VSS),.VDD(VDD),.Y(I17111),.A(g13809));
  NOT NOT1_2203(.VSS(VSS),.VDD(VDD),.Y(g16123),.A(g13530));
  NOT NOT1_2204(.VSS(VSS),.VDD(VDD),.Y(g24046),.A(g21256));
  NOT NOT1_2205(.VSS(VSS),.VDD(VDD),.Y(g17871),.A(I18845));
  NOT NOT1_2206(.VSS(VSS),.VDD(VDD),.Y(g16814),.A(g14058));
  NOT NOT1_2207(.VSS(VSS),.VDD(VDD),.Y(g21414),.A(g17929));
  NOT NOT1_2208(.VSS(VSS),.VDD(VDD),.Y(g32600),.A(g31542));
  NOT NOT1_2209(.VSS(VSS),.VDD(VDD),.Y(g7704),.A(I12167));
  NOT NOT1_2210(.VSS(VSS),.VDD(VDD),.Y(I16663),.A(g10981));
  NOT NOT1_2211(.VSS(VSS),.VDD(VDD),.Y(g23515),.A(g20785));
  NOT NOT1_2212(.VSS(VSS),.VDD(VDD),.Y(g28604),.A(g27759));
  NOT NOT1_2213(.VSS(VSS),.VDD(VDD),.Y(g23882),.A(g19277));
  NOT NOT1_2214(.VSS(VSS),.VDD(VDD),.Y(g23414),.A(I22525));
  NOT NOT1_2215(.VSS(VSS),.VDD(VDD),.Y(g32781),.A(g31376));
  NOT NOT1_2216(.VSS(VSS),.VDD(VDD),.Y(I23099),.A(g20682));
  NOT NOT1_2217(.VSS(VSS),.VDD(VDD),.Y(g31596),.A(I29204));
  NOT NOT1_2218(.VSS(VSS),.VDD(VDD),.Y(g8106),.A(g3133));
  NOT NOT1_2219(.VSS(VSS),.VDD(VDD),.Y(g14173),.A(g12076));
  NOT NOT1_2220(.VSS(VSS),.VDD(VDD),.Y(I23324),.A(g21697));
  NOT NOT1_2221(.VSS(VSS),.VDD(VDD),.Y(g20113),.A(g16826));
  NOT NOT1_2222(.VSS(VSS),.VDD(VDD),.Y(g21407),.A(g15171));
  NOT NOT1_2223(.VSS(VSS),.VDD(VDD),.Y(g31243),.A(g29933));
  NOT NOT1_2224(.VSS(VSS),.VDD(VDD),.Y(I17590),.A(g14591));
  NOT NOT1_2225(.VSS(VSS),.VDD(VDD),.Y(g19353),.A(I19831));
  NOT NOT1_2226(.VSS(VSS),.VDD(VDD),.Y(g24113),.A(g19984));
  NOT NOT1_2227(.VSS(VSS),.VDD(VDD),.Y(I32929),.A(g34649));
  NOT NOT1_2228(.VSS(VSS),.VDD(VDD),.Y(g32952),.A(g30937));
  NOT NOT1_2229(.VSS(VSS),.VDD(VDD),.Y(g19144),.A(g16031));
  NOT NOT1_2230(.VSS(VSS),.VDD(VDD),.Y(g12811),.A(g10319));
  NOT NOT1_2231(.VSS(VSS),.VDD(VDD),.Y(g27971),.A(g26673));
  NOT NOT1_2232(.VSS(VSS),.VDD(VDD),.Y(g8187),.A(g1657));
  NOT NOT1_2233(.VSS(VSS),.VDD(VDD),.Y(g32821),.A(g31021));
  NOT NOT1_2234(.VSS(VSS),.VDD(VDD),.Y(g8387),.A(g3080));
  NOT NOT1_2235(.VSS(VSS),.VDD(VDD),.Y(g25036),.A(g23733));
  NOT NOT1_2236(.VSS(VSS),.VDD(VDD),.Y(I31523),.A(g33187));
  NOT NOT1_2237(.VSS(VSS),.VDD(VDD),.Y(g7163),.A(g4593));
  NOT NOT1_2238(.VSS(VSS),.VDD(VDD),.Y(g29597),.A(g28444));
  NOT NOT1_2239(.VSS(VSS),.VDD(VDD),.Y(g25101),.A(g22384));
  NOT NOT1_2240(.VSS(VSS),.VDD(VDD),.Y(g20105),.A(g17433));
  NOT NOT1_2241(.VSS(VSS),.VDD(VDD),.Y(g24357),.A(g22325));
  NOT NOT1_2242(.VSS(VSS),.VDD(VDD),.Y(g25560),.A(g22550));
  NOT NOT1_2243(.VSS(VSS),.VDD(VDD),.Y(g10029),.A(I13548));
  NOT NOT1_2244(.VSS(VSS),.VDD(VDD),.Y(g8756),.A(g4049));
  NOT NOT1_2245(.VSS(VSS),.VDD(VDD),.Y(g22220),.A(I21802));
  NOT NOT1_2246(.VSS(VSS),.VDD(VDD),.Y(g13303),.A(I15869));
  NOT NOT1_2247(.VSS(VSS),.VDD(VDD),.Y(g24105),.A(g19935));
  NOT NOT1_2248(.VSS(VSS),.VDD(VDD),.Y(I17094),.A(g14331));
  NOT NOT1_2249(.VSS(VSS),.VDD(VDD),.Y(I18031),.A(g13680));
  NOT NOT1_2250(.VSS(VSS),.VDD(VDD),.Y(g29689),.A(I27954));
  NOT NOT1_2251(.VSS(VSS),.VDD(VDD),.Y(g14029),.A(g11283));
  NOT NOT1_2252(.VSS(VSS),.VDD(VDD),.Y(g29923),.A(g28874));
  NOT NOT1_2253(.VSS(VSS),.VDD(VDD),.Y(g25642),.A(I24787));
  NOT NOT1_2254(.VSS(VSS),.VDD(VDD),.Y(g32790),.A(g30825));
  NOT NOT1_2255(.VSS(VSS),.VDD(VDD),.Y(g9648),.A(g2177));
  NOT NOT1_2256(.VSS(VSS),.VDD(VDD),.Y(g32137),.A(g31134));
  NOT NOT1_2257(.VSS(VSS),.VDD(VDD),.Y(g10028),.A(g8));
  NOT NOT1_2258(.VSS(VSS),.VDD(VDD),.Y(g9875),.A(g5747));
  NOT NOT1_2259(.VSS(VSS),.VDD(VDD),.Y(g32516),.A(g31070));
  NOT NOT1_2260(.VSS(VSS),.VDD(VDD),.Y(g31655),.A(I29233));
  NOT NOT1_2261(.VSS(VSS),.VDD(VDD),.Y(I29579),.A(g30565));
  NOT NOT1_2262(.VSS(VSS),.VDD(VDD),.Y(g28262),.A(I26785));
  NOT NOT1_2263(.VSS(VSS),.VDD(VDD),.Y(I24445),.A(g22923));
  NOT NOT1_2264(.VSS(VSS),.VDD(VDD),.Y(g20640),.A(g15426));
  NOT NOT1_2265(.VSS(VSS),.VDD(VDD),.Y(I17801),.A(g14936));
  NOT NOT1_2266(.VSS(VSS),.VDD(VDD),.Y(g20769),.A(g17955));
  NOT NOT1_2267(.VSS(VSS),.VDD(VDD),.Y(g17472),.A(g14656));
  NOT NOT1_2268(.VSS(VSS),.VDD(VDD),.Y(I26406),.A(g26187));
  NOT NOT1_2269(.VSS(VSS),.VDD(VDD),.Y(g12368),.A(I15208));
  NOT NOT1_2270(.VSS(VSS),.VDD(VDD),.Y(I16040),.A(g10430));
  NOT NOT1_2271(.VSS(VSS),.VDD(VDD),.Y(I20499),.A(g16224));
  NOT NOT1_2272(.VSS(VSS),.VDD(VDD),.Y(I12086),.A(g622));
  NOT NOT1_2273(.VSS(VSS),.VDD(VDD),.Y(g33670),.A(I31504));
  NOT NOT1_2274(.VSS(VSS),.VDD(VDD),.Y(I31727),.A(g33076));
  NOT NOT1_2275(.VSS(VSS),.VDD(VDD),.Y(g32873),.A(g30614));
  NOT NOT1_2276(.VSS(VSS),.VDD(VDD),.Y(g8046),.A(g528));
  NOT NOT1_2277(.VSS(VSS),.VDD(VDD),.Y(g25064),.A(I24228));
  NOT NOT1_2278(.VSS(VSS),.VDD(VDD),.Y(g16510),.A(g14008));
  NOT NOT1_2279(.VSS(VSS),.VDD(VDD),.Y(g19364),.A(g15825));
  NOT NOT1_2280(.VSS(VSS),.VDD(VDD),.Y(g20768),.A(g17955));
  NOT NOT1_2281(.VSS(VSS),.VDD(VDD),.Y(g28633),.A(g27687));
  NOT NOT1_2282(.VSS(VSS),.VDD(VDD),.Y(g8514),.A(g4258));
  NOT NOT1_2283(.VSS(VSS),.VDD(VDD),.Y(I19238),.A(g15079));
  NOT NOT1_2284(.VSS(VSS),.VDD(VDD),.Y(g34570),.A(g34392));
  NOT NOT1_2285(.VSS(VSS),.VDD(VDD),.Y(g34712),.A(I32868));
  NOT NOT1_2286(.VSS(VSS),.VDD(VDD),.Y(g21725),.A(I21294));
  NOT NOT1_2287(.VSS(VSS),.VDD(VDD),.Y(g11796),.A(g7985));
  NOT NOT1_2288(.VSS(VSS),.VDD(VDD),.Y(g16579),.A(g13267));
  NOT NOT1_2289(.VSS(VSS),.VDD(VDD),.Y(g33335),.A(I30861));
  NOT NOT1_2290(.VSS(VSS),.VDD(VDD),.Y(g8403),.A(I12568));
  NOT NOT1_2291(.VSS(VSS),.VDD(VDD),.Y(g23759),.A(I22886));
  NOT NOT1_2292(.VSS(VSS),.VDD(VDD),.Y(g13174),.A(g10741));
  NOT NOT1_2293(.VSS(VSS),.VDD(VDD),.Y(I21766),.A(g19620));
  NOT NOT1_2294(.VSS(VSS),.VDD(VDD),.Y(I17695),.A(g14330));
  NOT NOT1_2295(.VSS(VSS),.VDD(VDD),.Y(g26941),.A(I25689));
  NOT NOT1_2296(.VSS(VSS),.VDD(VDD),.Y(g34914),.A(I33134));
  NOT NOT1_2297(.VSS(VSS),.VDD(VDD),.Y(g31839),.A(g29385));
  NOT NOT1_2298(.VSS(VSS),.VDD(VDD),.Y(g33839),.A(I31686));
  NOT NOT1_2299(.VSS(VSS),.VDD(VDD),.Y(I32827),.A(g34477));
  NOT NOT1_2300(.VSS(VSS),.VDD(VDD),.Y(g8345),.A(g3794));
  NOT NOT1_2301(.VSS(VSS),.VDD(VDD),.Y(g8841),.A(I12823));
  NOT NOT1_2302(.VSS(VSS),.VDD(VDD),.Y(I14671),.A(g7717));
  NOT NOT1_2303(.VSS(VSS),.VDD(VDD),.Y(g7157),.A(g5706));
  NOT NOT1_2304(.VSS(VSS),.VDD(VDD),.Y(I12159),.A(g608));
  NOT NOT1_2305(.VSS(VSS),.VDD(VDD),.Y(g22147),.A(g18997));
  NOT NOT1_2306(.VSS(VSS),.VDD(VDD),.Y(g26519),.A(I25380));
  NOT NOT1_2307(.VSS(VSS),.VDD(VDD),.Y(g16578),.A(I17750));
  NOT NOT1_2308(.VSS(VSS),.VDD(VDD),.Y(g15569),.A(I17148));
  NOT NOT1_2309(.VSS(VSS),.VDD(VDD),.Y(g8763),.A(I12749));
  NOT NOT1_2310(.VSS(VSS),.VDD(VDD),.Y(I16564),.A(g10429));
  NOT NOT1_2311(.VSS(VSS),.VDD(VDD),.Y(g23435),.A(g18833));
  NOT NOT1_2312(.VSS(VSS),.VDD(VDD),.Y(g31667),.A(g30142));
  NOT NOT1_2313(.VSS(VSS),.VDD(VDD),.Y(g31838),.A(g29385));
  NOT NOT1_2314(.VSS(VSS),.VDD(VDD),.Y(g23082),.A(g21024));
  NOT NOT1_2315(.VSS(VSS),.VDD(VDD),.Y(g32834),.A(g31672));
  NOT NOT1_2316(.VSS(VSS),.VDD(VDD),.Y(g9839),.A(g2724));
  NOT NOT1_2317(.VSS(VSS),.VDD(VDD),.Y(g30074),.A(g29046));
  NOT NOT1_2318(.VSS(VSS),.VDD(VDD),.Y(g26518),.A(g25233));
  NOT NOT1_2319(.VSS(VSS),.VDD(VDD),.Y(g17591),.A(I18526));
  NOT NOT1_2320(.VSS(VSS),.VDD(VDD),.Y(g12896),.A(g10402));
  NOT NOT1_2321(.VSS(VSS),.VDD(VDD),.Y(g17776),.A(g14905));
  NOT NOT1_2322(.VSS(VSS),.VDD(VDD),.Y(g27011),.A(g25917));
  NOT NOT1_2323(.VSS(VSS),.VDD(VDD),.Y(I27561),.A(g28163));
  NOT NOT1_2324(.VSS(VSS),.VDD(VDD),.Y(g15568),.A(g14984));
  NOT NOT1_2325(.VSS(VSS),.VDD(VDD),.Y(g15747),.A(g13307));
  NOT NOT1_2326(.VSS(VSS),.VDD(VDD),.Y(g25009),.A(g22472));
  NOT NOT1_2327(.VSS(VSS),.VDD(VDD),.Y(I13723),.A(g3167));
  NOT NOT1_2328(.VSS(VSS),.VDD(VDD),.Y(I26004),.A(g26818));
  NOT NOT1_2329(.VSS(VSS),.VDD(VDD),.Y(I18868),.A(g14315));
  NOT NOT1_2330(.VSS(VSS),.VDD(VDD),.Y(I23360),.A(g23360));
  NOT NOT1_2331(.VSS(VSS),.VDD(VDD),.Y(g18945),.A(g16100));
  NOT NOT1_2332(.VSS(VSS),.VDD(VDD),.Y(g30567),.A(g29930));
  NOT NOT1_2333(.VSS(VSS),.VDD(VDD),.Y(I30962),.A(g32021));
  NOT NOT1_2334(.VSS(VSS),.VDD(VDD),.Y(g17147),.A(g14321));
  NOT NOT1_2335(.VSS(VSS),.VDD(VDD),.Y(g22858),.A(g20751));
  NOT NOT1_2336(.VSS(VSS),.VDD(VDD),.Y(g34594),.A(I32690));
  NOT NOT1_2337(.VSS(VSS),.VDD(VDD),.Y(I13149),.A(g6745));
  NOT NOT1_2338(.VSS(VSS),.VDD(VDD),.Y(g17754),.A(g14262));
  NOT NOT1_2339(.VSS(VSS),.VDD(VDD),.Y(I16847),.A(g6329));
  NOT NOT1_2340(.VSS(VSS),.VDD(VDD),.Y(g26935),.A(I25677));
  NOT NOT1_2341(.VSS(VSS),.VDD(VDD),.Y(g25008),.A(g22432));
  NOT NOT1_2342(.VSS(VSS),.VDD(VDD),.Y(g32542),.A(g31554));
  NOT NOT1_2343(.VSS(VSS),.VDD(VDD),.Y(g8107),.A(g3179));
  NOT NOT1_2344(.VSS(VSS),.VDD(VDD),.Y(I32803),.A(g34584));
  NOT NOT1_2345(.VSS(VSS),.VDD(VDD),.Y(I25399),.A(g24489));
  NOT NOT1_2346(.VSS(VSS),.VDD(VDD),.Y(g31487),.A(I29149));
  NOT NOT1_2347(.VSS(VSS),.VDD(VDD),.Y(g32021),.A(I29579));
  NOT NOT1_2348(.VSS(VSS),.VDD(VDD),.Y(g32453),.A(I29981));
  NOT NOT1_2349(.VSS(VSS),.VDD(VDD),.Y(I29720),.A(g30931));
  NOT NOT1_2350(.VSS(VSS),.VDD(VDD),.Y(g11192),.A(g8038));
  NOT NOT1_2351(.VSS(VSS),.VDD(VDD),.Y(g22151),.A(I21734));
  NOT NOT1_2352(.VSS(VSS),.VDD(VDD),.Y(I11620),.A(g1));
  NOT NOT1_2353(.VSS(VSS),.VDD(VDD),.Y(I21162),.A(g17292));
  NOT NOT1_2354(.VSS(VSS),.VDD(VDD),.Y(I12144),.A(g554));
  NOT NOT1_2355(.VSS(VSS),.VDD(VDD),.Y(I12823),.A(g4311));
  NOT NOT1_2356(.VSS(VSS),.VDD(VDD),.Y(I18709),.A(g6668));
  NOT NOT1_2357(.VSS(VSS),.VDD(VDD),.Y(g20662),.A(g15171));
  NOT NOT1_2358(.VSS(VSS),.VDD(VDD),.Y(g21399),.A(g15224));
  NOT NOT1_2359(.VSS(VSS),.VDD(VDD),.Y(g23849),.A(g19277));
  NOT NOT1_2360(.VSS(VSS),.VDD(VDD),.Y(g22996),.A(g20330));
  NOT NOT1_2361(.VSS(VSS),.VDD(VDD),.Y(g23940),.A(g19074));
  NOT NOT1_2362(.VSS(VSS),.VDD(VDD),.Y(g25892),.A(g24528));
  NOT NOT1_2363(.VSS(VSS),.VDD(VDD),.Y(I20753),.A(g16677));
  NOT NOT1_2364(.VSS(VSS),.VDD(VDD),.Y(I15663),.A(g5308));
  NOT NOT1_2365(.VSS(VSS),.VDD(VDD),.Y(g23399),.A(g21514));
  NOT NOT1_2366(.VSS(VSS),.VDD(VDD),.Y(g32726),.A(g31672));
  NOT NOT1_2367(.VSS(VSS),.VDD(VDD),.Y(g32913),.A(g30825));
  NOT NOT1_2368(.VSS(VSS),.VDD(VDD),.Y(g24027),.A(g20014));
  NOT NOT1_2369(.VSS(VSS),.VDD(VDD),.Y(I18259),.A(g12946));
  NOT NOT1_2370(.VSS(VSS),.VDD(VDD),.Y(g9618),.A(g5794));
  NOT NOT1_2371(.VSS(VSS),.VDD(VDD),.Y(g11663),.A(g6905));
  NOT NOT1_2372(.VSS(VSS),.VDD(VDD),.Y(g16615),.A(I17801));
  NOT NOT1_2373(.VSS(VSS),.VDD(VDD),.Y(g22844),.A(g21163));
  NOT NOT1_2374(.VSS(VSS),.VDD(VDD),.Y(g13522),.A(g10981));
  NOT NOT1_2375(.VSS(VSS),.VDD(VDD),.Y(g34941),.A(g34926));
  NOT NOT1_2376(.VSS(VSS),.VDD(VDD),.Y(g13663),.A(g10971));
  NOT NOT1_2377(.VSS(VSS),.VDD(VDD),.Y(g21398),.A(g18008));
  NOT NOT1_2378(.VSS(VSS),.VDD(VDD),.Y(g23848),.A(g19210));
  NOT NOT1_2379(.VSS(VSS),.VDD(VDD),.Y(g25555),.A(g22550));
  NOT NOT1_2380(.VSS(VSS),.VDD(VDD),.Y(g32614),.A(g31542));
  NOT NOT1_2381(.VSS(VSS),.VDD(VDD),.Y(g7626),.A(I12112));
  NOT NOT1_2382(.VSS(VSS),.VDD(VDD),.Y(I12336),.A(g52));
  NOT NOT1_2383(.VSS(VSS),.VDD(VDD),.Y(g23398),.A(g21468));
  NOT NOT1_2384(.VSS(VSS),.VDD(VDD),.Y(I32881),.A(g34688));
  NOT NOT1_2385(.VSS(VSS),.VDD(VDD),.Y(g8858),.A(g671));
  NOT NOT1_2386(.VSS(VSS),.VDD(VDD),.Y(g33443),.A(I30971));
  NOT NOT1_2387(.VSS(VSS),.VDD(VDD),.Y(g16720),.A(g14234));
  NOT NOT1_2388(.VSS(VSS),.VDD(VDD),.Y(g9282),.A(g723));
  NOT NOT1_2389(.VSS(VSS),.VDD(VDD),.Y(g34675),.A(I32809));
  NOT NOT1_2390(.VSS(VSS),.VDD(VDD),.Y(I20650),.A(g17010));
  NOT NOT1_2391(.VSS(VSS),.VDD(VDD),.Y(g23652),.A(I22785));
  NOT NOT1_2392(.VSS(VSS),.VDD(VDD),.Y(g32607),.A(g31542));
  NOT NOT1_2393(.VSS(VSS),.VDD(VDD),.Y(g8016),.A(g3391));
  NOT NOT1_2394(.VSS(VSS),.VDD(VDD),.Y(g10981),.A(I14119));
  NOT NOT1_2395(.VSS(VSS),.VDD(VDD),.Y(g8757),.A(I12746));
  NOT NOT1_2396(.VSS(VSS),.VDD(VDD),.Y(g32905),.A(g30825));
  NOT NOT1_2397(.VSS(VSS),.VDD(VDD),.Y(g14563),.A(I16676));
  NOT NOT1_2398(.VSS(VSS),.VDD(VDD),.Y(g8416),.A(I12580));
  NOT NOT1_2399(.VSS(VSS),.VDD(VDD),.Y(g27112),.A(g26793));
  NOT NOT1_2400(.VSS(VSS),.VDD(VDD),.Y(g20710),.A(g15509));
  NOT NOT1_2401(.VSS(VSS),.VDD(VDD),.Y(g16746),.A(g14258));
  NOT NOT1_2402(.VSS(VSS),.VDD(VDD),.Y(I20529),.A(g16309));
  NOT NOT1_2403(.VSS(VSS),.VDD(VDD),.Y(I21911),.A(g21278));
  NOT NOT1_2404(.VSS(VSS),.VDD(VDD),.Y(g17844),.A(I18832));
  NOT NOT1_2405(.VSS(VSS),.VDD(VDD),.Y(g20552),.A(g17847));
  NOT NOT1_2406(.VSS(VSS),.VDD(VDD),.Y(g32530),.A(g30825));
  NOT NOT1_2407(.VSS(VSS),.VDD(VDD),.Y(g9693),.A(g1886));
  NOT NOT1_2408(.VSS(VSS),.VDD(VDD),.Y(g13483),.A(g11270));
  NOT NOT1_2409(.VSS(VSS),.VDD(VDD),.Y(I33264),.A(g34978));
  NOT NOT1_2410(.VSS(VSS),.VDD(VDD),.Y(I15862),.A(g11215));
  NOT NOT1_2411(.VSS(VSS),.VDD(VDD),.Y(g17367),.A(I18320));
  NOT NOT1_2412(.VSS(VSS),.VDD(VDD),.Y(g32593),.A(g31542));
  NOT NOT1_2413(.VSS(VSS),.VDD(VDD),.Y(g18932),.A(g16136));
  NOT NOT1_2414(.VSS(VSS),.VDD(VDD),.Y(g6985),.A(g4669));
  NOT NOT1_2415(.VSS(VSS),.VDD(VDD),.Y(I33137),.A(g34884));
  NOT NOT1_2416(.VSS(VSS),.VDD(VDD),.Y(g20204),.A(g16578));
  NOT NOT1_2417(.VSS(VSS),.VDD(VDD),.Y(g19687),.A(g17096));
  NOT NOT1_2418(.VSS(VSS),.VDD(VDD),.Y(I21246),.A(g16540));
  NOT NOT1_2419(.VSS(VSS),.VDD(VDD),.Y(g24003),.A(g21514));
  NOT NOT1_2420(.VSS(VSS),.VDD(VDD),.Y(g23263),.A(I22366));
  NOT NOT1_2421(.VSS(VSS),.VDD(VDD),.Y(I12631),.A(g1242));
  NOT NOT1_2422(.VSS(VSS),.VDD(VDD),.Y(g8522),.A(g298));
  NOT NOT1_2423(.VSS(VSS),.VDD(VDD),.Y(g20779),.A(g15509));
  NOT NOT1_2424(.VSS(VSS),.VDD(VDD),.Y(g22319),.A(I21831));
  NOT NOT1_2425(.VSS(VSS),.VDD(VDD),.Y(g12378),.A(g9417));
  NOT NOT1_2426(.VSS(VSS),.VDD(VDD),.Y(g34935),.A(I33189));
  NOT NOT1_2427(.VSS(VSS),.VDD(VDD),.Y(g23332),.A(g20785));
  NOT NOT1_2428(.VSS(VSS),.VDD(VDD),.Y(g32565),.A(g30735));
  NOT NOT1_2429(.VSS(VSS),.VDD(VDD),.Y(g32464),.A(g30735));
  NOT NOT1_2430(.VSS(VSS),.VDD(VDD),.Y(g25239),.A(g23972));
  NOT NOT1_2431(.VSS(VSS),.VDD(VDD),.Y(g19954),.A(g16540));
  NOT NOT1_2432(.VSS(VSS),.VDD(VDD),.Y(g11949),.A(I14773));
  NOT NOT1_2433(.VSS(VSS),.VDD(VDD),.Y(I24393),.A(g23453));
  NOT NOT1_2434(.VSS(VSS),.VDD(VDD),.Y(g19374),.A(g16047));
  NOT NOT1_2435(.VSS(VSS),.VDD(VDD),.Y(g20778),.A(g15224));
  NOT NOT1_2436(.VSS(VSS),.VDD(VDD),.Y(g34883),.A(g34852));
  NOT NOT1_2437(.VSS(VSS),.VDD(VDD),.Y(g10794),.A(g8470));
  NOT NOT1_2438(.VSS(VSS),.VDD(VDD),.Y(g9555),.A(I13206));
  NOT NOT1_2439(.VSS(VSS),.VDD(VDD),.Y(g18897),.A(g15509));
  NOT NOT1_2440(.VSS(VSS),.VDD(VDD),.Y(I15536),.A(g1227));
  NOT NOT1_2441(.VSS(VSS),.VDD(VDD),.Y(g10395),.A(g6995));
  NOT NOT1_2442(.VSS(VSS),.VDD(VDD),.Y(g22227),.A(g19801));
  NOT NOT1_2443(.VSS(VSS),.VDD(VDD),.Y(g24778),.A(g23286));
  NOT NOT1_2444(.VSS(VSS),.VDD(VDD),.Y(g9804),.A(g5456));
  NOT NOT1_2445(.VSS(VSS),.VDD(VDD),.Y(g10262),.A(g586));
  NOT NOT1_2446(.VSS(VSS),.VDD(VDD),.Y(g24081),.A(g21209));
  NOT NOT1_2447(.VSS(VSS),.VDD(VDD),.Y(g21406),.A(g17955));
  NOT NOT1_2448(.VSS(VSS),.VDD(VDD),.Y(g16684),.A(g14223));
  NOT NOT1_2449(.VSS(VSS),.VDD(VDD),.Y(g11948),.A(g10224));
  NOT NOT1_2450(.VSS(VSS),.VDD(VDD),.Y(I21776),.A(g21308));
  NOT NOT1_2451(.VSS(VSS),.VDD(VDD),.Y(I15702),.A(g12217));
  NOT NOT1_2452(.VSS(VSS),.VDD(VDD),.Y(g14262),.A(g10838));
  NOT NOT1_2453(.VSS(VSS),.VDD(VDD),.Y(g12944),.A(g12659));
  NOT NOT1_2454(.VSS(VSS),.VDD(VDD),.Y(I18810),.A(g13716));
  NOT NOT1_2455(.VSS(VSS),.VDD(VDD),.Y(g23406),.A(g20330));
  NOT NOT1_2456(.VSS(VSS),.VDD(VDD),.Y(g9792),.A(g5401));
  NOT NOT1_2457(.VSS(VSS),.VDD(VDD),.Y(g32641),.A(g30614));
  NOT NOT1_2458(.VSS(VSS),.VDD(VDD),.Y(g6832),.A(I11665));
  NOT NOT1_2459(.VSS(VSS),.VDD(VDD),.Y(g32797),.A(g30825));
  NOT NOT1_2460(.VSS(VSS),.VDD(VDD),.Y(g23962),.A(g19147));
  NOT NOT1_2461(.VSS(VSS),.VDD(VDD),.Y(g31815),.A(g29385));
  NOT NOT1_2462(.VSS(VSS),.VDD(VDD),.Y(g23361),.A(I22464));
  NOT NOT1_2463(.VSS(VSS),.VDD(VDD),.Y(g28032),.A(g26365));
  NOT NOT1_2464(.VSS(VSS),.VDD(VDD),.Y(I32482),.A(g34304));
  NOT NOT1_2465(.VSS(VSS),.VDD(VDD),.Y(g11702),.A(g6928));
  NOT NOT1_2466(.VSS(VSS),.VDD(VDD),.Y(g7778),.A(g1339));
  NOT NOT1_2467(.VSS(VSS),.VDD(VDD),.Y(g15579),.A(I17159));
  NOT NOT1_2468(.VSS(VSS),.VDD(VDD),.Y(g31601),.A(I29207));
  NOT NOT1_2469(.VSS(VSS),.VDD(VDD),.Y(g8654),.A(g1087));
  NOT NOT1_2470(.VSS(VSS),.VDD(VDD),.Y(I16452),.A(g11182));
  NOT NOT1_2471(.VSS(VSS),.VDD(VDD),.Y(I18879),.A(g13267));
  NOT NOT1_2472(.VSS(VSS),.VDD(VDD),.Y(g9621),.A(g6423));
  NOT NOT1_2473(.VSS(VSS),.VDD(VDD),.Y(g10191),.A(g6386));
  NOT NOT1_2474(.VSS(VSS),.VDD(VDD),.Y(g23500),.A(g20924));
  NOT NOT1_2475(.VSS(VSS),.VDD(VDD),.Y(g24356),.A(g22594));
  NOT NOT1_2476(.VSS(VSS),.VDD(VDD),.Y(g13621),.A(g10573));
  NOT NOT1_2477(.VSS(VSS),.VDD(VDD),.Y(g21049),.A(g17433));
  NOT NOT1_2478(.VSS(VSS),.VDD(VDD),.Y(I11896),.A(g4446));
  NOT NOT1_2479(.VSS(VSS),.VDD(VDD),.Y(g25185),.A(g22228));
  NOT NOT1_2480(.VSS(VSS),.VDD(VDD),.Y(g17059),.A(I18151));
  NOT NOT1_2481(.VSS(VSS),.VDD(VDD),.Y(g20380),.A(g17955));
  NOT NOT1_2482(.VSS(VSS),.VDD(VDD),.Y(g26083),.A(g24809));
  NOT NOT1_2483(.VSS(VSS),.VDD(VDD),.Y(g14191),.A(g12381));
  NOT NOT1_2484(.VSS(VSS),.VDD(VDD),.Y(g30729),.A(I28883));
  NOT NOT1_2485(.VSS(VSS),.VDD(VDD),.Y(I15564),.A(g11949));
  NOT NOT1_2486(.VSS(VSS),.VDD(VDD),.Y(g25092),.A(g23666));
  NOT NOT1_2487(.VSS(VSS),.VDD(VDD),.Y(g24999),.A(g23626));
  NOT NOT1_2488(.VSS(VSS),.VDD(VDD),.Y(g26284),.A(g24875));
  NOT NOT1_2489(.VSS(VSS),.VDD(VDD),.Y(I18337),.A(g1422));
  NOT NOT1_2490(.VSS(VSS),.VDD(VDD),.Y(g34501),.A(g34400));
  NOT NOT1_2491(.VSS(VSS),.VDD(VDD),.Y(g27730),.A(g26424));
  NOT NOT1_2492(.VSS(VSS),.VDD(VDD),.Y(g10521),.A(I13889));
  NOT NOT1_2493(.VSS(VSS),.VDD(VDD),.Y(g12857),.A(I15474));
  NOT NOT1_2494(.VSS(VSS),.VDD(VDD),.Y(I19348),.A(g15084));
  NOT NOT1_2495(.VSS(VSS),.VDD(VDD),.Y(g21048),.A(g17533));
  NOT NOT1_2496(.VSS(VSS),.VDD(VDD),.Y(g25154),.A(g22457));
  NOT NOT1_2497(.VSS(VSS),.VDD(VDD),.Y(g20090),.A(g17433));
  NOT NOT1_2498(.VSS(VSS),.VDD(VDD),.Y(g17058),.A(I18148));
  NOT NOT1_2499(.VSS(VSS),.VDD(VDD),.Y(g32635),.A(g31542));
  NOT NOT1_2500(.VSS(VSS),.VDD(VDD),.Y(g8880),.A(I12861));
  NOT NOT1_2501(.VSS(VSS),.VDD(VDD),.Y(g31937),.A(g30991));
  NOT NOT1_2502(.VSS(VSS),.VDD(VDD),.Y(g8595),.A(I12666));
  NOT NOT1_2503(.VSS(VSS),.VDD(VDD),.Y(g24090),.A(g19935));
  NOT NOT1_2504(.VSS(VSS),.VDD(VDD),.Y(g19489),.A(g16449));
  NOT NOT1_2505(.VSS(VSS),.VDD(VDD),.Y(g20233),.A(g17873));
  NOT NOT1_2506(.VSS(VSS),.VDD(VDD),.Y(g33937),.A(I31823));
  NOT NOT1_2507(.VSS(VSS),.VDD(VDD),.Y(g12793),.A(g10287));
  NOT NOT1_2508(.VSS(VSS),.VDD(VDD),.Y(I11716),.A(g4054));
  NOT NOT1_2509(.VSS(VSS),.VDD(VDD),.Y(g20182),.A(g16897));
  NOT NOT1_2510(.VSS(VSS),.VDD(VDD),.Y(g20651),.A(g15483));
  NOT NOT1_2511(.VSS(VSS),.VDD(VDD),.Y(g20672),.A(g15277));
  NOT NOT1_2512(.VSS(VSS),.VDD(VDD),.Y(I17876),.A(g13070));
  NOT NOT1_2513(.VSS(VSS),.VDD(VDD),.Y(g23004),.A(g20283));
  NOT NOT1_2514(.VSS(VSS),.VDD(VDD),.Y(I27495),.A(g27961));
  NOT NOT1_2515(.VSS(VSS),.VDD(VDD),.Y(g7475),.A(g896));
  NOT NOT1_2516(.VSS(VSS),.VDD(VDD),.Y(g21221),.A(g15680));
  NOT NOT1_2517(.VSS(VSS),.VDD(VDD),.Y(g24182),.A(I23390));
  NOT NOT1_2518(.VSS(VSS),.VDD(VDD),.Y(g19559),.A(g16129));
  NOT NOT1_2519(.VSS(VSS),.VDD(VDD),.Y(g23221),.A(g20785));
  NOT NOT1_2520(.VSS(VSS),.VDD(VDD),.Y(I14644),.A(g7717));
  NOT NOT1_2521(.VSS(VSS),.VDD(VDD),.Y(g11183),.A(g8135));
  NOT NOT1_2522(.VSS(VSS),.VDD(VDD),.Y(g29942),.A(g28867));
  NOT NOT1_2523(.VSS(VSS),.VDD(VDD),.Y(g22957),.A(I22143));
  NOT NOT1_2524(.VSS(VSS),.VDD(VDD),.Y(g31791),.A(I29363));
  NOT NOT1_2525(.VSS(VSS),.VDD(VDD),.Y(g7627),.A(g4311));
  NOT NOT1_2526(.VSS(VSS),.VDD(VDD),.Y(g19558),.A(g15938));
  NOT NOT1_2527(.VSS(VSS),.VDD(VDD),.Y(g6905),.A(I11708));
  NOT NOT1_2528(.VSS(VSS),.VDD(VDD),.Y(g16523),.A(g14041));
  NOT NOT1_2529(.VSS(VSS),.VDD(VDD),.Y(g8612),.A(g2775));
  NOT NOT1_2530(.VSS(VSS),.VDD(VDD),.Y(g23613),.A(I22748));
  NOT NOT1_2531(.VSS(VSS),.VDD(VDD),.Y(g9518),.A(g6219));
  NOT NOT1_2532(.VSS(VSS),.VDD(VDD),.Y(g15615),.A(I17181));
  NOT NOT1_2533(.VSS(VSS),.VDD(VDD),.Y(I17763),.A(g13191));
  NOT NOT1_2534(.VSS(VSS),.VDD(VDD),.Y(I31607),.A(g33164));
  NOT NOT1_2535(.VSS(VSS),.VDD(VDD),.Y(g13062),.A(g10981));
  NOT NOT1_2536(.VSS(VSS),.VDD(VDD),.Y(g7526),.A(I12013));
  NOT NOT1_2537(.VSS(VSS),.VDD(VDD),.Y(g7998),.A(g392));
  NOT NOT1_2538(.VSS(VSS),.VDD(VDD),.Y(g11509),.A(g7632));
  NOT NOT1_2539(.VSS(VSS),.VDD(VDD),.Y(g22146),.A(g18997));
  NOT NOT1_2540(.VSS(VSS),.VDD(VDD),.Y(g26653),.A(g25337));
  NOT NOT1_2541(.VSS(VSS),.VDD(VDD),.Y(g20513),.A(g18065));
  NOT NOT1_2542(.VSS(VSS),.VDD(VDD),.Y(g17301),.A(g14454));
  NOT NOT1_2543(.VSS(VSS),.VDD(VDD),.Y(g20449),.A(g15277));
  NOT NOT1_2544(.VSS(VSS),.VDD(VDD),.Y(g28162),.A(I26679));
  NOT NOT1_2545(.VSS(VSS),.VDD(VDD),.Y(g10389),.A(g6986));
  NOT NOT1_2546(.VSS(VSS),.VDD(VDD),.Y(g32891),.A(g30825));
  NOT NOT1_2547(.VSS(VSS),.VDD(VDD),.Y(I15872),.A(g11236));
  NOT NOT1_2548(.VSS(VSS),.VDD(VDD),.Y(g13933),.A(g11419));
  NOT NOT1_2549(.VSS(VSS),.VDD(VDD),.Y(g23947),.A(g19210));
  NOT NOT1_2550(.VSS(VSS),.VDD(VDD),.Y(g31479),.A(I29139));
  NOT NOT1_2551(.VSS(VSS),.VDD(VDD),.Y(g31666),.A(I29248));
  NOT NOT1_2552(.VSS(VSS),.VDD(VDD),.Y(I27954),.A(g28803));
  NOT NOT1_2553(.VSS(VSS),.VDD(VDD),.Y(g18097),.A(I18897));
  NOT NOT1_2554(.VSS(VSS),.VDD(VDD),.Y(g21273),.A(I21006));
  NOT NOT1_2555(.VSS(VSS),.VDD(VDD),.Y(g17120),.A(g14262));
  NOT NOT1_2556(.VSS(VSS),.VDD(VDD),.Y(g19544),.A(g16349));
  NOT NOT1_2557(.VSS(VSS),.VDD(VDD),.Y(g23273),.A(g21070));
  NOT NOT1_2558(.VSS(VSS),.VDD(VDD),.Y(g19865),.A(g15885));
  NOT NOT1_2559(.VSS(VSS),.VDD(VDD),.Y(g17739),.A(I18728));
  NOT NOT1_2560(.VSS(VSS),.VDD(VDD),.Y(g10612),.A(g10233));
  NOT NOT1_2561(.VSS(VSS),.VDD(VDD),.Y(g11872),.A(I14684));
  NOT NOT1_2562(.VSS(VSS),.VDD(VDD),.Y(g23605),.A(g20739));
  NOT NOT1_2563(.VSS(VSS),.VDD(VDD),.Y(g9776),.A(g5073));
  NOT NOT1_2564(.VSS(VSS),.VDD(VDD),.Y(g10099),.A(g6682));
  NOT NOT1_2565(.VSS(VSS),.VDD(VDD),.Y(g15746),.A(g13121));
  NOT NOT1_2566(.VSS(VSS),.VDD(VDD),.Y(g16475),.A(g14107));
  NOT NOT1_2567(.VSS(VSS),.VDD(VDD),.Y(g20448),.A(g15509));
  NOT NOT1_2568(.VSS(VSS),.VDD(VDD),.Y(g34304),.A(I32309));
  NOT NOT1_2569(.VSS(VSS),.VDD(VDD),.Y(I12954),.A(g4358));
  NOT NOT1_2570(.VSS(VSS),.VDD(VDD),.Y(g10388),.A(g6983));
  NOT NOT1_2571(.VSS(VSS),.VDD(VDD),.Y(I32651),.A(g34375));
  NOT NOT1_2572(.VSS(VSS),.VDD(VDD),.Y(g32575),.A(g31170));
  NOT NOT1_2573(.VSS(VSS),.VDD(VDD),.Y(g32474),.A(g31194));
  NOT NOT1_2574(.VSS(VSS),.VDD(VDD),.Y(g19713),.A(g16816));
  NOT NOT1_2575(.VSS(VSS),.VDD(VDD),.Y(g7439),.A(g6351));
  NOT NOT1_2576(.VSS(VSS),.VDD(VDD),.Y(g29930),.A(I28162));
  NOT NOT1_2577(.VSS(VSS),.VDD(VDD),.Y(g22698),.A(I22009));
  NOT NOT1_2578(.VSS(VSS),.VDD(VDD),.Y(g29993),.A(g29018));
  NOT NOT1_2579(.VSS(VSS),.VDD(VDD),.Y(g16727),.A(g14454));
  NOT NOT1_2580(.VSS(VSS),.VDD(VDD),.Y(g17738),.A(g14813));
  NOT NOT1_2581(.VSS(VSS),.VDD(VDD),.Y(g17645),.A(g15018));
  NOT NOT1_2582(.VSS(VSS),.VDD(VDD),.Y(g20505),.A(g15426));
  NOT NOT1_2583(.VSS(VSS),.VDD(VDD),.Y(g21463),.A(g15588));
  NOT NOT1_2584(.VSS(VSS),.VDD(VDD),.Y(g23812),.A(g18997));
  NOT NOT1_2585(.VSS(VSS),.VDD(VDD),.Y(g32711),.A(g31070));
  NOT NOT1_2586(.VSS(VSS),.VDD(VDD),.Y(g8130),.A(g4515));
  NOT NOT1_2587(.VSS(VSS),.VDD(VDD),.Y(g14701),.A(g12351));
  NOT NOT1_2588(.VSS(VSS),.VDD(VDD),.Y(I17456),.A(g13680));
  NOT NOT1_2589(.VSS(VSS),.VDD(VDD),.Y(I23318),.A(g21689));
  NOT NOT1_2590(.VSS(VSS),.VDD(VDD),.Y(g8542),.A(I12644));
  NOT NOT1_2591(.VSS(VSS),.VDD(VDD),.Y(g24505),.A(g22689));
  NOT NOT1_2592(.VSS(VSS),.VDD(VDD),.Y(g8330),.A(g2587));
  NOT NOT1_2593(.VSS(VSS),.VDD(VDD),.Y(g24404),.A(g22908));
  NOT NOT1_2594(.VSS(VSS),.VDD(VDD),.Y(g10272),.A(I13705));
  NOT NOT1_2595(.VSS(VSS),.VDD(VDD),.Y(g9965),.A(g127));
  NOT NOT1_2596(.VSS(VSS),.VDD(VDD),.Y(g29965),.A(g28903));
  NOT NOT1_2597(.VSS(VSS),.VDD(VDD),.Y(I33034),.A(g34769));
  NOT NOT1_2598(.VSS(VSS),.VDD(VDD),.Y(g14251),.A(g12308));
  NOT NOT1_2599(.VSS(VSS),.VDD(VDD),.Y(I17916),.A(g13087));
  NOT NOT1_2600(.VSS(VSS),.VDD(VDD),.Y(g20026),.A(g17271));
  NOT NOT1_2601(.VSS(VSS),.VDD(VDD),.Y(g32537),.A(g30825));
  NOT NOT1_2602(.VSS(VSS),.VDD(VDD),.Y(I18078),.A(g13350));
  NOT NOT1_2603(.VSS(VSS),.VDD(VDD),.Y(g20212),.A(g17194));
  NOT NOT1_2604(.VSS(VSS),.VDD(VDD),.Y(g23234),.A(g20375));
  NOT NOT1_2605(.VSS(VSS),.VDD(VDD),.Y(g24026),.A(g19919));
  NOT NOT1_2606(.VSS(VSS),.VDD(VDD),.Y(g9264),.A(g5396));
  NOT NOT1_2607(.VSS(VSS),.VDD(VDD),.Y(g15806),.A(I17302));
  NOT NOT1_2608(.VSS(VSS),.VDD(VDD),.Y(I21058),.A(g17747));
  NOT NOT1_2609(.VSS(VSS),.VDD(VDD),.Y(g25438),.A(g22763));
  NOT NOT1_2610(.VSS(VSS),.VDD(VDD),.Y(g6973),.A(I11743));
  NOT NOT1_2611(.VSS(VSS),.VDD(VDD),.Y(I17314),.A(g14078));
  NOT NOT1_2612(.VSS(VSS),.VDD(VDD),.Y(I32449),.A(g34127));
  NOT NOT1_2613(.VSS(VSS),.VDD(VDD),.Y(g19679),.A(g16782));
  NOT NOT1_2614(.VSS(VSS),.VDD(VDD),.Y(I18086),.A(g13856));
  NOT NOT1_2615(.VSS(VSS),.VDD(VDD),.Y(g27245),.A(g26209));
  NOT NOT1_2616(.VSS(VSS),.VDD(VDD),.Y(g34653),.A(I32763));
  NOT NOT1_2617(.VSS(VSS),.VDD(VDD),.Y(g9360),.A(g3372));
  NOT NOT1_2618(.VSS(VSS),.VDD(VDD),.Y(g9933),.A(g5759));
  NOT NOT1_2619(.VSS(VSS),.VDD(VDD),.Y(g32606),.A(g30673));
  NOT NOT1_2620(.VSS(VSS),.VDD(VDD),.Y(g10032),.A(g562));
  NOT NOT1_2621(.VSS(VSS),.VDD(VDD),.Y(I29236),.A(g29498));
  NOT NOT1_2622(.VSS(VSS),.VDD(VDD),.Y(g32492),.A(g31376));
  NOT NOT1_2623(.VSS(VSS),.VDD(VDD),.Y(g19678),.A(g16752));
  NOT NOT1_2624(.VSS(VSS),.VDD(VDD),.Y(I15205),.A(g10139));
  NOT NOT1_2625(.VSS(VSS),.VDD(VDD),.Y(g14032),.A(g11048));
  NOT NOT1_2626(.VSS(VSS),.VDD(VDD),.Y(g10140),.A(g19));
  NOT NOT1_2627(.VSS(VSS),.VDD(VDD),.Y(g29210),.A(I27546));
  NOT NOT1_2628(.VSS(VSS),.VDD(VDD),.Y(g9050),.A(g1087));
  NOT NOT1_2629(.VSS(VSS),.VDD(VDD),.Y(g17427),.A(I18364));
  NOT NOT1_2630(.VSS(VSS),.VDD(VDD),.Y(I13802),.A(g6971));
  NOT NOT1_2631(.VSS(VSS),.VDD(VDD),.Y(g13574),.A(I16024));
  NOT NOT1_2632(.VSS(VSS),.VDD(VDD),.Y(I25514),.A(g25073));
  NOT NOT1_2633(.VSS(VSS),.VDD(VDD),.Y(I13857),.A(g9780));
  NOT NOT1_2634(.VSS(VSS),.VDD(VDD),.Y(g17366),.A(g14454));
  NOT NOT1_2635(.VSS(VSS),.VDD(VDD),.Y(g7952),.A(g3774));
  NOT NOT1_2636(.VSS(VSS),.VDD(VDD),.Y(g25083),.A(g23782));
  NOT NOT1_2637(.VSS(VSS),.VDD(VDD),.Y(g25348),.A(g22763));
  NOT NOT1_2638(.VSS(VSS),.VDD(VDD),.Y(g9450),.A(g5817));
  NOT NOT1_2639(.VSS(VSS),.VDD(VDD),.Y(I14450),.A(g4191));
  NOT NOT1_2640(.VSS(VSS),.VDD(VDD),.Y(g16600),.A(I17780));
  NOT NOT1_2641(.VSS(VSS),.VDD(VDD),.Y(g19686),.A(g17062));
  NOT NOT1_2642(.VSS(VSS),.VDD(VDD),.Y(g25284),.A(I24474));
  NOT NOT1_2643(.VSS(VSS),.VDD(VDD),.Y(g21514),.A(I21189));
  NOT NOT1_2644(.VSS(VSS),.VDD(VDD),.Y(I11793),.A(g6049));
  NOT NOT1_2645(.VSS(VSS),.VDD(VDD),.Y(g11912),.A(g8989));
  NOT NOT1_2646(.VSS(VSS),.VDD(VDD),.Y(g26576),.A(I25399));
  NOT NOT1_2647(.VSS(VSS),.VDD(VDD),.Y(I26682),.A(g27774));
  NOT NOT1_2648(.VSS(VSS),.VDD(VDD),.Y(g28147),.A(I26654));
  NOT NOT1_2649(.VSS(VSS),.VDD(VDD),.Y(I27558),.A(g28155));
  NOT NOT1_2650(.VSS(VSS),.VDD(VDD),.Y(g32750),.A(g30937));
  NOT NOT1_2651(.VSS(VSS),.VDD(VDD),.Y(I12016),.A(g772));
  NOT NOT1_2652(.VSS(VSS),.VDD(VDD),.Y(I18125),.A(g13191));
  NOT NOT1_2653(.VSS(VSS),.VDD(VDD),.Y(g10061),.A(I13581));
  NOT NOT1_2654(.VSS(VSS),.VDD(VDD),.Y(g13311),.A(I15878));
  NOT NOT1_2655(.VSS(VSS),.VDD(VDD),.Y(g28754),.A(I27238));
  NOT NOT1_2656(.VSS(VSS),.VDD(VDD),.Y(g32381),.A(I29909));
  NOT NOT1_2657(.VSS(VSS),.VDD(VDD),.Y(g7616),.A(I12086));
  NOT NOT1_2658(.VSS(VSS),.VDD(VDD),.Y(I19484),.A(g15122));
  NOT NOT1_2659(.VSS(VSS),.VDD(VDD),.Y(g23507),.A(g21562));
  NOT NOT1_2660(.VSS(VSS),.VDD(VDD),.Y(g34852),.A(g34845));
  NOT NOT1_2661(.VSS(VSS),.VDD(VDD),.Y(g20433),.A(g17929));
  NOT NOT1_2662(.VSS(VSS),.VDD(VDD),.Y(g25566),.A(g22550));
  NOT NOT1_2663(.VSS(VSS),.VDD(VDD),.Y(g18896),.A(g16031));
  NOT NOT1_2664(.VSS(VSS),.VDD(VDD),.Y(g24149),.A(g19338));
  NOT NOT1_2665(.VSS(VSS),.VDD(VDD),.Y(g20387),.A(g15426));
  NOT NOT1_2666(.VSS(VSS),.VDD(VDD),.Y(g28370),.A(g27528));
  NOT NOT1_2667(.VSS(VSS),.VDD(VDD),.Y(I28866),.A(g29730));
  NOT NOT1_2668(.VSS(VSS),.VDD(VDD),.Y(I22180),.A(g21366));
  NOT NOT1_2669(.VSS(VSS),.VDD(VDD),.Y(g16821),.A(I18031));
  NOT NOT1_2670(.VSS(VSS),.VDD(VDD),.Y(g21421),.A(g15171));
  NOT NOT1_2671(.VSS(VSS),.VDD(VDD),.Y(g27737),.A(g26718));
  NOT NOT1_2672(.VSS(VSS),.VDD(VDD),.Y(I12893),.A(g4226));
  NOT NOT1_2673(.VSS(VSS),.VDD(VDD),.Y(g7004),.A(I11777));
  NOT NOT1_2674(.VSS(VSS),.VDD(VDD),.Y(g9379),.A(g5424));
  NOT NOT1_2675(.VSS(VSS),.VDD(VDD),.Y(g23421),.A(g21562));
  NOT NOT1_2676(.VSS(VSS),.VDD(VDD),.Y(g13051),.A(g11964));
  NOT NOT1_2677(.VSS(VSS),.VDD(VDD),.Y(g20097),.A(g17691));
  NOT NOT1_2678(.VSS(VSS),.VDD(VDD),.Y(g32796),.A(g31376));
  NOT NOT1_2679(.VSS(VSS),.VDD(VDD),.Y(g7527),.A(I12016));
  NOT NOT1_2680(.VSS(VSS),.VDD(VDD),.Y(I33164),.A(g34894));
  NOT NOT1_2681(.VSS(VSS),.VDD(VDD),.Y(g24097),.A(g19935));
  NOT NOT1_2682(.VSS(VSS),.VDD(VDD),.Y(g26608),.A(g25334));
  NOT NOT1_2683(.VSS(VSS),.VDD(VDD),.Y(g11592),.A(I14537));
  NOT NOT1_2684(.VSS(VSS),.VDD(VDD),.Y(g20104),.A(g17433));
  NOT NOT1_2685(.VSS(VSS),.VDD(VDD),.Y(g7647),.A(I12132));
  NOT NOT1_2686(.VSS(VSS),.VDD(VDD),.Y(g34664),.A(I32782));
  NOT NOT1_2687(.VSS(VSS),.VDD(VDD),.Y(I27713),.A(g28224));
  NOT NOT1_2688(.VSS(VSS),.VDD(VDD),.Y(I13548),.A(g94));
  NOT NOT1_2689(.VSS(VSS),.VDD(VDD),.Y(g10360),.A(g6836));
  NOT NOT1_2690(.VSS(VSS),.VDD(VDD),.Y(g23012),.A(g20330));
  NOT NOT1_2691(.VSS(VSS),.VDD(VDD),.Y(g24104),.A(g19890));
  NOT NOT1_2692(.VSS(VSS),.VDD(VDD),.Y(g17226),.A(I18252));
  NOT NOT1_2693(.VSS(VSS),.VDD(VDD),.Y(g25139),.A(g22472));
  NOT NOT1_2694(.VSS(VSS),.VDD(VDD),.Y(g17715),.A(I18700));
  NOT NOT1_2695(.VSS(VSS),.VDD(VDD),.Y(g6875),.A(I11697));
  NOT NOT1_2696(.VSS(VSS),.VDD(VDD),.Y(g9777),.A(g5112));
  NOT NOT1_2697(.VSS(VSS),.VDD(VDD),.Y(g17481),.A(g15005));
  NOT NOT1_2698(.VSS(VSS),.VDD(VDD),.Y(I25541),.A(g25180));
  NOT NOT1_2699(.VSS(VSS),.VDD(VDD),.Y(g32840),.A(g30825));
  NOT NOT1_2700(.VSS(VSS),.VDD(VDD),.Y(I28597),.A(g29374));
  NOT NOT1_2701(.VSS(VSS),.VDD(VDD),.Y(g28367),.A(I26880));
  NOT NOT1_2702(.VSS(VSS),.VDD(VDD),.Y(I31474),.A(g33212));
  NOT NOT1_2703(.VSS(VSS),.VDD(VDD),.Y(g24971),.A(g23590));
  NOT NOT1_2704(.VSS(VSS),.VDD(VDD),.Y(g27880),.A(I26427));
  NOT NOT1_2705(.VSS(VSS),.VDD(VDD),.Y(g25138),.A(g22472));
  NOT NOT1_2706(.VSS(VSS),.VDD(VDD),.Y(g34576),.A(I32654));
  NOT NOT1_2707(.VSS(VSS),.VDD(VDD),.Y(g16873),.A(I18063));
  NOT NOT1_2708(.VSS(VSS),.VDD(VDD),.Y(g23541),.A(g21514));
  NOT NOT1_2709(.VSS(VSS),.VDD(VDD),.Y(g31800),.A(g29385));
  NOT NOT1_2710(.VSS(VSS),.VDD(VDD),.Y(g12995),.A(g11820));
  NOT NOT1_2711(.VSS(VSS),.VDD(VDD),.Y(g7503),.A(g1351));
  NOT NOT1_2712(.VSS(VSS),.VDD(VDD),.Y(g7970),.A(g4688));
  NOT NOT1_2713(.VSS(VSS),.VDD(VDD),.Y(g13350),.A(I15906));
  NOT NOT1_2714(.VSS(VSS),.VDD(VDD),.Y(g23473),.A(g20785));
  NOT NOT1_2715(.VSS(VSS),.VDD(VDD),.Y(g33800),.A(I31642));
  NOT NOT1_2716(.VSS(VSS),.VDD(VDD),.Y(g8056),.A(g1246));
  NOT NOT1_2717(.VSS(VSS),.VDD(VDD),.Y(I13317),.A(g6144));
  NOT NOT1_2718(.VSS(VSS),.VDD(VDD),.Y(g11820),.A(I14644));
  NOT NOT1_2719(.VSS(VSS),.VDD(VDD),.Y(g33936),.A(I31820));
  NOT NOT1_2720(.VSS(VSS),.VDD(VDD),.Y(g8456),.A(g56));
  NOT NOT1_2721(.VSS(VSS),.VDD(VDD),.Y(g12880),.A(g10387));
  NOT NOT1_2722(.VSS(VSS),.VDD(VDD),.Y(I22131),.A(g19984));
  NOT NOT1_2723(.VSS(VSS),.VDD(VDD),.Y(I24078),.A(g22360));
  NOT NOT1_2724(.VSS(VSS),.VDD(VDD),.Y(g23789),.A(g21308));
  NOT NOT1_2725(.VSS(VSS),.VDD(VDD),.Y(I17839),.A(g13412));
  NOT NOT1_2726(.VSS(VSS),.VDD(VDD),.Y(g32192),.A(g31262));
  NOT NOT1_2727(.VSS(VSS),.VDD(VDD),.Y(I33109),.A(g34851));
  NOT NOT1_2728(.VSS(VSS),.VDD(VDD),.Y(I15846),.A(g11183));
  NOT NOT1_2729(.VSS(VSS),.VDD(VDD),.Y(I16357),.A(g884));
  NOT NOT1_2730(.VSS(VSS),.VDD(VDD),.Y(I25359),.A(g24715));
  NOT NOT1_2731(.VSS(VSS),.VDD(VDD),.Y(I19799),.A(g17817));
  NOT NOT1_2732(.VSS(VSS),.VDD(VDD),.Y(g30312),.A(g28970));
  NOT NOT1_2733(.VSS(VSS),.VDD(VDD),.Y(I12189),.A(g5869));
  NOT NOT1_2734(.VSS(VSS),.VDD(VDD),.Y(I19813),.A(g17952));
  NOT NOT1_2735(.VSS(VSS),.VDD(VDD),.Y(g24368),.A(g22228));
  NOT NOT1_2736(.VSS(VSS),.VDD(VDD),.Y(g21724),.A(I21291));
  NOT NOT1_2737(.VSS(VSS),.VDD(VDD),.Y(g23788),.A(g18997));
  NOT NOT1_2738(.VSS(VSS),.VDD(VDD),.Y(g8155),.A(g3380));
  NOT NOT1_2739(.VSS(VSS),.VDD(VDD),.Y(g34312),.A(g34098));
  NOT NOT1_2740(.VSS(VSS),.VDD(VDD),.Y(g26973),.A(g26105));
  NOT NOT1_2741(.VSS(VSS),.VDD(VDD),.Y(g34200),.A(g33895));
  NOT NOT1_2742(.VSS(VSS),.VDD(VDD),.Y(g7224),.A(g4601));
  NOT NOT1_2743(.VSS(VSS),.VDD(VDD),.Y(g32522),.A(g30735));
  NOT NOT1_2744(.VSS(VSS),.VDD(VDD),.Y(g23359),.A(I22458));
  NOT NOT1_2745(.VSS(VSS),.VDD(VDD),.Y(g32663),.A(g30673));
  NOT NOT1_2746(.VSS(VSS),.VDD(VDD),.Y(g8355),.A(I12534));
  NOT NOT1_2747(.VSS(VSS),.VDD(VDD),.Y(g8851),.A(g590));
  NOT NOT1_2748(.VSS(VSS),.VDD(VDD),.Y(I13057),.A(g112));
  NOT NOT1_2749(.VSS(VSS),.VDD(VDD),.Y(g14451),.A(I16606));
  NOT NOT1_2750(.VSS(VSS),.VDD(VDD),.Y(I23366),.A(g23321));
  NOT NOT1_2751(.VSS(VSS),.VDD(VDD),.Y(I18364),.A(g13009));
  NOT NOT1_2752(.VSS(VSS),.VDD(VDD),.Y(I22619),.A(g21193));
  NOT NOT1_2753(.VSS(VSS),.VDD(VDD),.Y(I17131),.A(g14384));
  NOT NOT1_2754(.VSS(VSS),.VDD(VDD),.Y(I22502),.A(g19376));
  NOT NOT1_2755(.VSS(VSS),.VDD(VDD),.Y(g22980),.A(I22153));
  NOT NOT1_2756(.VSS(VSS),.VDD(VDD),.Y(g21434),.A(g17248));
  NOT NOT1_2757(.VSS(VSS),.VDD(VDD),.Y(I22557),.A(g20695));
  NOT NOT1_2758(.VSS(VSS),.VDD(VDD),.Y(g21358),.A(g16307));
  NOT NOT1_2759(.VSS(VSS),.VDD(VDD),.Y(g6839),.A(g1858));
  NOT NOT1_2760(.VSS(VSS),.VDD(VDD),.Y(g23434),.A(g21611));
  NOT NOT1_2761(.VSS(VSS),.VDD(VDD),.Y(g24850),.A(I24022));
  NOT NOT1_2762(.VSS(VSS),.VDD(VDD),.Y(g30052),.A(g29018));
  NOT NOT1_2763(.VSS(VSS),.VDD(VDD),.Y(I19674),.A(g15932));
  NOT NOT1_2764(.VSS(VSS),.VDD(VDD),.Y(g8964),.A(g4269));
  NOT NOT1_2765(.VSS(VSS),.VDD(VDD),.Y(I29913),.A(g30605));
  NOT NOT1_2766(.VSS(VSS),.VDD(VDD),.Y(g27831),.A(I26406));
  NOT NOT1_2767(.VSS(VSS),.VDD(VDD),.Y(I11626),.A(g31));
  NOT NOT1_2768(.VSS(VSS),.VDD(VDD),.Y(g11413),.A(g9100));
  NOT NOT1_2769(.VSS(VSS),.VDD(VDD),.Y(g34921),.A(I33155));
  NOT NOT1_2770(.VSS(VSS),.VDD(VDD),.Y(g13413),.A(g11737));
  NOT NOT1_2771(.VSS(VSS),.VDD(VDD),.Y(g34052),.A(g33635));
  NOT NOT1_2772(.VSS(VSS),.VDD(VDD),.Y(g23946),.A(g19210));
  NOT NOT1_2773(.VSS(VSS),.VDD(VDD),.Y(g24133),.A(g19935));
  NOT NOT1_2774(.VSS(VSS),.VDD(VDD),.Y(g29169),.A(g27886));
  NOT NOT1_2775(.VSS(VSS),.VDD(VDD),.Y(g18096),.A(I18894));
  NOT NOT1_2776(.VSS(VSS),.VDD(VDD),.Y(g18944),.A(g15938));
  NOT NOT1_2777(.VSS(VSS),.VDD(VDD),.Y(g20229),.A(g17015));
  NOT NOT1_2778(.VSS(VSS),.VDD(VDD),.Y(g32483),.A(g30673));
  NOT NOT1_2779(.VSS(VSS),.VDD(VDD),.Y(g19617),.A(g16349));
  NOT NOT1_2780(.VSS(VSS),.VDD(VDD),.Y(g19470),.A(g16000));
  NOT NOT1_2781(.VSS(VSS),.VDD(VDD),.Y(g22181),.A(g19277));
  NOT NOT1_2782(.VSS(VSS),.VDD(VDD),.Y(g11691),.A(I14570));
  NOT NOT1_2783(.VSS(VSS),.VDD(VDD),.Y(g19915),.A(g16349));
  NOT NOT1_2784(.VSS(VSS),.VDD(VDD),.Y(g12831),.A(g9569));
  NOT NOT1_2785(.VSS(VSS),.VDD(VDD),.Y(g26732),.A(g25389));
  NOT NOT1_2786(.VSS(VSS),.VDD(VDD),.Y(I16803),.A(g6369));
  NOT NOT1_2787(.VSS(VSS),.VDD(VDD),.Y(I12030),.A(g595));
  NOT NOT1_2788(.VSS(VSS),.VDD(VDD),.Y(I17557),.A(g14510));
  NOT NOT1_2789(.VSS(VSS),.VDD(VDD),.Y(g9541),.A(g2012));
  NOT NOT1_2790(.VSS(VSS),.VDD(VDD),.Y(g32553),.A(g31170));
  NOT NOT1_2791(.VSS(VSS),.VDD(VDD),.Y(g32862),.A(g30825));
  NOT NOT1_2792(.VSS(VSS),.VDD(VDD),.Y(g7617),.A(I12089));
  NOT NOT1_2793(.VSS(VSS),.VDD(VDD),.Y(g16726),.A(g14454));
  NOT NOT1_2794(.VSS(VSS),.VDD(VDD),.Y(I26649),.A(g27675));
  NOT NOT1_2795(.VSS(VSS),.VDD(VDD),.Y(g34813),.A(I33027));
  NOT NOT1_2796(.VSS(VSS),.VDD(VDD),.Y(g10776),.A(I14033));
  NOT NOT1_2797(.VSS(VSS),.VDD(VDD),.Y(g19277),.A(I19813));
  NOT NOT1_2798(.VSS(VSS),.VDD(VDD),.Y(g32949),.A(g30825));
  NOT NOT1_2799(.VSS(VSS),.VDD(VDD),.Y(g9332),.A(g64));
  NOT NOT1_2800(.VSS(VSS),.VDD(VDD),.Y(g14591),.A(I16709));
  NOT NOT1_2801(.VSS(VSS),.VDD(VDD),.Y(g14785),.A(g12629));
  NOT NOT1_2802(.VSS(VSS),.VDD(VDD),.Y(I21226),.A(g16540));
  NOT NOT1_2803(.VSS(VSS),.VDD(VDD),.Y(I22286),.A(g19446));
  NOT NOT1_2804(.VSS(VSS),.VDD(VDD),.Y(g7516),.A(I12003));
  NOT NOT1_2805(.VSS(VSS),.VDD(VDD),.Y(g21682),.A(g16540));
  NOT NOT1_2806(.VSS(VSS),.VDD(VDD),.Y(I18224),.A(g13793));
  NOT NOT1_2807(.VSS(VSS),.VDD(VDD),.Y(g9680),.A(I13276));
  NOT NOT1_2808(.VSS(VSS),.VDD(VDD),.Y(g9153),.A(I12991));
  NOT NOT1_2809(.VSS(VSS),.VDD(VDD),.Y(g10147),.A(g728));
  NOT NOT1_2810(.VSS(VSS),.VDD(VDD),.Y(g20716),.A(g15277));
  NOT NOT1_2811(.VSS(VSS),.VDD(VDD),.Y(g27989),.A(g26759));
  NOT NOT1_2812(.VSS(VSS),.VDD(VDD),.Y(g29217),.A(I27567));
  NOT NOT1_2813(.VSS(VSS),.VDD(VDD),.Y(g34973),.A(I33235));
  NOT NOT1_2814(.VSS(VSS),.VDD(VDD),.Y(g25554),.A(g22550));
  NOT NOT1_2815(.VSS(VSS),.VDD(VDD),.Y(I15929),.A(g10430));
  NOT NOT1_2816(.VSS(VSS),.VDD(VDD),.Y(I18571),.A(g13074));
  NOT NOT1_2817(.VSS(VSS),.VDD(VDD),.Y(g21291),.A(g16620));
  NOT NOT1_2818(.VSS(VSS),.VDD(VDD),.Y(g32536),.A(g31376));
  NOT NOT1_2819(.VSS(VSS),.VDD(VDD),.Y(g14147),.A(I16357));
  NOT NOT1_2820(.VSS(VSS),.VDD(VDD),.Y(g30184),.A(g28144));
  NOT NOT1_2821(.VSS(VSS),.VDD(VDD),.Y(I31796),.A(g33176));
  NOT NOT1_2822(.VSS(VSS),.VDD(VDD),.Y(g10355),.A(g6816));
  NOT NOT1_2823(.VSS(VSS),.VDD(VDD),.Y(g32948),.A(g30735));
  NOT NOT1_2824(.VSS(VSS),.VDD(VDD),.Y(g23291),.A(g21070));
  NOT NOT1_2825(.VSS(VSS),.VDD(VDD),.Y(g16607),.A(g13960));
  NOT NOT1_2826(.VSS(VSS),.VDD(VDD),.Y(g19494),.A(g16349));
  NOT NOT1_2827(.VSS(VSS),.VDD(VDD),.Y(g11929),.A(I14745));
  NOT NOT1_2828(.VSS(VSS),.VDD(VDD),.Y(I11737),.A(g4467));
  NOT NOT1_2829(.VSS(VSS),.VDD(VDD),.Y(g34674),.A(I32806));
  NOT NOT1_2830(.VSS(VSS),.VDD(VDD),.Y(g8279),.A(I12487));
  NOT NOT1_2831(.VSS(VSS),.VDD(VDD),.Y(g16320),.A(g14454));
  NOT NOT1_2832(.VSS(VSS),.VDD(VDD),.Y(g20582),.A(g17873));
  NOT NOT1_2833(.VSS(VSS),.VDD(VDD),.Y(g32702),.A(g30735));
  NOT NOT1_2834(.VSS(VSS),.VDD(VDD),.Y(g9744),.A(g6486));
  NOT NOT1_2835(.VSS(VSS),.VDD(VDD),.Y(g10370),.A(g7095));
  NOT NOT1_2836(.VSS(VSS),.VDD(VDD),.Y(g31000),.A(g29737));
  NOT NOT1_2837(.VSS(VSS),.VDD(VDD),.Y(g32757),.A(g30937));
  NOT NOT1_2838(.VSS(VSS),.VDD(VDD),.Y(g32904),.A(g30735));
  NOT NOT1_2839(.VSS(VSS),.VDD(VDD),.Y(g6988),.A(g4765));
  NOT NOT1_2840(.VSS(VSS),.VDD(VDD),.Y(I14866),.A(g9748));
  NOT NOT1_2841(.VSS(VSS),.VDD(VDD),.Y(g16530),.A(g14454));
  NOT NOT1_2842(.VSS(VSS),.VDD(VDD),.Y(g26400),.A(I25351));
  NOT NOT1_2843(.VSS(VSS),.VDD(VDD),.Y(g11928),.A(I14742));
  NOT NOT1_2844(.VSS(VSS),.VDD(VDD),.Y(g25115),.A(I24281));
  NOT NOT1_2845(.VSS(VSS),.VDD(VDD),.Y(g13583),.A(I16028));
  NOT NOT1_2846(.VSS(VSS),.VDD(VDD),.Y(g32621),.A(g31542));
  NOT NOT1_2847(.VSS(VSS),.VDD(VDD),.Y(g8872),.A(g4258));
  NOT NOT1_2848(.VSS(VSS),.VDD(VDD),.Y(g22520),.A(g19801));
  NOT NOT1_2849(.VSS(VSS),.VDD(VDD),.Y(I22601),.A(g21127));
  NOT NOT1_2850(.VSS(VSS),.VDD(VDD),.Y(g10151),.A(g1992));
  NOT NOT1_2851(.VSS(VSS),.VDD(VDD),.Y(g28120),.A(g27108));
  NOT NOT1_2852(.VSS(VSS),.VDD(VDD),.Y(I32228),.A(g34122));
  NOT NOT1_2853(.VSS(VSS),.VDD(VDD),.Y(I11697),.A(g3352));
  NOT NOT1_2854(.VSS(VSS),.VDD(VDD),.Y(g10172),.A(g6459));
  NOT NOT1_2855(.VSS(VSS),.VDD(VDD),.Y(g20627),.A(g17433));
  NOT NOT1_2856(.VSS(VSS),.VDD(VDD),.Y(I12837),.A(g4222));
  NOT NOT1_2857(.VSS(VSS),.VDD(VDD),.Y(g7892),.A(g4801));
  NOT NOT1_2858(.VSS(VSS),.VDD(VDD),.Y(g34934),.A(g34918));
  NOT NOT1_2859(.VSS(VSS),.VDD(VDD),.Y(g9558),.A(g5841));
  NOT NOT1_2860(.VSS(VSS),.VDD(VDD),.Y(g20379),.A(g17821));
  NOT NOT1_2861(.VSS(VSS),.VDD(VDD),.Y(g8057),.A(g3068));
  NOT NOT1_2862(.VSS(VSS),.VDD(VDD),.Y(g32564),.A(g31376));
  NOT NOT1_2863(.VSS(VSS),.VDD(VDD),.Y(I13995),.A(g8744));
  NOT NOT1_2864(.VSS(VSS),.VDD(VDD),.Y(g24379),.A(g22550));
  NOT NOT1_2865(.VSS(VSS),.VDD(VDD),.Y(g8457),.A(g225));
  NOT NOT1_2866(.VSS(VSS),.VDD(VDD),.Y(g8989),.A(I12935));
  NOT NOT1_2867(.VSS(VSS),.VDD(VDD),.Y(g19352),.A(g15758));
  NOT NOT1_2868(.VSS(VSS),.VDD(VDD),.Y(g22546),.A(I21918));
  NOT NOT1_2869(.VSS(VSS),.VDD(VDD),.Y(g23760),.A(I22889));
  NOT NOT1_2870(.VSS(VSS),.VDD(VDD),.Y(g20050),.A(I20321));
  NOT NOT1_2871(.VSS(VSS),.VDD(VDD),.Y(g23029),.A(g20453));
  NOT NOT1_2872(.VSS(VSS),.VDD(VDD),.Y(g6804),.A(g490));
  NOT NOT1_2873(.VSS(VSS),.VDD(VDD),.Y(g24112),.A(g19935));
  NOT NOT1_2874(.VSS(VSS),.VDD(VDD),.Y(g10367),.A(g6870));
  NOT NOT1_2875(.VSS(VSS),.VDD(VDD),.Y(g10394),.A(g6994));
  NOT NOT1_2876(.VSS(VSS),.VDD(VDD),.Y(I25028),.A(g24484));
  NOT NOT1_2877(.VSS(VSS),.VDD(VDD),.Y(g24050),.A(g20841));
  NOT NOT1_2878(.VSS(VSS),.VDD(VDD),.Y(g9901),.A(g84));
  NOT NOT1_2879(.VSS(VSS),.VDD(VDD),.Y(g34692),.A(I32846));
  NOT NOT1_2880(.VSS(VSS),.VDD(VDD),.Y(I22143),.A(g20189));
  NOT NOT1_2881(.VSS(VSS),.VDD(VDD),.Y(I21784),.A(g19638));
  NOT NOT1_2882(.VSS(VSS),.VDD(VDD),.Y(g23506),.A(g21514));
  NOT NOT1_2883(.VSS(VSS),.VDD(VDD),.Y(g23028),.A(g20391));
  NOT NOT1_2884(.VSS(VSS),.VDD(VDD),.Y(I18752),.A(g6358));
  NOT NOT1_2885(.VSS(VSS),.VDD(VDD),.Y(I28480),.A(g28652));
  NOT NOT1_2886(.VSS(VSS),.VDD(VDD),.Y(g31814),.A(g29385));
  NOT NOT1_2887(.VSS(VSS),.VDD(VDD),.Y(g32673),.A(g31376));
  NOT NOT1_2888(.VSS(VSS),.VDD(VDD),.Y(g32847),.A(g30735));
  NOT NOT1_2889(.VSS(VSS),.VDD(VDD),.Y(g20386),.A(g15224));
  NOT NOT1_2890(.VSS(VSS),.VDD(VDD),.Y(I21297),.A(g18597));
  NOT NOT1_2891(.VSS(VSS),.VDD(VDD),.Y(g8971),.A(I12927));
  NOT NOT1_2892(.VSS(VSS),.VDD(VDD),.Y(g22860),.A(g20000));
  NOT NOT1_2893(.VSS(VSS),.VDD(VDD),.Y(g24386),.A(g22594));
  NOT NOT1_2894(.VSS(VSS),.VDD(VDD),.Y(g20603),.A(g17873));
  NOT NOT1_2895(.VSS(VSS),.VDD(VDD),.Y(g9511),.A(g5881));
  NOT NOT1_2896(.VSS(VSS),.VDD(VDD),.Y(g27736),.A(I26356));
  NOT NOT1_2897(.VSS(VSS),.VDD(VDD),.Y(g7738),.A(I12176));
  NOT NOT1_2898(.VSS(VSS),.VDD(VDD),.Y(g31807),.A(g29385));
  NOT NOT1_2899(.VSS(VSS),.VDD(VDD),.Y(g8686),.A(g2819));
  NOT NOT1_2900(.VSS(VSS),.VDD(VDD),.Y(g13302),.A(g12321));
  NOT NOT1_2901(.VSS(VSS),.VDD(VDD),.Y(g20096),.A(g16782));
  NOT NOT1_2902(.VSS(VSS),.VDD(VDD),.Y(g24603),.A(g23108));
  NOT NOT1_2903(.VSS(VSS),.VDD(VDD),.Y(g33772),.A(I31622));
  NOT NOT1_2904(.VSS(VSS),.VDD(VDD),.Y(g7991),.A(g4878));
  NOT NOT1_2905(.VSS(VSS),.VDD(VDD),.Y(I23354),.A(g23277));
  NOT NOT1_2906(.VSS(VSS),.VDD(VDD),.Y(g24096),.A(g19890));
  NOT NOT1_2907(.VSS(VSS),.VDD(VDD),.Y(g29922),.A(g28837));
  NOT NOT1_2908(.VSS(VSS),.VDD(VDD),.Y(g34400),.A(g34142));
  NOT NOT1_2909(.VSS(VSS),.VDD(VDD),.Y(g7244),.A(g4408));
  NOT NOT1_2910(.VSS(VSS),.VDD(VDD),.Y(g12887),.A(g10394));
  NOT NOT1_2911(.VSS(VSS),.VDD(VDD),.Y(g10420),.A(g9239));
  NOT NOT1_2912(.VSS(VSS),.VDD(VDD),.Y(I17143),.A(g14412));
  NOT NOT1_2913(.VSS(VSS),.VDD(VDD),.Y(g22497),.A(g19513));
  NOT NOT1_2914(.VSS(VSS),.VDD(VDD),.Y(g25184),.A(g22763));
  NOT NOT1_2915(.VSS(VSS),.VDD(VDD),.Y(g32509),.A(g31070));
  NOT NOT1_2916(.VSS(VSS),.VDD(VDD),.Y(g31639),.A(I29225));
  NOT NOT1_2917(.VSS(VSS),.VDD(VDD),.Y(g10319),.A(I13740));
  NOT NOT1_2918(.VSS(VSS),.VDD(VDD),.Y(g17088),.A(I18160));
  NOT NOT1_2919(.VSS(VSS),.VDD(VDD),.Y(g32933),.A(g31376));
  NOT NOT1_2920(.VSS(VSS),.VDD(VDD),.Y(g30329),.A(I28588));
  NOT NOT1_2921(.VSS(VSS),.VDD(VDD),.Y(g9492),.A(g2759));
  NOT NOT1_2922(.VSS(VSS),.VDD(VDD),.Y(I21181),.A(g17413));
  NOT NOT1_2923(.VSS(VSS),.VDD(VDD),.Y(g16136),.A(I17491));
  NOT NOT1_2924(.VSS(VSS),.VDD(VDD),.Y(g7340),.A(g4443));
  NOT NOT1_2925(.VSS(VSS),.VDD(VDD),.Y(g20681),.A(g15483));
  NOT NOT1_2926(.VSS(VSS),.VDD(VDD),.Y(g9600),.A(g3632));
  NOT NOT1_2927(.VSS(VSS),.VDD(VDD),.Y(I23671),.A(g23202));
  NOT NOT1_2928(.VSS(VSS),.VDD(VDD),.Y(g32508),.A(g30825));
  NOT NOT1_2929(.VSS(VSS),.VDD(VDD),.Y(g9574),.A(g6462));
  NOT NOT1_2930(.VSS(VSS),.VDD(VDD),.Y(g31638),.A(g29689));
  NOT NOT1_2931(.VSS(VSS),.VDD(VDD),.Y(g9864),.A(I13424));
  NOT NOT1_2932(.VSS(VSS),.VDD(VDD),.Y(g32634),.A(g30673));
  NOT NOT1_2933(.VSS(VSS),.VDD(VDD),.Y(g32851),.A(g31327));
  NOT NOT1_2934(.VSS(VSS),.VDD(VDD),.Y(g32872),.A(g31327));
  NOT NOT1_2935(.VSS(VSS),.VDD(VDD),.Y(g33638),.A(I31469));
  NOT NOT1_2936(.VSS(VSS),.VDD(VDD),.Y(g35001),.A(I33297));
  NOT NOT1_2937(.VSS(VSS),.VDD(VDD),.Y(g30328),.A(I28585));
  NOT NOT1_2938(.VSS(VSS),.VDD(VDD),.Y(g7907),.A(g3072));
  NOT NOT1_2939(.VSS(VSS),.VDD(VDD),.Y(g11640),.A(I14550));
  NOT NOT1_2940(.VSS(VSS),.VDD(VDD),.Y(g11769),.A(g8626));
  NOT NOT1_2941(.VSS(VSS),.VDD(VDD),.Y(g34539),.A(g34354));
  NOT NOT1_2942(.VSS(VSS),.VDD(VDD),.Y(g9714),.A(g4012));
  NOT NOT1_2943(.VSS(VSS),.VDD(VDD),.Y(g12843),.A(g10359));
  NOT NOT1_2944(.VSS(VSS),.VDD(VDD),.Y(g17497),.A(g14879));
  NOT NOT1_2945(.VSS(VSS),.VDD(VDD),.Y(g22987),.A(g20391));
  NOT NOT1_2946(.VSS(VSS),.VDD(VDD),.Y(g34328),.A(g34096));
  NOT NOT1_2947(.VSS(VSS),.VDD(VDD),.Y(g10059),.A(g6451));
  NOT NOT1_2948(.VSS(VSS),.VDD(VDD),.Y(g23927),.A(g19074));
  NOT NOT1_2949(.VSS(VSS),.VDD(VDD),.Y(I18842),.A(g13809));
  NOT NOT1_2950(.VSS(VSS),.VDD(VDD),.Y(g24429),.A(g22722));
  NOT NOT1_2951(.VSS(VSS),.VDD(VDD),.Y(g19524),.A(g15695));
  NOT NOT1_2952(.VSS(VSS),.VDD(VDD),.Y(I29891),.A(g31578));
  NOT NOT1_2953(.VSS(VSS),.VDD(VDD),.Y(g7517),.A(g962));
  NOT NOT1_2954(.VSS(VSS),.VDD(VDD),.Y(g22658),.A(I21969));
  NOT NOT1_2955(.VSS(VSS),.VDD(VDD),.Y(g29953),.A(g28907));
  NOT NOT1_2956(.VSS(VSS),.VDD(VDD),.Y(g10540),.A(g9392));
  NOT NOT1_2957(.VSS(VSS),.VDD(VDD),.Y(g10058),.A(g6497));
  NOT NOT1_2958(.VSS(VSS),.VDD(VDD),.Y(g31841),.A(g29385));
  NOT NOT1_2959(.VSS(VSS),.VDD(VDD),.Y(g24428),.A(g22722));
  NOT NOT1_2960(.VSS(VSS),.VDD(VDD),.Y(I32096),.A(g33641));
  NOT NOT1_2961(.VSS(VSS),.VDD(VDD),.Y(g33391),.A(g32384));
  NOT NOT1_2962(.VSS(VSS),.VDD(VDD),.Y(g19477),.A(g16431));
  NOT NOT1_2963(.VSS(VSS),.VDD(VDD),.Y(g12869),.A(g10376));
  NOT NOT1_2964(.VSS(VSS),.VDD(VDD),.Y(g16164),.A(I17507));
  NOT NOT1_2965(.VSS(VSS),.VDD(VDD),.Y(g23649),.A(g18833));
  NOT NOT1_2966(.VSS(VSS),.VDD(VDD),.Y(g26683),.A(g25514));
  NOT NOT1_2967(.VSS(VSS),.VDD(VDD),.Y(g7876),.A(g1495));
  NOT NOT1_2968(.VSS(VSS),.VDD(VDD),.Y(g25692),.A(I24839));
  NOT NOT1_2969(.VSS(VSS),.VDD(VDD),.Y(g15614),.A(g14914));
  NOT NOT1_2970(.VSS(VSS),.VDD(VDD),.Y(g22339),.A(g19801));
  NOT NOT1_2971(.VSS(VSS),.VDD(VDD),.Y(g20765),.A(g17748));
  NOT NOT1_2972(.VSS(VSS),.VDD(VDD),.Y(g8938),.A(g4899));
  NOT NOT1_2973(.VSS(VSS),.VDD(VDD),.Y(I19235),.A(g15078));
  NOT NOT1_2974(.VSS(VSS),.VDD(VDD),.Y(I20495),.A(g16283));
  NOT NOT1_2975(.VSS(VSS),.VDD(VDD),.Y(g29800),.A(g28363));
  NOT NOT1_2976(.VSS(VSS),.VDD(VDD),.Y(g10203),.A(g2393));
  NOT NOT1_2977(.VSS(VSS),.VDD(VDD),.Y(g12868),.A(g10377));
  NOT NOT1_2978(.VSS(VSS),.VDD(VDD),.Y(g21903),.A(I21480));
  NOT NOT1_2979(.VSS(VSS),.VDD(VDD),.Y(g14203),.A(g12381));
  NOT NOT1_2980(.VSS(VSS),.VDD(VDD),.Y(g20549),.A(g15277));
  NOT NOT1_2981(.VSS(VSS),.VDD(VDD),.Y(g23648),.A(g18833));
  NOT NOT1_2982(.VSS(VSS),.VDD(VDD),.Y(g13881),.A(I16181));
  NOT NOT1_2983(.VSS(VSS),.VDD(VDD),.Y(I16090),.A(g10430));
  NOT NOT1_2984(.VSS(VSS),.VDD(VDD),.Y(g22338),.A(g19801));
  NOT NOT1_2985(.VSS(VSS),.VDD(VDD),.Y(g23491),.A(g21514));
  NOT NOT1_2986(.VSS(VSS),.VDD(VDD),.Y(I20816),.A(g17088));
  NOT NOT1_2987(.VSS(VSS),.VDD(VDD),.Y(g23903),.A(g18997));
  NOT NOT1_2988(.VSS(VSS),.VDD(VDD),.Y(I33252),.A(g34974));
  NOT NOT1_2989(.VSS(VSS),.VDD(VDD),.Y(I32681),.A(g34429));
  NOT NOT1_2990(.VSS(VSS),.VDD(VDD),.Y(g10044),.A(g5357));
  NOT NOT1_2991(.VSS(VSS),.VDD(VDD),.Y(g34241),.A(I32222));
  NOT NOT1_2992(.VSS(VSS),.VDD(VDD),.Y(g27709),.A(I26337));
  NOT NOT1_2993(.VSS(VSS),.VDD(VDD),.Y(g21604),.A(g15938));
  NOT NOT1_2994(.VSS(VSS),.VDD(VDD),.Y(I22580),.A(g20982));
  NOT NOT1_2995(.VSS(VSS),.VDD(VDD),.Y(I16651),.A(g10542));
  NOT NOT1_2996(.VSS(VSS),.VDD(VDD),.Y(g20548),.A(g15426));
  NOT NOT1_2997(.VSS(VSS),.VDD(VDD),.Y(g8519),.A(g287));
  NOT NOT1_2998(.VSS(VSS),.VDD(VDD),.Y(g8740),.A(I12735));
  NOT NOT1_2999(.VSS(VSS),.VDD(VDD),.Y(g31578),.A(I29199));
  NOT NOT1_3000(.VSS(VSS),.VDD(VDD),.Y(g25013),.A(g23599));
  NOT NOT1_3001(.VSS(VSS),.VDD(VDD),.Y(g31835),.A(g29385));
  NOT NOT1_3002(.VSS(VSS),.VDD(VDD),.Y(g32574),.A(g31070));
  NOT NOT1_3003(.VSS(VSS),.VDD(VDD),.Y(I20985),.A(g16300));
  NOT NOT1_3004(.VSS(VSS),.VDD(VDD),.Y(g24548),.A(g22942));
  NOT NOT1_3005(.VSS(VSS),.VDD(VDD),.Y(I31564),.A(g33204));
  NOT NOT1_3006(.VSS(VSS),.VDD(VDD),.Y(g17296),.A(I18280));
  NOT NOT1_3007(.VSS(VSS),.VDD(VDD),.Y(g25214),.A(g22228));
  NOT NOT1_3008(.VSS(VSS),.VDD(VDD),.Y(g27708),.A(I26334));
  NOT NOT1_3009(.VSS(VSS),.VDD(VDD),.Y(I12418),.A(g55));
  NOT NOT1_3010(.VSS(VSS),.VDD(VDD),.Y(g17644),.A(g15002));
  NOT NOT1_3011(.VSS(VSS),.VDD(VDD),.Y(g20504),.A(g18008));
  NOT NOT1_3012(.VSS(VSS),.VDD(VDD),.Y(g30100),.A(g29131));
  NOT NOT1_3013(.VSS(VSS),.VDD(VDD),.Y(g23563),.A(g20682));
  NOT NOT1_3014(.VSS(VSS),.VDD(VDD),.Y(g10377),.A(g6940));
  NOT NOT1_3015(.VSS(VSS),.VDD(VDD),.Y(g32912),.A(g30735));
  NOT NOT1_3016(.VSS(VSS),.VDD(VDD),.Y(g8606),.A(g4653));
  NOT NOT1_3017(.VSS(VSS),.VDD(VDD),.Y(I18865),.A(g14314));
  NOT NOT1_3018(.VSS(VSS),.VDD(VDD),.Y(I20954),.A(g16228));
  NOT NOT1_3019(.VSS(VSS),.VDD(VDD),.Y(g19748),.A(g17015));
  NOT NOT1_3020(.VSS(VSS),.VDD(VDD),.Y(g10120),.A(g1902));
  NOT NOT1_3021(.VSS(VSS),.VDD(VDD),.Y(g22197),.A(g19074));
  NOT NOT1_3022(.VSS(VSS),.VDD(VDD),.Y(g14377),.A(g12201));
  NOT NOT1_3023(.VSS(VSS),.VDD(VDD),.Y(I11753),.A(g4492));
  NOT NOT1_3024(.VSS(VSS),.VDD(VDD),.Y(g22855),.A(g20391));
  NOT NOT1_3025(.VSS(VSS),.VDD(VDD),.Y(g19276),.A(g17367));
  NOT NOT1_3026(.VSS(VSS),.VDD(VDD),.Y(g9889),.A(g6128));
  NOT NOT1_3027(.VSS(VSS),.VDD(VDD),.Y(g13027),.A(I15647));
  NOT NOT1_3028(.VSS(VSS),.VDD(VDD),.Y(g7110),.A(g6682));
  NOT NOT1_3029(.VSS(VSS),.VDD(VDD),.Y(I14660),.A(g9746));
  NOT NOT1_3030(.VSS(VSS),.VDD(VDD),.Y(g33442),.A(g31937));
  NOT NOT1_3031(.VSS(VSS),.VDD(VDD),.Y(g22870),.A(g20887));
  NOT NOT1_3032(.VSS(VSS),.VDD(VDD),.Y(g22527),.A(g19546));
  NOT NOT1_3033(.VSS(VSS),.VDD(VDD),.Y(I21860),.A(g19638));
  NOT NOT1_3034(.VSS(VSS),.VDD(VDD),.Y(g34683),.A(I32827));
  NOT NOT1_3035(.VSS(VSS),.VDD(VDD),.Y(g28127),.A(g27102));
  NOT NOT1_3036(.VSS(VSS),.VDD(VDD),.Y(g25538),.A(g22594));
  NOT NOT1_3037(.VSS(VSS),.VDD(VDD),.Y(g29216),.A(I27564));
  NOT NOT1_3038(.VSS(VSS),.VDD(VDD),.Y(I32690),.A(g34432));
  NOT NOT1_3039(.VSS(VSS),.VDD(VDD),.Y(g11249),.A(g8405));
  NOT NOT1_3040(.VSS(VSS),.VDD(VDD),.Y(I28838),.A(g29372));
  NOT NOT1_3041(.VSS(VSS),.VDD(VDD),.Y(I13031),.A(g6747));
  NOT NOT1_3042(.VSS(VSS),.VDD(VDD),.Y(g14738),.A(I16821));
  NOT NOT1_3043(.VSS(VSS),.VDD(VDD),.Y(g13249),.A(g10590));
  NOT NOT1_3044(.VSS(VSS),.VDD(VDD),.Y(g14562),.A(g12036));
  NOT NOT1_3045(.VSS(VSS),.VDD(VDD),.Y(g14645),.A(I16755));
  NOT NOT1_3046(.VSS(VSS),.VDD(VDD),.Y(I30861),.A(g32383));
  NOT NOT1_3047(.VSS(VSS),.VDD(VDD),.Y(g20129),.A(g17328));
  NOT NOT1_3048(.VSS(VSS),.VDD(VDD),.Y(g16606),.A(g14110));
  NOT NOT1_3049(.VSS(VSS),.VDD(VDD),.Y(g17197),.A(I18233));
  NOT NOT1_3050(.VSS(VSS),.VDD(VDD),.Y(g18880),.A(g15656));
  NOT NOT1_3051(.VSS(VSS),.VDD(VDD),.Y(g23767),.A(g18997));
  NOT NOT1_3052(.VSS(VSS),.VDD(VDD),.Y(g23794),.A(g19147));
  NOT NOT1_3053(.VSS(VSS),.VDD(VDD),.Y(g21395),.A(g17873));
  NOT NOT1_3054(.VSS(VSS),.VDD(VDD),.Y(g24129),.A(g20857));
  NOT NOT1_3055(.VSS(VSS),.VDD(VDD),.Y(g32592),.A(g30673));
  NOT NOT1_3056(.VSS(VSS),.VDD(VDD),.Y(g20057),.A(g16349));
  NOT NOT1_3057(.VSS(VSS),.VDD(VDD),.Y(g32756),.A(g31021));
  NOT NOT1_3058(.VSS(VSS),.VDD(VDD),.Y(g23395),.A(I22502));
  NOT NOT1_3059(.VSS(VSS),.VDD(VDD),.Y(g24057),.A(g20841));
  NOT NOT1_3060(.VSS(VSS),.VDD(VDD),.Y(g20128),.A(g17533));
  NOT NOT1_3061(.VSS(VSS),.VDD(VDD),.Y(I12167),.A(g5176));
  NOT NOT1_3062(.VSS(VSS),.VDD(VDD),.Y(g14290),.A(I16460));
  NOT NOT1_3063(.VSS(VSS),.VDD(VDD),.Y(g17870),.A(I18842));
  NOT NOT1_3064(.VSS(VSS),.VDD(VDD),.Y(g17411),.A(g14454));
  NOT NOT1_3065(.VSS(VSS),.VDD(VDD),.Y(g17527),.A(g14741));
  NOT NOT1_3066(.VSS(VSS),.VDD(VDD),.Y(g23899),.A(g19277));
  NOT NOT1_3067(.VSS(VSS),.VDD(VDD),.Y(g7002),.A(g5160));
  NOT NOT1_3068(.VSS(VSS),.VDD(VDD),.Y(g13003),.A(I15609));
  NOT NOT1_3069(.VSS(VSS),.VDD(VDD),.Y(g24128),.A(g20720));
  NOT NOT1_3070(.VSS(VSS),.VDD(VDD),.Y(g11204),.A(I14271));
  NOT NOT1_3071(.VSS(VSS),.VDD(VDD),.Y(I14550),.A(g10072));
  NOT NOT1_3072(.VSS(VSS),.VDD(VDD),.Y(g7824),.A(g4169));
  NOT NOT1_3073(.VSS(VSS),.VDD(VDD),.Y(g30991),.A(I28925));
  NOT NOT1_3074(.VSS(VSS),.VDD(VDD),.Y(g6996),.A(g4955));
  NOT NOT1_3075(.VSS(VSS),.VDD(VDD),.Y(g25241),.A(g23651));
  NOT NOT1_3076(.VSS(VSS),.VDD(VDD),.Y(g11779),.A(g9602));
  NOT NOT1_3077(.VSS(VSS),.VDD(VDD),.Y(I18270),.A(g13191));
  NOT NOT1_3078(.VSS(VSS),.VDD(VDD),.Y(g16750),.A(g14454));
  NOT NOT1_3079(.VSS(VSS),.VDD(VDD),.Y(g22867),.A(g20391));
  NOT NOT1_3080(.VSS(VSS),.VDD(VDD),.Y(g34991),.A(I33273));
  NOT NOT1_3081(.VSS(VSS),.VDD(VDD),.Y(g7236),.A(g4608));
  NOT NOT1_3082(.VSS(VSS),.VDD(VDD),.Y(g9285),.A(g2715));
  NOT NOT1_3083(.VSS(VSS),.VDD(VDD),.Y(g20626),.A(g15483));
  NOT NOT1_3084(.VSS(VSS),.VDD(VDD),.Y(g27774),.A(I26381));
  NOT NOT1_3085(.VSS(VSS),.VDD(VDD),.Y(I27401),.A(g27051));
  NOT NOT1_3086(.VSS(VSS),.VDD(VDD),.Y(I11843),.A(g111));
  NOT NOT1_3087(.VSS(VSS),.VDD(VDD),.Y(g23898),.A(g19277));
  NOT NOT1_3088(.VSS(VSS),.VDD(VDD),.Y(g9500),.A(g5495));
  NOT NOT1_3089(.VSS(VSS),.VDD(VDD),.Y(g20323),.A(g17873));
  NOT NOT1_3090(.VSS(VSS),.VDD(VDD),.Y(I21250),.A(g16540));
  NOT NOT1_3091(.VSS(VSS),.VDD(VDD),.Y(g29117),.A(g27886));
  NOT NOT1_3092(.VSS(VSS),.VDD(VDD),.Y(g24626),.A(g23139));
  NOT NOT1_3093(.VSS(VSS),.VDD(VDD),.Y(g33430),.A(g32421));
  NOT NOT1_3094(.VSS(VSS),.VDD(VDD),.Y(g23191),.A(I22289));
  NOT NOT1_3095(.VSS(VSS),.VDD(VDD),.Y(g20533),.A(g17271));
  NOT NOT1_3096(.VSS(VSS),.VDD(VDD),.Y(g10427),.A(g10053));
  NOT NOT1_3097(.VSS(VSS),.VDD(VDD),.Y(g12955),.A(I15577));
  NOT NOT1_3098(.VSS(VSS),.VDD(VDD),.Y(g32820),.A(g31672));
  NOT NOT1_3099(.VSS(VSS),.VDD(VDD),.Y(I18460),.A(g5276));
  NOT NOT1_3100(.VSS(VSS),.VDD(VDD),.Y(g8341),.A(g3119));
  NOT NOT1_3101(.VSS(VSS),.VDD(VDD),.Y(g10366),.A(g6895));
  NOT NOT1_3102(.VSS(VSS),.VDD(VDD),.Y(g24533),.A(g22876));
  NOT NOT1_3103(.VSS(VSS),.VDD(VDD),.Y(g25100),.A(g22384));
  NOT NOT1_3104(.VSS(VSS),.VDD(VDD),.Y(g12879),.A(g10381));
  NOT NOT1_3105(.VSS(VSS),.VDD(VDD),.Y(g22714),.A(g20436));
  NOT NOT1_3106(.VSS(VSS),.VDD(VDD),.Y(g11786),.A(g7549));
  NOT NOT1_3107(.VSS(VSS),.VDD(VDD),.Y(g14366),.A(I16526));
  NOT NOT1_3108(.VSS(VSS),.VDD(VDD),.Y(g17503),.A(g14892));
  NOT NOT1_3109(.VSS(VSS),.VDD(VDD),.Y(I14054),.A(g10028));
  NOT NOT1_3110(.VSS(VSS),.VDD(VDD),.Y(g9184),.A(g6120));
  NOT NOT1_3111(.VSS(VSS),.VDD(VDD),.Y(g23521),.A(g21468));
  NOT NOT1_3112(.VSS(VSS),.VDD(VDD),.Y(g28181),.A(I26700));
  NOT NOT1_3113(.VSS(VSS),.VDD(VDD),.Y(g25771),.A(I24920));
  NOT NOT1_3114(.VSS(VSS),.VDD(VDD),.Y(g20775),.A(g18008));
  NOT NOT1_3115(.VSS(VSS),.VDD(VDD),.Y(g18831),.A(g15224));
  NOT NOT1_3116(.VSS(VSS),.VDD(VDD),.Y(I15647),.A(g12109));
  NOT NOT1_3117(.VSS(VSS),.VDD(VDD),.Y(I23339),.A(g23232));
  NOT NOT1_3118(.VSS(VSS),.VDD(VDD),.Y(g32846),.A(g31376));
  NOT NOT1_3119(.VSS(VSS),.VDD(VDD),.Y(g9339),.A(g2295));
  NOT NOT1_3120(.VSS(VSS),.VDD(VDD),.Y(I19759),.A(g17767));
  NOT NOT1_3121(.VSS(VSS),.VDD(VDD),.Y(g19733),.A(g16856));
  NOT NOT1_3122(.VSS(VSS),.VDD(VDD),.Y(I24558),.A(g23777));
  NOT NOT1_3123(.VSS(VSS),.VDD(VDD),.Y(g12878),.A(g10386));
  NOT NOT1_3124(.VSS(VSS),.VDD(VDD),.Y(g26758),.A(g25389));
  NOT NOT1_3125(.VSS(VSS),.VDD(VDD),.Y(I27749),.A(g28917));
  NOT NOT1_3126(.VSS(VSS),.VDD(VDD),.Y(I20830),.A(g17657));
  NOT NOT1_3127(.VSS(VSS),.VDD(VDD),.Y(g12337),.A(g9340));
  NOT NOT1_3128(.VSS(VSS),.VDD(VDD),.Y(g32731),.A(g31376));
  NOT NOT1_3129(.VSS(VSS),.VDD(VDD),.Y(g31806),.A(g29385));
  NOT NOT1_3130(.VSS(VSS),.VDD(VDD),.Y(g22202),.A(I21784));
  NOT NOT1_3131(.VSS(VSS),.VDD(VDD),.Y(g33806),.A(I31650));
  NOT NOT1_3132(.VSS(VSS),.VDD(VDD),.Y(g9024),.A(g4358));
  NOT NOT1_3133(.VSS(VSS),.VDD(VDD),.Y(I12749),.A(g4575));
  NOT NOT1_3134(.VSS(VSS),.VDD(VDD),.Y(g11826),.A(I14650));
  NOT NOT1_3135(.VSS(VSS),.VDD(VDD),.Y(g17714),.A(g14930));
  NOT NOT1_3136(.VSS(VSS),.VDD(VDD),.Y(g12886),.A(g10393));
  NOT NOT1_3137(.VSS(VSS),.VDD(VDD),.Y(g22979),.A(g20453));
  NOT NOT1_3138(.VSS(VSS),.VDD(VDD),.Y(g20737),.A(g15656));
  NOT NOT1_3139(.VSS(VSS),.VDD(VDD),.Y(g22496),.A(g19510));
  NOT NOT1_3140(.VSS(VSS),.VDD(VDD),.Y(g10403),.A(g7040));
  NOT NOT1_3141(.VSS(VSS),.VDD(VDD),.Y(I21969),.A(g21370));
  NOT NOT1_3142(.VSS(VSS),.VDD(VDD),.Y(g23440),.A(I22557));
  NOT NOT1_3143(.VSS(VSS),.VDD(VDD),.Y(g13999),.A(g11048));
  NOT NOT1_3144(.VSS(VSS),.VDD(VDD),.Y(g7222),.A(g4427));
  NOT NOT1_3145(.VSS(VSS),.VDD(VDD),.Y(g27967),.A(I26479));
  NOT NOT1_3146(.VSS(VSS),.VDD(VDD),.Y(g27994),.A(g26793));
  NOT NOT1_3147(.VSS(VSS),.VDD(VDD),.Y(g33142),.A(g32072));
  NOT NOT1_3148(.VSS(VSS),.VDD(VDD),.Y(g19630),.A(g16897));
  NOT NOT1_3149(.VSS(VSS),.VDD(VDD),.Y(g9809),.A(g6082));
  NOT NOT1_3150(.VSS(VSS),.VDD(VDD),.Y(g20232),.A(g16931));
  NOT NOT1_3151(.VSS(VSS),.VDD(VDD),.Y(I14773),.A(g9581));
  NOT NOT1_3152(.VSS(VSS),.VDD(VDD),.Y(g29814),.A(I28062));
  NOT NOT1_3153(.VSS(VSS),.VDD(VDD),.Y(g17819),.A(I18825));
  NOT NOT1_3154(.VSS(VSS),.VDD(VDD),.Y(g17707),.A(g14758));
  NOT NOT1_3155(.VSS(VSS),.VDD(VDD),.Y(I33047),.A(g34776));
  NOT NOT1_3156(.VSS(VSS),.VDD(VDD),.Y(g30206),.A(g28436));
  NOT NOT1_3157(.VSS(VSS),.VDD(VDD),.Y(g7928),.A(g4776));
  NOT NOT1_3158(.VSS(VSS),.VDD(VDD),.Y(g26744),.A(g25400));
  NOT NOT1_3159(.VSS(VSS),.VDD(VDD),.Y(g12967),.A(g11790));
  NOT NOT1_3160(.VSS(VSS),.VDD(VDD),.Y(g23861),.A(g19147));
  NOT NOT1_3161(.VSS(VSS),.VDD(VDD),.Y(g23573),.A(g20248));
  NOT NOT1_3162(.VSS(VSS),.VDD(VDD),.Y(g32691),.A(g30673));
  NOT NOT1_3163(.VSS(VSS),.VDD(VDD),.Y(g18989),.A(g16000));
  NOT NOT1_3164(.VSS(VSS),.VDD(VDD),.Y(g8879),.A(I12858));
  NOT NOT1_3165(.VSS(VSS),.VDD(VDD),.Y(g8607),.A(g37));
  NOT NOT1_3166(.VSS(VSS),.VDD(VDD),.Y(g11233),.A(g9664));
  NOT NOT1_3167(.VSS(VSS),.VDD(VDD),.Y(I18875),.A(g13782));
  NOT NOT1_3168(.VSS(VSS),.VDD(VDD),.Y(g21247),.A(g15171));
  NOT NOT1_3169(.VSS(VSS),.VDD(VDD),.Y(g23247),.A(g20924));
  NOT NOT1_3170(.VSS(VSS),.VDD(VDD),.Y(g11182),.A(I14241));
  NOT NOT1_3171(.VSS(VSS),.VDD(VDD),.Y(I11708),.A(g3703));
  NOT NOT1_3172(.VSS(VSS),.VDD(VDD),.Y(g7064),.A(g5990));
  NOT NOT1_3173(.VSS(VSS),.VDD(VDD),.Y(g17818),.A(I18822));
  NOT NOT1_3174(.VSS(VSS),.VDD(VDD),.Y(g9672),.A(g5390));
  NOT NOT1_3175(.VSS(VSS),.VDD(VDD),.Y(I13708),.A(g136));
  NOT NOT1_3176(.VSS(VSS),.VDD(VDD),.Y(g20697),.A(g17433));
  NOT NOT1_3177(.VSS(VSS),.VDD(VDD),.Y(g14226),.A(g11618));
  NOT NOT1_3178(.VSS(VSS),.VDD(VDD),.Y(g9077),.A(g504));
  NOT NOT1_3179(.VSS(VSS),.VDD(VDD),.Y(g17496),.A(g14683));
  NOT NOT1_3180(.VSS(VSS),.VDD(VDD),.Y(I19345),.A(g15083));
  NOT NOT1_3181(.VSS(VSS),.VDD(VDD),.Y(g22986),.A(g20330));
  NOT NOT1_3182(.VSS(VSS),.VDD(VDD),.Y(g8659),.A(g2815));
  NOT NOT1_3183(.VSS(VSS),.VDD(VDD),.Y(g25882),.A(g25026));
  NOT NOT1_3184(.VSS(VSS),.VDD(VDD),.Y(g23926),.A(g19074));
  NOT NOT1_3185(.VSS(VSS),.VDD(VDD),.Y(g8358),.A(I12541));
  NOT NOT1_3186(.VSS(VSS),.VDD(VDD),.Y(g18988),.A(g15979));
  NOT NOT1_3187(.VSS(VSS),.VDD(VDD),.Y(I32775),.A(g34512));
  NOT NOT1_3188(.VSS(VSS),.VDD(VDD),.Y(g9477),.A(I13149));
  NOT NOT1_3189(.VSS(VSS),.VDD(VDD),.Y(g8506),.A(g3782));
  NOT NOT1_3190(.VSS(VSS),.VDD(VDD),.Y(I30766),.A(g32363));
  NOT NOT1_3191(.VSS(VSS),.VDD(VDD),.Y(g9523),.A(g6419));
  NOT NOT1_3192(.VSS(VSS),.VDD(VDD),.Y(g24995),.A(g22763));
  NOT NOT1_3193(.VSS(VSS),.VDD(VDD),.Y(g34759),.A(I32935));
  NOT NOT1_3194(.VSS(VSS),.VDD(VDD),.Y(g7785),.A(g4621));
  NOT NOT1_3195(.VSS(VSS),.VDD(VDD),.Y(g16522),.A(g13889));
  NOT NOT1_3196(.VSS(VSS),.VDD(VDD),.Y(g23612),.A(I22745));
  NOT NOT1_3197(.VSS(VSS),.VDD(VDD),.Y(g10572),.A(g10233));
  NOT NOT1_3198(.VSS(VSS),.VDD(VDD),.Y(I25534),.A(g25448));
  NOT NOT1_3199(.VSS(VSS),.VDD(VDD),.Y(I17964),.A(g3661));
  NOT NOT1_3200(.VSS(VSS),.VDD(VDD),.Y(g23388),.A(g21070));
  NOT NOT1_3201(.VSS(VSS),.VDD(VDD),.Y(I15932),.A(g12381));
  NOT NOT1_3202(.VSS(VSS),.VDD(VDD),.Y(g17590),.A(I18523));
  NOT NOT1_3203(.VSS(VSS),.VDD(VDD),.Y(g19476),.A(g16326));
  NOT NOT1_3204(.VSS(VSS),.VDD(VDD),.Y(g12919),.A(I15536));
  NOT NOT1_3205(.VSS(VSS),.VDD(VDD),.Y(I12808),.A(g4322));
  NOT NOT1_3206(.VSS(VSS),.VDD(VDD),.Y(g6799),.A(g199));
  NOT NOT1_3207(.VSS(VSS),.VDD(VDD),.Y(g26804),.A(g25400));
  NOT NOT1_3208(.VSS(VSS),.VDD(VDD),.Y(g20512),.A(g18062));
  NOT NOT1_3209(.VSS(VSS),.VDD(VDD),.Y(g34435),.A(I32476));
  NOT NOT1_3210(.VSS(VSS),.VDD(VDD),.Y(g23777),.A(I22918));
  NOT NOT1_3211(.VSS(VSS),.VDD(VDD),.Y(g23534),.A(I22665));
  NOT NOT1_3212(.VSS(VSS),.VDD(VDD),.Y(I26451),.A(g26862));
  NOT NOT1_3213(.VSS(VSS),.VDD(VDD),.Y(g13932),.A(g11534));
  NOT NOT1_3214(.VSS(VSS),.VDD(VDD),.Y(g32929),.A(g31710));
  NOT NOT1_3215(.VSS(VSS),.VDD(VDD),.Y(g8587),.A(g3689));
  NOT NOT1_3216(.VSS(VSS),.VDD(VDD),.Y(I14839),.A(g9689));
  NOT NOT1_3217(.VSS(VSS),.VDD(VDD),.Y(g23272),.A(g20924));
  NOT NOT1_3218(.VSS(VSS),.VDD(VDD),.Y(g11513),.A(g7948));
  NOT NOT1_3219(.VSS(VSS),.VDD(VDD),.Y(g19454),.A(g16349));
  NOT NOT1_3220(.VSS(VSS),.VDD(VDD),.Y(g7563),.A(g6322));
  NOT NOT1_3221(.VSS(VSS),.VDD(VDD),.Y(g17741),.A(g12972));
  NOT NOT1_3222(.VSS(VSS),.VDD(VDD),.Y(g12918),.A(I15533));
  NOT NOT1_3223(.VSS(VSS),.VDD(VDD),.Y(I18160),.A(g14441));
  NOT NOT1_3224(.VSS(VSS),.VDD(VDD),.Y(I15448),.A(g10877));
  NOT NOT1_3225(.VSS(VSS),.VDD(VDD),.Y(g17384),.A(I18323));
  NOT NOT1_3226(.VSS(VSS),.VDD(VDD),.Y(g32583),.A(g30614));
  NOT NOT1_3227(.VSS(VSS),.VDD(VDD),.Y(g32928),.A(g31672));
  NOT NOT1_3228(.VSS(VSS),.VDD(VDD),.Y(g19570),.A(g16349));
  NOT NOT1_3229(.VSS(VSS),.VDD(VDD),.Y(g19712),.A(g17096));
  NOT NOT1_3230(.VSS(VSS),.VDD(VDD),.Y(g6997),.A(g4578));
  NOT NOT1_3231(.VSS(VSS),.VDD(VDD),.Y(g22150),.A(g21280));
  NOT NOT1_3232(.VSS(VSS),.VDD(VDD),.Y(g11897),.A(I14705));
  NOT NOT1_3233(.VSS(VSS),.VDD(VDD),.Y(I22000),.A(g20277));
  NOT NOT1_3234(.VSS(VSS),.VDD(VDD),.Y(g10490),.A(g9274));
  NOT NOT1_3235(.VSS(VSS),.VDD(VDD),.Y(g9551),.A(g3281));
  NOT NOT1_3236(.VSS(VSS),.VDD(VDD),.Y(g9742),.A(g6144));
  NOT NOT1_3237(.VSS(VSS),.VDD(VDD),.Y(g9104),.A(I12987));
  NOT NOT1_3238(.VSS(VSS),.VDD(VDD),.Y(g23462),.A(I22589));
  NOT NOT1_3239(.VSS(VSS),.VDD(VDD),.Y(g9099),.A(g3706));
  NOT NOT1_3240(.VSS(VSS),.VDD(VDD),.Y(g34345),.A(I32352));
  NOT NOT1_3241(.VSS(VSS),.VDD(VDD),.Y(g9499),.A(g5152));
  NOT NOT1_3242(.VSS(VSS),.VDD(VDD),.Y(g11404),.A(g7596));
  NOT NOT1_3243(.VSS(VSS),.VDD(VDD),.Y(g15750),.A(g13291));
  NOT NOT1_3244(.VSS(VSS),.VDD(VDD),.Y(g34940),.A(g34924));
  NOT NOT1_3245(.VSS(VSS),.VDD(VDD),.Y(g13505),.A(g10981));
  NOT NOT1_3246(.VSS(VSS),.VDD(VDD),.Y(I15717),.A(g6346));
  NOT NOT1_3247(.VSS(VSS),.VDD(VDD),.Y(g16326),.A(I17658));
  NOT NOT1_3248(.VSS(VSS),.VDD(VDD),.Y(g18887),.A(g15373));
  NOT NOT1_3249(.VSS(VSS),.VDD(VDD),.Y(g20445),.A(g15224));
  NOT NOT1_3250(.VSS(VSS),.VDD(VDD),.Y(I31820),.A(g33323));
  NOT NOT1_3251(.VSS(VSS),.VDD(VDD),.Y(I12064),.A(g617));
  NOT NOT1_3252(.VSS(VSS),.VDD(VDD),.Y(g23032),.A(I22211));
  NOT NOT1_3253(.VSS(VSS),.VDD(VDD),.Y(g10376),.A(g6923));
  NOT NOT1_3254(.VSS(VSS),.VDD(VDD),.Y(g10385),.A(I13805));
  NOT NOT1_3255(.VSS(VSS),.VDD(VDD),.Y(g25206),.A(g23613));
  NOT NOT1_3256(.VSS(VSS),.VDD(VDD),.Y(g12598),.A(g7004));
  NOT NOT1_3257(.VSS(VSS),.VDD(VDD),.Y(g14376),.A(g12126));
  NOT NOT1_3258(.VSS(VSS),.VDD(VDD),.Y(g14385),.A(I16541));
  NOT NOT1_3259(.VSS(VSS),.VDD(VDD),.Y(g34848),.A(I33070));
  NOT NOT1_3260(.VSS(VSS),.VDD(VDD),.Y(g19074),.A(I19772));
  NOT NOT1_3261(.VSS(VSS),.VDD(VDD),.Y(g17735),.A(g14807));
  NOT NOT1_3262(.VSS(VSS),.VDD(VDD),.Y(g14297),.A(g10869));
  NOT NOT1_3263(.VSS(VSS),.VDD(VDD),.Y(g20499),.A(g15483));
  NOT NOT1_3264(.VSS(VSS),.VDD(VDD),.Y(g7394),.A(g5637));
  NOT NOT1_3265(.VSS(VSS),.VDD(VDD),.Y(g10980),.A(g9051));
  NOT NOT1_3266(.VSS(VSS),.VDD(VDD),.Y(g11026),.A(g8434));
  NOT NOT1_3267(.VSS(VSS),.VDD(VDD),.Y(I26785),.A(g27013));
  NOT NOT1_3268(.VSS(VSS),.VDD(VDD),.Y(g12086),.A(g9654));
  NOT NOT1_3269(.VSS(VSS),.VDD(VDD),.Y(g32787),.A(g30937));
  NOT NOT1_3270(.VSS(VSS),.VDD(VDD),.Y(g13026),.A(g11018));
  NOT NOT1_3271(.VSS(VSS),.VDD(VDD),.Y(g31863),.A(I29447));
  NOT NOT1_3272(.VSS(VSS),.VDD(VDD),.Y(I14619),.A(g4185));
  NOT NOT1_3273(.VSS(VSS),.VDD(VDD),.Y(g10354),.A(g6811));
  NOT NOT1_3274(.VSS(VSS),.VDD(VDD),.Y(I23315),.A(g21685));
  NOT NOT1_3275(.VSS(VSS),.VDD(VDD),.Y(I33152),.A(g34900));
  NOT NOT1_3276(.VSS(VSS),.VDD(VDD),.Y(g19567),.A(g16164));
  NOT NOT1_3277(.VSS(VSS),.VDD(VDD),.Y(g14095),.A(g11326));
  NOT NOT1_3278(.VSS(VSS),.VDD(VDD),.Y(g29014),.A(g27742));
  NOT NOT1_3279(.VSS(VSS),.VDD(VDD),.Y(g22526),.A(g19801));
  NOT NOT1_3280(.VSS(VSS),.VDD(VDD),.Y(I17569),.A(g14564));
  NOT NOT1_3281(.VSS(VSS),.VDD(VDD),.Y(g9754),.A(g2020));
  NOT NOT1_3282(.VSS(VSS),.VDD(VDD),.Y(g21061),.A(I20929));
  NOT NOT1_3283(.VSS(VSS),.VDD(VDD),.Y(g28126),.A(g27122));
  NOT NOT1_3284(.VSS(VSS),.VDD(VDD),.Y(g18528),.A(I19348));
  NOT NOT1_3285(.VSS(VSS),.VDD(VDD),.Y(g20498),.A(g15348));
  NOT NOT1_3286(.VSS(VSS),.VDD(VDD),.Y(g6802),.A(g468));
  NOT NOT1_3287(.VSS(VSS),.VDD(VDD),.Y(g8284),.A(g5002));
  NOT NOT1_3288(.VSS(VSS),.VDD(VDD),.Y(g23061),.A(g20283));
  NOT NOT1_3289(.VSS(VSS),.VDD(VDD),.Y(g8239),.A(g1056));
  NOT NOT1_3290(.VSS(VSS),.VDD(VDD),.Y(g28250),.A(g27074));
  NOT NOT1_3291(.VSS(VSS),.VDD(VDD),.Y(g10181),.A(g2551));
  NOT NOT1_3292(.VSS(VSS),.VDD(VDD),.Y(g25114),.A(I24278));
  NOT NOT1_3293(.VSS(VSS),.VDD(VDD),.Y(g7557),.A(g1500));
  NOT NOT1_3294(.VSS(VSS),.VDD(VDD),.Y(g8180),.A(g262));
  NOT NOT1_3295(.VSS(VSS),.VDD(VDD),.Y(I17747),.A(g13298));
  NOT NOT1_3296(.VSS(VSS),.VDD(VDD),.Y(g12322),.A(I15162));
  NOT NOT1_3297(.VSS(VSS),.VDD(VDD),.Y(g27977),.A(g26105));
  NOT NOT1_3298(.VSS(VSS),.VDD(VDD),.Y(g32743),.A(g30937));
  NOT NOT1_3299(.VSS(VSS),.VDD(VDD),.Y(g32827),.A(g31672));
  NOT NOT1_3300(.VSS(VSS),.VDD(VDD),.Y(g25082),.A(g22342));
  NOT NOT1_3301(.VSS(VSS),.VDD(VDD),.Y(g8591),.A(g3763));
  NOT NOT1_3302(.VSS(VSS),.VDD(VDD),.Y(g30332),.A(I28597));
  NOT NOT1_3303(.VSS(VSS),.VDD(VDD),.Y(g24056),.A(g20014));
  NOT NOT1_3304(.VSS(VSS),.VDD(VDD),.Y(g9613),.A(g5062));
  NOT NOT1_3305(.VSS(VSS),.VDD(VDD),.Y(g12901),.A(g10404));
  NOT NOT1_3306(.VSS(VSS),.VDD(VDD),.Y(g20611),.A(g18008));
  NOT NOT1_3307(.VSS(VSS),.VDD(VDD),.Y(g17526),.A(I18469));
  NOT NOT1_3308(.VSS(VSS),.VDD(VDD),.Y(g12977),.A(I15590));
  NOT NOT1_3309(.VSS(VSS),.VDD(VDD),.Y(g20080),.A(g17328));
  NOT NOT1_3310(.VSS(VSS),.VDD(VDD),.Y(g7471),.A(g6012));
  NOT NOT1_3311(.VSS(VSS),.VDD(VDD),.Y(g9044),.A(g604));
  NOT NOT1_3312(.VSS(VSS),.VDD(VDD),.Y(g20924),.A(I20895));
  NOT NOT1_3313(.VSS(VSS),.VDD(VDD),.Y(g19519),.A(g16795));
  NOT NOT1_3314(.VSS(VSS),.VDD(VDD),.Y(g24080),.A(g21143));
  NOT NOT1_3315(.VSS(VSS),.VDD(VDD),.Y(g19675),.A(g16987));
  NOT NOT1_3316(.VSS(VSS),.VDD(VDD),.Y(g9444),.A(g5535));
  NOT NOT1_3317(.VSS(VSS),.VDD(VDD),.Y(g9269),.A(g5517));
  NOT NOT1_3318(.VSS(VSS),.VDD(VDD),.Y(g22866),.A(g20330));
  NOT NOT1_3319(.VSS(VSS),.VDD(VDD),.Y(I17814),.A(g3274));
  NOT NOT1_3320(.VSS(VSS),.VDD(VDD),.Y(g32640),.A(g31154));
  NOT NOT1_3321(.VSS(VSS),.VDD(VDD),.Y(g20432),.A(g17847));
  NOT NOT1_3322(.VSS(VSS),.VDD(VDD),.Y(g32769),.A(g31672));
  NOT NOT1_3323(.VSS(VSS),.VDD(VDD),.Y(g23360),.A(I22461));
  NOT NOT1_3324(.VSS(VSS),.VDD(VDD),.Y(g29116),.A(g27837));
  NOT NOT1_3325(.VSS(VSS),.VDD(VDD),.Y(g19518),.A(g16239));
  NOT NOT1_3326(.VSS(VSS),.VDD(VDD),.Y(g8507),.A(g3712));
  NOT NOT1_3327(.VSS(VSS),.VDD(VDD),.Y(g9983),.A(g4239));
  NOT NOT1_3328(.VSS(VSS),.VDD(VDD),.Y(g12656),.A(g7028));
  NOT NOT1_3329(.VSS(VSS),.VDD(VDD),.Y(I15620),.A(g12038));
  NOT NOT1_3330(.VSS(VSS),.VDD(VDD),.Y(I17772),.A(g14888));
  NOT NOT1_3331(.VSS(VSS),.VDD(VDD),.Y(g25849),.A(g24491));
  NOT NOT1_3332(.VSS(VSS),.VDD(VDD),.Y(g9862),.A(g5413));
  NOT NOT1_3333(.VSS(VSS),.VDD(VDD),.Y(I27555),.A(g28142));
  NOT NOT1_3334(.VSS(VSS),.VDD(VDD),.Y(g23447),.A(g21562));
  NOT NOT1_3335(.VSS(VSS),.VDD(VDD),.Y(g32768),.A(g30825));
  NOT NOT1_3336(.VSS(VSS),.VDD(VDD),.Y(g32803),.A(g31376));
  NOT NOT1_3337(.VSS(VSS),.VDD(VDD),.Y(g25399),.A(g22763));
  NOT NOT1_3338(.VSS(VSS),.VDD(VDD),.Y(g12295),.A(g7139));
  NOT NOT1_3339(.VSS(VSS),.VDD(VDD),.Y(I23384),.A(g23362));
  NOT NOT1_3340(.VSS(VSS),.VDD(VDD),.Y(g10190),.A(g6044));
  NOT NOT1_3341(.VSS(VSS),.VDD(VDD),.Y(g29041),.A(I27385));
  NOT NOT1_3342(.VSS(VSS),.VDD(VDD),.Y(g13620),.A(g10556));
  NOT NOT1_3343(.VSS(VSS),.VDD(VDD),.Y(g12823),.A(g9206));
  NOT NOT1_3344(.VSS(VSS),.VDD(VDD),.Y(I17639),.A(g13350));
  NOT NOT1_3345(.VSS(VSS),.VDD(VDD),.Y(I27570),.A(g28262));
  NOT NOT1_3346(.VSS(VSS),.VDD(VDD),.Y(I15811),.A(g11128));
  NOT NOT1_3347(.VSS(VSS),.VDD(VDD),.Y(I21067),.A(g15573));
  NOT NOT1_3348(.VSS(VSS),.VDD(VDD),.Y(I18822),.A(g13745));
  NOT NOT1_3349(.VSS(VSS),.VDD(VDD),.Y(g16509),.A(g13873));
  NOT NOT1_3350(.VSS(VSS),.VDD(VDD),.Y(I32056),.A(g33641));
  NOT NOT1_3351(.VSS(VSS),.VDD(VDD),.Y(g11811),.A(g9724));
  NOT NOT1_3352(.VSS(VSS),.VDD(VDD),.Y(I12712),.A(g59));
  NOT NOT1_3353(.VSS(VSS),.VDD(VDD),.Y(g20145),.A(g17533));
  NOT NOT1_3354(.VSS(VSS),.VDD(VDD),.Y(g34833),.A(I33047));
  NOT NOT1_3355(.VSS(VSS),.VDD(VDD),.Y(g34049),.A(g33678));
  NOT NOT1_3356(.VSS(VSS),.VDD(VDD),.Y(I13010),.A(g6749));
  NOT NOT1_3357(.VSS(VSS),.VDD(VDD),.Y(g31821),.A(g29385));
  NOT NOT1_3358(.VSS(VSS),.VDD(VDD),.Y(g32881),.A(g30673));
  NOT NOT1_3359(.VSS(VSS),.VDD(VDD),.Y(I32988),.A(g34755));
  NOT NOT1_3360(.VSS(VSS),.VDD(VDD),.Y(g24031),.A(g21193));
  NOT NOT1_3361(.VSS(VSS),.VDD(VDD),.Y(I33020),.A(g34781));
  NOT NOT1_3362(.VSS(VSS),.VDD(VDD),.Y(g16508),.A(I17704));
  NOT NOT1_3363(.VSS(VSS),.VDD(VDD),.Y(I24455),.A(g22541));
  NOT NOT1_3364(.VSS(VSS),.VDD(VDD),.Y(g26605),.A(g25293));
  NOT NOT1_3365(.VSS(VSS),.VDD(VDD),.Y(g20650),.A(g15348));
  NOT NOT1_3366(.VSS(VSS),.VDD(VDD),.Y(g23629),.A(g21514));
  NOT NOT1_3367(.VSS(VSS),.VDD(VDD),.Y(g21451),.A(I21162));
  NOT NOT1_3368(.VSS(VSS),.VDD(VDD),.Y(g16872),.A(I18060));
  NOT NOT1_3369(.VSS(VSS),.VDD(VDD),.Y(I12907),.A(g4322));
  NOT NOT1_3370(.VSS(VSS),.VDD(VDD),.Y(g22923),.A(I22124));
  NOT NOT1_3371(.VSS(VSS),.VDD(VDD),.Y(I17416),.A(g13806));
  NOT NOT1_3372(.VSS(VSS),.VDD(VDD),.Y(g23472),.A(g21062));
  NOT NOT1_3373(.VSS(VSS),.VDD(VDD),.Y(g15483),.A(I17128));
  NOT NOT1_3374(.VSS(VSS),.VDD(VDD),.Y(g9534),.A(g90));
  NOT NOT1_3375(.VSS(VSS),.VDD(VDD),.Y(g9729),.A(g5138));
  NOT NOT1_3376(.VSS(VSS),.VDD(VDD),.Y(g9961),.A(g6404));
  NOT NOT1_3377(.VSS(VSS),.VDD(VDD),.Y(g7438),.A(g5983));
  NOT NOT1_3378(.VSS(VSS),.VDD(VDD),.Y(g25263),.A(g22763));
  NOT NOT1_3379(.VSS(VSS),.VDD(VDD),.Y(g29983),.A(g28977));
  NOT NOT1_3380(.VSS(VSS),.VDD(VDD),.Y(g20529),.A(g15509));
  NOT NOT1_3381(.VSS(VSS),.VDD(VDD),.Y(g22300),.A(I21815));
  NOT NOT1_3382(.VSS(VSS),.VDD(VDD),.Y(g26812),.A(g25439));
  NOT NOT1_3383(.VSS(VSS),.VDD(VDD),.Y(I21019),.A(g17325));
  NOT NOT1_3384(.VSS(VSS),.VDD(VDD),.Y(g27017),.A(g25895));
  NOT NOT1_3385(.VSS(VSS),.VDD(VDD),.Y(I27567),.A(g28181));
  NOT NOT1_3386(.VSS(VSS),.VDD(VDD),.Y(g15862),.A(I17355));
  NOT NOT1_3387(.VSS(VSS),.VDD(VDD),.Y(g8515),.A(I12631));
  NOT NOT1_3388(.VSS(VSS),.VDD(VDD),.Y(g34221),.A(I32192));
  NOT NOT1_3389(.VSS(VSS),.VDD(VDD),.Y(g8630),.A(g4843));
  NOT NOT1_3390(.VSS(VSS),.VDD(VDD),.Y(g21246),.A(I20985));
  NOT NOT1_3391(.VSS(VSS),.VDD(VDD),.Y(I27238),.A(g27320));
  NOT NOT1_3392(.VSS(VSS),.VDD(VDD),.Y(g23246),.A(g20785));
  NOT NOT1_3393(.VSS(VSS),.VDD(VDD),.Y(g20528),.A(g15224));
  NOT NOT1_3394(.VSS(VSS),.VDD(VDD),.Y(g20696),.A(g17533));
  NOT NOT1_3395(.VSS(VSS),.VDD(VDD),.Y(g25135),.A(g22457));
  NOT NOT1_3396(.VSS(VSS),.VDD(VDD),.Y(g20330),.A(I20542));
  NOT NOT1_3397(.VSS(VSS),.VDD(VDD),.Y(g9927),.A(g5689));
  NOT NOT1_3398(.VSS(VSS),.VDD(VDD),.Y(g32662),.A(g30614));
  NOT NOT1_3399(.VSS(VSS),.VDD(VDD),.Y(g8300),.A(g1242));
  NOT NOT1_3400(.VSS(VSS),.VDD(VDD),.Y(g32027),.A(I29585));
  NOT NOT1_3401(.VSS(VSS),.VDD(VDD),.Y(I32461),.A(g34244));
  NOT NOT1_3402(.VSS(VSS),.VDD(VDD),.Y(g19577),.A(g16129));
  NOT NOT1_3403(.VSS(VSS),.VDD(VDD),.Y(g17688),.A(I18667));
  NOT NOT1_3404(.VSS(VSS),.VDD(VDD),.Y(g9014),.A(g3004));
  NOT NOT1_3405(.VSS(VSS),.VDD(VDD),.Y(g20764),.A(I20819));
  NOT NOT1_3406(.VSS(VSS),.VDD(VDD),.Y(g10497),.A(g10102));
  NOT NOT1_3407(.VSS(VSS),.VDD(VDD),.Y(I25591),.A(g25380));
  NOT NOT1_3408(.VSS(VSS),.VDD(VDD),.Y(g32890),.A(g30735));
  NOT NOT1_3409(.VSS(VSS),.VDD(VDD),.Y(I33282),.A(g34987));
  NOT NOT1_3410(.VSS(VSS),.VDD(VDD),.Y(I27941),.A(g28803));
  NOT NOT1_3411(.VSS(VSS),.VDD(VDD),.Y(g9414),.A(g2004));
  NOT NOT1_3412(.VSS(VSS),.VDD(VDD),.Y(g7212),.A(g6411));
  NOT NOT1_3413(.VSS(VSS),.VDD(VDD),.Y(g19439),.A(g15885));
  NOT NOT1_3414(.VSS(VSS),.VDD(VDD),.Y(g9660),.A(g3267));
  NOT NOT1_3415(.VSS(VSS),.VDD(VDD),.Y(g9946),.A(g6093));
  NOT NOT1_3416(.VSS(VSS),.VDD(VDD),.Y(g20132),.A(g16931));
  NOT NOT1_3417(.VSS(VSS),.VDD(VDD),.Y(g24365),.A(g22594));
  NOT NOT1_3418(.VSS(VSS),.VDD(VDD),.Y(g20869),.A(g15615));
  NOT NOT1_3419(.VSS(VSS),.VDD(VDD),.Y(g13412),.A(g11963));
  NOT NOT1_3420(.VSS(VSS),.VDD(VDD),.Y(g23776),.A(g21177));
  NOT NOT1_3421(.VSS(VSS),.VDD(VDD),.Y(g34947),.A(g34938));
  NOT NOT1_3422(.VSS(VSS),.VDD(VDD),.Y(I12382),.A(g47));
  NOT NOT1_3423(.VSS(VSS),.VDD(VDD),.Y(g24132),.A(g19890));
  NOT NOT1_3424(.VSS(VSS),.VDD(VDD),.Y(g32482),.A(g30614));
  NOT NOT1_3425(.VSS(VSS),.VDD(VDD),.Y(g24869),.A(I24041));
  NOT NOT1_3426(.VSS(VSS),.VDD(VDD),.Y(g24960),.A(g23716));
  NOT NOT1_3427(.VSS(VSS),.VDD(VDD),.Y(g19438),.A(g16249));
  NOT NOT1_3428(.VSS(VSS),.VDD(VDD),.Y(I12519),.A(g3447));
  NOT NOT1_3429(.VSS(VSS),.VDD(VDD),.Y(g17157),.A(g13350));
  NOT NOT1_3430(.VSS(VSS),.VDD(VDD),.Y(I12176),.A(g5523));
  NOT NOT1_3431(.VSS(VSS),.VDD(VDD),.Y(g9903),.A(g681));
  NOT NOT1_3432(.VSS(VSS),.VDD(VDD),.Y(g13133),.A(g11330));
  NOT NOT1_3433(.VSS(VSS),.VDD(VDD),.Y(g32710),.A(g30825));
  NOT NOT1_3434(.VSS(VSS),.VDD(VDD),.Y(I12092),.A(g790));
  NOT NOT1_3435(.VSS(VSS),.VDD(VDD),.Y(g14700),.A(g12512));
  NOT NOT1_3436(.VSS(VSS),.VDD(VDD),.Y(g21355),.A(g17821));
  NOT NOT1_3437(.VSS(VSS),.VDD(VDD),.Y(g32552),.A(g30825));
  NOT NOT1_3438(.VSS(VSS),.VDD(VDD),.Y(g31834),.A(g29385));
  NOT NOT1_3439(.VSS(VSS),.VDD(VDD),.Y(g23355),.A(g21070));
  NOT NOT1_3440(.VSS(VSS),.VDD(VDD),.Y(g34812),.A(I33024));
  NOT NOT1_3441(.VSS(VSS),.VDD(VDD),.Y(g10658),.A(I13979));
  NOT NOT1_3442(.VSS(VSS),.VDD(VDD),.Y(g21370),.A(g16323));
  NOT NOT1_3443(.VSS(VSS),.VDD(VDD),.Y(g23859),.A(g19074));
  NOT NOT1_3444(.VSS(VSS),.VDD(VDD),.Y(g28819),.A(I27271));
  NOT NOT1_3445(.VSS(VSS),.VDD(VDD),.Y(g16311),.A(g13273));
  NOT NOT1_3446(.VSS(VSS),.VDD(VDD),.Y(g32779),.A(g30937));
  NOT NOT1_3447(.VSS(VSS),.VDD(VDD),.Y(I17442),.A(g13638));
  NOT NOT1_3448(.VSS(VSS),.VDD(VDD),.Y(g18878),.A(g15426));
  NOT NOT1_3449(.VSS(VSS),.VDD(VDD),.Y(g24161),.A(I23327));
  NOT NOT1_3450(.VSS(VSS),.VDD(VDD),.Y(g29130),.A(g27907));
  NOT NOT1_3451(.VSS(VSS),.VDD(VDD),.Y(I32696),.A(g34434));
  NOT NOT1_3452(.VSS(VSS),.VDD(VDD),.Y(I32843),.A(g34499));
  NOT NOT1_3453(.VSS(VSS),.VDD(VDD),.Y(g7993),.A(I12333));
  NOT NOT1_3454(.VSS(VSS),.VDD(VDD),.Y(g20709),.A(g15426));
  NOT NOT1_3455(.VSS(VSS),.VDD(VDD),.Y(g11011),.A(g10274));
  NOT NOT1_3456(.VSS(VSS),.VDD(VDD),.Y(g22854),.A(g20330));
  NOT NOT1_3457(.VSS(VSS),.VDD(VDD),.Y(g34951),.A(g34941));
  NOT NOT1_3458(.VSS(VSS),.VDD(VDD),.Y(g34972),.A(I33232));
  NOT NOT1_3459(.VSS(VSS),.VDD(VDD),.Y(g23858),.A(g18997));
  NOT NOT1_3460(.VSS(VSS),.VDD(VDD),.Y(g13011),.A(I15623));
  NOT NOT1_3461(.VSS(VSS),.VDD(VDD),.Y(I12935),.A(g6753));
  NOT NOT1_3462(.VSS(VSS),.VDD(VDD),.Y(g32778),.A(g31021));
  NOT NOT1_3463(.VSS(VSS),.VDD(VDD),.Y(g18886),.A(g16000));
  NOT NOT1_3464(.VSS(VSS),.VDD(VDD),.Y(I31803),.A(g33176));
  NOT NOT1_3465(.VSS(VSS),.VDD(VDD),.Y(g9036),.A(g5084));
  NOT NOT1_3466(.VSS(VSS),.VDD(VDD),.Y(I18313),.A(g13350));
  NOT NOT1_3467(.VSS(VSS),.VDD(VDD),.Y(g25221),.A(g23653));
  NOT NOT1_3468(.VSS(VSS),.VDD(VDD),.Y(I22275),.A(g20127));
  NOT NOT1_3469(.VSS(VSS),.VDD(VDD),.Y(g8440),.A(g3431));
  NOT NOT1_3470(.VSS(VSS),.VDD(VDD),.Y(g20708),.A(g15426));
  NOT NOT1_3471(.VSS(VSS),.VDD(VDD),.Y(g22763),.A(I22046));
  NOT NOT1_3472(.VSS(VSS),.VDD(VDD),.Y(g9679),.A(g5475));
  NOT NOT1_3473(.VSS(VSS),.VDD(VDD),.Y(g23172),.A(I22275));
  NOT NOT1_3474(.VSS(VSS),.VDD(VDD),.Y(g13716),.A(I16090));
  NOT NOT1_3475(.VSS(VSS),.VDD(VDD),.Y(I17615),.A(g13251));
  NOT NOT1_3476(.VSS(VSS),.VDD(VDD),.Y(g20087),.A(g17249));
  NOT NOT1_3477(.VSS(VSS),.VDD(VDD),.Y(g32786),.A(g31021));
  NOT NOT1_3478(.VSS(VSS),.VDD(VDD),.Y(g33726),.A(I31581));
  NOT NOT1_3479(.VSS(VSS),.VDD(VDD),.Y(I32960),.A(g34653));
  NOT NOT1_3480(.VSS(VSS),.VDD(VDD),.Y(g8123),.A(g3808));
  NOT NOT1_3481(.VSS(VSS),.VDD(VDD),.Y(g19566),.A(g16136));
  NOT NOT1_3482(.VSS(VSS),.VDD(VDD),.Y(g14338),.A(I16502));
  NOT NOT1_3483(.VSS(VSS),.VDD(VDD),.Y(g24087),.A(g21143));
  NOT NOT1_3484(.VSS(VSS),.VDD(VDD),.Y(I18276),.A(g1075));
  NOT NOT1_3485(.VSS(VSS),.VDD(VDD),.Y(I18285),.A(g13638));
  NOT NOT1_3486(.VSS(VSS),.VDD(VDD),.Y(g28590),.A(g27724));
  NOT NOT1_3487(.VSS(VSS),.VDD(VDD),.Y(g23844),.A(g21308));
  NOT NOT1_3488(.VSS(VSS),.VDD(VDD),.Y(g32647),.A(g31154));
  NOT NOT1_3489(.VSS(VSS),.VDD(VDD),.Y(g23394),.A(I22499));
  NOT NOT1_3490(.VSS(VSS),.VDD(VDD),.Y(I32868),.A(g34579));
  NOT NOT1_3491(.VSS(VSS),.VDD(VDD),.Y(g9831),.A(g2269));
  NOT NOT1_3492(.VSS(VSS),.VDD(VDD),.Y(g32945),.A(g30937));
  NOT NOT1_3493(.VSS(VSS),.VDD(VDD),.Y(g33436),.A(I30962));
  NOT NOT1_3494(.VSS(VSS),.VDD(VDD),.Y(g22660),.A(g19140));
  NOT NOT1_3495(.VSS(VSS),.VDD(VDD),.Y(g15509),.A(I17136));
  NOT NOT1_3496(.VSS(VSS),.VDD(VDD),.Y(I19012),.A(g15060));
  NOT NOT1_3497(.VSS(VSS),.VDD(VDD),.Y(g17763),.A(g15011));
  NOT NOT1_3498(.VSS(VSS),.VDD(VDD),.Y(g8666),.A(g3703));
  NOT NOT1_3499(.VSS(VSS),.VDD(VDD),.Y(g10060),.A(g6541));
  NOT NOT1_3500(.VSS(VSS),.VDD(VDD),.Y(I18900),.A(g16767));
  NOT NOT1_3501(.VSS(VSS),.VDD(VDD),.Y(g27976),.A(g26703));
  NOT NOT1_3502(.VSS(VSS),.VDD(VDD),.Y(g27985),.A(g26131));
  NOT NOT1_3503(.VSS(VSS),.VDD(VDD),.Y(I32161),.A(g33791));
  NOT NOT1_3504(.VSS(VSS),.VDD(VDD),.Y(g32826),.A(g30825));
  NOT NOT1_3505(.VSS(VSS),.VDD(VDD),.Y(g25273),.A(g23978));
  NOT NOT1_3506(.VSS(VSS),.VDD(VDD),.Y(g29863),.A(g28410));
  NOT NOT1_3507(.VSS(VSS),.VDD(VDD),.Y(g24043),.A(g20982));
  NOT NOT1_3508(.VSS(VSS),.VDD(VDD),.Y(g10197),.A(g31));
  NOT NOT1_3509(.VSS(VSS),.VDD(VDD),.Y(I21300),.A(g18598));
  NOT NOT1_3510(.VSS(VSS),.VDD(VDD),.Y(g22456),.A(g19801));
  NOT NOT1_3511(.VSS(VSS),.VDD(VDD),.Y(g12976),.A(I15587));
  NOT NOT1_3512(.VSS(VSS),.VDD(VDD),.Y(g15634),.A(I17188));
  NOT NOT1_3513(.VSS(VSS),.VDD(VDD),.Y(I23688),.A(g23244));
  NOT NOT1_3514(.VSS(VSS),.VDD(VDD),.Y(I23300),.A(g21665));
  NOT NOT1_3515(.VSS(VSS),.VDD(VDD),.Y(g14197),.A(g12160));
  NOT NOT1_3516(.VSS(VSS),.VDD(VDD),.Y(g32090),.A(g31003));
  NOT NOT1_3517(.VSS(VSS),.VDD(VDD),.Y(g9805),.A(g5485));
  NOT NOT1_3518(.VSS(VSS),.VDD(VDD),.Y(g9916),.A(g3625));
  NOT NOT1_3519(.VSS(VSS),.VDD(VDD),.Y(g19653),.A(g16897));
  NOT NOT1_3520(.VSS(VSS),.VDD(VDD),.Y(g33346),.A(g32132));
  NOT NOT1_3521(.VSS(VSS),.VDD(VDD),.Y(I18101),.A(g13416));
  NOT NOT1_3522(.VSS(VSS),.VDD(VDD),.Y(I32225),.A(g34121));
  NOT NOT1_3523(.VSS(VSS),.VDD(VDD),.Y(g10527),.A(I13892));
  NOT NOT1_3524(.VSS(VSS),.VDD(VDD),.Y(I12577),.A(g1227));
  NOT NOT1_3525(.VSS(VSS),.VDD(VDD),.Y(g10411),.A(g7086));
  NOT NOT1_3526(.VSS(VSS),.VDD(VDD),.Y(g23420),.A(g21514));
  NOT NOT1_3527(.VSS(VSS),.VDD(VDD),.Y(g9749),.A(g1691));
  NOT NOT1_3528(.VSS(VSS),.VDD(VDD),.Y(I18177),.A(g13191));
  NOT NOT1_3529(.VSS(VSS),.VDD(VDD),.Y(I18560),.A(g5969));
  NOT NOT1_3530(.VSS(VSS),.VDD(VDD),.Y(g32651),.A(g31376));
  NOT NOT1_3531(.VSS(VSS),.VDD(VDD),.Y(g18918),.A(I19704));
  NOT NOT1_3532(.VSS(VSS),.VDD(VDD),.Y(g32672),.A(g31579));
  NOT NOT1_3533(.VSS(VSS),.VDD(VDD),.Y(I19789),.A(g17793));
  NOT NOT1_3534(.VSS(VSS),.VDD(VDD),.Y(g24069),.A(g19968));
  NOT NOT1_3535(.VSS(VSS),.VDD(VDD),.Y(g22550),.A(I21922));
  NOT NOT1_3536(.VSS(VSS),.VDD(VDD),.Y(I33027),.A(g34767));
  NOT NOT1_3537(.VSS(VSS),.VDD(VDD),.Y(g26788),.A(g25349));
  NOT NOT1_3538(.VSS(VSS),.VDD(VDD),.Y(g26724),.A(g25341));
  NOT NOT1_3539(.VSS(VSS),.VDD(VDD),.Y(g20657),.A(g17433));
  NOT NOT1_3540(.VSS(VSS),.VDD(VDD),.Y(g20774),.A(g18008));
  NOT NOT1_3541(.VSS(VSS),.VDD(VDD),.Y(I26427),.A(g26859));
  NOT NOT1_3542(.VSS(VSS),.VDD(VDD),.Y(g8655),.A(g2787));
  NOT NOT1_3543(.VSS(VSS),.VDD(VDD),.Y(g23446),.A(g21562));
  NOT NOT1_3544(.VSS(VSS),.VDD(VDD),.Y(I16057),.A(g10430));
  NOT NOT1_3545(.VSS(VSS),.VDD(VDD),.Y(I28908),.A(g30182));
  NOT NOT1_3546(.VSS(VSS),.VDD(VDD),.Y(g19636),.A(g16987));
  NOT NOT1_3547(.VSS(VSS),.VDD(VDD),.Y(g23227),.A(g20924));
  NOT NOT1_3548(.VSS(VSS),.VDD(VDD),.Y(g30012),.A(I28241));
  NOT NOT1_3549(.VSS(VSS),.VDD(VDD),.Y(g19415),.A(g15758));
  NOT NOT1_3550(.VSS(VSS),.VDD(VDD),.Y(g24068),.A(g19919));
  NOT NOT1_3551(.VSS(VSS),.VDD(VDD),.Y(g24375),.A(g22722));
  NOT NOT1_3552(.VSS(VSS),.VDD(VDD),.Y(g21059),.A(g15509));
  NOT NOT1_3553(.VSS(VSS),.VDD(VDD),.Y(I33249),.A(g34971));
  NOT NOT1_3554(.VSS(VSS),.VDD(VDD),.Y(g7462),.A(g2599));
  NOT NOT1_3555(.VSS(VSS),.VDD(VDD),.Y(g23059),.A(g20453));
  NOT NOT1_3556(.VSS(VSS),.VDD(VDD),.Y(g31797),.A(g29385));
  NOT NOT1_3557(.VSS(VSS),.VDD(VDD),.Y(g6838),.A(g1724));
  NOT NOT1_3558(.VSS(VSS),.VDD(VDD),.Y(g13096),.A(I15727));
  NOT NOT1_3559(.VSS(VSS),.VDD(VDD),.Y(g33641),.A(I31474));
  NOT NOT1_3560(.VSS(VSS),.VDD(VDD),.Y(g32932),.A(g31327));
  NOT NOT1_3561(.VSS(VSS),.VDD(VDD),.Y(g33797),.A(g33306));
  NOT NOT1_3562(.VSS(VSS),.VDD(VDD),.Y(I31482),.A(g33204));
  NOT NOT1_3563(.VSS(VSS),.VDD(VDD),.Y(g19852),.A(g17015));
  NOT NOT1_3564(.VSS(VSS),.VDD(VDD),.Y(g22721),.A(I22028));
  NOT NOT1_3565(.VSS(VSS),.VDD(VDD),.Y(g10503),.A(g8879));
  NOT NOT1_3566(.VSS(VSS),.VDD(VDD),.Y(I16626),.A(g11986));
  NOT NOT1_3567(.VSS(VSS),.VDD(VDD),.Y(g21058),.A(g15426));
  NOT NOT1_3568(.VSS(VSS),.VDD(VDD),.Y(g6809),.A(g341));
  NOT NOT1_3569(.VSS(VSS),.VDD(VDD),.Y(g32513),.A(g31376));
  NOT NOT1_3570(.VSS(VSS),.VDD(VDD),.Y(I20864),.A(g16960));
  NOT NOT1_3571(.VSS(VSS),.VDD(VDD),.Y(g23058),.A(g20453));
  NOT NOT1_3572(.VSS(VSS),.VDD(VDD),.Y(g32449),.A(I29977));
  NOT NOT1_3573(.VSS(VSS),.VDD(VDD),.Y(g14503),.A(g12256));
  NOT NOT1_3574(.VSS(VSS),.VDD(VDD),.Y(g16691),.A(g14160));
  NOT NOT1_3575(.VSS(VSS),.VDD(VDD),.Y(I24022),.A(g22182));
  NOT NOT1_3576(.VSS(VSS),.VDD(VDD),.Y(g19963),.A(g16326));
  NOT NOT1_3577(.VSS(VSS),.VDD(VDD),.Y(g12842),.A(g10355));
  NOT NOT1_3578(.VSS(VSS),.VDD(VDD),.Y(g34473),.A(g34426));
  NOT NOT1_3579(.VSS(VSS),.VDD(VDD),.Y(I12083),.A(g568));
  NOT NOT1_3580(.VSS(VSS),.VDD(VDD),.Y(g17085),.A(g14238));
  NOT NOT1_3581(.VSS(VSS),.VDD(VDD),.Y(I31779),.A(g33212));
  NOT NOT1_3582(.VSS(VSS),.VDD(VDD),.Y(g24171),.A(I23357));
  NOT NOT1_3583(.VSS(VSS),.VDD(VDD),.Y(g32897),.A(g30735));
  NOT NOT1_3584(.VSS(VSS),.VDD(VDD),.Y(g32961),.A(g31376));
  NOT NOT1_3585(.VSS(VSS),.VDD(VDD),.Y(g23203),.A(g20073));
  NOT NOT1_3586(.VSS(VSS),.VDD(VDD),.Y(g8839),.A(I12819));
  NOT NOT1_3587(.VSS(VSS),.VDD(VDD),.Y(g34789),.A(I32997));
  NOT NOT1_3588(.VSS(VSS),.VDD(VDD),.Y(g7788),.A(g4674));
  NOT NOT1_3589(.VSS(VSS),.VDD(VDD),.Y(g11429),.A(g7616));
  NOT NOT1_3590(.VSS(VSS),.VDD(VDD),.Y(g17721),.A(g12915));
  NOT NOT1_3591(.VSS(VSS),.VDD(VDD),.Y(g29372),.A(I27738));
  NOT NOT1_3592(.VSS(VSS),.VDD(VDD),.Y(g10581),.A(g9529));
  NOT NOT1_3593(.VSS(VSS),.VDD(VDD),.Y(I16775),.A(g12183));
  NOT NOT1_3594(.VSS(VSS),.VDD(VDD),.Y(g13857),.A(I16163));
  NOT NOT1_3595(.VSS(VSS),.VDD(VDD),.Y(g32505),.A(g31566));
  NOT NOT1_3596(.VSS(VSS),.VDD(VDD),.Y(g20994),.A(g15615));
  NOT NOT1_3597(.VSS(VSS),.VDD(VDD),.Y(g9095),.A(g3368));
  NOT NOT1_3598(.VSS(VSS),.VDD(VDD),.Y(g32404),.A(I29936));
  NOT NOT1_3599(.VSS(VSS),.VDD(VDD),.Y(I14800),.A(g10107));
  NOT NOT1_3600(.VSS(VSS),.VDD(VDD),.Y(g33136),.A(g32057));
  NOT NOT1_3601(.VSS(VSS),.VDD(VDD),.Y(g9037),.A(g164));
  NOT NOT1_3602(.VSS(VSS),.VDD(VDD),.Y(g14714),.A(g11405));
  NOT NOT1_3603(.VSS(VSS),.VDD(VDD),.Y(g33635),.A(g33436));
  NOT NOT1_3604(.VSS(VSS),.VDD(VDD),.Y(g24994),.A(g22432));
  NOT NOT1_3605(.VSS(VSS),.VDD(VDD),.Y(g14315),.A(I16479));
  NOT NOT1_3606(.VSS(VSS),.VDD(VDD),.Y(g30325),.A(I28576));
  NOT NOT1_3607(.VSS(VSS),.VDD(VDD),.Y(g34788),.A(I32994));
  NOT NOT1_3608(.VSS(VSS),.VDD(VDD),.Y(g11793),.A(I14633));
  NOT NOT1_3609(.VSS(VSS),.VDD(VDD),.Y(g11428),.A(g7615));
  NOT NOT1_3610(.VSS(VSS),.VDD(VDD),.Y(g26682),.A(g25309));
  NOT NOT1_3611(.VSS(VSS),.VDD(VDD),.Y(g9653),.A(g2441));
  NOT NOT1_3612(.VSS(VSS),.VDD(VDD),.Y(g17431),.A(I18376));
  NOT NOT1_3613(.VSS(VSS),.VDD(VDD),.Y(g13793),.A(I16120));
  NOT NOT1_3614(.VSS(VSS),.VDD(VDD),.Y(g22341),.A(g19801));
  NOT NOT1_3615(.VSS(VSS),.VDD(VDD),.Y(g32717),.A(g30735));
  NOT NOT1_3616(.VSS(VSS),.VDD(VDD),.Y(g34325),.A(g34092));
  NOT NOT1_3617(.VSS(VSS),.VDD(VDD),.Y(I15765),.A(g10823));
  NOT NOT1_3618(.VSS(VSS),.VDD(VDD),.Y(I18009),.A(g13680));
  NOT NOT1_3619(.VSS(VSS),.VDD(VDD),.Y(g21281),.A(g16286));
  NOT NOT1_3620(.VSS(VSS),.VDD(VDD),.Y(g18977),.A(g16100));
  NOT NOT1_3621(.VSS(VSS),.VDD(VDD),.Y(I31786),.A(g33197));
  NOT NOT1_3622(.VSS(VSS),.VDD(VDD),.Y(I32970),.A(g34716));
  NOT NOT1_3623(.VSS(VSS),.VDD(VDD),.Y(g22156),.A(g19147));
  NOT NOT1_3624(.VSS(VSS),.VDD(VDD),.Y(g27830),.A(g26802));
  NOT NOT1_3625(.VSS(VSS),.VDD(VDD),.Y(g21902),.A(I21477));
  NOT NOT1_3626(.VSS(VSS),.VDD(VDD),.Y(g34920),.A(I33152));
  NOT NOT1_3627(.VSS(VSS),.VDD(VDD),.Y(g8172),.A(g3873));
  NOT NOT1_3628(.VSS(VSS),.VDD(VDD),.Y(g8278),.A(g3096));
  NOT NOT1_3629(.VSS(VSS),.VDD(VDD),.Y(g34434),.A(I32473));
  NOT NOT1_3630(.VSS(VSS),.VDD(VDD),.Y(g23902),.A(g21468));
  NOT NOT1_3631(.VSS(VSS),.VDD(VDD),.Y(g23301),.A(g21037));
  NOT NOT1_3632(.VSS(VSS),.VDD(VDD),.Y(g34358),.A(I32364));
  NOT NOT1_3633(.VSS(VSS),.VDD(VDD),.Y(g28917),.A(I27314));
  NOT NOT1_3634(.VSS(VSS),.VDD(VDD),.Y(g23377),.A(g21070));
  NOT NOT1_3635(.VSS(VSS),.VDD(VDD),.Y(I32878),.A(g34501));
  NOT NOT1_3636(.VSS(VSS),.VDD(VDD),.Y(g22180),.A(g19210));
  NOT NOT1_3637(.VSS(VSS),.VDD(VDD),.Y(g24425),.A(g22722));
  NOT NOT1_3638(.VSS(VSS),.VDD(VDD),.Y(g19554),.A(g16861));
  NOT NOT1_3639(.VSS(VSS),.VDD(VDD),.Y(g10111),.A(g1858));
  NOT NOT1_3640(.VSS(VSS),.VDD(VDD),.Y(g12830),.A(g9995));
  NOT NOT1_3641(.VSS(VSS),.VDD(VDD),.Y(g12893),.A(g10391));
  NOT NOT1_3642(.VSS(VSS),.VDD(VDD),.Y(I11816),.A(g93));
  NOT NOT1_3643(.VSS(VSS),.VDD(VDD),.Y(g16583),.A(g14069));
  NOT NOT1_3644(.VSS(VSS),.VDD(VDD),.Y(g7392),.A(g4438));
  NOT NOT1_3645(.VSS(VSS),.VDD(VDD),.Y(g20919),.A(g15224));
  NOT NOT1_3646(.VSS(VSS),.VDD(VDD),.Y(g15756),.A(g13315));
  NOT NOT1_3647(.VSS(VSS),.VDD(VDD),.Y(I25146),.A(g24911));
  NOT NOT1_3648(.VSS(VSS),.VDD(VDD),.Y(g34946),.A(g34934));
  NOT NOT1_3649(.VSS(VSS),.VDD(VDD),.Y(I25562),.A(g25250));
  NOT NOT1_3650(.VSS(VSS),.VDD(VDD),.Y(g19609),.A(g16264));
  NOT NOT1_3651(.VSS(VSS),.VDD(VDD),.Y(g8235),.A(I12463));
  NOT NOT1_3652(.VSS(VSS),.VDD(VDD),.Y(g8343),.A(g3447));
  NOT NOT1_3653(.VSS(VSS),.VDD(VDD),.Y(I18476),.A(g14031));
  NOT NOT1_3654(.VSS(VSS),.VDD(VDD),.Y(g34121),.A(I32056));
  NOT NOT1_3655(.VSS(VSS),.VDD(VDD),.Y(I14964),.A(g10230));
  NOT NOT1_3656(.VSS(VSS),.VDD(VDD),.Y(g19200),.A(I19789));
  NOT NOT1_3657(.VSS(VSS),.VDD(VDD),.Y(g21562),.A(I21199));
  NOT NOT1_3658(.VSS(VSS),.VDD(VDD),.Y(g9752),.A(g1840));
  NOT NOT1_3659(.VSS(VSS),.VDD(VDD),.Y(g12865),.A(g10372));
  NOT NOT1_3660(.VSS(VSS),.VDD(VDD),.Y(g20010),.A(g17226));
  NOT NOT1_3661(.VSS(VSS),.VDD(VDD),.Y(g8282),.A(g3841));
  NOT NOT1_3662(.VSS(VSS),.VDD(VDD),.Y(g20918),.A(g15224));
  NOT NOT1_3663(.VSS(VSS),.VDD(VDD),.Y(g23645),.A(g20875));
  NOT NOT1_3664(.VSS(VSS),.VDD(VDD),.Y(g8566),.A(g3831));
  NOT NOT1_3665(.VSS(VSS),.VDD(VDD),.Y(I18555),.A(g5630));
  NOT NOT1_3666(.VSS(VSS),.VDD(VDD),.Y(g24010),.A(g21562));
  NOT NOT1_3667(.VSS(VSS),.VDD(VDD),.Y(g9917),.A(I13473));
  NOT NOT1_3668(.VSS(VSS),.VDD(VDD),.Y(I32967),.A(g34648));
  NOT NOT1_3669(.VSS(VSS),.VDD(VDD),.Y(I32994),.A(g34739));
  NOT NOT1_3670(.VSS(VSS),.VDD(VDD),.Y(g10741),.A(g8411));
  NOT NOT1_3671(.VSS(VSS),.VDD(VDD),.Y(I21480),.A(g18696));
  NOT NOT1_3672(.VSS(VSS),.VDD(VDD),.Y(g7854),.A(g1152));
  NOT NOT1_3673(.VSS(VSS),.VDD(VDD),.Y(g13504),.A(g11303));
  NOT NOT1_3674(.VSS(VSS),.VDD(VDD),.Y(g25541),.A(g22763));
  NOT NOT1_3675(.VSS(VSS),.VDD(VDD),.Y(g20545),.A(g15373));
  NOT NOT1_3676(.VSS(VSS),.VDD(VDD),.Y(g20079),.A(g17328));
  NOT NOT1_3677(.VSS(VSS),.VDD(VDD),.Y(g20444),.A(g15373));
  NOT NOT1_3678(.VSS(VSS),.VDD(VDD),.Y(g21290),.A(I21029));
  NOT NOT1_3679(.VSS(VSS),.VDD(VDD),.Y(g32723),.A(g31327));
  NOT NOT1_3680(.VSS(VSS),.VDD(VDD),.Y(I31672),.A(g33149));
  NOT NOT1_3681(.VSS(VSS),.VDD(VDD),.Y(g10384),.A(I13802));
  NOT NOT1_3682(.VSS(VSS),.VDD(VDD),.Y(g8134),.A(I12415));
  NOT NOT1_3683(.VSS(VSS),.VDD(VDD),.Y(g23290),.A(g20924));
  NOT NOT1_3684(.VSS(VSS),.VDD(VDD),.Y(I33182),.A(g34910));
  NOT NOT1_3685(.VSS(VSS),.VDD(VDD),.Y(I13374),.A(g6490));
  NOT NOT1_3686(.VSS(VSS),.VDD(VDD),.Y(g8334),.A(g3034));
  NOT NOT1_3687(.VSS(VSS),.VDD(VDD),.Y(g24079),.A(g20998));
  NOT NOT1_3688(.VSS(VSS),.VDD(VDD),.Y(g21698),.A(g18562));
  NOT NOT1_3689(.VSS(VSS),.VDD(VDD),.Y(g14384),.A(I16538));
  NOT NOT1_3690(.VSS(VSS),.VDD(VDD),.Y(g22667),.A(g21156));
  NOT NOT1_3691(.VSS(VSS),.VDD(VDD),.Y(g34682),.A(I32824));
  NOT NOT1_3692(.VSS(VSS),.VDD(VDD),.Y(g29209),.A(I27543));
  NOT NOT1_3693(.VSS(VSS),.VDD(VDD),.Y(g20599),.A(g18065));
  NOT NOT1_3694(.VSS(VSS),.VDD(VDD),.Y(g6926),.A(g3853));
  NOT NOT1_3695(.VSS(VSS),.VDD(VDD),.Y(I16512),.A(g12811));
  NOT NOT1_3696(.VSS(VSS),.VDD(VDD),.Y(g23698),.A(g21611));
  NOT NOT1_3697(.VSS(VSS),.VDD(VDD),.Y(I12415),.A(g48));
  NOT NOT1_3698(.VSS(VSS),.VDD(VDD),.Y(g11317),.A(I14346));
  NOT NOT1_3699(.VSS(VSS),.VDD(VDD),.Y(g20078),.A(g16846));
  NOT NOT1_3700(.VSS(VSS),.VDD(VDD),.Y(I12333),.A(g45));
  NOT NOT1_3701(.VSS(VSS),.VDD(VDD),.Y(g32433),.A(I29961));
  NOT NOT1_3702(.VSS(VSS),.VDD(VDD),.Y(g19745),.A(g16877));
  NOT NOT1_3703(.VSS(VSS),.VDD(VDD),.Y(g24078),.A(g20857));
  NOT NOT1_3704(.VSS(VSS),.VDD(VDD),.Y(g6754),.A(I11617));
  NOT NOT1_3705(.VSS(VSS),.VDD(VDD),.Y(g12705),.A(g7051));
  NOT NOT1_3706(.VSS(VSS),.VDD(VDD),.Y(g20598),.A(g17929));
  NOT NOT1_3707(.VSS(VSS),.VDD(VDD),.Y(g32620),.A(g30673));
  NOT NOT1_3708(.VSS(VSS),.VDD(VDD),.Y(I28579),.A(g29474));
  NOT NOT1_3709(.VSS(VSS),.VDD(VDD),.Y(g20086),.A(I20355));
  NOT NOT1_3710(.VSS(VSS),.VDD(VDD),.Y(g19799),.A(g17062));
  NOT NOT1_3711(.VSS(VSS),.VDD(VDD),.Y(g25325),.A(g22228));
  NOT NOT1_3712(.VSS(VSS),.VDD(VDD),.Y(I32458),.A(g34243));
  NOT NOT1_3713(.VSS(VSS),.VDD(VDD),.Y(g11129),.A(g7994));
  NOT NOT1_3714(.VSS(VSS),.VDD(VDD),.Y(I25366),.A(g24477));
  NOT NOT1_3715(.VSS(VSS),.VDD(VDD),.Y(g8804),.A(g4035));
  NOT NOT1_3716(.VSS(VSS),.VDD(VDD),.Y(g10150),.A(g1700));
  NOT NOT1_3717(.VSS(VSS),.VDD(VDD),.Y(g24086),.A(g20998));
  NOT NOT1_3718(.VSS(VSS),.VDD(VDD),.Y(g16743),.A(g13986));
  NOT NOT1_3719(.VSS(VSS),.VDD(VDD),.Y(g21427),.A(g17367));
  NOT NOT1_3720(.VSS(VSS),.VDD(VDD),.Y(g15731),.A(g13326));
  NOT NOT1_3721(.VSS(VSS),.VDD(VDD),.Y(g9364),.A(g5041));
  NOT NOT1_3722(.VSS(VSS),.VDD(VDD),.Y(g10877),.A(I14079));
  NOT NOT1_3723(.VSS(VSS),.VDD(VDD),.Y(g23427),.A(I22542));
  NOT NOT1_3724(.VSS(VSS),.VDD(VDD),.Y(g25535),.A(g22763));
  NOT NOT1_3725(.VSS(VSS),.VDD(VDD),.Y(g32811),.A(g30735));
  NOT NOT1_3726(.VSS(VSS),.VDD(VDD),.Y(I12963),.A(g640));
  NOT NOT1_3727(.VSS(VSS),.VDD(VDD),.Y(g14150),.A(g12381));
  NOT NOT1_3728(.VSS(VSS),.VDD(VDD),.Y(g21366),.A(I21100));
  NOT NOT1_3729(.VSS(VSS),.VDD(VDD),.Y(g32646),.A(g31070));
  NOT NOT1_3730(.VSS(VSS),.VDD(VDD),.Y(g8792),.A(I12790));
  NOT NOT1_3731(.VSS(VSS),.VDD(VDD),.Y(g7219),.A(g4405));
  NOT NOT1_3732(.VSS(VSS),.VDD(VDD),.Y(g19798),.A(g17200));
  NOT NOT1_3733(.VSS(VSS),.VDD(VDD),.Y(I28014),.A(g28158));
  NOT NOT1_3734(.VSS(VSS),.VDD(VDD),.Y(g11128),.A(g7993));
  NOT NOT1_3735(.VSS(VSS),.VDD(VDD),.Y(g7640),.A(I12128));
  NOT NOT1_3736(.VSS(VSS),.VDD(VDD),.Y(I18238),.A(g13144));
  NOT NOT1_3737(.VSS(VSS),.VDD(VDD),.Y(g10019),.A(g6479));
  NOT NOT1_3738(.VSS(VSS),.VDD(VDD),.Y(g28157),.A(I26670));
  NOT NOT1_3739(.VSS(VSS),.VDD(VDD),.Y(I15626),.A(g12041));
  NOT NOT1_3740(.VSS(VSS),.VDD(VDD),.Y(g22210),.A(I21792));
  NOT NOT1_3741(.VSS(VSS),.VDD(VDD),.Y(g20322),.A(g17873));
  NOT NOT1_3742(.VSS(VSS),.VDD(VDD),.Y(g32971),.A(g31672));
  NOT NOT1_3743(.VSS(VSS),.VDD(VDD),.Y(g7431),.A(g2555));
  NOT NOT1_3744(.VSS(VSS),.VDD(VDD),.Y(I32079),.A(g33937));
  NOT NOT1_3745(.VSS(VSS),.VDD(VDD),.Y(g7252),.A(g1592));
  NOT NOT1_3746(.VSS(VSS),.VDD(VDD),.Y(g16640),.A(I17834));
  NOT NOT1_3747(.VSS(VSS),.VDD(VDD),.Y(g29913),.A(g28840));
  NOT NOT1_3748(.VSS(VSS),.VDD(VDD),.Y(g34760),.A(I32938));
  NOT NOT1_3749(.VSS(VSS),.VDD(VDD),.Y(g7812),.A(I12214));
  NOT NOT1_3750(.VSS(VSS),.VDD(VDD),.Y(g16769),.A(g13530));
  NOT NOT1_3751(.VSS(VSS),.VDD(VDD),.Y(g20159),.A(g17533));
  NOT NOT1_3752(.VSS(VSS),.VDD(VDD),.Y(g34134),.A(I32079));
  NOT NOT1_3753(.VSS(VSS),.VDD(VDD),.Y(g25121),.A(g22432));
  NOT NOT1_3754(.VSS(VSS),.VDD(VDD),.Y(g20901),.A(I20867));
  NOT NOT1_3755(.VSS(VSS),.VDD(VDD),.Y(g13626),.A(g11273));
  NOT NOT1_3756(.VSS(VSS),.VDD(VDD),.Y(g20532),.A(g15277));
  NOT NOT1_3757(.VSS(VSS),.VDD(VDD),.Y(g17487),.A(I18414));
  NOT NOT1_3758(.VSS(VSS),.VDD(VDD),.Y(I27576),.A(g28173));
  NOT NOT1_3759(.VSS(VSS),.VDD(VDD),.Y(I15533),.A(g11867));
  NOT NOT1_3760(.VSS(VSS),.VDD(VDD),.Y(g24159),.A(I23321));
  NOT NOT1_3761(.VSS(VSS),.VDD(VDD),.Y(g13323),.A(g11048));
  NOT NOT1_3762(.VSS(VSS),.VDD(VDD),.Y(g24125),.A(g19890));
  NOT NOT1_3763(.VSS(VSS),.VDD(VDD),.Y(g6983),.A(g4698));
  NOT NOT1_3764(.VSS(VSS),.VDD(VDD),.Y(I18382),.A(g13350));
  NOT NOT1_3765(.VSS(VSS),.VDD(VDD),.Y(g21661),.A(I21222));
  NOT NOT1_3766(.VSS(VSS),.VDD(VDD),.Y(g17502),.A(g14697));
  NOT NOT1_3767(.VSS(VSS),.VDD(VDD),.Y(g16768),.A(g13223));
  NOT NOT1_3768(.VSS(VSS),.VDD(VDD),.Y(I19927),.A(g17408));
  NOT NOT1_3769(.VSS(VSS),.VDD(VDD),.Y(g20158),.A(g16971));
  NOT NOT1_3770(.VSS(VSS),.VDD(VDD),.Y(g8113),.A(g3466));
  NOT NOT1_3771(.VSS(VSS),.VDD(VDD),.Y(g12938),.A(I15556));
  NOT NOT1_3772(.VSS(VSS),.VDD(VDD),.Y(I16498),.A(g10430));
  NOT NOT1_3773(.VSS(VSS),.VDD(VDD),.Y(g23403),.A(I22512));
  NOT NOT1_3774(.VSS(VSS),.VDD(VDD),.Y(g23547),.A(g21611));
  NOT NOT1_3775(.VSS(VSS),.VDD(VDD),.Y(g23895),.A(g19147));
  NOT NOT1_3776(.VSS(VSS),.VDD(VDD),.Y(I13424),.A(g5689));
  NOT NOT1_3777(.VSS(VSS),.VDD(VDD),.Y(g24158),.A(I23318));
  NOT NOT1_3778(.VSS(VSS),.VDD(VDD),.Y(g33750),.A(I31607));
  NOT NOT1_3779(.VSS(VSS),.VDD(VDD),.Y(I18092),.A(g3668));
  NOT NOT1_3780(.VSS(VSS),.VDD(VDD),.Y(g7405),.A(g1936));
  NOT NOT1_3781(.VSS(VSS),.VDD(VDD),.Y(g13298),.A(I15862));
  NOT NOT1_3782(.VSS(VSS),.VDD(VDD),.Y(g19732),.A(g17096));
  NOT NOT1_3783(.VSS(VSS),.VDD(VDD),.Y(I22264),.A(g20100));
  NOT NOT1_3784(.VSS(VSS),.VDD(VDD),.Y(I30980),.A(g32132));
  NOT NOT1_3785(.VSS(VSS),.VDD(VDD),.Y(I24008),.A(g22182));
  NOT NOT1_3786(.VSS(VSS),.VDD(VDD),.Y(g29905),.A(g28783));
  NOT NOT1_3787(.VSS(VSS),.VDD(VDD),.Y(g20561),.A(g17873));
  NOT NOT1_3788(.VSS(VSS),.VDD(VDD),.Y(g20656),.A(g17249));
  NOT NOT1_3789(.VSS(VSS),.VDD(VDD),.Y(g9553),.A(I13202));
  NOT NOT1_3790(.VSS(VSS),.VDD(VDD),.Y(I18518),.A(g13835));
  NOT NOT1_3791(.VSS(VSS),.VDD(VDD),.Y(I18154),.A(g13177));
  NOT NOT1_3792(.VSS(VSS),.VDD(VDD),.Y(g23226),.A(g20924));
  NOT NOT1_3793(.VSS(VSS),.VDD(VDD),.Y(g7765),.A(g4165));
  NOT NOT1_3794(.VSS(VSS),.VDD(VDD),.Y(g20680),.A(g15348));
  NOT NOT1_3795(.VSS(VSS),.VDD(VDD),.Y(g26648),.A(g25115));
  NOT NOT1_3796(.VSS(VSS),.VDD(VDD),.Y(g20144),.A(g17533));
  NOT NOT1_3797(.VSS(VSS),.VDD(VDD),.Y(g10402),.A(g7023));
  NOT NOT1_3798(.VSS(VSS),.VDD(VDD),.Y(g23715),.A(g20764));
  NOT NOT1_3799(.VSS(VSS),.VDD(VDD),.Y(g23481),.A(I22604));
  NOT NOT1_3800(.VSS(VSS),.VDD(VDD),.Y(g32850),.A(g30937));
  NOT NOT1_3801(.VSS(VSS),.VDD(VDD),.Y(g31796),.A(g29385));
  NOT NOT1_3802(.VSS(VSS),.VDD(VDD),.Y(g19761),.A(g17015));
  NOT NOT1_3803(.VSS(VSS),.VDD(VDD),.Y(I12608),.A(g1582));
  NOT NOT1_3804(.VSS(VSS),.VDD(VDD),.Y(g12875),.A(I15494));
  NOT NOT1_3805(.VSS(VSS),.VDD(VDD),.Y(I21734),.A(g19268));
  NOT NOT1_3806(.VSS(VSS),.VDD(VDD),.Y(g6961),.A(I11734));
  NOT NOT1_3807(.VSS(VSS),.VDD(VDD),.Y(g8567),.A(g4082));
  NOT NOT1_3808(.VSS(VSS),.VDD(VDD),.Y(I21930),.A(g21297));
  NOT NOT1_3809(.VSS(VSS),.VDD(VDD),.Y(g34927),.A(I33173));
  NOT NOT1_3810(.VSS(VSS),.VDD(VDD),.Y(g7733),.A(g4093));
  NOT NOT1_3811(.VSS(VSS),.VDD(VDD),.Y(I22422),.A(g19330));
  NOT NOT1_3812(.VSS(VSS),.VDD(VDD),.Y(I15697),.A(g6000));
  NOT NOT1_3813(.VSS(VSS),.VDD(VDD),.Y(I17873),.A(g15017));
  NOT NOT1_3814(.VSS(VSS),.VDD(VDD),.Y(g31840),.A(g29385));
  NOT NOT1_3815(.VSS(VSS),.VDD(VDD),.Y(I32158),.A(g33791));
  NOT NOT1_3816(.VSS(VSS),.VDD(VDD),.Y(g12218),.A(I15073));
  NOT NOT1_3817(.VSS(VSS),.VDD(VDD),.Y(g32896),.A(g31376));
  NOT NOT1_3818(.VSS(VSS),.VDD(VDD),.Y(g12837),.A(g10354));
  NOT NOT1_3819(.VSS(VSS),.VDD(VDD),.Y(g23127),.A(g21163));
  NOT NOT1_3820(.VSS(VSS),.VDD(VDD),.Y(g6927),.A(g3845));
  NOT NOT1_3821(.VSS(VSS),.VDD(VDD),.Y(I21838),.A(g19263));
  NOT NOT1_3822(.VSS(VSS),.VDD(VDD),.Y(g25134),.A(g22417));
  NOT NOT1_3823(.VSS(VSS),.VDD(VDD),.Y(g10001),.A(g6105));
  NOT NOT1_3824(.VSS(VSS),.VDD(VDD),.Y(g22975),.A(g20391));
  NOT NOT1_3825(.VSS(VSS),.VDD(VDD),.Y(g13856),.A(I16160));
  NOT NOT1_3826(.VSS(VSS),.VDD(VDD),.Y(I23694),.A(g23252));
  NOT NOT1_3827(.VSS(VSS),.VDD(VDD),.Y(I29248),.A(g29491));
  NOT NOT1_3828(.VSS(VSS),.VDD(VDD),.Y(g9888),.A(g5831));
  NOT NOT1_3829(.VSS(VSS),.VDD(VDD),.Y(g10077),.A(g1724));
  NOT NOT1_3830(.VSS(VSS),.VDD(VDD),.Y(g13995),.A(g11261));
  NOT NOT1_3831(.VSS(VSS),.VDD(VDD),.Y(I33149),.A(g34900));
  NOT NOT1_3832(.VSS(VSS),.VDD(VDD),.Y(g8593),.A(g3759));
  NOT NOT1_3833(.VSS(VSS),.VDD(VDD),.Y(g29153),.A(g27937));
  NOT NOT1_3834(.VSS(VSS),.VDD(VDD),.Y(g24966),.A(g22763));
  NOT NOT1_3835(.VSS(VSS),.VDD(VDD),.Y(g7073),.A(g6191));
  NOT NOT1_3836(.VSS(VSS),.VDD(VDD),.Y(I12799),.A(g59));
  NOT NOT1_3837(.VSS(VSS),.VDD(VDD),.Y(g20631),.A(g15171));
  NOT NOT1_3838(.VSS(VSS),.VDD(VDD),.Y(g17815),.A(g14348));
  NOT NOT1_3839(.VSS(VSS),.VDD(VDD),.Y(g10597),.A(g10233));
  NOT NOT1_3840(.VSS(VSS),.VDD(VDD),.Y(g23490),.A(g21514));
  NOT NOT1_3841(.VSS(VSS),.VDD(VDD),.Y(g25506),.A(g22228));
  NOT NOT1_3842(.VSS(VSS),.VDD(VDD),.Y(g9429),.A(g3723));
  NOT NOT1_3843(.VSS(VSS),.VDD(VDD),.Y(I13705),.A(g63));
  NOT NOT1_3844(.VSS(VSS),.VDD(VDD),.Y(I29204),.A(g29505));
  NOT NOT1_3845(.VSS(VSS),.VDD(VDD),.Y(g32716),.A(g31376));
  NOT NOT1_3846(.VSS(VSS),.VDD(VDD),.Y(g7473),.A(g6697));
  NOT NOT1_3847(.VSS(VSS),.VDD(VDD),.Y(g16249),.A(I17590));
  NOT NOT1_3848(.VSS(VSS),.VDD(VDD),.Y(g18976),.A(g16100));
  NOT NOT1_3849(.VSS(VSS),.VDD(VDD),.Y(g14597),.A(I16713));
  NOT NOT1_3850(.VSS(VSS),.VDD(VDD),.Y(g19539),.A(g16129));
  NOT NOT1_3851(.VSS(VSS),.VDD(VDD),.Y(g6946),.A(I11721));
  NOT NOT1_3852(.VSS(VSS),.VDD(VDD),.Y(g24017),.A(g18833));
  NOT NOT1_3853(.VSS(VSS),.VDD(VDD),.Y(g11512),.A(g7634));
  NOT NOT1_3854(.VSS(VSS),.VDD(VDD),.Y(g34648),.A(I32752));
  NOT NOT1_3855(.VSS(VSS),.VDD(VDD),.Y(g24364),.A(g22722));
  NOT NOT1_3856(.VSS(VSS),.VDD(VDD),.Y(g17677),.A(g14882));
  NOT NOT1_3857(.VSS(VSS),.VDD(VDD),.Y(g34491),.A(I32550));
  NOT NOT1_3858(.VSS(VSS),.VDD(VDD),.Y(I22542),.A(g19773));
  NOT NOT1_3859(.VSS(VSS),.VDD(VDD),.Y(g16482),.A(g13464));
  NOT NOT1_3860(.VSS(VSS),.VDD(VDD),.Y(I17834),.A(g14977));
  NOT NOT1_3861(.VSS(VSS),.VDD(VDD),.Y(g31522),.A(I29185));
  NOT NOT1_3862(.VSS(VSS),.VDD(VDD),.Y(g32582),.A(g31170));
  NOT NOT1_3863(.VSS(VSS),.VDD(VDD),.Y(g7980),.A(g3161));
  NOT NOT1_3864(.VSS(VSS),.VDD(VDD),.Y(g21297),.A(I21042));
  NOT NOT1_3865(.VSS(VSS),.VDD(VDD),.Y(g18954),.A(g17427));
  NOT NOT1_3866(.VSS(VSS),.VDD(VDD),.Y(g23376),.A(g21070));
  NOT NOT1_3867(.VSS(VSS),.VDD(VDD),.Y(g23385),.A(I22488));
  NOT NOT1_3868(.VSS(VSS),.VDD(VDD),.Y(I25095),.A(g25265));
  NOT NOT1_3869(.VSS(VSS),.VDD(VDD),.Y(g19538),.A(g16100));
  NOT NOT1_3870(.VSS(VSS),.VDD(VDD),.Y(g6903),.A(g3502));
  NOT NOT1_3871(.VSS(VSS),.VDD(VDD),.Y(g7069),.A(g6137));
  NOT NOT1_3872(.VSS(VSS),.VDD(VDD),.Y(g9281),.A(I13057));
  NOT NOT1_3873(.VSS(VSS),.VDD(VDD),.Y(I12805),.A(g4098));
  NOT NOT1_3874(.VSS(VSS),.VDD(VDD),.Y(g26990),.A(g26105));
  NOT NOT1_3875(.VSS(VSS),.VDD(VDD),.Y(g34755),.A(I32929));
  NOT NOT1_3876(.VSS(VSS),.VDD(VDD),.Y(g23889),.A(g20682));
  NOT NOT1_3877(.VSS(VSS),.VDD(VDD),.Y(I13124),.A(g2729));
  NOT NOT1_3878(.VSS(VSS),.VDD(VDD),.Y(I18728),.A(g6012));
  NOT NOT1_3879(.VSS(VSS),.VDD(VDD),.Y(I21210),.A(g17526));
  NOT NOT1_3880(.VSS(VSS),.VDD(VDD),.Y(g23354),.A(g20453));
  NOT NOT1_3881(.VSS(VSS),.VDD(VDD),.Y(I14579),.A(g8792));
  NOT NOT1_3882(.VSS(VSS),.VDD(VDD),.Y(g22169),.A(g19147));
  NOT NOT1_3883(.VSS(VSS),.VDD(VDD),.Y(I26700),.A(g27956));
  NOT NOT1_3884(.VSS(VSS),.VDD(VDD),.Y(g34770),.A(I32956));
  NOT NOT1_3885(.VSS(VSS),.VDD(VDD),.Y(g12470),.A(I15284));
  NOT NOT1_3886(.VSS(VSS),.VDD(VDD),.Y(g7540),.A(I12026));
  NOT NOT1_3887(.VSS(VSS),.VDD(VDD),.Y(g8160),.A(g3423));
  NOT NOT1_3888(.VSS(VSS),.VDD(VDD),.Y(g22884),.A(g20453));
  NOT NOT1_3889(.VSS(VSS),.VDD(VDD),.Y(g34981),.A(g34973));
  NOT NOT1_3890(.VSS(VSS),.VDD(VDD),.Y(g23888),.A(g18997));
  NOT NOT1_3891(.VSS(VSS),.VDD(VDD),.Y(g23824),.A(g21271));
  NOT NOT1_3892(.VSS(VSS),.VDD(VDD),.Y(I15831),.A(g10416));
  NOT NOT1_3893(.VSS(VSS),.VDD(VDD),.Y(g32627),.A(g30673));
  NOT NOT1_3894(.VSS(VSS),.VDD(VDD),.Y(g28307),.A(g27306));
  NOT NOT1_3895(.VSS(VSS),.VDD(VDD),.Y(g32959),.A(g30937));
  NOT NOT1_3896(.VSS(VSS),.VDD(VDD),.Y(g32925),.A(g31327));
  NOT NOT1_3897(.VSS(VSS),.VDD(VDD),.Y(g21181),.A(g15426));
  NOT NOT1_3898(.VSS(VSS),.VDD(VDD),.Y(g22168),.A(g19147));
  NOT NOT1_3899(.VSS(VSS),.VDD(VDD),.Y(g10102),.A(g6727));
  NOT NOT1_3900(.VSS(VSS),.VDD(VDD),.Y(g10157),.A(g2036));
  NOT NOT1_3901(.VSS(VSS),.VDD(VDD),.Y(g31862),.A(I29444));
  NOT NOT1_3902(.VSS(VSS),.VDD(VDD),.Y(g32958),.A(g31710));
  NOT NOT1_3903(.VSS(VSS),.VDD(VDD),.Y(I15316),.A(g10087));
  NOT NOT1_3904(.VSS(VSS),.VDD(VDD),.Y(I19719),.A(g17431));
  NOT NOT1_3905(.VSS(VSS),.VDD(VDD),.Y(g8450),.A(g3821));
  NOT NOT1_3906(.VSS(VSS),.VDD(VDD),.Y(g24023),.A(g21127));
  NOT NOT1_3907(.VSS(VSS),.VDD(VDD),.Y(g26718),.A(g25168));
  NOT NOT1_3908(.VSS(VSS),.VDD(VDD),.Y(I32364),.A(g34208));
  NOT NOT1_3909(.VSS(VSS),.VDD(VDD),.Y(g17791),.A(g14950));
  NOT NOT1_3910(.VSS(VSS),.VDD(VDD),.Y(g20571),.A(g15277));
  NOT NOT1_3911(.VSS(VSS),.VDD(VDD),.Y(g9684),.A(g6191));
  NOT NOT1_3912(.VSS(VSS),.VDD(VDD),.Y(g11316),.A(g8967));
  NOT NOT1_3913(.VSS(VSS),.VDD(VDD),.Y(g9745),.A(g6537));
  NOT NOT1_3914(.VSS(VSS),.VDD(VDD),.Y(g12075),.A(I14935));
  NOT NOT1_3915(.VSS(VSS),.VDD(VDD),.Y(I17436),.A(g13416));
  NOT NOT1_3916(.VSS(VSS),.VDD(VDD),.Y(g28431),.A(I26925));
  NOT NOT1_3917(.VSS(VSS),.VDD(VDD),.Y(g9639),.A(g1752));
  NOT NOT1_3918(.VSS(VSS),.VDD(VDD),.Y(I18906),.A(g16963));
  NOT NOT1_3919(.VSS(VSS),.VDD(VDD),.Y(g9338),.A(g1870));
  NOT NOT1_3920(.VSS(VSS),.VDD(VDD),.Y(g24571),.A(g22942));
  NOT NOT1_3921(.VSS(VSS),.VDD(VDD),.Y(g10231),.A(g2661));
  NOT NOT1_3922(.VSS(VSS),.VDD(VDD),.Y(I18083),.A(g13394));
  NOT NOT1_3923(.VSS(VSS),.VDD(VDD),.Y(g9963),.A(g7));
  NOT NOT1_3924(.VSS(VSS),.VDD(VDD),.Y(I26296),.A(g26820));
  NOT NOT1_3925(.VSS(VSS),.VDD(VDD),.Y(g33326),.A(g32318));
  NOT NOT1_3926(.VSS(VSS),.VDD(VDD),.Y(g17410),.A(g12955));
  NOT NOT1_3927(.VSS(VSS),.VDD(VDD),.Y(I12761),.A(g4188));
  NOT NOT1_3928(.VSS(VSS),.VDD(VDD),.Y(g11498),.A(I14475));
  NOT NOT1_3929(.VSS(VSS),.VDD(VDD),.Y(g34767),.A(I32947));
  NOT NOT1_3930(.VSS(VSS),.VDD(VDD),.Y(g14231),.A(g12246));
  NOT NOT1_3931(.VSS(VSS),.VDD(VDD),.Y(g26832),.A(g24850));
  NOT NOT1_3932(.VSS(VSS),.VDD(VDD),.Y(g34845),.A(g34773));
  NOT NOT1_3933(.VSS(VSS),.VDD(VDD),.Y(g32603),.A(g31070));
  NOT NOT1_3934(.VSS(VSS),.VDD(VDD),.Y(g6831),.A(g1413));
  NOT NOT1_3935(.VSS(VSS),.VDD(VDD),.Y(I22464),.A(g21222));
  NOT NOT1_3936(.VSS(VSS),.VDD(VDD),.Y(g23931),.A(g20875));
  NOT NOT1_3937(.VSS(VSS),.VDD(VDD),.Y(g32742),.A(g31021));
  NOT NOT1_3938(.VSS(VSS),.VDD(VDD),.Y(I29233),.A(g30295));
  NOT NOT1_3939(.VSS(VSS),.VDD(VDD),.Y(g9309),.A(g5462));
  NOT NOT1_3940(.VSS(VSS),.VDD(VDD),.Y(I23306),.A(g21673));
  NOT NOT1_3941(.VSS(VSS),.VDD(VDD),.Y(g30990),.A(g29676));
  NOT NOT1_3942(.VSS(VSS),.VDD(VDD),.Y(I18304),.A(g14790));
  NOT NOT1_3943(.VSS(VSS),.VDD(VDD),.Y(g19771),.A(g17096));
  NOT NOT1_3944(.VSS(VSS),.VDD(VDD),.Y(g25240),.A(g23650));
  NOT NOT1_3945(.VSS(VSS),.VDD(VDD),.Y(g32944),.A(g31021));
  NOT NOT1_3946(.VSS(VSS),.VDD(VDD),.Y(I29182),.A(g30012));
  NOT NOT1_3947(.VSS(VSS),.VDD(VDD),.Y(g29474),.A(I27758));
  NOT NOT1_3948(.VSS(VSS),.VDD(VDD),.Y(g34990),.A(I33270));
  NOT NOT1_3949(.VSS(VSS),.VDD(VDD),.Y(g11989),.A(I14839));
  NOT NOT1_3950(.VSS(VSS),.VDD(VDD),.Y(I25190),.A(g25423));
  NOT NOT1_3951(.VSS(VSS),.VDD(VDD),.Y(g16826),.A(I18034));
  NOT NOT1_3952(.VSS(VSS),.VDD(VDD),.Y(g17479),.A(g14855));
  NOT NOT1_3953(.VSS(VSS),.VDD(VDD),.Y(g21426),.A(g15277));
  NOT NOT1_3954(.VSS(VSS),.VDD(VDD),.Y(g8179),.A(g4999));
  NOT NOT1_3955(.VSS(VSS),.VDD(VDD),.Y(g12037),.A(I14893));
  NOT NOT1_3956(.VSS(VSS),.VDD(VDD),.Y(g20495),.A(g17926));
  NOT NOT1_3957(.VSS(VSS),.VDD(VDD),.Y(g23426),.A(I22539));
  NOT NOT1_3958(.VSS(VSS),.VDD(VDD),.Y(g25903),.A(I25005));
  NOT NOT1_3959(.VSS(VSS),.VDD(VDD),.Y(g27984),.A(g26737));
  NOT NOT1_3960(.VSS(VSS),.VDD(VDD),.Y(I13875),.A(g1233));
  NOT NOT1_3961(.VSS(VSS),.VDD(VDD),.Y(g33702),.A(I31545));
  NOT NOT1_3962(.VSS(VSS),.VDD(VDD),.Y(g9808),.A(g5827));
  NOT NOT1_3963(.VSS(VSS),.VDD(VDD),.Y(g19683),.A(g16931));
  NOT NOT1_3964(.VSS(VSS),.VDD(VDD),.Y(g23190),.A(I22286));
  NOT NOT1_3965(.VSS(VSS),.VDD(VDD),.Y(I16709),.A(g10430));
  NOT NOT1_3966(.VSS(VSS),.VDD(VDD),.Y(g11988),.A(I14836));
  NOT NOT1_3967(.VSS(VSS),.VDD(VDD),.Y(I21815),.A(g21308));
  NOT NOT1_3968(.VSS(VSS),.VDD(VDD),.Y(g17478),.A(g14996));
  NOT NOT1_3969(.VSS(VSS),.VDD(VDD),.Y(g28156),.A(I26667));
  NOT NOT1_3970(.VSS(VSS),.VDD(VDD),.Y(I12013),.A(g590));
  NOT NOT1_3971(.VSS(VSS),.VDD(VDD),.Y(g17015),.A(I18143));
  NOT NOT1_3972(.VSS(VSS),.VDD(VDD),.Y(g32681),.A(g30735));
  NOT NOT1_3973(.VSS(VSS),.VDD(VDD),.Y(I32309),.A(g34210));
  NOT NOT1_3974(.VSS(VSS),.VDD(VDD),.Y(I12214),.A(g6561));
  NOT NOT1_3975(.VSS(VSS),.VDD(VDD),.Y(g16182),.A(g13846));
  NOT NOT1_3976(.VSS(VSS),.VDD(VDD),.Y(g16651),.A(g14005));
  NOT NOT1_3977(.VSS(VSS),.VDD(VDD),.Y(I22153),.A(g20014));
  NOT NOT1_3978(.VSS(VSS),.VDD(VDD),.Y(g23520),.A(g21468));
  NOT NOT1_3979(.VSS(VSS),.VDD(VDD),.Y(g27155),.A(g26131));
  NOT NOT1_3980(.VSS(VSS),.VDD(VDD),.Y(g9759),.A(g2265));
  NOT NOT1_3981(.VSS(VSS),.VDD(VDD),.Y(g18830),.A(g18008));
  NOT NOT1_3982(.VSS(VSS),.VDD(VDD),.Y(I16471),.A(g12367));
  NOT NOT1_3983(.VSS(VSS),.VDD(VDD),.Y(g17486),.A(I18411));
  NOT NOT1_3984(.VSS(VSS),.VDD(VDD),.Y(g7898),.A(g4991));
  NOT NOT1_3985(.VSS(VSS),.VDD(VDD),.Y(g25563),.A(g22594));
  NOT NOT1_3986(.VSS(VSS),.VDD(VDD),.Y(g32802),.A(g31327));
  NOT NOT1_3987(.VSS(VSS),.VDD(VDD),.Y(g32857),.A(g30937));
  NOT NOT1_3988(.VSS(VSS),.VDD(VDD),.Y(g22223),.A(g19210));
  NOT NOT1_3989(.VSS(VSS),.VDD(VDD),.Y(g13271),.A(I15834));
  NOT NOT1_3990(.VSS(VSS),.VDD(VDD),.Y(g34718),.A(I32884));
  NOT NOT1_3991(.VSS(VSS),.VDD(VDD),.Y(g24985),.A(g23586));
  NOT NOT1_3992(.VSS(VSS),.VDD(VDD),.Y(g34521),.A(g34270));
  NOT NOT1_3993(.VSS(VSS),.VDD(VDD),.Y(g32730),.A(g31327));
  NOT NOT1_3994(.VSS(VSS),.VDD(VDD),.Y(g23546),.A(g21611));
  NOT NOT1_3995(.VSS(VSS),.VDD(VDD),.Y(I24215),.A(g22360));
  NOT NOT1_3996(.VSS(VSS),.VDD(VDD),.Y(g32793),.A(g31021));
  NOT NOT1_3997(.VSS(VSS),.VDD(VDD),.Y(I18653),.A(g5681));
  NOT NOT1_3998(.VSS(VSS),.VDD(VDD),.Y(g20374),.A(g18065));
  NOT NOT1_3999(.VSS(VSS),.VDD(VDD),.Y(g23211),.A(g21308));
  NOT NOT1_4000(.VSS(VSS),.VDD(VDD),.Y(I30644),.A(g32024));
  NOT NOT1_4001(.VSS(VSS),.VDD(VDD),.Y(g19882),.A(g16540));
  NOT NOT1_4002(.VSS(VSS),.VDD(VDD),.Y(g19414),.A(g16349));
  NOT NOT1_4003(.VSS(VSS),.VDD(VDD),.Y(g26701),.A(g25341));
  NOT NOT1_4004(.VSS(VSS),.VDD(VDD),.Y(g7245),.A(I11896));
  NOT NOT1_4005(.VSS(VSS),.VDD(VDD),.Y(g17580),.A(I18509));
  NOT NOT1_4006(.VSS(VSS),.VDD(VDD),.Y(g11753),.A(g8587));
  NOT NOT1_4007(.VSS(VSS),.VDD(VDD),.Y(I29961),.A(g30984));
  NOT NOT1_4008(.VSS(VSS),.VDD(VDD),.Y(I12538),.A(g58));
  NOT NOT1_4009(.VSS(VSS),.VDD(VDD),.Y(g26777),.A(g25439));
  NOT NOT1_4010(.VSS(VSS),.VDD(VDD),.Y(g20643),.A(g15962));
  NOT NOT1_4011(.VSS(VSS),.VDD(VDD),.Y(I18138),.A(g14277));
  NOT NOT1_4012(.VSS(VSS),.VDD(VDD),.Y(g9049),.A(g640));
  NOT NOT1_4013(.VSS(VSS),.VDD(VDD),.Y(g23088),.A(I22240));
  NOT NOT1_4014(.VSS(VSS),.VDD(VDD),.Y(g31847),.A(g29385));
  NOT NOT1_4015(.VSS(VSS),.VDD(VDD),.Y(g32765),.A(g31327));
  NOT NOT1_4016(.VSS(VSS),.VDD(VDD),.Y(g19407),.A(g16268));
  NOT NOT1_4017(.VSS(VSS),.VDD(VDD),.Y(g9449),.A(g5770));
  NOT NOT1_4018(.VSS(VSS),.VDD(VDD),.Y(g16449),.A(I17679));
  NOT NOT1_4019(.VSS(VSS),.VDD(VDD),.Y(g11031),.A(g8609));
  NOT NOT1_4020(.VSS(VSS),.VDD(VDD),.Y(g22922),.A(g20330));
  NOT NOT1_4021(.VSS(VSS),.VDD(VDD),.Y(g23860),.A(g19074));
  NOT NOT1_4022(.VSS(VSS),.VDD(VDD),.Y(I15650),.A(g12110));
  NOT NOT1_4023(.VSS(VSS),.VDD(VDD),.Y(g32690),.A(g31070));
  NOT NOT1_4024(.VSS(VSS),.VDD(VDD),.Y(g9575),.A(g6509));
  NOT NOT1_4025(.VSS(VSS),.VDD(VDD),.Y(g32549),.A(g31554));
  NOT NOT1_4026(.VSS(VSS),.VDD(VDD),.Y(I15736),.A(g12322));
  NOT NOT1_4027(.VSS(VSS),.VDD(VDD),.Y(I14684),.A(g7717));
  NOT NOT1_4028(.VSS(VSS),.VDD(VDD),.Y(I18333),.A(g1083));
  NOT NOT1_4029(.VSS(VSS),.VDD(VDD),.Y(g22179),.A(g19210));
  NOT NOT1_4030(.VSS(VSS),.VDD(VDD),.Y(I29717),.A(g30931));
  NOT NOT1_4031(.VSS(VSS),.VDD(VDD),.Y(g25262),.A(g22763));
  NOT NOT1_4032(.VSS(VSS),.VDD(VDD),.Y(I11617),.A(g1));
  NOT NOT1_4033(.VSS(VSS),.VDD(VDD),.Y(g11736),.A(g8165));
  NOT NOT1_4034(.VSS(VSS),.VDD(VDD),.Y(g20669),.A(g15426));
  NOT NOT1_4035(.VSS(VSS),.VDD(VDD),.Y(I17136),.A(g14398));
  NOT NOT1_4036(.VSS(VSS),.VDD(VDD),.Y(g16897),.A(I18083));
  NOT NOT1_4037(.VSS(VSS),.VDD(VDD),.Y(I26503),.A(g26811));
  NOT NOT1_4038(.VSS(VSS),.VDD(VDD),.Y(g34573),.A(I32645));
  NOT NOT1_4039(.VSS(VSS),.VDD(VDD),.Y(g7344),.A(g5659));
  NOT NOT1_4040(.VSS(VSS),.VDD(VDD),.Y(g25899),.A(g24997));
  NOT NOT1_4041(.VSS(VSS),.VDD(VDD),.Y(g13736),.A(g11313));
  NOT NOT1_4042(.VSS(VSS),.VDD(VDD),.Y(g32548),.A(g30673));
  NOT NOT1_4043(.VSS(VSS),.VDD(VDD),.Y(I18852),.A(g13716));
  NOT NOT1_4044(.VSS(VSS),.VDD(VDD),.Y(I32687),.A(g34431));
  NOT NOT1_4045(.VSS(VSS),.VDD(VDD),.Y(g34247),.A(I32240));
  NOT NOT1_4046(.VSS(VSS),.VDD(VDD),.Y(I32976),.A(g34699));
  NOT NOT1_4047(.VSS(VSS),.VDD(VDD),.Y(I32985),.A(g34736));
  NOT NOT1_4048(.VSS(VSS),.VDD(VDD),.Y(g22178),.A(g19147));
  NOT NOT1_4049(.VSS(VSS),.VDD(VDD),.Y(g9498),.A(g5101));
  NOT NOT1_4050(.VSS(VSS),.VDD(VDD),.Y(g6873),.A(g3151));
  NOT NOT1_4051(.VSS(VSS),.VDD(VDD),.Y(g20668),.A(g15426));
  NOT NOT1_4052(.VSS(VSS),.VDD(VDD),.Y(g34926),.A(I33170));
  NOT NOT1_4053(.VSS(VSS),.VDD(VDD),.Y(g32504),.A(g30673));
  NOT NOT1_4054(.VSS(VSS),.VDD(VDD),.Y(g31851),.A(g29385));
  NOT NOT1_4055(.VSS(VSS),.VDD(VDD),.Y(I15843),.A(g11181));
  NOT NOT1_4056(.VSS(VSS),.VDD(VDD),.Y(I32752),.A(g34510));
  NOT NOT1_4057(.VSS(VSS),.VDD(VDD),.Y(g9833),.A(g2449));
  NOT NOT1_4058(.VSS(VSS),.VDD(VDD),.Y(g10287),.A(I13715));
  NOT NOT1_4059(.VSS(VSS),.VDD(VDD),.Y(g7259),.A(g4375));
  NOT NOT1_4060(.VSS(VSS),.VDD(VDD),.Y(g21659),.A(g17727));
  NOT NOT1_4061(.VSS(VSS),.VDD(VDD),.Y(I33050),.A(g34777));
  NOT NOT1_4062(.VSS(VSS),.VDD(VDD),.Y(g14314),.A(I16476));
  NOT NOT1_4063(.VSS(VSS),.VDD(VDD),.Y(g16717),.A(g13951));
  NOT NOT1_4064(.VSS(VSS),.VDD(VDD),.Y(g17531),.A(I18476));
  NOT NOT1_4065(.VSS(VSS),.VDD(VDD),.Y(g12836),.A(g10351));
  NOT NOT1_4066(.VSS(VSS),.VDD(VDD),.Y(g20195),.A(g16931));
  NOT NOT1_4067(.VSS(VSS),.VDD(VDD),.Y(I26581),.A(g26942));
  NOT NOT1_4068(.VSS(VSS),.VDD(VDD),.Y(g8997),.A(g577));
  NOT NOT1_4069(.VSS(VSS),.VDD(VDD),.Y(g23987),.A(g19277));
  NOT NOT1_4070(.VSS(VSS),.VDD(VDD),.Y(g10085),.A(g1768));
  NOT NOT1_4071(.VSS(VSS),.VDD(VDD),.Y(g8541),.A(g3498));
  NOT NOT1_4072(.VSS(VSS),.VDD(VDD),.Y(g23250),.A(g21070));
  NOT NOT1_4073(.VSS(VSS),.VDD(VDD),.Y(g24489),.A(I23694));
  NOT NOT1_4074(.VSS(VSS),.VDD(VDD),.Y(I23363),.A(g23385));
  NOT NOT1_4075(.VSS(VSS),.VDD(VDD),.Y(g14307),.A(I16468));
  NOT NOT1_4076(.VSS(VSS),.VDD(VDD),.Y(I27235),.A(g27320));
  NOT NOT1_4077(.VSS(VSS),.VDD(VDD),.Y(g17178),.A(I18214));
  NOT NOT1_4078(.VSS(VSS),.VDD(VDD),.Y(g6869),.A(I11691));
  NOT NOT1_4079(.VSS(VSS),.VDD(VDD),.Y(g34777),.A(I32973));
  NOT NOT1_4080(.VSS(VSS),.VDD(VDD),.Y(g12477),.A(I15295));
  NOT NOT1_4081(.VSS(VSS),.VDD(VDD),.Y(g20525),.A(g17955));
  NOT NOT1_4082(.VSS(VSS),.VDD(VDD),.Y(I15869),.A(g11234));
  NOT NOT1_4083(.VSS(VSS),.VDD(VDD),.Y(g18939),.A(g16077));
  NOT NOT1_4084(.VSS(VSS),.VDD(VDD),.Y(g8132),.A(I12411));
  NOT NOT1_4085(.VSS(VSS),.VDD(VDD),.Y(g28443),.A(I26936));
  NOT NOT1_4086(.VSS(VSS),.VDD(VDD),.Y(g34272),.A(g34229));
  NOT NOT1_4087(.VSS(VSS),.VDD(VDD),.Y(g24525),.A(g22670));
  NOT NOT1_4088(.VSS(VSS),.VDD(VDD),.Y(g24424),.A(g22722));
  NOT NOT1_4089(.VSS(VSS),.VDD(VDD),.Y(I11623),.A(g28));
  NOT NOT1_4090(.VSS(VSS),.VDD(VDD),.Y(g13132),.A(g10632));
  NOT NOT1_4091(.VSS(VSS),.VDD(VDD),.Y(g17685),.A(I18662));
  NOT NOT1_4092(.VSS(VSS),.VDD(VDD),.Y(g17676),.A(g12941));
  NOT NOT1_4093(.VSS(VSS),.VDD(VDD),.Y(g13869),.A(g10831));
  NOT NOT1_4094(.VSS(VSS),.VDD(VDD),.Y(g20558),.A(I20650));
  NOT NOT1_4095(.VSS(VSS),.VDD(VDD),.Y(g8680),.A(g686));
  NOT NOT1_4096(.VSS(VSS),.VDD(VDD),.Y(g22936),.A(g20283));
  NOT NOT1_4097(.VSS(VSS),.VDD(VDD),.Y(I13623),.A(g4294));
  NOT NOT1_4098(.VSS(VSS),.VDD(VDD),.Y(I21486),.A(g18727));
  NOT NOT1_4099(.VSS(VSS),.VDD(VDD),.Y(g17953),.A(I18861));
  NOT NOT1_4100(.VSS(VSS),.VDD(VDD),.Y(I22327),.A(g19367));
  NOT NOT1_4101(.VSS(VSS),.VDD(VDD),.Y(g23339),.A(g21070));
  NOT NOT1_4102(.VSS(VSS),.VDD(VDD),.Y(g8353),.A(I12530));
  NOT NOT1_4103(.VSS(VSS),.VDD(VDD),.Y(g18938),.A(g16053));
  NOT NOT1_4104(.VSS(VSS),.VDD(VDD),.Y(g23943),.A(g19147));
  NOT NOT1_4105(.VSS(VSS),.VDD(VDD),.Y(g18093),.A(I18885));
  NOT NOT1_4106(.VSS(VSS),.VDD(VDD),.Y(I13037),.A(g4304));
  NOT NOT1_4107(.VSS(VSS),.VDD(VDD),.Y(I29149),.A(g29384));
  NOT NOT1_4108(.VSS(VSS),.VDD(VDD),.Y(g14431),.A(g12208));
  NOT NOT1_4109(.VSS(VSS),.VDD(VDD),.Y(g31213),.A(I29013));
  NOT NOT1_4110(.VSS(VSS),.VDD(VDD),.Y(g11868),.A(g9185));
  NOT NOT1_4111(.VSS(VSS),.VDD(VDD),.Y(g12864),.A(g10373));
  NOT NOT1_4112(.VSS(VSS),.VDD(VDD),.Y(g13868),.A(g11493));
  NOT NOT1_4113(.VSS(VSS),.VDD(VDD),.Y(g6917),.A(g3684));
  NOT NOT1_4114(.VSS(VSS),.VDD(VDD),.Y(g8744),.A(g691));
  NOT NOT1_4115(.VSS(VSS),.VDD(VDD),.Y(g23338),.A(g20453));
  NOT NOT1_4116(.VSS(VSS),.VDD(VDD),.Y(g18065),.A(I18875));
  NOT NOT1_4117(.VSS(VSS),.VDD(VDD),.Y(g24893),.A(I24060));
  NOT NOT1_4118(.VSS(VSS),.VDD(VDD),.Y(g12749),.A(g7074));
  NOT NOT1_4119(.VSS(VSS),.VDD(VDD),.Y(g19435),.A(g16449));
  NOT NOT1_4120(.VSS(VSS),.VDD(VDD),.Y(g9162),.A(g622));
  NOT NOT1_4121(.VSS(VSS),.VDD(VDD),.Y(g9019),.A(I12950));
  NOT NOT1_4122(.VSS(VSS),.VDD(VDD),.Y(g17417),.A(g14804));
  NOT NOT1_4123(.VSS(VSS),.VDD(VDD),.Y(I18609),.A(g5976));
  NOT NOT1_4124(.VSS(VSS),.VDD(VDD),.Y(g7886),.A(g1442));
  NOT NOT1_4125(.VSS(VSS),.VDD(VDD),.Y(g20544),.A(g15171));
  NOT NOT1_4126(.VSS(VSS),.VDD(VDD),.Y(g23969),.A(g19277));
  NOT NOT1_4127(.VSS(VSS),.VDD(VDD),.Y(g32626),.A(g30614));
  NOT NOT1_4128(.VSS(VSS),.VDD(VDD),.Y(g28039),.A(g26365));
  NOT NOT1_4129(.VSS(VSS),.VDD(VDD),.Y(I32195),.A(g33628));
  NOT NOT1_4130(.VSS(VSS),.VDD(VDD),.Y(I13352),.A(g4146));
  NOT NOT1_4131(.VSS(VSS),.VDD(VDD),.Y(g11709),.A(I14584));
  NOT NOT1_4132(.VSS(VSS),.VDD(VDD),.Y(g30997),.A(g29702));
  NOT NOT1_4133(.VSS(VSS),.VDD(VDD),.Y(g10156),.A(g2675));
  NOT NOT1_4134(.VSS(VSS),.VDD(VDD),.Y(g20713),.A(g15277));
  NOT NOT1_4135(.VSS(VSS),.VDD(VDD),.Y(g21060),.A(g15509));
  NOT NOT1_4136(.VSS(VSS),.VDD(VDD),.Y(g34997),.A(I33291));
  NOT NOT1_4137(.VSS(VSS),.VDD(VDD),.Y(I12991),.A(g6752));
  NOT NOT1_4138(.VSS(VSS),.VDD(VDD),.Y(g23060),.A(g19908));
  NOT NOT1_4139(.VSS(VSS),.VDD(VDD),.Y(g23968),.A(g18833));
  NOT NOT1_4140(.VSS(VSS),.VDD(VDD),.Y(g18875),.A(g15171));
  NOT NOT1_4141(.VSS(VSS),.VDD(VDD),.Y(g32533),.A(g30614));
  NOT NOT1_4142(.VSS(VSS),.VDD(VDD),.Y(g8558),.A(g3787));
  NOT NOT1_4143(.VSS(VSS),.VDD(VDD),.Y(g28038),.A(g26365));
  NOT NOT1_4144(.VSS(VSS),.VDD(VDD),.Y(I32525),.A(g34285));
  NOT NOT1_4145(.VSS(VSS),.VDD(VDD),.Y(g13259),.A(I15824));
  NOT NOT1_4146(.VSS(VSS),.VDD(VDD),.Y(g33912),.A(I31770));
  NOT NOT1_4147(.VSS(VSS),.VDD(VDD),.Y(g19744),.A(g15885));
  NOT NOT1_4148(.VSS(VSS),.VDD(VDD),.Y(g16620),.A(I17808));
  NOT NOT1_4149(.VSS(VSS),.VDD(VDD),.Y(g7314),.A(g1740));
  NOT NOT1_4150(.VSS(VSS),.VDD(VDD),.Y(g10180),.A(g2259));
  NOT NOT1_4151(.VSS(VSS),.VDD(VDD),.Y(I14006),.A(g9104));
  NOT NOT1_4152(.VSS(VSS),.VDD(VDD),.Y(I17108),.A(g13782));
  NOT NOT1_4153(.VSS(VSS),.VDD(VDD),.Y(I14475),.A(g10175));
  NOT NOT1_4154(.VSS(VSS),.VDD(VDD),.Y(g11471),.A(g7626));
  NOT NOT1_4155(.VSS(VSS),.VDD(VDD),.Y(g19345),.A(g17591));
  NOT NOT1_4156(.VSS(VSS),.VDD(VDD),.Y(g25099),.A(g22369));
  NOT NOT1_4157(.VSS(VSS),.VDD(VDD),.Y(g13087),.A(g12012));
  NOT NOT1_4158(.VSS(VSS),.VDD(VDD),.Y(g32775),.A(g30825));
  NOT NOT1_4159(.VSS(VSS),.VDD(VDD),.Y(g25388),.A(g22763));
  NOT NOT1_4160(.VSS(VSS),.VDD(VDD),.Y(g25324),.A(g22228));
  NOT NOT1_4161(.VSS(VSS),.VDD(VDD),.Y(I14727),.A(g7753));
  NOT NOT1_4162(.VSS(VSS),.VDD(VDD),.Y(g13258),.A(I15821));
  NOT NOT1_4163(.VSS(VSS),.VDD(VDD),.Y(g12900),.A(g10406));
  NOT NOT1_4164(.VSS(VSS),.VDD(VDD),.Y(g19399),.A(g16489));
  NOT NOT1_4165(.VSS(VSS),.VDD(VDD),.Y(g20610),.A(g18008));
  NOT NOT1_4166(.VSS(VSS),.VDD(VDD),.Y(g7870),.A(g1193));
  NOT NOT1_4167(.VSS(VSS),.VDD(VDD),.Y(g21411),.A(g15426));
  NOT NOT1_4168(.VSS(VSS),.VDD(VDD),.Y(g17762),.A(g13000));
  NOT NOT1_4169(.VSS(VSS),.VDD(VDD),.Y(g20705),.A(I20793));
  NOT NOT1_4170(.VSS(VSS),.VDD(VDD),.Y(g34766),.A(g34703));
  NOT NOT1_4171(.VSS(VSS),.VDD(VDD),.Y(g23870),.A(g21293));
  NOT NOT1_4172(.VSS(VSS),.VDD(VDD),.Y(I16010),.A(g11148));
  NOT NOT1_4173(.VSS(VSS),.VDD(VDD),.Y(g23411),.A(g20734));
  NOT NOT1_4174(.VSS(VSS),.VDD(VDD),.Y(g23527),.A(g21611));
  NOT NOT1_4175(.VSS(VSS),.VDD(VDD),.Y(g28187),.A(I26710));
  NOT NOT1_4176(.VSS(VSS),.VDD(VDD),.Y(I14222),.A(g8286));
  NOT NOT1_4177(.VSS(VSS),.VDD(VDD),.Y(I21922),.A(g21335));
  NOT NOT1_4178(.VSS(VSS),.VDD(VDD),.Y(g25534),.A(g22763));
  NOT NOT1_4179(.VSS(VSS),.VDD(VDD),.Y(g15932),.A(I17395));
  NOT NOT1_4180(.VSS(VSS),.VDD(VDD),.Y(g25098),.A(g22369));
  NOT NOT1_4181(.VSS(VSS),.VDD(VDD),.Y(g10335),.A(g4483));
  NOT NOT1_4182(.VSS(VSS),.VDD(VDD),.Y(I23321),.A(g21693));
  NOT NOT1_4183(.VSS(VSS),.VDD(VDD),.Y(g7650),.A(g4064));
  NOT NOT1_4184(.VSS(VSS),.VDD(VDD),.Y(g27101),.A(g26770));
  NOT NOT1_4185(.VSS(VSS),.VDD(VDD),.Y(g25272),.A(g23715));
  NOT NOT1_4186(.VSS(VSS),.VDD(VDD),.Y(g29862),.A(g28406));
  NOT NOT1_4187(.VSS(VSS),.VDD(VDD),.Y(g24042),.A(g20014));
  NOT NOT1_4188(.VSS(VSS),.VDD(VDD),.Y(g33072),.A(g31945));
  NOT NOT1_4189(.VSS(VSS),.VDD(VDD),.Y(g20189),.A(I20447));
  NOT NOT1_4190(.VSS(VSS),.VDD(VDD),.Y(g19398),.A(g16489));
  NOT NOT1_4191(.VSS(VSS),.VDD(VDD),.Y(g20679),.A(g15634));
  NOT NOT1_4192(.VSS(VSS),.VDD(VDD),.Y(I29368),.A(g30321));
  NOT NOT1_4193(.VSS(VSS),.VDD(VDD),.Y(g17423),.A(I18360));
  NOT NOT1_4194(.VSS(VSS),.VDD(VDD),.Y(g16971),.A(I18131));
  NOT NOT1_4195(.VSS(VSS),.VDD(VDD),.Y(g11043),.A(g8561));
  NOT NOT1_4196(.VSS(VSS),.VDD(VDD),.Y(g12036),.A(g9245));
  NOT NOT1_4197(.VSS(VSS),.VDD(VDD),.Y(g9086),.A(g847));
  NOT NOT1_4198(.VSS(VSS),.VDD(VDD),.Y(g32737),.A(g31327));
  NOT NOT1_4199(.VSS(VSS),.VDD(VDD),.Y(I18813),.A(g5673));
  NOT NOT1_4200(.VSS(VSS),.VDD(VDD),.Y(g17216),.A(g14454));
  NOT NOT1_4201(.VSS(VSS),.VDD(VDD),.Y(g20270),.A(g15277));
  NOT NOT1_4202(.VSS(VSS),.VDD(VDD),.Y(g9728),.A(g5109));
  NOT NOT1_4203(.VSS(VSS),.VDD(VDD),.Y(g19652),.A(g16897));
  NOT NOT1_4204(.VSS(VSS),.VDD(VDD),.Y(I30986),.A(g32437));
  NOT NOT1_4205(.VSS(VSS),.VDD(VDD),.Y(I17750),.A(g14383));
  NOT NOT1_4206(.VSS(VSS),.VDD(VDD),.Y(g22543),.A(g19801));
  NOT NOT1_4207(.VSS(VSS),.VDD(VDD),.Y(g17587),.A(I18518));
  NOT NOT1_4208(.VSS(VSS),.VDD(VDD),.Y(g9730),.A(g5436));
  NOT NOT1_4209(.VSS(VSS),.VDD(VDD),.Y(I31504),.A(g33164));
  NOT NOT1_4210(.VSS(VSS),.VDD(VDD),.Y(g24124),.A(g21209));
  NOT NOT1_4211(.VSS(VSS),.VDD(VDD),.Y(g8092),.A(g1589));
  NOT NOT1_4212(.VSS(VSS),.VDD(VDD),.Y(g14694),.A(I16795));
  NOT NOT1_4213(.VSS(VSS),.VDD(VDD),.Y(g29948),.A(g28853));
  NOT NOT1_4214(.VSS(VSS),.VDD(VDD),.Y(g8492),.A(g3396));
  NOT NOT1_4215(.VSS(VSS),.VDD(VDD),.Y(g9185),.A(I13007));
  NOT NOT1_4216(.VSS(VSS),.VDD(VDD),.Y(g23503),.A(g21468));
  NOT NOT1_4217(.VSS(VSS),.VDD(VDD),.Y(g23894),.A(g19074));
  NOT NOT1_4218(.VSS(VSS),.VDD(VDD),.Y(g19263),.A(I19799));
  NOT NOT1_4219(.VSS(VSS),.VDD(VDD),.Y(g32697),.A(g31070));
  NOT NOT1_4220(.VSS(VSS),.VDD(VDD),.Y(g27064),.A(I25786));
  NOT NOT1_4221(.VSS(VSS),.VDD(VDD),.Y(I18674),.A(g13101));
  NOT NOT1_4222(.VSS(VSS),.VDD(VDD),.Y(g25032),.A(g23639));
  NOT NOT1_4223(.VSS(VSS),.VDD(VDD),.Y(g20383),.A(g15373));
  NOT NOT1_4224(.VSS(VSS),.VDD(VDD),.Y(g32856),.A(g31021));
  NOT NOT1_4225(.VSS(VSS),.VDD(VDD),.Y(I28913),.A(g30322));
  NOT NOT1_4226(.VSS(VSS),.VDD(VDD),.Y(g11810),.A(g9664));
  NOT NOT1_4227(.VSS(VSS),.VDD(VDD),.Y(g25140),.A(g22228));
  NOT NOT1_4228(.VSS(VSS),.VDD(VDD),.Y(g9070),.A(g5428));
  NOT NOT1_4229(.VSS(VSS),.VDD(VDD),.Y(g8714),.A(g4859));
  NOT NOT1_4230(.VSS(VSS),.VDD(VDD),.Y(g7594),.A(I12064));
  NOT NOT1_4231(.VSS(VSS),.VDD(VDD),.Y(g31820),.A(g29385));
  NOT NOT1_4232(.VSS(VSS),.VDD(VDD),.Y(g10487),.A(g10233));
  NOT NOT1_4233(.VSS(VSS),.VDD(VDD),.Y(g32880),.A(g30614));
  NOT NOT1_4234(.VSS(VSS),.VDD(VDD),.Y(g13068),.A(I15697));
  NOT NOT1_4235(.VSS(VSS),.VDD(VDD),.Y(g25997),.A(I25095));
  NOT NOT1_4236(.VSS(VSS),.VDD(VDD),.Y(g7972),.A(g1046));
  NOT NOT1_4237(.VSS(VSS),.VDD(VDD),.Y(g24030),.A(g21127));
  NOT NOT1_4238(.VSS(VSS),.VDD(VDD),.Y(g20267),.A(g17955));
  NOT NOT1_4239(.VSS(VSS),.VDD(VDD),.Y(g24093),.A(g20998));
  NOT NOT1_4240(.VSS(VSS),.VDD(VDD),.Y(g10502),.A(g8876));
  NOT NOT1_4241(.VSS(VSS),.VDD(VDD),.Y(g26776),.A(g25498));
  NOT NOT1_4242(.VSS(VSS),.VDD(VDD),.Y(g23714),.A(g20751));
  NOT NOT1_4243(.VSS(VSS),.VDD(VDD),.Y(I27758),.A(g28119));
  NOT NOT1_4244(.VSS(VSS),.VDD(VDD),.Y(g23450),.A(I22571));
  NOT NOT1_4245(.VSS(VSS),.VDD(VDD),.Y(I29228),.A(g30314));
  NOT NOT1_4246(.VSS(VSS),.VDD(VDD),.Y(g32512),.A(g31566));
  NOT NOT1_4247(.VSS(VSS),.VDD(VDD),.Y(g7806),.A(g4681));
  NOT NOT1_4248(.VSS(VSS),.VDD(VDD),.Y(I15878),.A(g11249));
  NOT NOT1_4249(.VSS(VSS),.VDD(VDD),.Y(g20065),.A(g16846));
  NOT NOT1_4250(.VSS(VSS),.VDD(VDD),.Y(g31846),.A(g29385));
  NOT NOT1_4251(.VSS(VSS),.VDD(VDD),.Y(g7943),.A(g1395));
  NOT NOT1_4252(.VSS(VSS),.VDD(VDD),.Y(g24065),.A(g20982));
  NOT NOT1_4253(.VSS(VSS),.VDD(VDD),.Y(g11878),.A(I14690));
  NOT NOT1_4254(.VSS(VSS),.VDD(VDD),.Y(g19361),.A(I19843));
  NOT NOT1_4255(.VSS(VSS),.VDD(VDD),.Y(I20609),.A(g16539));
  NOT NOT1_4256(.VSS(VSS),.VDD(VDD),.Y(I12758),.A(g4093));
  NOT NOT1_4257(.VSS(VSS),.VDD(VDD),.Y(g23819),.A(g19147));
  NOT NOT1_4258(.VSS(VSS),.VDD(VDD),.Y(g12874),.A(g10383));
  NOT NOT1_4259(.VSS(VSS),.VDD(VDD),.Y(g26754),.A(g25300));
  NOT NOT1_4260(.VSS(VSS),.VDD(VDD),.Y(g34472),.A(I32525));
  NOT NOT1_4261(.VSS(VSS),.VDD(VDD),.Y(g25766),.A(g24439));
  NOT NOT1_4262(.VSS(VSS),.VDD(VDD),.Y(g28479),.A(g27654));
  NOT NOT1_4263(.VSS(VSS),.VDD(VDD),.Y(I32678),.A(g34428));
  NOT NOT1_4264(.VSS(VSS),.VDD(VDD),.Y(g23202),.A(I22302));
  NOT NOT1_4265(.VSS(VSS),.VDD(VDD),.Y(g14443),.A(I16596));
  NOT NOT1_4266(.VSS(VSS),.VDD(VDD),.Y(g23257),.A(g20924));
  NOT NOT1_4267(.VSS(VSS),.VDD(VDD),.Y(g26859),.A(I25591));
  NOT NOT1_4268(.VSS(VSS),.VDD(VDD),.Y(g27009),.A(g25911));
  NOT NOT1_4269(.VSS(VSS),.VDD(VDD),.Y(g26825),.A(I25541));
  NOT NOT1_4270(.VSS(VSS),.VDD(VDD),.Y(g21055),.A(g15224));
  NOT NOT1_4271(.VSS(VSS),.VDD(VDD),.Y(g23496),.A(g20248));
  NOT NOT1_4272(.VSS(VSS),.VDD(VDD),.Y(g7322),.A(g1862));
  NOT NOT1_4273(.VSS(VSS),.VDD(VDD),.Y(g16228),.A(I17569));
  NOT NOT1_4274(.VSS(VSS),.VDD(VDD),.Y(g20219),.A(I20495));
  NOT NOT1_4275(.VSS(VSS),.VDD(VDD),.Y(g23055),.A(g20887));
  NOT NOT1_4276(.VSS(VSS),.VDD(VDD),.Y(g6990),.A(g4742));
  NOT NOT1_4277(.VSS(VSS),.VDD(VDD),.Y(g17242),.A(g14454));
  NOT NOT1_4278(.VSS(VSS),.VDD(VDD),.Y(g34246),.A(I32237));
  NOT NOT1_4279(.VSS(VSS),.VDD(VDD),.Y(g10278),.A(g4628));
  NOT NOT1_4280(.VSS(VSS),.VDD(VDD),.Y(g33413),.A(g31971));
  NOT NOT1_4281(.VSS(VSS),.VDD(VDD),.Y(g29847),.A(g28395));
  NOT NOT1_4282(.VSS(VSS),.VDD(VDD),.Y(I29582),.A(g30591));
  NOT NOT1_4283(.VSS(VSS),.VDD(VDD),.Y(g23111),.A(g20391));
  NOT NOT1_4284(.VSS(VSS),.VDD(VDD),.Y(g12009),.A(I14862));
  NOT NOT1_4285(.VSS(VSS),.VDD(VDD),.Y(g21070),.A(I20937));
  NOT NOT1_4286(.VSS(VSS),.VDD(VDD),.Y(g6888),.A(I11701));
  NOT NOT1_4287(.VSS(VSS),.VDD(VDD),.Y(g22974),.A(g20330));
  NOT NOT1_4288(.VSS(VSS),.VDD(VDD),.Y(g32831),.A(g31376));
  NOT NOT1_4289(.VSS(VSS),.VDD(VDD),.Y(g33691),.A(I31528));
  NOT NOT1_4290(.VSS(VSS),.VDD(VDD),.Y(g32445),.A(I29973));
  NOT NOT1_4291(.VSS(VSS),.VDD(VDD),.Y(I32938),.A(g34663));
  NOT NOT1_4292(.VSS(VSS),.VDD(VDD),.Y(I32093),.A(g33670));
  NOT NOT1_4293(.VSS(VSS),.VDD(VDD),.Y(I13276),.A(g5798));
  NOT NOT1_4294(.VSS(VSS),.VDD(VDD),.Y(g16716),.A(g13948));
  NOT NOT1_4295(.VSS(VSS),.VDD(VDD),.Y(g9678),.A(g5406));
  NOT NOT1_4296(.VSS(VSS),.VDD(VDD),.Y(g10039),.A(g2273));
  NOT NOT1_4297(.VSS(VSS),.VDD(VDD),.Y(g10306),.A(I13726));
  NOT NOT1_4298(.VSS(VSS),.VDD(VDD),.Y(g32499),.A(g31376));
  NOT NOT1_4299(.VSS(VSS),.VDD(VDD),.Y(g23986),.A(g18833));
  NOT NOT1_4300(.VSS(VSS),.VDD(VDD),.Y(g30591),.A(I28851));
  NOT NOT1_4301(.VSS(VSS),.VDD(VDD),.Y(g6956),.A(g4242));
  NOT NOT1_4302(.VSS(VSS),.VDD(VDD),.Y(g18984),.A(g17486));
  NOT NOT1_4303(.VSS(VSS),.VDD(VDD),.Y(g8623),.A(g3990));
  NOT NOT1_4304(.VSS(VSS),.VDD(VDD),.Y(I11809),.A(g6741));
  NOT NOT1_4305(.VSS(VSS),.VDD(VDD),.Y(g34591),.A(I32681));
  NOT NOT1_4306(.VSS(VSS),.VDD(VDD),.Y(I18214),.A(g12918));
  NOT NOT1_4307(.VSS(VSS),.VDD(VDD),.Y(g12892),.A(g10398));
  NOT NOT1_4308(.VSS(VSS),.VDD(VDD),.Y(g34785),.A(I32985));
  NOT NOT1_4309(.VSS(VSS),.VDD(VDD),.Y(g16582),.A(g13915));
  NOT NOT1_4310(.VSS(VSS),.VDD(VDD),.Y(g17772),.A(g14297));
  NOT NOT1_4311(.VSS(VSS),.VDD(VDD),.Y(g34776),.A(I32970));
  NOT NOT1_4312(.VSS(VSS),.VDD(VDD),.Y(g11425),.A(g7640));
  NOT NOT1_4313(.VSS(VSS),.VDD(VDD),.Y(g10038),.A(g2241));
  NOT NOT1_4314(.VSS(VSS),.VDD(VDD),.Y(g32498),.A(g31566));
  NOT NOT1_4315(.VSS(VSS),.VDD(VDD),.Y(g23384),.A(I22485));
  NOT NOT1_4316(.VSS(VSS),.VDD(VDD),.Y(g17639),.A(I18600));
  NOT NOT1_4317(.VSS(VSS),.VDD(VDD),.Y(I12141),.A(g599));
  NOT NOT1_4318(.VSS(VSS),.VDD(VDD),.Y(g34147),.A(g33823));
  NOT NOT1_4319(.VSS(VSS),.VDD(VDD),.Y(g9682),.A(I13280));
  NOT NOT1_4320(.VSS(VSS),.VDD(VDD),.Y(g9766),.A(g2748));
  NOT NOT1_4321(.VSS(VSS),.VDD(VDD),.Y(g15811),.A(g13125));
  NOT NOT1_4322(.VSS(VSS),.VDD(VDD),.Y(g16310),.A(g13223));
  NOT NOT1_4323(.VSS(VSS),.VDD(VDD),.Y(g7096),.A(g6537));
  NOT NOT1_4324(.VSS(VSS),.VDD(VDD),.Y(g10815),.A(g9917));
  NOT NOT1_4325(.VSS(VSS),.VDD(VDD),.Y(g13458),.A(g11048));
  NOT NOT1_4326(.VSS(VSS),.VDD(VDD),.Y(g24160),.A(I23324));
  NOT NOT1_4327(.VSS(VSS),.VDD(VDD),.Y(I15918),.A(g12381));
  NOT NOT1_4328(.VSS(VSS),.VDD(VDD),.Y(g9305),.A(g5381));
  NOT NOT1_4329(.VSS(VSS),.VDD(VDD),.Y(g7496),.A(g5969));
  NOT NOT1_4330(.VSS(VSS),.VDD(VDD),.Y(g33929),.A(I31803));
  NOT NOT1_4331(.VSS(VSS),.VDD(VDD),.Y(g16627),.A(I17819));
  NOT NOT1_4332(.VSS(VSS),.VDD(VDD),.Y(g17638),.A(g14838));
  NOT NOT1_4333(.VSS(VSS),.VDD(VDD),.Y(g22841),.A(g20391));
  NOT NOT1_4334(.VSS(VSS),.VDD(VDD),.Y(g34950),.A(g34940));
  NOT NOT1_4335(.VSS(VSS),.VDD(VDD),.Y(g12914),.A(g12235));
  NOT NOT1_4336(.VSS(VSS),.VDD(VDD),.Y(g13010),.A(I15620));
  NOT NOT1_4337(.VSS(VSS),.VDD(VDD),.Y(g32611),.A(g31154));
  NOT NOT1_4338(.VSS(VSS),.VDD(VDD),.Y(g7845),.A(g1146));
  NOT NOT1_4339(.VSS(VSS),.VDD(VDD),.Y(I33232),.A(g34957));
  NOT NOT1_4340(.VSS(VSS),.VDD(VDD),.Y(g25451),.A(g22228));
  NOT NOT1_4341(.VSS(VSS),.VDD(VDD),.Y(g32722),.A(g30937));
  NOT NOT1_4342(.VSS(VSS),.VDD(VDD),.Y(g25220),.A(I24396));
  NOT NOT1_4343(.VSS(VSS),.VDD(VDD),.Y(g32924),.A(g30937));
  NOT NOT1_4344(.VSS(VSS),.VDD(VDD),.Y(g33928),.A(I31800));
  NOT NOT1_4345(.VSS(VSS),.VDD(VDD),.Y(g19947),.A(g17226));
  NOT NOT1_4346(.VSS(VSS),.VDD(VDD),.Y(g7195),.A(g25));
  NOT NOT1_4347(.VSS(VSS),.VDD(VDD),.Y(g12907),.A(g10415));
  NOT NOT1_4348(.VSS(VSS),.VDD(VDD),.Y(g20617),.A(g15277));
  NOT NOT1_4349(.VSS(VSS),.VDD(VDD),.Y(g17416),.A(g14956));
  NOT NOT1_4350(.VSS(VSS),.VDD(VDD),.Y(g7395),.A(g6005));
  NOT NOT1_4351(.VSS(VSS),.VDD(VDD),.Y(g7891),.A(g2994));
  NOT NOT1_4352(.VSS(VSS),.VDD(VDD),.Y(g8651),.A(g758));
  NOT NOT1_4353(.VSS(VSS),.VDD(VDD),.Y(g16958),.A(g14238));
  NOT NOT1_4354(.VSS(VSS),.VDD(VDD),.Y(g9748),.A(g114));
  NOT NOT1_4355(.VSS(VSS),.VDD(VDD),.Y(g13545),.A(I16010));
  NOT NOT1_4356(.VSS(VSS),.VDD(VDD),.Y(g23877),.A(g19147));
  NOT NOT1_4357(.VSS(VSS),.VDD(VDD),.Y(g19273),.A(g16100));
  NOT NOT1_4358(.VSS(VSS),.VDD(VDD),.Y(g20915),.A(I20882));
  NOT NOT1_4359(.VSS(VSS),.VDD(VDD),.Y(g7913),.A(g1052));
  NOT NOT1_4360(.VSS(VSS),.VDD(VDD),.Y(g27074),.A(I25790));
  NOT NOT1_4361(.VSS(VSS),.VDD(VDD),.Y(g28321),.A(g27317));
  NOT NOT1_4362(.VSS(VSS),.VDD(VDD),.Y(I32837),.A(g34498));
  NOT NOT1_4363(.VSS(VSS),.VDD(VDD),.Y(g30996),.A(g29694));
  NOT NOT1_4364(.VSS(VSS),.VDD(VDD),.Y(g25246),.A(g23828));
  NOT NOT1_4365(.VSS(VSS),.VDD(VDD),.Y(g34151),.A(I32106));
  NOT NOT1_4366(.VSS(VSS),.VDD(VDD),.Y(I12135),.A(g807));
  NOT NOT1_4367(.VSS(VSS),.VDD(VDD),.Y(g10143),.A(g568));
  NOT NOT1_4368(.VSS(VSS),.VDD(VDD),.Y(g29213),.A(I27555));
  NOT NOT1_4369(.VSS(VSS),.VDD(VDD),.Y(g34996),.A(I33288));
  NOT NOT1_4370(.VSS(VSS),.VDD(VDD),.Y(g23019),.A(g19866));
  NOT NOT1_4371(.VSS(VSS),.VDD(VDD),.Y(I33261),.A(g34977));
  NOT NOT1_4372(.VSS(VSS),.VDD(VDD),.Y(g8285),.A(I12497));
  NOT NOT1_4373(.VSS(VSS),.VDD(VDD),.Y(g12074),.A(I14932));
  NOT NOT1_4374(.VSS(VSS),.VDD(VDD),.Y(I25695),.A(g25690));
  NOT NOT1_4375(.VSS(VSS),.VDD(VDD),.Y(g9226),.A(g1564));
  NOT NOT1_4376(.VSS(VSS),.VDD(VDD),.Y(g20277),.A(g16487));
  NOT NOT1_4377(.VSS(VSS),.VDD(VDD),.Y(g16603),.A(I17787));
  NOT NOT1_4378(.VSS(VSS),.VDD(VDD),.Y(g16742),.A(g13983));
  NOT NOT1_4379(.VSS(VSS),.VDD(VDD),.Y(g23196),.A(g20785));
  NOT NOT1_4380(.VSS(VSS),.VDD(VDD),.Y(g34844),.A(g34737));
  NOT NOT1_4381(.VSS(VSS),.VDD(VDD),.Y(I22564),.A(g20857));
  NOT NOT1_4382(.VSS(VSS),.VDD(VDD),.Y(g16096),.A(g13530));
  NOT NOT1_4383(.VSS(VSS),.VDD(VDD),.Y(g23018),.A(g19801));
  NOT NOT1_4384(.VSS(VSS),.VDD(VDD),.Y(g32753),.A(g30735));
  NOT NOT1_4385(.VSS(VSS),.VDD(VDD),.Y(g12238),.A(I15102));
  NOT NOT1_4386(.VSS(VSS),.VDD(VDD),.Y(g32461),.A(g30614));
  NOT NOT1_4387(.VSS(VSS),.VDD(VDD),.Y(I21242),.A(g16540));
  NOT NOT1_4388(.VSS(VSS),.VDD(VDD),.Y(g10169),.A(g6395));
  NOT NOT1_4389(.VSS(VSS),.VDD(VDD),.Y(g24075),.A(g19935));
  NOT NOT1_4390(.VSS(VSS),.VDD(VDD),.Y(g17579),.A(g14959));
  NOT NOT1_4391(.VSS(VSS),.VDD(VDD),.Y(g19371),.A(I19857));
  NOT NOT1_4392(.VSS(VSS),.VDD(VDD),.Y(g20595),.A(g15877));
  NOT NOT1_4393(.VSS(VSS),.VDD(VDD),.Y(g23526),.A(g21611));
  NOT NOT1_4394(.VSS(VSS),.VDD(VDD),.Y(g6808),.A(g554));
  NOT NOT1_4395(.VSS(VSS),.VDD(VDD),.Y(g20494),.A(g17847));
  NOT NOT1_4396(.VSS(VSS),.VDD(VDD),.Y(g14169),.A(g12381));
  NOT NOT1_4397(.VSS(VSS),.VDD(VDD),.Y(g8139),.A(g1648));
  NOT NOT1_4398(.VSS(VSS),.VDD(VDD),.Y(I16289),.A(g12107));
  NOT NOT1_4399(.VSS(VSS),.VDD(VDD),.Y(I32455),.A(g34242));
  NOT NOT1_4400(.VSS(VSS),.VDD(VDD),.Y(g7266),.A(g35));
  NOT NOT1_4401(.VSS(VSS),.VDD(VDD),.Y(g29912),.A(g28827));
  NOT NOT1_4402(.VSS(VSS),.VDD(VDD),.Y(g29311),.A(g28998));
  NOT NOT1_4403(.VSS(VSS),.VDD(VDD),.Y(g10410),.A(g7069));
  NOT NOT1_4404(.VSS(VSS),.VDD(VDD),.Y(g20623),.A(g17929));
  NOT NOT1_4405(.VSS(VSS),.VDD(VDD),.Y(g27675),.A(I26309));
  NOT NOT1_4406(.VSS(VSS),.VDD(VDD),.Y(I12049),.A(g781));
  NOT NOT1_4407(.VSS(VSS),.VDD(VDD),.Y(g9373),.A(g5142));
  NOT NOT1_4408(.VSS(VSS),.VDD(VDD),.Y(g17014),.A(g14297));
  NOT NOT1_4409(.VSS(VSS),.VDD(VDD),.Y(g27092),.A(g26737));
  NOT NOT1_4410(.VSS(VSS),.VDD(VDD),.Y(g9091),.A(g1430));
  NOT NOT1_4411(.VSS(VSS),.VDD(VDD),.Y(g20037),.A(g17328));
  NOT NOT1_4412(.VSS(VSS),.VDD(VDD),.Y(g31827),.A(g29385));
  NOT NOT1_4413(.VSS(VSS),.VDD(VDD),.Y(g32736),.A(g30937));
  NOT NOT1_4414(.VSS(VSS),.VDD(VDD),.Y(I32617),.A(g34333));
  NOT NOT1_4415(.VSS(VSS),.VDD(VDD),.Y(g13322),.A(g10918));
  NOT NOT1_4416(.VSS(VSS),.VDD(VDD),.Y(g32887),.A(g30614));
  NOT NOT1_4417(.VSS(VSS),.VDD(VDD),.Y(I32470),.A(g34247));
  NOT NOT1_4418(.VSS(VSS),.VDD(VDD),.Y(g24623),.A(g23076));
  NOT NOT1_4419(.VSS(VSS),.VDD(VDD),.Y(g33827),.A(I31672));
  NOT NOT1_4420(.VSS(VSS),.VDD(VDD),.Y(g9491),.A(g2729));
  NOT NOT1_4421(.VSS(VSS),.VDD(VDD),.Y(I14905),.A(g9822));
  NOT NOT1_4422(.VSS(VSS),.VDD(VDD),.Y(g24037),.A(g21127));
  NOT NOT1_4423(.VSS(VSS),.VDD(VDD),.Y(g34420),.A(g34152));
  NOT NOT1_4424(.VSS(VSS),.VDD(VDD),.Y(g16429),.A(I17671));
  NOT NOT1_4425(.VSS(VSS),.VDD(VDD),.Y(I11665),.A(g1589));
  NOT NOT1_4426(.VSS(VSS),.VDD(VDD),.Y(g20782),.A(g15853));
  NOT NOT1_4427(.VSS(VSS),.VDD(VDD),.Y(g21457),.A(g17367));
  NOT NOT1_4428(.VSS(VSS),.VDD(VDD),.Y(g13901),.A(g11480));
  NOT NOT1_4429(.VSS(VSS),.VDD(VDD),.Y(g23402),.A(g20875));
  NOT NOT1_4430(.VSS(VSS),.VDD(VDD),.Y(I13166),.A(g5101));
  NOT NOT1_4431(.VSS(VSS),.VDD(VDD),.Y(g32529),.A(g30735));
  NOT NOT1_4432(.VSS(VSS),.VDD(VDD),.Y(g23457),.A(I22580));
  NOT NOT1_4433(.VSS(VSS),.VDD(VDD),.Y(g25370),.A(g22228));
  NOT NOT1_4434(.VSS(VSS),.VDD(VDD),.Y(g8795),.A(I12793));
  NOT NOT1_4435(.VSS(VSS),.VDD(VDD),.Y(g10363),.A(I13779));
  NOT NOT1_4436(.VSS(VSS),.VDD(VDD),.Y(I24400),.A(g23954));
  NOT NOT1_4437(.VSS(VSS),.VDD(VDD),.Y(g10217),.A(g2102));
  NOT NOT1_4438(.VSS(VSS),.VDD(VDD),.Y(I14593),.A(g9978));
  NOT NOT1_4439(.VSS(VSS),.VDD(VDD),.Y(g30318),.A(g28274));
  NOT NOT1_4440(.VSS(VSS),.VDD(VDD),.Y(g14363),.A(I16521));
  NOT NOT1_4441(.VSS(VSS),.VDD(VDD),.Y(g14217),.A(I16417));
  NOT NOT1_4442(.VSS(VSS),.VDD(VDD),.Y(g9283),.A(g1736));
  NOT NOT1_4443(.VSS(VSS),.VDD(VDD),.Y(I14346),.A(g10233));
  NOT NOT1_4444(.VSS(VSS),.VDD(VDD),.Y(g16428),.A(I17668));
  NOT NOT1_4445(.VSS(VSS),.VDD(VDD),.Y(g9369),.A(g5084));
  NOT NOT1_4446(.VSS(VSS),.VDD(VDD),.Y(g32528),.A(g31554));
  NOT NOT1_4447(.VSS(VSS),.VDD(VDD),.Y(g32696),.A(g30825));
  NOT NOT1_4448(.VSS(VSS),.VDD(VDD),.Y(g9007),.A(g1083));
  NOT NOT1_4449(.VSS(VSS),.VDD(VDD),.Y(I21230),.A(g16540));
  NOT NOT1_4450(.VSS(VSS),.VDD(VDD),.Y(g32843),.A(g31021));
  NOT NOT1_4451(.VSS(VSS),.VDD(VDD),.Y(g6957),.A(g2932));
  NOT NOT1_4452(.VSS(VSS),.VDD(VDD),.Y(g24419),.A(g22722));
  NOT NOT1_4453(.VSS(VSS),.VDD(VDD),.Y(g32393),.A(g30922));
  NOT NOT1_4454(.VSS(VSS),.VDD(VDD),.Y(g9407),.A(g6549));
  NOT NOT1_4455(.VSS(VSS),.VDD(VDD),.Y(I15295),.A(g8515));
  NOT NOT1_4456(.VSS(VSS),.VDD(VDD),.Y(I11892),.A(g4408));
  NOT NOT1_4457(.VSS(VSS),.VDD(VDD),.Y(g34059),.A(g33658));
  NOT NOT1_4458(.VSS(VSS),.VDD(VDD),.Y(g8672),.A(g4669));
  NOT NOT1_4459(.VSS(VSS),.VDD(VDD),.Y(g9920),.A(g4322));
  NOT NOT1_4460(.VSS(VSS),.VDD(VDD),.Y(I15144),.A(g5659));
  NOT NOT1_4461(.VSS(VSS),.VDD(VDD),.Y(I13892),.A(g1576));
  NOT NOT1_4462(.VSS(VSS),.VDD(VDD),.Y(g31803),.A(g29385));
  NOT NOT1_4463(.VSS(VSS),.VDD(VDD),.Y(g32764),.A(g30937));
  NOT NOT1_4464(.VSS(VSS),.VDD(VDD),.Y(g24155),.A(I23309));
  NOT NOT1_4465(.VSS(VSS),.VDD(VDD),.Y(g24418),.A(g22722));
  NOT NOT1_4466(.VSS(VSS),.VDD(VDD),.Y(I32467),.A(g34246));
  NOT NOT1_4467(.VSS(VSS),.VDD(VDD),.Y(g20266),.A(g17873));
  NOT NOT1_4468(.VSS(VSS),.VDD(VDD),.Y(g8477),.A(g3061));
  NOT NOT1_4469(.VSS(VSS),.VDD(VDD),.Y(g34540),.A(I32607));
  NOT NOT1_4470(.VSS(VSS),.VDD(VDD),.Y(g11823),.A(I14647));
  NOT NOT1_4471(.VSS(VSS),.VDD(VDD),.Y(g13680),.A(I16077));
  NOT NOT1_4472(.VSS(VSS),.VDD(VDD),.Y(g17615),.A(I18574));
  NOT NOT1_4473(.VSS(VSS),.VDD(VDD),.Y(g12883),.A(g10390));
  NOT NOT1_4474(.VSS(VSS),.VDD(VDD),.Y(g13144),.A(I15773));
  NOT NOT1_4475(.VSS(VSS),.VDD(VDD),.Y(g22493),.A(g19801));
  NOT NOT1_4476(.VSS(VSS),.VDD(VDD),.Y(g7097),.A(I11809));
  NOT NOT1_4477(.VSS(VSS),.VDD(VDD),.Y(g23001),.A(g19801));
  NOT NOT1_4478(.VSS(VSS),.VDD(VDD),.Y(g34058),.A(g33660));
  NOT NOT1_4479(.VSS(VSS),.VDD(VDD),.Y(g24170),.A(I23354));
  NOT NOT1_4480(.VSS(VSS),.VDD(VDD),.Y(g32869),.A(g30735));
  NOT NOT1_4481(.VSS(VSS),.VDD(VDD),.Y(I18882),.A(g16580));
  NOT NOT1_4482(.VSS(VSS),.VDD(VDD),.Y(g32960),.A(g31327));
  NOT NOT1_4483(.VSS(VSS),.VDD(VDD),.Y(I18414),.A(g14359));
  NOT NOT1_4484(.VSS(VSS),.VDD(VDD),.Y(g7497),.A(g6358));
  NOT NOT1_4485(.VSS(VSS),.VDD(VDD),.Y(I14797),.A(g9636));
  NOT NOT1_4486(.VSS(VSS),.VDD(VDD),.Y(g19421),.A(g16326));
  NOT NOT1_4487(.VSS(VSS),.VDD(VDD),.Y(g17720),.A(g15045));
  NOT NOT1_4488(.VSS(VSS),.VDD(VDD),.Y(I33056),.A(g34778));
  NOT NOT1_4489(.VSS(VSS),.VDD(VDD),.Y(I25689),.A(g25688));
  NOT NOT1_4490(.VSS(VSS),.VDD(VDD),.Y(g9582),.A(g703));
  NOT NOT1_4491(.VSS(VSS),.VDD(VDD),.Y(g11336),.A(g7620));
  NOT NOT1_4492(.VSS(VSS),.VDD(VDD),.Y(g7960),.A(g1404));
  NOT NOT1_4493(.VSS(VSS),.VDD(VDD),.Y(g32868),.A(g31376));
  NOT NOT1_4494(.VSS(VSS),.VDD(VDD),.Y(g8205),.A(g2208));
  NOT NOT1_4495(.VSS(VSS),.VDD(VDD),.Y(I32782),.A(g34571));
  NOT NOT1_4496(.VSS(VSS),.VDD(VDD),.Y(g10223),.A(g4561));
  NOT NOT1_4497(.VSS(VSS),.VDD(VDD),.Y(g21689),.A(I21250));
  NOT NOT1_4498(.VSS(VSS),.VDD(VDD),.Y(g23256),.A(g20785));
  NOT NOT1_4499(.VSS(VSS),.VDD(VDD),.Y(I12106),.A(g626));
  NOT NOT1_4500(.VSS(VSS),.VDD(VDD),.Y(I12605),.A(g1570));
  NOT NOT1_4501(.VSS(VSS),.VDD(VDD),.Y(g17430),.A(I18373));
  NOT NOT1_4502(.VSS(VSS),.VDD(VDD),.Y(g17746),.A(g14825));
  NOT NOT1_4503(.VSS(VSS),.VDD(VDD),.Y(g20853),.A(g15595));
  NOT NOT1_4504(.VSS(VSS),.VDD(VDD),.Y(g34044),.A(g33675));
  NOT NOT1_4505(.VSS(VSS),.VDD(VDD),.Y(g21280),.A(g16601));
  NOT NOT1_4506(.VSS(VSS),.VDD(VDD),.Y(g23923),.A(g18997));
  NOT NOT1_4507(.VSS(VSS),.VDD(VDD),.Y(I14409),.A(g8364));
  NOT NOT1_4508(.VSS(VSS),.VDD(VDD),.Y(g29152),.A(g27907));
  NOT NOT1_4509(.VSS(VSS),.VDD(VDD),.Y(g29846),.A(g28391));
  NOT NOT1_4510(.VSS(VSS),.VDD(VDD),.Y(I32352),.A(g34169));
  NOT NOT1_4511(.VSS(VSS),.VDD(VDD),.Y(I29002),.A(g29675));
  NOT NOT1_4512(.VSS(VSS),.VDD(VDD),.Y(g21300),.A(I21047));
  NOT NOT1_4513(.VSS(VSS),.VDD(VDD),.Y(g20167),.A(g16971));
  NOT NOT1_4514(.VSS(VSS),.VDD(VDD),.Y(g20194),.A(g16897));
  NOT NOT1_4515(.VSS(VSS),.VDD(VDD),.Y(g20589),.A(g15224));
  NOT NOT1_4516(.VSS(VSS),.VDD(VDD),.Y(g32709),.A(g30735));
  NOT NOT1_4517(.VSS(VSS),.VDD(VDD),.Y(g11966),.A(I14800));
  NOT NOT1_4518(.VSS(VSS),.VDD(VDD),.Y(g23300),.A(g20283));
  NOT NOT1_4519(.VSS(VSS),.VDD(VDD),.Y(I12463),.A(g4812));
  NOT NOT1_4520(.VSS(VSS),.VDD(VDD),.Y(g17465),.A(g12955));
  NOT NOT1_4521(.VSS(VSS),.VDD(VDD),.Y(g8742),.A(g4035));
  NOT NOT1_4522(.VSS(VSS),.VDD(VDD),.Y(g13966),.A(I16246));
  NOT NOT1_4523(.VSS(VSS),.VDD(VDD),.Y(g10084),.A(g2837));
  NOT NOT1_4524(.VSS(VSS),.VDD(VDD),.Y(g24167),.A(I23345));
  NOT NOT1_4525(.VSS(VSS),.VDD(VDD),.Y(g9415),.A(g2169));
  NOT NOT1_4526(.VSS(VSS),.VDD(VDD),.Y(g19541),.A(g16136));
  NOT NOT1_4527(.VSS(VSS),.VDD(VDD),.Y(g30301),.A(I28548));
  NOT NOT1_4528(.VSS(VSS),.VDD(VDD),.Y(g10110),.A(g661));
  NOT NOT1_4529(.VSS(VSS),.VDD(VDD),.Y(g11631),.A(g8595));
  NOT NOT1_4530(.VSS(VSS),.VDD(VDD),.Y(g19473),.A(g16349));
  NOT NOT1_4531(.VSS(VSS),.VDD(VDD),.Y(g18101),.A(I18909));
  NOT NOT1_4532(.VSS(VSS),.VDD(VDD),.Y(g11017),.A(g10289));
  NOT NOT1_4533(.VSS(VSS),.VDD(VDD),.Y(g20588),.A(g18008));
  NOT NOT1_4534(.VSS(VSS),.VDD(VDD),.Y(g20524),.A(g17873));
  NOT NOT1_4535(.VSS(VSS),.VDD(VDD),.Y(g32708),.A(g31376));
  NOT NOT1_4536(.VSS(VSS),.VDD(VDD),.Y(I32170),.A(g33638));
  NOT NOT1_4537(.VSS(VSS),.VDD(VDD),.Y(I12033),.A(g776));
  NOT NOT1_4538(.VSS(VSS),.VDD(VDD),.Y(g13017),.A(I15633));
  NOT NOT1_4539(.VSS(VSS),.VDD(VDD),.Y(I28174),.A(g28803));
  NOT NOT1_4540(.VSS(VSS),.VDD(VDD),.Y(I29245),.A(g29491));
  NOT NOT1_4541(.VSS(VSS),.VDD(VDD),.Y(g32471),.A(g31376));
  NOT NOT1_4542(.VSS(VSS),.VDD(VDD),.Y(g19789),.A(g17015));
  NOT NOT1_4543(.VSS(VSS),.VDD(VDD),.Y(g24524),.A(g22876));
  NOT NOT1_4544(.VSS(VSS),.VDD(VDD),.Y(g24836),.A(I24008));
  NOT NOT1_4545(.VSS(VSS),.VDD(VDD),.Y(g16129),.A(I17488));
  NOT NOT1_4546(.VSS(VSS),.VDD(VDD),.Y(g25227),.A(g22763));
  NOT NOT1_4547(.VSS(VSS),.VDD(VDD),.Y(g14321),.A(g10874));
  NOT NOT1_4548(.VSS(VSS),.VDD(VDD),.Y(g34739),.A(I32909));
  NOT NOT1_4549(.VSS(VSS),.VDD(VDD),.Y(g10531),.A(g8925));
  NOT NOT1_4550(.VSS(VSS),.VDD(VDD),.Y(g17684),.A(g15036));
  NOT NOT1_4551(.VSS(VSS),.VDD(VDD),.Y(g27438),.A(I26130));
  NOT NOT1_4552(.VSS(VSS),.VDD(VDD),.Y(g14179),.A(g11048));
  NOT NOT1_4553(.VSS(VSS),.VDD(VDD),.Y(g25025),.A(g22498));
  NOT NOT1_4554(.VSS(VSS),.VDD(VDD),.Y(g7267),.A(g1604));
  NOT NOT1_4555(.VSS(VSS),.VDD(VDD),.Y(g24477),.A(I23680));
  NOT NOT1_4556(.VSS(VSS),.VDD(VDD),.Y(g10178),.A(g2126));
  NOT NOT1_4557(.VSS(VSS),.VDD(VDD),.Y(g26632),.A(g25473));
  NOT NOT1_4558(.VSS(VSS),.VDD(VDD),.Y(g24119),.A(g19935));
  NOT NOT1_4559(.VSS(VSS),.VDD(VDD),.Y(g27349),.A(g26352));
  NOT NOT1_4560(.VSS(VSS),.VDD(VDD),.Y(I31650),.A(g33212));
  NOT NOT1_4561(.VSS(VSS),.VDD(VDD),.Y(g23066),.A(g20330));
  NOT NOT1_4562(.VSS(VSS),.VDD(VDD),.Y(I28390),.A(g29185));
  NOT NOT1_4563(.VSS(VSS),.VDD(VDD),.Y(g9721),.A(g5097));
  NOT NOT1_4564(.VSS(VSS),.VDD(VDD),.Y(g23231),.A(g20050));
  NOT NOT1_4565(.VSS(VSS),.VDD(VDD),.Y(g34699),.A(I32855));
  NOT NOT1_4566(.VSS(VSS),.VDD(VDD),.Y(g19434),.A(g16326));
  NOT NOT1_4567(.VSS(VSS),.VDD(VDD),.Y(g16626),.A(g14133));
  NOT NOT1_4568(.VSS(VSS),.VDD(VDD),.Y(g8273),.A(g2453));
  NOT NOT1_4569(.VSS(VSS),.VDD(VDD),.Y(g10685),.A(I13995));
  NOT NOT1_4570(.VSS(VSS),.VDD(VDD),.Y(I16489),.A(g12793));
  NOT NOT1_4571(.VSS(VSS),.VDD(VDD),.Y(g16323),.A(I17653));
  NOT NOT1_4572(.VSS(VSS),.VDD(VDD),.Y(g24118),.A(g19890));
  NOT NOT1_4573(.VSS(VSS),.VDD(VDD),.Y(g10373),.A(g6917));
  NOT NOT1_4574(.VSS(VSS),.VDD(VDD),.Y(g14186),.A(g11346));
  NOT NOT1_4575(.VSS(VSS),.VDD(VDD),.Y(g14676),.A(I16775));
  NOT NOT1_4576(.VSS(VSS),.VDD(VDD),.Y(g24022),.A(g20982));
  NOT NOT1_4577(.VSS(VSS),.VDD(VDD),.Y(g34698),.A(g34550));
  NOT NOT1_4578(.VSS(VSS),.VDD(VDD),.Y(g7293),.A(g4452));
  NOT NOT1_4579(.VSS(VSS),.VDD(VDD),.Y(g12906),.A(g10413));
  NOT NOT1_4580(.VSS(VSS),.VDD(VDD),.Y(g16533),.A(I17733));
  NOT NOT1_4581(.VSS(VSS),.VDD(VDD),.Y(g20616),.A(g15277));
  NOT NOT1_4582(.VSS(VSS),.VDD(VDD),.Y(I18114),.A(g14509));
  NOT NOT1_4583(.VSS(VSS),.VDD(VDD),.Y(g23876),.A(g19074));
  NOT NOT1_4584(.VSS(VSS),.VDD(VDD),.Y(I18758),.A(g6719));
  NOT NOT1_4585(.VSS(VSS),.VDD(VDD),.Y(g13023),.A(g11897));
  NOT NOT1_4586(.VSS(VSS),.VDD(VDD),.Y(g18874),.A(g15938));
  NOT NOT1_4587(.VSS(VSS),.VDD(VDD),.Y(I31528),.A(g33219));
  NOT NOT1_4588(.VSS(VSS),.VDD(VDD),.Y(g25044),.A(g23675));
  NOT NOT1_4589(.VSS(VSS),.VDD(VDD),.Y(I19661),.A(g17587));
  NOT NOT1_4590(.VSS(VSS),.VDD(VDD),.Y(g29929),.A(g28914));
  NOT NOT1_4591(.VSS(VSS),.VDD(VDD),.Y(g16775),.A(I17999));
  NOT NOT1_4592(.VSS(VSS),.VDD(VDD),.Y(I18107),.A(g4019));
  NOT NOT1_4593(.VSS(VSS),.VDD(VDD),.Y(g10417),.A(g7117));
  NOT NOT1_4594(.VSS(VSS),.VDD(VDD),.Y(I25511),.A(g25073));
  NOT NOT1_4595(.VSS(VSS),.VDD(VDD),.Y(g32602),.A(g30825));
  NOT NOT1_4596(.VSS(VSS),.VDD(VDD),.Y(g32810),.A(g31376));
  NOT NOT1_4597(.VSS(VSS),.VDD(VDD),.Y(I13637),.A(g102));
  NOT NOT1_4598(.VSS(VSS),.VDD(VDD),.Y(I20882),.A(g17619));
  NOT NOT1_4599(.VSS(VSS),.VDD(VDD),.Y(g32657),.A(g31528));
  NOT NOT1_4600(.VSS(VSS),.VDD(VDD),.Y(g32774),.A(g30735));
  NOT NOT1_4601(.VSS(VSS),.VDD(VDD),.Y(g33778),.A(I31625));
  NOT NOT1_4602(.VSS(VSS),.VDD(VDD),.Y(g7828),.A(g4871));
  NOT NOT1_4603(.VSS(VSS),.VDD(VDD),.Y(g32955),.A(g30735));
  NOT NOT1_4604(.VSS(VSS),.VDD(VDD),.Y(g21511),.A(g15483));
  NOT NOT1_4605(.VSS(VSS),.VDD(VDD),.Y(g29928),.A(g28871));
  NOT NOT1_4606(.VSS(VSS),.VDD(VDD),.Y(I26670),.A(g27709));
  NOT NOT1_4607(.VSS(VSS),.VDD(VDD),.Y(g20704),.A(g15373));
  NOT NOT1_4608(.VSS(VSS),.VDD(VDD),.Y(g23511),.A(I22640));
  NOT NOT1_4609(.VSS(VSS),.VDD(VDD),.Y(g34427),.A(I32452));
  NOT NOT1_4610(.VSS(VSS),.VDD(VDD),.Y(I32119),.A(g33648));
  NOT NOT1_4611(.VSS(VSS),.VDD(VDD),.Y(g32879),.A(g31327));
  NOT NOT1_4612(.VSS(VSS),.VDD(VDD),.Y(g8572),.A(I12654));
  NOT NOT1_4613(.VSS(VSS),.VDD(VDD),.Y(g20053),.A(g17328));
  NOT NOT1_4614(.VSS(VSS),.VDD(VDD),.Y(g32970),.A(g30825));
  NOT NOT1_4615(.VSS(VSS),.VDD(VDD),.Y(g10334),.A(g4420));
  NOT NOT1_4616(.VSS(VSS),.VDD(VDD),.Y(g19682),.A(g17015));
  NOT NOT1_4617(.VSS(VSS),.VDD(VDD),.Y(I14537),.A(g10106));
  NOT NOT1_4618(.VSS(VSS),.VDD(VDD),.Y(g24053),.A(g21256));
  NOT NOT1_4619(.VSS(VSS),.VDD(VDD),.Y(g25120),.A(g22432));
  NOT NOT1_4620(.VSS(VSS),.VDD(VDD),.Y(I17780),.A(g13303));
  NOT NOT1_4621(.VSS(VSS),.VDD(VDD),.Y(g17523),.A(g14732));
  NOT NOT1_4622(.VSS(VSS),.VDD(VDD),.Y(g20900),.A(I20864));
  NOT NOT1_4623(.VSS(VSS),.VDD(VDD),.Y(g8712),.A(I12712));
  NOT NOT1_4624(.VSS(VSS),.VDD(VDD),.Y(g7592),.A(g347));
  NOT NOT1_4625(.VSS(VSS),.VDD(VDD),.Y(I16544),.A(g11931));
  NOT NOT1_4626(.VSS(VSS),.VDD(VDD),.Y(I18849),.A(g14290));
  NOT NOT1_4627(.VSS(VSS),.VDD(VDD),.Y(g18008),.A(I18868));
  NOT NOT1_4628(.VSS(VSS),.VDD(VDD),.Y(g32878),.A(g30937));
  NOT NOT1_4629(.VSS(VSS),.VDD(VDD),.Y(g31945),.A(g31189));
  NOT NOT1_4630(.VSS(VSS),.VDD(VDD),.Y(g21660),.A(g17694));
  NOT NOT1_4631(.VSS(VSS),.VDD(VDD),.Y(g24466),.A(I23671));
  NOT NOT1_4632(.VSS(VSS),.VDD(VDD),.Y(I16713),.A(g5331));
  NOT NOT1_4633(.VSS(VSS),.VDD(VDD),.Y(g9689),.A(g124));
  NOT NOT1_4634(.VSS(VSS),.VDD(VDD),.Y(g10762),.A(g8470));
  NOT NOT1_4635(.VSS(VSS),.VDD(VDD),.Y(g25562),.A(g22763));
  NOT NOT1_4636(.VSS(VSS),.VDD(VDD),.Y(g18892),.A(g15680));
  NOT NOT1_4637(.VSS(VSS),.VDD(VDD),.Y(g20036),.A(g17433));
  NOT NOT1_4638(.VSS(VSS),.VDD(VDD),.Y(g31826),.A(g29385));
  NOT NOT1_4639(.VSS(VSS),.VDD(VDD),.Y(g32886),.A(g31327));
  NOT NOT1_4640(.VSS(VSS),.VDD(VDD),.Y(I33161),.A(g34894));
  NOT NOT1_4641(.VSS(VSS),.VDD(VDD),.Y(I18398),.A(g13745));
  NOT NOT1_4642(.VSS(VSS),.VDD(VDD),.Y(g20101),.A(g17533));
  NOT NOT1_4643(.VSS(VSS),.VDD(VDD),.Y(g24036),.A(g20982));
  NOT NOT1_4644(.VSS(VSS),.VDD(VDD),.Y(I12541),.A(g194));
  NOT NOT1_4645(.VSS(VSS),.VDD(VDD),.Y(g20560),.A(g17328));
  NOT NOT1_4646(.VSS(VSS),.VDD(VDD),.Y(g16856),.A(I18048));
  NOT NOT1_4647(.VSS(VSS),.VDD(VDD),.Y(g21456),.A(g15509));
  NOT NOT1_4648(.VSS(VSS),.VDD(VDD),.Y(I26667),.A(g27585));
  NOT NOT1_4649(.VSS(VSS),.VDD(VDD),.Y(g11985),.A(I14827));
  NOT NOT1_4650(.VSS(VSS),.VDD(VDD),.Y(g17475),.A(I18398));
  NOT NOT1_4651(.VSS(VSS),.VDD(VDD),.Y(g24101),.A(g20998));
  NOT NOT1_4652(.VSS(VSS),.VDD(VDD),.Y(I23684),.A(g23230));
  NOT NOT1_4653(.VSS(VSS),.VDD(VDD),.Y(g32792),.A(g31710));
  NOT NOT1_4654(.VSS(VSS),.VDD(VDD),.Y(g23456),.A(g21514));
  NOT NOT1_4655(.VSS(VSS),.VDD(VDD),.Y(g13976),.A(g11130));
  NOT NOT1_4656(.VSS(VSS),.VDD(VDD),.Y(g24177),.A(I23375));
  NOT NOT1_4657(.VSS(VSS),.VDD(VDD),.Y(g24560),.A(g22942));
  NOT NOT1_4658(.VSS(VSS),.VDD(VDD),.Y(I15954),.A(g12381));
  NOT NOT1_4659(.VSS(VSS),.VDD(VDD),.Y(g32967),.A(g31327));
  NOT NOT1_4660(.VSS(VSS),.VDD(VDD),.Y(g10216),.A(I13684));
  NOT NOT1_4661(.VSS(VSS),.VDD(VDD),.Y(g14423),.A(I16579));
  NOT NOT1_4662(.VSS(VSS),.VDD(VDD),.Y(g8534),.A(g3338));
  NOT NOT1_4663(.VSS(VSS),.VDD(VDD),.Y(I16610),.A(g10981));
  NOT NOT1_4664(.VSS(VSS),.VDD(VDD),.Y(g9671),.A(g5134));
  NOT NOT1_4665(.VSS(VSS),.VDD(VDD),.Y(g20642),.A(g15277));
  NOT NOT1_4666(.VSS(VSS),.VDD(VDD),.Y(g23480),.A(I22601));
  NOT NOT1_4667(.VSS(VSS),.VDD(VDD),.Y(g27415),.A(g26382));
  NOT NOT1_4668(.VSS(VSS),.VDD(VDD),.Y(I20584),.A(g16587));
  NOT NOT1_4669(.VSS(VSS),.VDD(VDD),.Y(g23916),.A(g19277));
  NOT NOT1_4670(.VSS(VSS),.VDD(VDD),.Y(g9030),.A(g4793));
  NOT NOT1_4671(.VSS(VSS),.VDD(VDD),.Y(g19760),.A(g17015));
  NOT NOT1_4672(.VSS(VSS),.VDD(VDD),.Y(I32305),.A(g34209));
  NOT NOT1_4673(.VSS(VSS),.VDD(VDD),.Y(I14381),.A(g8300));
  NOT NOT1_4674(.VSS(VSS),.VDD(VDD),.Y(g16512),.A(g14015));
  NOT NOT1_4675(.VSS(VSS),.VDD(VDD),.Y(I16679),.A(g12039));
  NOT NOT1_4676(.VSS(VSS),.VDD(VDD),.Y(g23550),.A(g20248));
  NOT NOT1_4677(.VSS(VSS),.VDD(VDD),.Y(g26784),.A(g25341));
  NOT NOT1_4678(.VSS(VSS),.VDD(VDD),.Y(g9247),.A(g1559));
  NOT NOT1_4679(.VSS(VSS),.VDD(VDD),.Y(I33258),.A(g34976));
  NOT NOT1_4680(.VSS(VSS),.VDD(VDD),.Y(I32809),.A(g34586));
  NOT NOT1_4681(.VSS(VSS),.VDD(VDD),.Y(g18907),.A(g15979));
  NOT NOT1_4682(.VSS(VSS),.VDD(VDD),.Y(g7624),.A(I12106));
  NOT NOT1_4683(.VSS(VSS),.VDD(VDD),.Y(g32459),.A(g31070));
  NOT NOT1_4684(.VSS(VSS),.VDD(VDD),.Y(g20064),.A(g17533));
  NOT NOT1_4685(.VSS(VSS),.VDD(VDD),.Y(g7953),.A(g4966));
  NOT NOT1_4686(.VSS(VSS),.VDD(VDD),.Y(g30572),.A(g29945));
  NOT NOT1_4687(.VSS(VSS),.VDD(VDD),.Y(g24064),.A(g20841));
  NOT NOT1_4688(.VSS(VSS),.VDD(VDD),.Y(g28579),.A(g27714));
  NOT NOT1_4689(.VSS(VSS),.VDD(VDD),.Y(g9564),.A(g6120));
  NOT NOT1_4690(.VSS(VSS),.VDD(VDD),.Y(I18135),.A(g13144));
  NOT NOT1_4691(.VSS(VSS),.VDD(VDD),.Y(g23307),.A(g20924));
  NOT NOT1_4692(.VSS(VSS),.VDD(VDD),.Y(g32919),.A(g30735));
  NOT NOT1_4693(.VSS(VSS),.VDD(VDD),.Y(g23085),.A(g19957));
  NOT NOT1_4694(.VSS(VSS),.VDD(VDD),.Y(g32458),.A(g30825));
  NOT NOT1_4695(.VSS(VSS),.VDD(VDD),.Y(I24759),.A(g24229));
  NOT NOT1_4696(.VSS(VSS),.VDD(VDD),.Y(g14543),.A(I16660));
  NOT NOT1_4697(.VSS(VSS),.VDD(VDD),.Y(g33932),.A(I31810));
  NOT NOT1_4698(.VSS(VSS),.VDD(VDD),.Y(g9826),.A(g1844));
  NOT NOT1_4699(.VSS(VSS),.VDD(VDD),.Y(g10117),.A(g2509));
  NOT NOT1_4700(.VSS(VSS),.VDD(VDD),.Y(g10000),.A(g6151));
  NOT NOT1_4701(.VSS(VSS),.VDD(VDD),.Y(g26824),.A(g25298));
  NOT NOT1_4702(.VSS(VSS),.VDD(VDD),.Y(I16460),.A(g10430));
  NOT NOT1_4703(.VSS(VSS),.VDD(VDD),.Y(g20874),.A(g15680));
  NOT NOT1_4704(.VSS(VSS),.VDD(VDD),.Y(g21054),.A(g15373));
  NOT NOT1_4705(.VSS(VSS),.VDD(VDD),.Y(g32918),.A(g31327));
  NOT NOT1_4706(.VSS(VSS),.VDD(VDD),.Y(g23243),.A(g21070));
  NOT NOT1_4707(.VSS(VSS),.VDD(VDD),.Y(g20630),.A(g17955));
  NOT NOT1_4708(.VSS(VSS),.VDD(VDD),.Y(g11842),.A(I14660));
  NOT NOT1_4709(.VSS(VSS),.VDD(VDD),.Y(g21431),.A(g18065));
  NOT NOT1_4710(.VSS(VSS),.VDD(VDD),.Y(g9741),.A(I13317));
  NOT NOT1_4711(.VSS(VSS),.VDD(VDD),.Y(g8903),.A(g1075));
  NOT NOT1_4712(.VSS(VSS),.VDD(VDD),.Y(g23431),.A(g21514));
  NOT NOT1_4713(.VSS(VSS),.VDD(VDD),.Y(I13906),.A(g7620));
  NOT NOT1_4714(.VSS(VSS),.VDD(VDD),.Y(g32545),.A(g31070));
  NOT NOT1_4715(.VSS(VSS),.VDD(VDD),.Y(g9910),.A(g2108));
  NOT NOT1_4716(.VSS(VSS),.VDD(VDD),.Y(g17600),.A(g14659));
  NOT NOT1_4717(.VSS(VSS),.VDD(VDD),.Y(I19671),.A(g15932));
  NOT NOT1_4718(.VSS(VSS),.VDD(VDD),.Y(g34490),.A(I32547));
  NOT NOT1_4719(.VSS(VSS),.VDD(VDD),.Y(g20166),.A(g16886));
  NOT NOT1_4720(.VSS(VSS),.VDD(VDD),.Y(g20009),.A(g16349));
  NOT NOT1_4721(.VSS(VSS),.VDD(VDD),.Y(I22583),.A(g20998));
  NOT NOT1_4722(.VSS(VSS),.VDD(VDD),.Y(g27576),.A(g26081));
  NOT NOT1_4723(.VSS(VSS),.VDD(VDD),.Y(g27585),.A(g25994));
  NOT NOT1_4724(.VSS(VSS),.VDD(VDD),.Y(g20665),.A(g15373));
  NOT NOT1_4725(.VSS(VSS),.VDD(VDD),.Y(g25547),.A(g22550));
  NOT NOT1_4726(.VSS(VSS),.VDD(VDD),.Y(g32599),.A(g30673));
  NOT NOT1_4727(.VSS(VSS),.VDD(VDD),.Y(I20744),.A(g17141));
  NOT NOT1_4728(.VSS(VSS),.VDD(VDD),.Y(I31810),.A(g33164));
  NOT NOT1_4729(.VSS(VSS),.VDD(VDD),.Y(g9638),.A(g1620));
  NOT NOT1_4730(.VSS(VSS),.VDD(VDD),.Y(g21269),.A(g15506));
  NOT NOT1_4731(.VSS(VSS),.VDD(VDD),.Y(g24166),.A(I23342));
  NOT NOT1_4732(.VSS(VSS),.VDD(VDD),.Y(g24665),.A(g23067));
  NOT NOT1_4733(.VSS(VSS),.VDD(VDD),.Y(g7716),.A(g1199));
  NOT NOT1_4734(.VSS(VSS),.VDD(VDD),.Y(g7149),.A(g4564));
  NOT NOT1_4735(.VSS(VSS),.VDD(VDD),.Y(g34784),.A(I32982));
  NOT NOT1_4736(.VSS(VSS),.VDD(VDD),.Y(g7349),.A(g1270));
  NOT NOT1_4737(.VSS(VSS),.VDD(VDD),.Y(g30297),.A(g28758));
  NOT NOT1_4738(.VSS(VSS),.VDD(VDD),.Y(g27554),.A(g26625));
  NOT NOT1_4739(.VSS(VSS),.VDD(VDD),.Y(g20008),.A(g16449));
  NOT NOT1_4740(.VSS(VSS),.VDD(VDD),.Y(g34956),.A(I33214));
  NOT NOT1_4741(.VSS(VSS),.VDD(VDD),.Y(g17952),.A(I18858));
  NOT NOT1_4742(.VSS(VSS),.VDD(VDD),.Y(g32598),.A(g30614));
  NOT NOT1_4743(.VSS(VSS),.VDD(VDD),.Y(g13016),.A(g11878));
  NOT NOT1_4744(.VSS(VSS),.VDD(VDD),.Y(I22046),.A(g19330));
  NOT NOT1_4745(.VSS(VSS),.VDD(VDD),.Y(g23942),.A(g21562));
  NOT NOT1_4746(.VSS(VSS),.VDD(VDD),.Y(I20399),.A(g16205));
  NOT NOT1_4747(.VSS(VSS),.VDD(VDD),.Y(g23341),.A(g21163));
  NOT NOT1_4748(.VSS(VSS),.VDD(VDD),.Y(g18092),.A(I18882));
  NOT NOT1_4749(.VSS(VSS),.VDD(VDD),.Y(g21268),.A(g15680));
  NOT NOT1_4750(.VSS(VSS),.VDD(VDD),.Y(I14192),.A(g10233));
  NOT NOT1_4751(.VSS(VSS),.VDD(VDD),.Y(I18048),.A(g13638));
  NOT NOT1_4752(.VSS(VSS),.VDD(VDD),.Y(I28062),.A(g29194));
  NOT NOT1_4753(.VSS(VSS),.VDD(VDD),.Y(g25226),.A(g22763));
  NOT NOT1_4754(.VSS(VSS),.VDD(VDD),.Y(g22137),.A(g21370));
  NOT NOT1_4755(.VSS(VSS),.VDD(VDD),.Y(g21156),.A(g17247));
  NOT NOT1_4756(.VSS(VSS),.VDD(VDD),.Y(g17821),.A(I18829));
  NOT NOT1_4757(.VSS(VSS),.VDD(VDD),.Y(g8178),.A(I12437));
  NOT NOT1_4758(.VSS(VSS),.VDD(VDD),.Y(g6801),.A(g391));
  NOT NOT1_4759(.VSS(VSS),.VDD(VDD),.Y(I21006),.A(g15579));
  NOT NOT1_4760(.VSS(VSS),.VDD(VDD),.Y(g28615),.A(g27817));
  NOT NOT1_4761(.VSS(VSS),.VDD(VDD),.Y(I16875),.A(g6675));
  NOT NOT1_4762(.VSS(VSS),.VDD(VDD),.Y(g25481),.A(g22228));
  NOT NOT1_4763(.VSS(VSS),.VDD(VDD),.Y(I15893),.A(g10430));
  NOT NOT1_4764(.VSS(VSS),.VDD(VDD),.Y(I31878),.A(g33696));
  NOT NOT1_4765(.VSS(VSS),.VDD(VDD),.Y(g19649),.A(g17015));
  NOT NOT1_4766(.VSS(VSS),.VDD(VDD),.Y(I32874),.A(g34504));
  NOT NOT1_4767(.VSS(VSS),.VDD(VDD),.Y(g21180),.A(g18008));
  NOT NOT1_4768(.VSS(VSS),.VDD(VDD),.Y(I14663),.A(g9747));
  NOT NOT1_4769(.VSS(VSS),.VDD(VDD),.Y(g21670),.A(g16540));
  NOT NOT1_4770(.VSS(VSS),.VDD(VDD),.Y(I18221),.A(g13605));
  NOT NOT1_4771(.VSS(VSS),.VDD(VDD),.Y(g16722),.A(I17938));
  NOT NOT1_4772(.VSS(VSS),.VDD(VDD),.Y(g16924),.A(I18092));
  NOT NOT1_4773(.VSS(VSS),.VDD(VDD),.Y(g20555),.A(g15480));
  NOT NOT1_4774(.VSS(VSS),.VDD(VDD),.Y(g32817),.A(g31376));
  NOT NOT1_4775(.VSS(VSS),.VDD(VDD),.Y(I28851),.A(g29317));
  NOT NOT1_4776(.VSS(VSS),.VDD(VDD),.Y(I28872),.A(g30072));
  NOT NOT1_4777(.VSS(VSS),.VDD(VDD),.Y(I32693),.A(g34433));
  NOT NOT1_4778(.VSS(VSS),.VDD(VDD),.Y(g8135),.A(I12418));
  NOT NOT1_4779(.VSS(VSS),.VDD(VDD),.Y(I21222),.A(g18091));
  NOT NOT1_4780(.VSS(VSS),.VDD(VDD),.Y(g19491),.A(g16349));
  NOT NOT1_4781(.VSS(VSS),.VDD(VDD),.Y(g34181),.A(g33913));
  NOT NOT1_4782(.VSS(VSS),.VDD(VDD),.Y(g34671),.A(I32797));
  NOT NOT1_4783(.VSS(VSS),.VDD(VDD),.Y(g20570),.A(g15277));
  NOT NOT1_4784(.VSS(VSS),.VDD(VDD),.Y(g20712),.A(g15509));
  NOT NOT1_4785(.VSS(VSS),.VDD(VDD),.Y(g11865),.A(g10124));
  NOT NOT1_4786(.VSS(VSS),.VDD(VDD),.Y(I22302),.A(g19353));
  NOT NOT1_4787(.VSS(VSS),.VDD(VDD),.Y(g13865),.A(I16168));
  NOT NOT1_4788(.VSS(VSS),.VDD(VDD),.Y(g20914),.A(g15373));
  NOT NOT1_4789(.VSS(VSS),.VDD(VDD),.Y(g21335),.A(I21067));
  NOT NOT1_4790(.VSS(VSS),.VDD(VDD),.Y(g18883),.A(g15938));
  NOT NOT1_4791(.VSS(VSS),.VDD(VDD),.Y(g32532),.A(g31170));
  NOT NOT1_4792(.VSS(VSS),.VDD(VDD),.Y(g32901),.A(g31327));
  NOT NOT1_4793(.VSS(VSS),.VDD(VDD),.Y(g14639),.A(I16747));
  NOT NOT1_4794(.VSS(VSS),.VDD(VDD),.Y(g10230),.A(I13694));
  NOT NOT1_4795(.VSS(VSS),.VDD(VDD),.Y(g23335),.A(g20391));
  NOT NOT1_4796(.VSS(VSS),.VDD(VDD),.Y(I32665),.A(g34386));
  NOT NOT1_4797(.VSS(VSS),.VDD(VDD),.Y(g19755),.A(g15915));
  NOT NOT1_4798(.VSS(VSS),.VDD(VDD),.Y(g6755),.A(I11620));
  NOT NOT1_4799(.VSS(VSS),.VDD(VDD),.Y(g12921),.A(g12228));
  NOT NOT1_4800(.VSS(VSS),.VDD(VDD),.Y(g23839),.A(g18997));
  NOT NOT1_4801(.VSS(VSS),.VDD(VDD),.Y(I17787),.A(g3267));
  NOT NOT1_4802(.VSS(VSS),.VDD(VDD),.Y(g17873),.A(I18849));
  NOT NOT1_4803(.VSS(VSS),.VDD(VDD),.Y(g23930),.A(g19147));
  NOT NOT1_4804(.VSS(VSS),.VDD(VDD),.Y(g23993),.A(g19277));
  NOT NOT1_4805(.VSS(VSS),.VDD(VDD),.Y(g32783),.A(g30825));
  NOT NOT1_4806(.VSS(VSS),.VDD(VDD),.Y(g19770),.A(g17062));
  NOT NOT1_4807(.VSS(VSS),.VDD(VDD),.Y(I29199),.A(g30237));
  NOT NOT1_4808(.VSS(VSS),.VDD(VDD),.Y(g30931),.A(I28913));
  NOT NOT1_4809(.VSS(VSS),.VDD(VDD),.Y(g8805),.A(I12799));
  NOT NOT1_4810(.VSS(VSS),.VDD(VDD),.Y(I14862),.A(g8092));
  NOT NOT1_4811(.VSS(VSS),.VDD(VDD),.Y(g8916),.A(I12887));
  NOT NOT1_4812(.VSS(VSS),.VDD(VDD),.Y(I16160),.A(g11237));
  NOT NOT1_4813(.VSS(VSS),.VDD(VDD),.Y(g21694),.A(g16540));
  NOT NOT1_4814(.VSS(VSS),.VDD(VDD),.Y(g23838),.A(g18997));
  NOT NOT1_4815(.VSS(VSS),.VDD(VDD),.Y(g9861),.A(g5459));
  NOT NOT1_4816(.VSS(VSS),.VDD(VDD),.Y(g10416),.A(g10318));
  NOT NOT1_4817(.VSS(VSS),.VDD(VDD),.Y(I15705),.A(g12218));
  NOT NOT1_4818(.VSS(VSS),.VDD(VDD),.Y(g9048),.A(I12963));
  NOT NOT1_4819(.VSS(VSS),.VDD(VDD),.Y(I17302),.A(g14044));
  NOT NOT1_4820(.VSS(VSS),.VDD(VDD),.Y(g32561),.A(g30614));
  NOT NOT1_4821(.VSS(VSS),.VDD(VDD),.Y(g32656),.A(g30673));
  NOT NOT1_4822(.VSS(VSS),.VDD(VDD),.Y(g23965),.A(g21611));
  NOT NOT1_4823(.VSS(VSS),.VDD(VDD),.Y(I31459),.A(g33219));
  NOT NOT1_4824(.VSS(VSS),.VDD(VDD),.Y(g20239),.A(g17128));
  NOT NOT1_4825(.VSS(VSS),.VDD(VDD),.Y(I32476),.A(g34277));
  NOT NOT1_4826(.VSS(VSS),.VDD(VDD),.Y(g11705),.A(I14576));
  NOT NOT1_4827(.VSS(VSS),.VDD(VDD),.Y(I22640),.A(g21256));
  NOT NOT1_4828(.VSS(VSS),.VDD(VDD),.Y(g24074),.A(g21193));
  NOT NOT1_4829(.VSS(VSS),.VDD(VDD),.Y(I22769),.A(g21277));
  NOT NOT1_4830(.VSS(VSS),.VDD(VDD),.Y(g26860),.A(I25594));
  NOT NOT1_4831(.VSS(VSS),.VDD(VDD),.Y(I14326),.A(g8607));
  NOT NOT1_4832(.VSS(VSS),.VDD(VDD),.Y(g34426),.A(I32449));
  NOT NOT1_4833(.VSS(VSS),.VDD(VDD),.Y(g11042),.A(g8691));
  NOT NOT1_4834(.VSS(VSS),.VDD(VDD),.Y(g16031),.A(I17436));
  NOT NOT1_4835(.VSS(VSS),.VDD(VDD),.Y(g20567),.A(g15426));
  NOT NOT1_4836(.VSS(VSS),.VDD(VDD),.Y(g20594),.A(g15277));
  NOT NOT1_4837(.VSS(VSS),.VDD(VDD),.Y(g32680),.A(g31376));
  NOT NOT1_4838(.VSS(VSS),.VDD(VDD),.Y(g10391),.A(g6988));
  NOT NOT1_4839(.VSS(VSS),.VDD(VDD),.Y(I16455),.A(g11845));
  NOT NOT1_4840(.VSS(VSS),.VDD(VDD),.Y(g32823),.A(g31327));
  NOT NOT1_4841(.VSS(VSS),.VDD(VDD),.Y(g20238),.A(g17096));
  NOT NOT1_4842(.VSS(VSS),.VDD(VDD),.Y(g25297),.A(g23746));
  NOT NOT1_4843(.VSS(VSS),.VDD(VDD),.Y(g13255),.A(g10632));
  NOT NOT1_4844(.VSS(VSS),.VDD(VDD),.Y(g9827),.A(g1974));
  NOT NOT1_4845(.VSS(VSS),.VDD(VDD),.Y(g13189),.A(g10762));
  NOT NOT1_4846(.VSS(VSS),.VDD(VDD),.Y(g22542),.A(g19801));
  NOT NOT1_4847(.VSS(VSS),.VDD(VDD),.Y(g13679),.A(g10573));
  NOT NOT1_4848(.VSS(VSS),.VDD(VDD),.Y(g28142),.A(I26649));
  NOT NOT1_4849(.VSS(VSS),.VDD(VDD),.Y(g31811),.A(g29385));
  NOT NOT1_4850(.VSS(VSS),.VDD(VDD),.Y(g23487),.A(g20924));
  NOT NOT1_4851(.VSS(VSS),.VDD(VDD),.Y(g14510),.A(I16629));
  NOT NOT1_4852(.VSS(VSS),.VDD(VDD),.Y(g31646),.A(I29228));
  NOT NOT1_4853(.VSS(VSS),.VDD(VDD),.Y(g9333),.A(g417));
  NOT NOT1_4854(.VSS(VSS),.VDD(VDD),.Y(I14702),.A(g7717));
  NOT NOT1_4855(.VSS(VSS),.VDD(VDD),.Y(g19794),.A(g16489));
  NOT NOT1_4856(.VSS(VSS),.VDD(VDD),.Y(g11678),.A(I14563));
  NOT NOT1_4857(.VSS(VSS),.VDD(VDD),.Y(g12184),.A(I15036));
  NOT NOT1_4858(.VSS(VSS),.VDD(VDD),.Y(g16529),.A(g14055));
  NOT NOT1_4859(.VSS(VSS),.VDD(VDD),.Y(g29081),.A(g27837));
  NOT NOT1_4860(.VSS(VSS),.VDD(VDD),.Y(g12805),.A(g9511));
  NOT NOT1_4861(.VSS(VSS),.VDD(VDD),.Y(g13188),.A(g10909));
  NOT NOT1_4862(.VSS(VSS),.VDD(VDD),.Y(g19395),.A(g16431));
  NOT NOT1_4863(.VSS(VSS),.VDD(VDD),.Y(g23502),.A(g21070));
  NOT NOT1_4864(.VSS(VSS),.VDD(VDD),.Y(I27927),.A(g28803));
  NOT NOT1_4865(.VSS(VSS),.VDD(VDD),.Y(g20382),.A(g15171));
  NOT NOT1_4866(.VSS(VSS),.VDD(VDD),.Y(I16201),.A(g4023));
  NOT NOT1_4867(.VSS(VSS),.VDD(VDD),.Y(I23351),.A(g23263));
  NOT NOT1_4868(.VSS(VSS),.VDD(VDD),.Y(I31545),.A(g33219));
  NOT NOT1_4869(.VSS(VSS),.VDD(VDD),.Y(I23372),.A(g23361));
  NOT NOT1_4870(.VSS(VSS),.VDD(VDD),.Y(g26700),.A(g25429));
  NOT NOT1_4871(.VSS(VSS),.VDD(VDD),.Y(g7258),.A(g4414));
  NOT NOT1_4872(.VSS(VSS),.VDD(VDD),.Y(I33079),.A(g34809));
  NOT NOT1_4873(.VSS(VSS),.VDD(VDD),.Y(g11686),.A(I14567));
  NOT NOT1_4874(.VSS(VSS),.VDD(VDD),.Y(g16528),.A(g14154));
  NOT NOT1_4875(.VSS(VSS),.VDD(VDD),.Y(g7577),.A(g1263));
  NOT NOT1_4876(.VSS(VSS),.VDD(VDD),.Y(g7867),.A(g1489));
  NOT NOT1_4877(.VSS(VSS),.VDD(VDD),.Y(g13460),.A(I15942));
  NOT NOT1_4878(.VSS(VSS),.VDD(VDD),.Y(g15831),.A(g13385));
  NOT NOT1_4879(.VSS(VSS),.VDD(VDD),.Y(I26479),.A(g25771));
  NOT NOT1_4880(.VSS(VSS),.VDD(VDD),.Y(I12927),.A(g4332));
  NOT NOT1_4881(.VSS(VSS),.VDD(VDD),.Y(g26987),.A(g26131));
  NOT NOT1_4882(.VSS(VSS),.VDD(VDD),.Y(g11383),.A(g9061));
  NOT NOT1_4883(.VSS(VSS),.VDD(VDD),.Y(g10014),.A(g6439));
  NOT NOT1_4884(.VSS(VSS),.VDD(VDD),.Y(g23443),.A(g21468));
  NOT NOT1_4885(.VSS(VSS),.VDD(VDD),.Y(I15030),.A(g10073));
  NOT NOT1_4886(.VSS(VSS),.VDD(VDD),.Y(I18795),.A(g5327));
  NOT NOT1_4887(.VSS(VSS),.VDD(VDD),.Y(g21279),.A(g15680));
  NOT NOT1_4888(.VSS(VSS),.VDD(VDD),.Y(g24176),.A(I23372));
  NOT NOT1_4889(.VSS(VSS),.VDD(VDD),.Y(g24185),.A(I23399));
  NOT NOT1_4890(.VSS(VSS),.VDD(VDD),.Y(g23279),.A(g21037));
  NOT NOT1_4891(.VSS(VSS),.VDD(VDD),.Y(g32966),.A(g31021));
  NOT NOT1_4892(.VSS(VSS),.VDD(VDD),.Y(g19633),.A(g16931));
  NOT NOT1_4893(.VSS(VSS),.VDD(VDD),.Y(g7717),.A(I12172));
  NOT NOT1_4894(.VSS(VSS),.VDD(VDD),.Y(g30088),.A(g29094));
  NOT NOT1_4895(.VSS(VSS),.VDD(VDD),.Y(g24092),.A(g20857));
  NOT NOT1_4896(.VSS(VSS),.VDD(VDD),.Y(I32074),.A(g33670));
  NOT NOT1_4897(.VSS(VSS),.VDD(VDD),.Y(g29945),.A(I28174));
  NOT NOT1_4898(.VSS(VSS),.VDD(VDD),.Y(g6868),.A(I11688));
  NOT NOT1_4899(.VSS(VSS),.VDD(VDD),.Y(g11030),.A(g8292));
  NOT NOT1_4900(.VSS(VSS),.VDD(VDD),.Y(g20154),.A(I20412));
  NOT NOT1_4901(.VSS(VSS),.VDD(VDD),.Y(g22905),.A(I22114));
  NOT NOT1_4902(.VSS(VSS),.VDD(VDD),.Y(g32631),.A(g30825));
  NOT NOT1_4903(.VSS(VSS),.VDD(VDD),.Y(g19719),.A(g16897));
  NOT NOT1_4904(.VSS(VSS),.VDD(VDD),.Y(g21278),.A(I21013));
  NOT NOT1_4905(.VSS(VSS),.VDD(VDD),.Y(g11294),.A(g7598));
  NOT NOT1_4906(.VSS(VSS),.VDD(VDD),.Y(g24154),.A(I23306));
  NOT NOT1_4907(.VSS(VSS),.VDD(VDD),.Y(I32594),.A(g34298));
  NOT NOT1_4908(.VSS(VSS),.VDD(VDD),.Y(g8037),.A(g405));
  NOT NOT1_4909(.VSS(VSS),.VDD(VDD),.Y(g23278),.A(g20283));
  NOT NOT1_4910(.VSS(VSS),.VDD(VDD),.Y(g13267),.A(I15831));
  NOT NOT1_4911(.VSS(VSS),.VDD(VDD),.Y(g29999),.A(g28973));
  NOT NOT1_4912(.VSS(VSS),.VDD(VDD),.Y(g32364),.A(I29894));
  NOT NOT1_4913(.VSS(VSS),.VDD(VDD),.Y(g6767),.A(I11626));
  NOT NOT1_4914(.VSS(VSS),.VDD(VDD),.Y(g17614),.A(I18571));
  NOT NOT1_4915(.VSS(VSS),.VDD(VDD),.Y(g22593),.A(g19801));
  NOT NOT1_4916(.VSS(VSS),.VDD(VDD),.Y(g9780),.A(I13360));
  NOT NOT1_4917(.VSS(VSS),.VDD(VDD),.Y(g16960),.A(I18114));
  NOT NOT1_4918(.VSS(VSS),.VDD(VDD),.Y(g20637),.A(g15224));
  NOT NOT1_4919(.VSS(VSS),.VDD(VDD),.Y(g26943),.A(I25695));
  NOT NOT1_4920(.VSS(VSS),.VDD(VDD),.Y(g8102),.A(g3072));
  NOT NOT1_4921(.VSS(VSS),.VDD(VDD),.Y(g13065),.A(g10476));
  NOT NOT1_4922(.VSS(VSS),.VDD(VDD),.Y(g19718),.A(g17015));
  NOT NOT1_4923(.VSS(VSS),.VDD(VDD),.Y(g21286),.A(g15509));
  NOT NOT1_4924(.VSS(VSS),.VDD(VDD),.Y(g8302),.A(g1926));
  NOT NOT1_4925(.VSS(VSS),.VDD(VDD),.Y(g14442),.A(I16593));
  NOT NOT1_4926(.VSS(VSS),.VDD(VDD),.Y(g29998),.A(g28966));
  NOT NOT1_4927(.VSS(VSS),.VDD(VDD),.Y(g17607),.A(I18560));
  NOT NOT1_4928(.VSS(VSS),.VDD(VDD),.Y(g21468),.A(I21181));
  NOT NOT1_4929(.VSS(VSS),.VDD(VDD),.Y(g17320),.A(I18297));
  NOT NOT1_4930(.VSS(VSS),.VDD(VDD),.Y(g21306),.A(g15582));
  NOT NOT1_4931(.VSS(VSS),.VDD(VDD),.Y(g31850),.A(g29385));
  NOT NOT1_4932(.VSS(VSS),.VDD(VDD),.Y(g8579),.A(g2771));
  NOT NOT1_4933(.VSS(VSS),.VDD(VDD),.Y(g23306),.A(g20924));
  NOT NOT1_4934(.VSS(VSS),.VDD(VDD),.Y(I29225),.A(g30311));
  NOT NOT1_4935(.VSS(VSS),.VDD(VDD),.Y(I31817),.A(g33323));
  NOT NOT1_4936(.VSS(VSS),.VDD(VDD),.Y(g7975),.A(g3040));
  NOT NOT1_4937(.VSS(VSS),.VDD(VDD),.Y(g33850),.A(I31701));
  NOT NOT1_4938(.VSS(VSS),.VDD(VDD),.Y(g17530),.A(g14947));
  NOT NOT1_4939(.VSS(VSS),.VDD(VDD),.Y(g10116),.A(g2413));
  NOT NOT1_4940(.VSS(VSS),.VDD(VDD),.Y(g9662),.A(g3983));
  NOT NOT1_4941(.VSS(VSS),.VDD(VDD),.Y(g9018),.A(g4273));
  NOT NOT1_4942(.VSS(VSS),.VDD(VDD),.Y(g11875),.A(I14687));
  NOT NOT1_4943(.VSS(VSS),.VDD(VDD),.Y(g8719),.A(I12719));
  NOT NOT1_4944(.VSS(VSS),.VDD(VDD),.Y(g27013),.A(I25743));
  NOT NOT1_4945(.VSS(VSS),.VDD(VDD),.Y(g7026),.A(g5507));
  NOT NOT1_4946(.VSS(VSS),.VDD(VDD),.Y(I32675),.A(g34427));
  NOT NOT1_4947(.VSS(VSS),.VDD(VDD),.Y(g9467),.A(g6434));
  NOT NOT1_4948(.VSS(VSS),.VDD(VDD),.Y(g19440),.A(g15915));
  NOT NOT1_4949(.VSS(VSS),.VDD(VDD),.Y(g16709),.A(I17919));
  NOT NOT1_4950(.VSS(VSS),.VDD(VDD),.Y(g17122),.A(g14348));
  NOT NOT1_4951(.VSS(VSS),.VDD(VDD),.Y(g34126),.A(I32067));
  NOT NOT1_4952(.VSS(VSS),.VDD(VDD),.Y(g34659),.A(I32775));
  NOT NOT1_4953(.VSS(VSS),.VDD(VDD),.Y(I12770),.A(g4200));
  NOT NOT1_4954(.VSS(VSS),.VDD(VDD),.Y(I12563),.A(g3798));
  NOT NOT1_4955(.VSS(VSS),.VDD(VDD),.Y(g12013),.A(I14866));
  NOT NOT1_4956(.VSS(VSS),.VDD(VDD),.Y(g23815),.A(g19074));
  NOT NOT1_4957(.VSS(VSS),.VDD(VDD),.Y(g34987),.A(I33261));
  NOT NOT1_4958(.VSS(VSS),.VDD(VDD),.Y(I25677),.A(g25640));
  NOT NOT1_4959(.VSS(VSS),.VDD(VDD),.Y(I15837),.A(g1459));
  NOT NOT1_4960(.VSS(VSS),.VDD(VDD),.Y(I33158),.A(g34897));
  NOT NOT1_4961(.VSS(VSS),.VDD(VDD),.Y(g7170),.A(g5719));
  NOT NOT1_4962(.VSS(VSS),.VDD(VDD),.Y(g19861),.A(g17096));
  NOT NOT1_4963(.VSS(VSS),.VDD(VDD),.Y(g10275),.A(g4584));
  NOT NOT1_4964(.VSS(VSS),.VDD(VDD),.Y(g19573),.A(g16877));
  NOT NOT1_4965(.VSS(VSS),.VDD(VDD),.Y(g8917),.A(I12890));
  NOT NOT1_4966(.VSS(VSS),.VDD(VDD),.Y(g16708),.A(I17916));
  NOT NOT1_4967(.VSS(VSS),.VDD(VDD),.Y(g22153),.A(g18997));
  NOT NOT1_4968(.VSS(VSS),.VDD(VDD),.Y(g21677),.A(I21238));
  NOT NOT1_4969(.VSS(VSS),.VDD(VDD),.Y(g33228),.A(I30766));
  NOT NOT1_4970(.VSS(VSS),.VDD(VDD),.Y(g10430),.A(I13847));
  NOT NOT1_4971(.VSS(VSS),.VDD(VDD),.Y(g14275),.A(g12358));
  NOT NOT1_4972(.VSS(VSS),.VDD(VDD),.Y(g25546),.A(g22550));
  NOT NOT1_4973(.VSS(VSS),.VDD(VDD),.Y(g32571),.A(g31376));
  NOT NOT1_4974(.VSS(VSS),.VDD(VDD),.Y(I31561),.A(g33197));
  NOT NOT1_4975(.VSS(VSS),.VDD(VDD),.Y(I17249),.A(g13605));
  NOT NOT1_4976(.VSS(VSS),.VDD(VDD),.Y(g25211),.A(g22763));
  NOT NOT1_4977(.VSS(VSS),.VDD(VDD),.Y(I32935),.A(g34657));
  NOT NOT1_4978(.VSS(VSS),.VDD(VDD),.Y(g22409),.A(I21860));
  NOT NOT1_4979(.VSS(VSS),.VDD(VDD),.Y(g19389),.A(g17532));
  NOT NOT1_4980(.VSS(VSS),.VDD(VDD),.Y(g17641),.A(g14845));
  NOT NOT1_4981(.VSS(VSS),.VDD(VDD),.Y(g20501),.A(g17955));
  NOT NOT1_4982(.VSS(VSS),.VDD(VDD),.Y(g26870),.A(I25606));
  NOT NOT1_4983(.VSS(VSS),.VDD(VDD),.Y(g30296),.A(g28889));
  NOT NOT1_4984(.VSS(VSS),.VDD(VDD),.Y(g20577),.A(g15483));
  NOT NOT1_4985(.VSS(VSS),.VDD(VDD),.Y(g34339),.A(g34077));
  NOT NOT1_4986(.VSS(VSS),.VDD(VDD),.Y(g9816),.A(g6167));
  NOT NOT1_4987(.VSS(VSS),.VDD(VDD),.Y(g34943),.A(I33197));
  NOT NOT1_4988(.VSS(VSS),.VDD(VDD),.Y(I20951),.A(g17782));
  NOT NOT1_4989(.VSS(VSS),.VDD(VDD),.Y(g25024),.A(g22472));
  NOT NOT1_4990(.VSS(VSS),.VDD(VDD),.Y(g33716),.A(I31569));
  NOT NOT1_4991(.VSS(VSS),.VDD(VDD),.Y(I31823),.A(g33149));
  NOT NOT1_4992(.VSS(VSS),.VDD(VDD),.Y(g19612),.A(g16897));
  NOT NOT1_4993(.VSS(VSS),.VDD(VDD),.Y(g34296),.A(I32297));
  NOT NOT1_4994(.VSS(VSS),.VDD(VDD),.Y(g7280),.A(g2153));
  NOT NOT1_4995(.VSS(VSS),.VDD(VDD),.Y(g29897),.A(I28128));
  NOT NOT1_4996(.VSS(VSS),.VDD(VDD),.Y(g7939),.A(g1280));
  NOT NOT1_4997(.VSS(VSS),.VDD(VDD),.Y(g22136),.A(g20277));
  NOT NOT1_4998(.VSS(VSS),.VDD(VDD),.Y(g29961),.A(g28892));
  NOT NOT1_4999(.VSS(VSS),.VDD(VDD),.Y(g8442),.A(g3476));
  NOT NOT1_5000(.VSS(VSS),.VDD(VDD),.Y(g22408),.A(g19483));
  NOT NOT1_5001(.VSS(VSS),.VDD(VDD),.Y(g22635),.A(g19801));
  NOT NOT1_5002(.VSS(VSS),.VDD(VDD),.Y(I12767),.A(g4197));
  NOT NOT1_5003(.VSS(VSS),.VDD(VDD),.Y(g14237),.A(g11666));
  NOT NOT1_5004(.VSS(VSS),.VDD(VDD),.Y(g8786),.A(I12770));
  NOT NOT1_5005(.VSS(VSS),.VDD(VDD),.Y(g23937),.A(g19277));
  NOT NOT1_5006(.VSS(VSS),.VDD(VDD),.Y(g10035),.A(g1720));
  NOT NOT1_5007(.VSS(VSS),.VDD(VDD),.Y(g32495),.A(g31070));
  NOT NOT1_5008(.VSS(VSS),.VDD(VDD),.Y(g29505),.A(g29186));
  NOT NOT1_5009(.VSS(VSS),.VDD(VDD),.Y(g19777),.A(g17015));
  NOT NOT1_5010(.VSS(VSS),.VDD(VDD),.Y(g17409),.A(I18344));
  NOT NOT1_5011(.VSS(VSS),.VDD(VDD),.Y(I12899),.A(g4232));
  NOT NOT1_5012(.VSS(VSS),.VDD(VDD),.Y(g7544),.A(g918));
  NOT NOT1_5013(.VSS(VSS),.VDD(VDD),.Y(g8164),.A(g3484));
  NOT NOT1_5014(.VSS(VSS),.VDD(VDD),.Y(g9381),.A(g5527));
  NOT NOT1_5015(.VSS(VSS),.VDD(VDD),.Y(I15617),.A(g12037));
  NOT NOT1_5016(.VSS(VSS),.VDD(VDD),.Y(I13805),.A(g6976));
  NOT NOT1_5017(.VSS(VSS),.VDD(VDD),.Y(I18788),.A(g13138));
  NOT NOT1_5018(.VSS(VSS),.VDD(VDD),.Y(g8364),.A(g1585));
  NOT NOT1_5019(.VSS(VSS),.VDD(VDD),.Y(g32816),.A(g31327));
  NOT NOT1_5020(.VSS(VSS),.VDD(VDD),.Y(I15915),.A(g10430));
  NOT NOT1_5021(.VSS(VSS),.VDD(VDD),.Y(g24438),.A(g22722));
  NOT NOT1_5022(.VSS(VSS),.VDD(VDD),.Y(g11470),.A(g7625));
  NOT NOT1_5023(.VSS(VSS),.VDD(VDD),.Y(g17136),.A(g14348));
  NOT NOT1_5024(.VSS(VSS),.VDD(VDD),.Y(g10142),.A(I13637));
  NOT NOT1_5025(.VSS(VSS),.VDD(VDD),.Y(g17408),.A(I18341));
  NOT NOT1_5026(.VSS(VSS),.VDD(VDD),.Y(g34060),.A(g33704));
  NOT NOT1_5027(.VSS(VSS),.VDD(VDD),.Y(g29212),.A(I27552));
  NOT NOT1_5028(.VSS(VSS),.VDD(VDD),.Y(g7636),.A(g4098));
  NOT NOT1_5029(.VSS(VSS),.VDD(VDD),.Y(g9685),.A(g6533));
  NOT NOT1_5030(.VSS(VSS),.VDD(VDD),.Y(I26676),.A(g27736));
  NOT NOT1_5031(.VSS(VSS),.VDD(VDD),.Y(g9197),.A(g1221));
  NOT NOT1_5032(.VSS(VSS),.VDD(VDD),.Y(I18829),.A(g13350));
  NOT NOT1_5033(.VSS(VSS),.VDD(VDD),.Y(g32687),.A(g31376));
  NOT NOT1_5034(.VSS(VSS),.VDD(VDD),.Y(g9397),.A(g6088));
  NOT NOT1_5035(.VSS(VSS),.VDD(VDD),.Y(I18434),.A(g13782));
  NOT NOT1_5036(.VSS(VSS),.VDD(VDD),.Y(g33959),.A(I31878));
  NOT NOT1_5037(.VSS(VSS),.VDD(VDD),.Y(g9021),.A(I12954));
  NOT NOT1_5038(.VSS(VSS),.VDD(VDD),.Y(I12719),.A(g365));
  NOT NOT1_5039(.VSS(VSS),.VDD(VDD),.Y(g16602),.A(g14101));
  NOT NOT1_5040(.VSS(VSS),.VDD(VDD),.Y(g21410),.A(g15224));
  NOT NOT1_5041(.VSS(VSS),.VDD(VDD),.Y(g34197),.A(g33812));
  NOT NOT1_5042(.VSS(VSS),.VDD(VDD),.Y(I27718),.A(g28231));
  NOT NOT1_5043(.VSS(VSS),.VDD(VDD),.Y(I16401),.A(g869));
  NOT NOT1_5044(.VSS(VSS),.VDD(VDD),.Y(g16774),.A(g14024));
  NOT NOT1_5045(.VSS(VSS),.VDD(VDD),.Y(g23410),.A(g21562));
  NOT NOT1_5046(.VSS(VSS),.VDD(VDD),.Y(g8770),.A(g749));
  NOT NOT1_5047(.VSS(VSS),.VDD(VDD),.Y(I29337),.A(g30286));
  NOT NOT1_5048(.VSS(VSS),.VDD(VDD),.Y(g34855),.A(I33079));
  NOT NOT1_5049(.VSS(VSS),.VDD(VDD),.Y(I26654),.A(g27576));
  NOT NOT1_5050(.VSS(VSS),.VDD(VDD),.Y(I22380),.A(g21156));
  NOT NOT1_5051(.VSS(VSS),.VDD(VDD),.Y(g16955),.A(I18107));
  NOT NOT1_5052(.VSS(VSS),.VDD(VDD),.Y(g32752),.A(g31376));
  NOT NOT1_5053(.VSS(VSS),.VDD(VDD),.Y(g8296),.A(g246));
  NOT NOT1_5054(.VSS(VSS),.VDD(VDD),.Y(g25250),.A(I24434));
  NOT NOT1_5055(.VSS(VSS),.VDD(VDD),.Y(g27100),.A(g26759));
  NOT NOT1_5056(.VSS(VSS),.VDD(VDD),.Y(g32954),.A(g31376));
  NOT NOT1_5057(.VSS(VSS),.VDD(VDD),.Y(g8725),.A(g739));
  NOT NOT1_5058(.VSS(VSS),.VDD(VDD),.Y(g24083),.A(g19984));
  NOT NOT1_5059(.VSS(VSS),.VDD(VDD),.Y(g33378),.A(I30904));
  NOT NOT1_5060(.VSS(VSS),.VDD(VDD),.Y(g21666),.A(g16540));
  NOT NOT1_5061(.VSS(VSS),.VDD(VDD),.Y(g23479),.A(g21562));
  NOT NOT1_5062(.VSS(VSS),.VDD(VDD),.Y(I26936),.A(g27599));
  NOT NOT1_5063(.VSS(VSS),.VDD(VDD),.Y(g32643),.A(g31376));
  NOT NOT1_5064(.VSS(VSS),.VDD(VDD),.Y(g6940),.A(g4035));
  NOT NOT1_5065(.VSS(VSS),.VDD(VDD),.Y(I15494),.A(g10385));
  NOT NOT1_5066(.VSS(VSS),.VDD(VDD),.Y(g13075),.A(I15705));
  NOT NOT1_5067(.VSS(VSS),.VDD(VDD),.Y(g23363),.A(I22470));
  NOT NOT1_5068(.VSS(VSS),.VDD(VDD),.Y(I18344),.A(g13003));
  NOT NOT1_5069(.VSS(VSS),.VDD(VDD),.Y(g7187),.A(g6065));
  NOT NOT1_5070(.VSS(VSS),.VDD(VDD),.Y(g7387),.A(g2421));
  NOT NOT1_5071(.VSS(VSS),.VDD(VDD),.Y(g20622),.A(g15595));
  NOT NOT1_5072(.VSS(VSS),.VDD(VDD),.Y(g11467),.A(g7623));
  NOT NOT1_5073(.VSS(VSS),.VDD(VDD),.Y(g13595),.A(g10951));
  NOT NOT1_5074(.VSS(VSS),.VDD(VDD),.Y(I17999),.A(g4012));
  NOT NOT1_5075(.VSS(VSS),.VDD(VDD),.Y(g20566),.A(g15224));
  NOT NOT1_5076(.VSS(VSS),.VDD(VDD),.Y(g7461),.A(g2567));
  NOT NOT1_5077(.VSS(VSS),.VDD(VDD),.Y(I15623),.A(g12040));
  NOT NOT1_5078(.VSS(VSS),.VDD(VDD),.Y(g23478),.A(g21514));
  NOT NOT1_5079(.VSS(VSS),.VDD(VDD),.Y(g13494),.A(g11912));
  NOT NOT1_5080(.VSS(VSS),.VDD(VDD),.Y(g23015),.A(g20391));
  NOT NOT1_5081(.VSS(VSS),.VDD(VDD),.Y(g8553),.A(g3747));
  NOT NOT1_5082(.VSS(VSS),.VDD(VDD),.Y(I26334),.A(g26834));
  NOT NOT1_5083(.VSS(VSS),.VDD(VDD),.Y(I19707),.A(g17590));
  NOT NOT1_5084(.VSS(VSS),.VDD(VDD),.Y(g25296),.A(g23745));
  NOT NOT1_5085(.VSS(VSS),.VDD(VDD),.Y(g10130),.A(g5694));
  NOT NOT1_5086(.VSS(VSS),.VDD(VDD),.Y(g16171),.A(g13530));
  NOT NOT1_5087(.VSS(VSS),.VDD(VDD),.Y(g33944),.A(I31829));
  NOT NOT1_5088(.VSS(VSS),.VDD(VDD),.Y(g19061),.A(I19762));
  NOT NOT1_5089(.VSS(VSS),.VDD(VDD),.Y(g26818),.A(I25530));
  NOT NOT1_5090(.VSS(VSS),.VDD(VDD),.Y(g16886),.A(I18078));
  NOT NOT1_5091(.VSS(VSS),.VDD(VDD),.Y(I27573),.A(g28157));
  NOT NOT1_5092(.VSS(VSS),.VDD(VDD),.Y(g32669),.A(g30614));
  NOT NOT1_5093(.VSS(VSS),.VDD(VDD),.Y(I15782),.A(g10430));
  NOT NOT1_5094(.VSS(VSS),.VDD(VDD),.Y(g23486),.A(g20785));
  NOT NOT1_5095(.VSS(VSS),.VDD(VDD),.Y(g26055),.A(I25115));
  NOT NOT1_5096(.VSS(VSS),.VDD(VDD),.Y(g13037),.A(g10981));
  NOT NOT1_5097(.VSS(VSS),.VDD(VDD),.Y(g10362),.A(g6850));
  NOT NOT1_5098(.VSS(VSS),.VDD(VDD),.Y(g29149),.A(g27837));
  NOT NOT1_5099(.VSS(VSS),.VDD(VDD),.Y(g7027),.A(g5499));
  NOT NOT1_5100(.VSS(VSS),.VDD(VDD),.Y(I19818),.A(g1056));
  NOT NOT1_5101(.VSS(VSS),.VDD(VDD),.Y(g19766),.A(g16449));
  NOT NOT1_5102(.VSS(VSS),.VDD(VDD),.Y(g21556),.A(g15669));
  NOT NOT1_5103(.VSS(VSS),.VDD(VDD),.Y(I12861),.A(g4372));
  NOT NOT1_5104(.VSS(VSS),.VDD(VDD),.Y(g10165),.A(g5698));
  NOT NOT1_5105(.VSS(VSS),.VDD(VDD),.Y(g13782),.A(I16117));
  NOT NOT1_5106(.VSS(VSS),.VDD(VDD),.Y(g17575),.A(g14921));
  NOT NOT1_5107(.VSS(VSS),.VDD(VDD),.Y(g28137),.A(I26638));
  NOT NOT1_5108(.VSS(VSS),.VDD(VDD),.Y(g11984),.A(g9186));
  NOT NOT1_5109(.VSS(VSS),.VDD(VDD),.Y(g16967),.A(I18125));
  NOT NOT1_5110(.VSS(VSS),.VDD(VDD),.Y(I22331),.A(g19417));
  NOT NOT1_5111(.VSS(VSS),.VDD(VDD),.Y(g32668),.A(g31070));
  NOT NOT1_5112(.VSS(VSS),.VDD(VDD),.Y(g32842),.A(g31710));
  NOT NOT1_5113(.VSS(VSS),.VDD(VDD),.Y(g17711),.A(I18694));
  NOT NOT1_5114(.VSS(VSS),.VDD(VDD),.Y(g7046),.A(g5791));
  NOT NOT1_5115(.VSS(VSS),.VDD(VDD),.Y(I32284),.A(g34052));
  NOT NOT1_5116(.VSS(VSS),.VDD(VDD),.Y(g20653),.A(I20747));
  NOT NOT1_5117(.VSS(VSS),.VDD(VDD),.Y(g27991),.A(g25852));
  NOT NOT1_5118(.VSS(VSS),.VDD(VDD),.Y(I33288),.A(g34989));
  NOT NOT1_5119(.VSS(VSS),.VDD(VDD),.Y(g31802),.A(g29385));
  NOT NOT1_5120(.VSS(VSS),.VDD(VDD),.Y(g9631),.A(g6573));
  NOT NOT1_5121(.VSS(VSS),.VDD(VDD),.Y(g17327),.A(I18310));
  NOT NOT1_5122(.VSS(VSS),.VDD(VDD),.Y(g25060),.A(g23708));
  NOT NOT1_5123(.VSS(VSS),.VDD(VDD),.Y(g32489),.A(g30614));
  NOT NOT1_5124(.VSS(VSS),.VDD(VDD),.Y(g8389),.A(g3125));
  NOT NOT1_5125(.VSS(VSS),.VDD(VDD),.Y(I13329),.A(g86));
  NOT NOT1_5126(.VSS(VSS),.VDD(VDD),.Y(I27388),.A(g27698));
  NOT NOT1_5127(.VSS(VSS),.VDD(VDD),.Y(g31857),.A(g29385));
  NOT NOT1_5128(.VSS(VSS),.VDD(VDD),.Y(g7446),.A(g1256));
  NOT NOT1_5129(.VSS(VSS),.VDD(VDD),.Y(g18200),.A(I19012));
  NOT NOT1_5130(.VSS(VSS),.VDD(VDD),.Y(g29811),.A(g28376));
  NOT NOT1_5131(.VSS(VSS),.VDD(VDD),.Y(g23223),.A(g21308));
  NOT NOT1_5132(.VSS(VSS),.VDD(VDD),.Y(g7514),.A(g6704));
  NOT NOT1_5133(.VSS(VSS),.VDD(VDD),.Y(g19360),.A(g16249));
  NOT NOT1_5134(.VSS(VSS),.VDD(VDD),.Y(g11418),.A(I14424));
  NOT NOT1_5135(.VSS(VSS),.VDD(VDD),.Y(g34714),.A(I32874));
  NOT NOT1_5136(.VSS(VSS),.VDD(VDD),.Y(g8990),.A(g146));
  NOT NOT1_5137(.VSS(VSS),.VDD(VDD),.Y(g12882),.A(g10389));
  NOT NOT1_5138(.VSS(VSS),.VDD(VDD),.Y(g9257),.A(g5115));
  NOT NOT1_5139(.VSS(VSS),.VDD(VDD),.Y(g22492),.A(g19614));
  NOT NOT1_5140(.VSS(VSS),.VDD(VDD),.Y(g25197),.A(g23958));
  NOT NOT1_5141(.VSS(VSS),.VDD(VDD),.Y(g29343),.A(g28174));
  NOT NOT1_5142(.VSS(VSS),.VDD(VDD),.Y(g7003),.A(g5152));
  NOT NOT1_5143(.VSS(VSS),.VDD(VDD),.Y(I13539),.A(g6381));
  NOT NOT1_5144(.VSS(VSS),.VDD(VDD),.Y(g22303),.A(g19277));
  NOT NOT1_5145(.VSS(VSS),.VDD(VDD),.Y(I27777),.A(g29043));
  NOT NOT1_5146(.VSS(VSS),.VDD(VDD),.Y(g9817),.A(I13374));
  NOT NOT1_5147(.VSS(VSS),.VDD(VDD),.Y(g32559),.A(g30825));
  NOT NOT1_5148(.VSS(VSS),.VDD(VDD),.Y(g34315),.A(g34085));
  NOT NOT1_5149(.VSS(VSS),.VDD(VDD),.Y(g10475),.A(g8844));
  NOT NOT1_5150(.VSS(VSS),.VDD(VDD),.Y(I17932),.A(g3310));
  NOT NOT1_5151(.VSS(VSS),.VDD(VDD),.Y(g24138),.A(g21143));
  NOT NOT1_5152(.VSS(VSS),.VDD(VDD),.Y(g32525),.A(g31170));
  NOT NOT1_5153(.VSS(VSS),.VDD(VDD),.Y(g32488),.A(g31194));
  NOT NOT1_5154(.VSS(VSS),.VDD(VDD),.Y(g11170),.A(g8476));
  NOT NOT1_5155(.VSS(VSS),.VDD(VDD),.Y(g34910),.A(g34864));
  NOT NOT1_5156(.VSS(VSS),.VDD(VDD),.Y(I29444),.A(g30928));
  NOT NOT1_5157(.VSS(VSS),.VDD(VDD),.Y(g8171),.A(g3817));
  NOT NOT1_5158(.VSS(VSS),.VDD(VDD),.Y(g10727),.A(I14016));
  NOT NOT1_5159(.VSS(VSS),.VDD(VDD),.Y(g7345),.A(g6415));
  NOT NOT1_5160(.VSS(VSS),.VDD(VDD),.Y(g7841),.A(g904));
  NOT NOT1_5161(.VSS(VSS),.VDD(VDD),.Y(I12534),.A(g50));
  NOT NOT1_5162(.VSS(VSS),.VDD(VDD),.Y(g20636),.A(g18008));
  NOT NOT1_5163(.VSS(VSS),.VDD(VDD),.Y(I19384),.A(g15085));
  NOT NOT1_5164(.VSS(VSS),.VDD(VDD),.Y(g8787),.A(I12773));
  NOT NOT1_5165(.VSS(VSS),.VDD(VDD),.Y(g32558),.A(g30735));
  NOT NOT1_5166(.VSS(VSS),.VDD(VDD),.Y(g34202),.A(I32161));
  NOT NOT1_5167(.VSS(VSS),.VDD(VDD),.Y(g23084),.A(g19954));
  NOT NOT1_5168(.VSS(VSS),.VDD(VDD),.Y(g24636),.A(g23121));
  NOT NOT1_5169(.VSS(VSS),.VDD(VDD),.Y(g6826),.A(g218));
  NOT NOT1_5170(.VSS(VSS),.VDD(VDD),.Y(g10222),.A(g4492));
  NOT NOT1_5171(.VSS(VSS),.VDD(VDD),.Y(g7191),.A(g6398));
  NOT NOT1_5172(.VSS(VSS),.VDD(VDD),.Y(g30055),.A(g29157));
  NOT NOT1_5173(.VSS(VSS),.VDD(VDD),.Y(g17606),.A(g14999));
  NOT NOT1_5174(.VSS(VSS),.VDD(VDD),.Y(g20852),.A(g15595));
  NOT NOT1_5175(.VSS(VSS),.VDD(VDD),.Y(g32830),.A(g31327));
  NOT NOT1_5176(.VSS(VSS),.VDD(VDD),.Y(g23922),.A(g18997));
  NOT NOT1_5177(.VSS(VSS),.VDD(VDD),.Y(g23321),.A(I22422));
  NOT NOT1_5178(.VSS(VSS),.VDD(VDD),.Y(g32893),.A(g30937));
  NOT NOT1_5179(.VSS(VSS),.VDD(VDD),.Y(I18028),.A(g13638));
  NOT NOT1_5180(.VSS(VSS),.VDD(VDD),.Y(g21179),.A(g15373));
  NOT NOT1_5181(.VSS(VSS),.VDD(VDD),.Y(I24920),.A(g25513));
  NOT NOT1_5182(.VSS(VSS),.VDD(VDD),.Y(g26801),.A(I25511));
  NOT NOT1_5183(.VSS(VSS),.VDD(VDD),.Y(I24434),.A(g22763));
  NOT NOT1_5184(.VSS(VSS),.VDD(VDD),.Y(g29368),.A(I27730));
  NOT NOT1_5185(.VSS(VSS),.VDD(VDD),.Y(g9751),.A(g1710));
  NOT NOT1_5186(.VSS(VSS),.VDD(VDD),.Y(g34070),.A(g33725));
  NOT NOT1_5187(.VSS(VSS),.VDD(VDD),.Y(g8281),.A(g3494));
  NOT NOT1_5188(.VSS(VSS),.VDD(VDD),.Y(g32544),.A(g30735));
  NOT NOT1_5189(.VSS(VSS),.VDD(VDD),.Y(g19629),.A(g17015));
  NOT NOT1_5190(.VSS(VSS),.VDD(VDD),.Y(g32865),.A(g31327));
  NOT NOT1_5191(.VSS(VSS),.VDD(VDD),.Y(g19451),.A(g15938));
  NOT NOT1_5192(.VSS(VSS),.VDD(VDD),.Y(g21178),.A(g17955));
  NOT NOT1_5193(.VSS(VSS),.VDD(VDD),.Y(g34590),.A(I32678));
  NOT NOT1_5194(.VSS(VSS),.VDD(VDD),.Y(g19472),.A(g16349));
  NOT NOT1_5195(.VSS(VSS),.VDD(VDD),.Y(g24963),.A(g22342));
  NOT NOT1_5196(.VSS(VSS),.VDD(VDD),.Y(g20664),.A(g15373));
  NOT NOT1_5197(.VSS(VSS),.VDD(VDD),.Y(g34986),.A(I33258));
  NOT NOT1_5198(.VSS(VSS),.VDD(VDD),.Y(g32713),.A(g30673));
  NOT NOT1_5199(.VSS(VSS),.VDD(VDD),.Y(g7536),.A(g5976));
  NOT NOT1_5200(.VSS(VSS),.VDD(VDD),.Y(g9585),.A(g1616));
  NOT NOT1_5201(.VSS(VSS),.VDD(VDD),.Y(g8297),.A(g142));
  NOT NOT1_5202(.VSS(VSS),.VDD(VDD),.Y(g10347),.A(I13759));
  NOT NOT1_5203(.VSS(VSS),.VDD(VDD),.Y(g21685),.A(I21246));
  NOT NOT1_5204(.VSS(VSS),.VDD(VDD),.Y(I16733),.A(g12026));
  NOT NOT1_5205(.VSS(VSS),.VDD(VDD),.Y(I12997),.A(g351));
  NOT NOT1_5206(.VSS(VSS),.VDD(VDD),.Y(g28726),.A(g27937));
  NOT NOT1_5207(.VSS(VSS),.VDD(VDD),.Y(g34384),.A(I32391));
  NOT NOT1_5208(.VSS(VSS),.VDD(VDD),.Y(g23953),.A(g19277));
  NOT NOT1_5209(.VSS(VSS),.VDD(VDD),.Y(g30067),.A(g29060));
  NOT NOT1_5210(.VSS(VSS),.VDD(VDD),.Y(g11401),.A(g7593));
  NOT NOT1_5211(.VSS(VSS),.VDD(VDD),.Y(g22840),.A(g20330));
  NOT NOT1_5212(.VSS(VSS),.VDD(VDD),.Y(g21654),.A(g17619));
  NOT NOT1_5213(.VSS(VSS),.VDD(VDD),.Y(I29977),.A(g31596));
  NOT NOT1_5214(.VSS(VSS),.VDD(VDD),.Y(g7858),.A(g947));
  NOT NOT1_5215(.VSS(VSS),.VDD(VDD),.Y(g32610),.A(g31070));
  NOT NOT1_5216(.VSS(VSS),.VDD(VDD),.Y(g20576),.A(g18065));
  NOT NOT1_5217(.VSS(VSS),.VDD(VDD),.Y(g20585),.A(g17955));
  NOT NOT1_5218(.VSS(VSS),.VDD(VDD),.Y(g23654),.A(g20248));
  NOT NOT1_5219(.VSS(VSS),.VDD(VDD),.Y(I12061),.A(g562));
  NOT NOT1_5220(.VSS(VSS),.VDD(VDD),.Y(g32705),.A(g30614));
  NOT NOT1_5221(.VSS(VSS),.VDD(VDD),.Y(g34094),.A(g33772));
  NOT NOT1_5222(.VSS(VSS),.VDD(VDD),.Y(g13477),.A(I15954));
  NOT NOT1_5223(.VSS(VSS),.VDD(VDD),.Y(g8745),.A(g744));
  NOT NOT1_5224(.VSS(VSS),.VDD(VDD),.Y(g28436),.A(I26929));
  NOT NOT1_5225(.VSS(VSS),.VDD(VDD),.Y(g8138),.A(g1500));
  NOT NOT1_5226(.VSS(VSS),.VDD(VDD),.Y(g8639),.A(g2807));
  NOT NOT1_5227(.VSS(VSS),.VDD(VDD),.Y(g24585),.A(g23063));
  NOT NOT1_5228(.VSS(VSS),.VDD(VDD),.Y(I22149),.A(g21036));
  NOT NOT1_5229(.VSS(VSS),.VDD(VDD),.Y(g19071),.A(g15591));
  NOT NOT1_5230(.VSS(VSS),.VDD(VDD),.Y(g23800),.A(g21246));
  NOT NOT1_5231(.VSS(VSS),.VDD(VDD),.Y(I23711),.A(g23192));
  NOT NOT1_5232(.VSS(VSS),.VDD(VDD),.Y(g20554),.A(g15348));
  NOT NOT1_5233(.VSS(VSS),.VDD(VDD),.Y(g23417),.A(g20391));
  NOT NOT1_5234(.VSS(VSS),.VDD(VDD),.Y(g32679),.A(g31579));
  NOT NOT1_5235(.VSS(VSS),.VDD(VDD),.Y(g16322),.A(I17650));
  NOT NOT1_5236(.VSS(VSS),.VDD(VDD),.Y(g8791),.A(I12787));
  NOT NOT1_5237(.VSS(VSS),.VDD(VDD),.Y(g10351),.A(g6802));
  NOT NOT1_5238(.VSS(VSS),.VDD(VDD),.Y(g23936),.A(g19210));
  NOT NOT1_5239(.VSS(VSS),.VDD(VDD),.Y(g10372),.A(g6900));
  NOT NOT1_5240(.VSS(VSS),.VDD(VDD),.Y(I23327),.A(g22647));
  NOT NOT1_5241(.VSS(VSS),.VDD(VDD),.Y(g25202),.A(g23932));
  NOT NOT1_5242(.VSS(VSS),.VDD(VDD),.Y(g19776),.A(g17015));
  NOT NOT1_5243(.VSS(VSS),.VDD(VDD),.Y(g19785),.A(g16987));
  NOT NOT1_5244(.VSS(VSS),.VDD(VDD),.Y(g34150),.A(I32103));
  NOT NOT1_5245(.VSS(VSS),.VDD(VDD),.Y(I32963),.A(g34650));
  NOT NOT1_5246(.VSS(VSS),.VDD(VDD),.Y(g16159),.A(g13584));
  NOT NOT1_5247(.VSS(VSS),.VDD(VDD),.Y(g22192),.A(g19801));
  NOT NOT1_5248(.VSS(VSS),.VDD(VDD),.Y(g20609),.A(g15373));
  NOT NOT1_5249(.VSS(VSS),.VDD(VDD),.Y(g28274),.A(I26799));
  NOT NOT1_5250(.VSS(VSS),.VDD(VDD),.Y(g15171),.A(I17098));
  NOT NOT1_5251(.VSS(VSS),.VDD(VDD),.Y(g34877),.A(I33103));
  NOT NOT1_5252(.VSS(VSS),.VDD(VDD),.Y(g10175),.A(g28));
  NOT NOT1_5253(.VSS(VSS),.VDD(VDD),.Y(I17723),.A(g13177));
  NOT NOT1_5254(.VSS(VSS),.VDD(VDD),.Y(g12082),.A(g9645));
  NOT NOT1_5255(.VSS(VSS),.VDD(VDD),.Y(g17390),.A(g14755));
  NOT NOT1_5256(.VSS(VSS),.VDD(VDD),.Y(g28593),.A(g27727));
  NOT NOT1_5257(.VSS(VSS),.VDD(VDD),.Y(g32678),.A(g31528));
  NOT NOT1_5258(.VSS(VSS),.VDD(VDD),.Y(g13022),.A(g11894));
  NOT NOT1_5259(.VSS(VSS),.VDD(VDD),.Y(g7522),.A(g6661));
  NOT NOT1_5260(.VSS(VSS),.VDD(VDD),.Y(g23334),.A(g20785));
  NOT NOT1_5261(.VSS(VSS),.VDD(VDD),.Y(g25055),.A(g23590));
  NOT NOT1_5262(.VSS(VSS),.VDD(VDD),.Y(g19147),.A(I19786));
  NOT NOT1_5263(.VSS(VSS),.VDD(VDD),.Y(g30019),.A(g29060));
  NOT NOT1_5264(.VSS(VSS),.VDD(VDD),.Y(g7115),.A(g12));
  NOT NOT1_5265(.VSS(VSS),.VDD(VDD),.Y(g12107),.A(g9687));
  NOT NOT1_5266(.VSS(VSS),.VDD(VDD),.Y(g8808),.A(g595));
  NOT NOT1_5267(.VSS(VSS),.VDD(VDD),.Y(g19754),.A(g17062));
  NOT NOT1_5268(.VSS(VSS),.VDD(VDD),.Y(g7315),.A(g1772));
  NOT NOT1_5269(.VSS(VSS),.VDD(VDD),.Y(g16158),.A(g13555));
  NOT NOT1_5270(.VSS(VSS),.VDD(VDD),.Y(g20608),.A(g15171));
  NOT NOT1_5271(.VSS(VSS),.VDD(VDD),.Y(g25111),.A(g23699));
  NOT NOT1_5272(.VSS(VSS),.VDD(VDD),.Y(g9669),.A(g5092));
  NOT NOT1_5273(.VSS(VSS),.VDD(VDD),.Y(g19355),.A(g16027));
  NOT NOT1_5274(.VSS(VSS),.VDD(VDD),.Y(I12360),.A(g528));
  NOT NOT1_5275(.VSS(VSS),.VDD(VDD),.Y(g25070),.A(g23590));
  NOT NOT1_5276(.VSS(VSS),.VDD(VDD),.Y(g32460),.A(g31194));
  NOT NOT1_5277(.VSS(VSS),.VDD(VDD),.Y(g32686),.A(g31579));
  NOT NOT1_5278(.VSS(VSS),.VDD(VDD),.Y(I22343),.A(g19371));
  NOT NOT1_5279(.VSS(VSS),.VDD(VDD),.Y(g24115),.A(g20998));
  NOT NOT1_5280(.VSS(VSS),.VDD(VDD),.Y(g32939),.A(g31327));
  NOT NOT1_5281(.VSS(VSS),.VDD(VDD),.Y(I18903),.A(g16872));
  NOT NOT1_5282(.VSS(VSS),.VDD(VDD),.Y(g30018),.A(g28987));
  NOT NOT1_5283(.VSS(VSS),.VDD(VDD),.Y(g32383),.A(I29913));
  NOT NOT1_5284(.VSS(VSS),.VDD(VDD),.Y(g19950),.A(g15885));
  NOT NOT1_5285(.VSS(VSS),.VDD(VDD),.Y(g14063),.A(g11048));
  NOT NOT1_5286(.VSS(VSS),.VDD(VDD),.Y(g19370),.A(g15915));
  NOT NOT1_5287(.VSS(VSS),.VDD(VDD),.Y(I19917),.A(g18088));
  NOT NOT1_5288(.VSS(VSS),.VDD(VDD),.Y(I14046),.A(g9900));
  NOT NOT1_5289(.VSS(VSS),.VDD(VDD),.Y(I17148),.A(g14442));
  NOT NOT1_5290(.VSS(VSS),.VDD(VDD),.Y(g16656),.A(I17852));
  NOT NOT1_5291(.VSS(VSS),.VDD(VDD),.Y(g9772),.A(I13352));
  NOT NOT1_5292(.VSS(VSS),.VDD(VDD),.Y(I26638),.A(g27965));
  NOT NOT1_5293(.VSS(VSS),.VDD(VDD),.Y(g20921),.A(g15426));
  NOT NOT1_5294(.VSS(VSS),.VDD(VDD),.Y(g12345),.A(g7158));
  NOT NOT1_5295(.VSS(VSS),.VDD(VDD),.Y(I16476),.A(g10430));
  NOT NOT1_5296(.VSS(VSS),.VDD(VDD),.Y(g14790),.A(I16855));
  NOT NOT1_5297(.VSS(VSS),.VDD(VDD),.Y(g20052),.A(g17533));
  NOT NOT1_5298(.VSS(VSS),.VDD(VDD),.Y(g23964),.A(g19147));
  NOT NOT1_5299(.VSS(VSS),.VDD(VDD),.Y(I23303),.A(g21669));
  NOT NOT1_5300(.VSS(VSS),.VDD(VDD),.Y(g32938),.A(g30937));
  NOT NOT1_5301(.VSS(VSS),.VDD(VDD),.Y(g28034),.A(g26365));
  NOT NOT1_5302(.VSS(VSS),.VDD(VDD),.Y(g33533),.A(I31361));
  NOT NOT1_5303(.VSS(VSS),.VDD(VDD),.Y(g29310),.A(g28991));
  NOT NOT1_5304(.VSS(VSS),.VDD(VDD),.Y(g16680),.A(g13223));
  NOT NOT1_5305(.VSS(VSS),.VDD(VDD),.Y(g24052),.A(g21193));
  NOT NOT1_5306(.VSS(VSS),.VDD(VDD),.Y(I17104),.A(g12932));
  NOT NOT1_5307(.VSS(VSS),.VDD(VDD),.Y(g12940),.A(g11744));
  NOT NOT1_5308(.VSS(VSS),.VDD(VDD),.Y(g17522),.A(g14927));
  NOT NOT1_5309(.VSS(VSS),.VDD(VDD),.Y(g21423),.A(g15224));
  NOT NOT1_5310(.VSS(VSS),.VDD(VDD),.Y(g12399),.A(g9920));
  NOT NOT1_5311(.VSS(VSS),.VDD(VDD),.Y(g9743),.A(I13321));
  NOT NOT1_5312(.VSS(VSS),.VDD(VDD),.Y(I16555),.A(g10430));
  NOT NOT1_5313(.VSS(VSS),.VDD(VDD),.Y(g23423),.A(g20871));
  NOT NOT1_5314(.VSS(VSS),.VDD(VDD),.Y(g8201),.A(g1894));
  NOT NOT1_5315(.VSS(VSS),.VDD(VDD),.Y(g9890),.A(g6058));
  NOT NOT1_5316(.VSS(VSS),.VDD(VDD),.Y(g13305),.A(g11048));
  NOT NOT1_5317(.VSS(VSS),.VDD(VDD),.Y(g6827),.A(g1277));
  NOT NOT1_5318(.VSS(VSS),.VDD(VDD),.Y(g14873),.A(I16898));
  NOT NOT1_5319(.VSS(VSS),.VDD(VDD),.Y(g23216),.A(g20924));
  NOT NOT1_5320(.VSS(VSS),.VDD(VDD),.Y(g11900),.A(I14708));
  NOT NOT1_5321(.VSS(VSS),.VDD(VDD),.Y(g19996),.A(g17271));
  NOT NOT1_5322(.VSS(VSS),.VDD(VDD),.Y(g29379),.A(I27749));
  NOT NOT1_5323(.VSS(VSS),.VDD(VDD),.Y(g29925),.A(g28820));
  NOT NOT1_5324(.VSS(VSS),.VDD(VDD),.Y(g13809),.A(I16135));
  NOT NOT1_5325(.VSS(VSS),.VDD(VDD),.Y(I23381),.A(g23322));
  NOT NOT1_5326(.VSS(VSS),.VDD(VDD),.Y(I15036),.A(g799));
  NOT NOT1_5327(.VSS(VSS),.VDD(VDD),.Y(g8449),.A(g3752));
  NOT NOT1_5328(.VSS(VSS),.VDD(VDD),.Y(g12804),.A(g9927));
  NOT NOT1_5329(.VSS(VSS),.VDD(VDD),.Y(g9011),.A(g1422));
  NOT NOT1_5330(.VSS(VSS),.VDD(VDD),.Y(g19367),.A(I19851));
  NOT NOT1_5331(.VSS(VSS),.VDD(VDD),.Y(g19394),.A(g16326));
  NOT NOT1_5332(.VSS(VSS),.VDD(VDD),.Y(I12451),.A(g3092));
  NOT NOT1_5333(.VSS(VSS),.VDD(VDD),.Y(g6846),.A(g2152));
  NOT NOT1_5334(.VSS(VSS),.VDD(VDD),.Y(g9856),.A(g5343));
  NOT NOT1_5335(.VSS(VSS),.VDD(VDD),.Y(g8575),.A(g291));
  NOT NOT1_5336(.VSS(VSS),.VDD(VDD),.Y(g13036),.A(g10981));
  NOT NOT1_5337(.VSS(VSS),.VDD(VDD),.Y(g32875),.A(g31376));
  NOT NOT1_5338(.VSS(VSS),.VDD(VDD),.Y(g30917),.A(I28897));
  NOT NOT1_5339(.VSS(VSS),.VDD(VDD),.Y(I14827),.A(g9686));
  NOT NOT1_5340(.VSS(VSS),.VDD(VDD),.Y(g11560),.A(g7647));
  NOT NOT1_5341(.VSS(VSS),.VDD(VDD),.Y(g13101),.A(I15736));
  NOT NOT1_5342(.VSS(VSS),.VDD(VDD),.Y(g14209),.A(g11415));
  NOT NOT1_5343(.VSS(VSS),.VDD(VDD),.Y(g7880),.A(g1291));
  NOT NOT1_5344(.VSS(VSS),.VDD(VDD),.Y(g13177),.A(I15782));
  NOT NOT1_5345(.VSS(VSS),.VDD(VDD),.Y(g34917),.A(I33143));
  NOT NOT1_5346(.VSS(VSS),.VDD(VDD),.Y(g8715),.A(g4927));
  NOT NOT1_5347(.VSS(VSS),.VDD(VDD),.Y(g20674),.A(g15277));
  NOT NOT1_5348(.VSS(VSS),.VDD(VDD),.Y(g7595),.A(I12067));
  NOT NOT1_5349(.VSS(VSS),.VDD(VDD),.Y(g23543),.A(g21514));
  NOT NOT1_5350(.VSS(VSS),.VDD(VDD),.Y(g6803),.A(g496));
  NOT NOT1_5351(.VSS(VSS),.VDD(VDD),.Y(g16966),.A(g14291));
  NOT NOT1_5352(.VSS(VSS),.VDD(VDD),.Y(g7537),.A(g311));
  NOT NOT1_5353(.VSS(VSS),.VDD(VDD),.Y(g24184),.A(I23396));
  NOT NOT1_5354(.VSS(VSS),.VDD(VDD),.Y(I18845),.A(g6711));
  NOT NOT1_5355(.VSS(VSS),.VDD(VDD),.Y(I32921),.A(g34650));
  NOT NOT1_5356(.VSS(VSS),.VDD(VDD),.Y(g16631),.A(g14454));
  NOT NOT1_5357(.VSS(VSS),.VDD(VDD),.Y(g14208),.A(g11563));
  NOT NOT1_5358(.VSS(VSS),.VDD(VDD),.Y(I18262),.A(g13857));
  NOT NOT1_5359(.VSS(VSS),.VDD(VDD),.Y(g29944),.A(g28911));
  NOT NOT1_5360(.VSS(VSS),.VDD(VDD),.Y(g22904),.A(I22111));
  NOT NOT1_5361(.VSS(VSS),.VDD(VDD),.Y(g23000),.A(g20453));
  NOT NOT1_5362(.VSS(VSS),.VDD(VDD),.Y(I26578),.A(g26941));
  NOT NOT1_5363(.VSS(VSS),.VDD(VDD),.Y(g23908),.A(g20739));
  NOT NOT1_5364(.VSS(VSS),.VDD(VDD),.Y(g17326),.A(I18307));
  NOT NOT1_5365(.VSS(VSS),.VDD(VDD),.Y(g32837),.A(g31327));
  NOT NOT1_5366(.VSS(VSS),.VDD(VDD),.Y(g31856),.A(g29385));
  NOT NOT1_5367(.VSS(VSS),.VDD(VDD),.Y(I13206),.A(g5448));
  NOT NOT1_5368(.VSS(VSS),.VDD(VDD),.Y(g8833),.A(g794));
  NOT NOT1_5369(.VSS(VSS),.VDD(VDD),.Y(g30077),.A(g29057));
  NOT NOT1_5370(.VSS(VSS),.VDD(VDD),.Y(g9992),.A(g5990));
  NOT NOT1_5371(.VSS(VSS),.VDD(VDD),.Y(g20732),.A(g15595));
  NOT NOT1_5372(.VSS(VSS),.VDD(VDD),.Y(g23569),.A(g21611));
  NOT NOT1_5373(.VSS(VSS),.VDD(VDD),.Y(g25196),.A(g22763));
  NOT NOT1_5374(.VSS(VSS),.VDD(VDD),.Y(g10542),.A(g7196));
  NOT NOT1_5375(.VSS(VSS),.VDD(VDD),.Y(I31610),.A(g33149));
  NOT NOT1_5376(.VSS(VSS),.VDD(VDD),.Y(I23390),.A(g23395));
  NOT NOT1_5377(.VSS(VSS),.VDD(VDD),.Y(g13064),.A(g11705));
  NOT NOT1_5378(.VSS(VSS),.VDD(VDD),.Y(g24732),.A(g23042));
  NOT NOT1_5379(.VSS(VSS),.VDD(VDD),.Y(g14453),.A(I16610));
  NOT NOT1_5380(.VSS(VSS),.VDD(VDD),.Y(g7017),.A(g128));
  NOT NOT1_5381(.VSS(VSS),.VDD(VDD),.Y(I30992),.A(g32445));
  NOT NOT1_5382(.VSS(VSS),.VDD(VDD),.Y(g7243),.A(I11892));
  NOT NOT1_5383(.VSS(VSS),.VDD(VDD),.Y(g19446),.A(I19917));
  NOT NOT1_5384(.VSS(VSS),.VDD(VDD),.Y(g34597),.A(I32699));
  NOT NOT1_5385(.VSS(VSS),.VDD(VDD),.Y(I12776),.A(g4207));
  NOT NOT1_5386(.VSS(VSS),.VDD(VDD),.Y(I13759),.A(g6754));
  NOT NOT1_5387(.VSS(VSS),.VDD(VDD),.Y(I18191),.A(g14385));
  NOT NOT1_5388(.VSS(VSS),.VDD(VDD),.Y(g23568),.A(g21611));
  NOT NOT1_5389(.VSS(VSS),.VDD(VDD),.Y(I33255),.A(g34975));
  NOT NOT1_5390(.VSS(VSS),.VDD(VDD),.Y(I33189),.A(g34929));
  NOT NOT1_5391(.VSS(VSS),.VDD(VDD),.Y(g8584),.A(g3639));
  NOT NOT1_5392(.VSS(VSS),.VDD(VDD),.Y(g8539),.A(g3454));
  NOT NOT1_5393(.VSS(VSS),.VDD(VDD),.Y(g23242),.A(g21070));
  NOT NOT1_5394(.VSS(VSS),.VDD(VDD),.Y(I32973),.A(g34714));
  NOT NOT1_5395(.VSS(VSS),.VDD(VDD),.Y(I29571),.A(g31783));
  NOT NOT1_5396(.VSS(VSS),.VDD(VDD),.Y(g34689),.A(I32837));
  NOT NOT1_5397(.VSS(VSS),.VDD(VDD),.Y(I33270),.A(g34982));
  NOT NOT1_5398(.VSS(VSS),.VDD(VDD),.Y(g34923),.A(I33161));
  NOT NOT1_5399(.VSS(VSS),.VDD(VDD),.Y(g9863),.A(g5503));
  NOT NOT1_5400(.VSS(VSS),.VDD(VDD),.Y(I12355),.A(g46));
  NOT NOT1_5401(.VSS(VSS),.VDD(VDD),.Y(g16289),.A(g13223));
  NOT NOT1_5402(.VSS(VSS),.VDD(VDD),.Y(g9480),.A(g559));
  NOT NOT1_5403(.VSS(VSS),.VDD(VDD),.Y(I17228),.A(g13350));
  NOT NOT1_5404(.VSS(VSS),.VDD(VDD),.Y(g6994),.A(g4933));
  NOT NOT1_5405(.VSS(VSS),.VDD(VDD),.Y(g21123),.A(g15615));
  NOT NOT1_5406(.VSS(VSS),.VDD(VDD),.Y(g18100),.A(I18906));
  NOT NOT1_5407(.VSS(VSS),.VDD(VDD),.Y(g34688),.A(I32834));
  NOT NOT1_5408(.VSS(VSS),.VDD(VDD),.Y(g9713),.A(g3618));
  NOT NOT1_5409(.VSS(VSS),.VDD(VDD),.Y(g10607),.A(g10233));
  NOT NOT1_5410(.VSS(VSS),.VDD(VDD),.Y(g12833),.A(I15448));
  NOT NOT1_5411(.VSS(VSS),.VDD(VDD),.Y(g22847),.A(g20283));
  NOT NOT1_5412(.VSS(VSS),.VDD(VDD),.Y(g16309),.A(I17639));
  NOT NOT1_5413(.VSS(VSS),.VDD(VDD),.Y(I12950),.A(g4287));
  NOT NOT1_5414(.VSS(VSS),.VDD(VDD),.Y(g23814),.A(g19074));
  NOT NOT1_5415(.VSS(VSS),.VDD(VDD),.Y(g10320),.A(g817));
  NOT NOT1_5416(.VSS(VSS),.VDD(VDD),.Y(g32617),.A(g30825));
  NOT NOT1_5417(.VSS(VSS),.VDD(VDD),.Y(g28575),.A(g27711));
  NOT NOT1_5418(.VSS(VSS),.VDD(VDD),.Y(g32470),.A(g31566));
  NOT NOT1_5419(.VSS(VSS),.VDD(VDD),.Y(g10073),.A(g134));
  NOT NOT1_5420(.VSS(VSS),.VDD(VDD),.Y(I18832),.A(g13782));
  NOT NOT1_5421(.VSS(VSS),.VDD(VDD),.Y(I31686),.A(g33164));
  NOT NOT1_5422(.VSS(VSS),.VDD(VDD),.Y(g7328),.A(g2197));
  NOT NOT1_5423(.VSS(VSS),.VDD(VDD),.Y(g32915),.A(g31710));
  NOT NOT1_5424(.VSS(VSS),.VDD(VDD),.Y(g10274),.A(g976));
  NOT NOT1_5425(.VSS(VSS),.VDD(VDD),.Y(g29765),.A(I28014));
  NOT NOT1_5426(.VSS(VSS),.VDD(VDD),.Y(g10530),.A(g8922));
  NOT NOT1_5427(.VSS(VSS),.VDD(VDD),.Y(g7542),.A(I12030));
  NOT NOT1_5428(.VSS(VSS),.VDD(VDD),.Y(I12858),.A(g4340));
  NOT NOT1_5429(.VSS(VSS),.VDD(VDD),.Y(g28711),.A(g27886));
  NOT NOT1_5430(.VSS(VSS),.VDD(VDD),.Y(g13009),.A(I15617));
  NOT NOT1_5431(.VSS(VSS),.VDD(VDD),.Y(g16308),.A(I17636));
  NOT NOT1_5432(.VSS(VSS),.VDD(VDD),.Y(g9569),.A(g6227));
  NOT NOT1_5433(.VSS(VSS),.VDD(VDD),.Y(g13665),.A(g11306));
  NOT NOT1_5434(.VSS(VSS),.VDD(VDD),.Y(g27004),.A(g26131));
  NOT NOT1_5435(.VSS(VSS),.VDD(VDD),.Y(g30102),.A(g29157));
  NOT NOT1_5436(.VSS(VSS),.VDD(VDD),.Y(g8362),.A(g194));
  NOT NOT1_5437(.VSS(VSS),.VDD(VDD),.Y(I13744),.A(g3518));
  NOT NOT1_5438(.VSS(VSS),.VDD(VDD),.Y(g31831),.A(g29385));
  NOT NOT1_5439(.VSS(VSS),.VDD(VDD),.Y(g32201),.A(g31509));
  NOT NOT1_5440(.VSS(VSS),.VDD(VDD),.Y(g24013),.A(g21611));
  NOT NOT1_5441(.VSS(VSS),.VDD(VDD),.Y(I33030),.A(g34768));
  NOT NOT1_5442(.VSS(VSS),.VDD(VDD),.Y(I12151),.A(g604));
  NOT NOT1_5443(.VSS(VSS),.VDD(VDD),.Y(g10122),.A(I13623));
  NOT NOT1_5444(.VSS(VSS),.VDD(VDD),.Y(g6816),.A(g933));
  NOT NOT1_5445(.VSS(VSS),.VDD(VDD),.Y(I12172),.A(g2715));
  NOT NOT1_5446(.VSS(VSS),.VDD(VDD),.Y(g17183),.A(I18221));
  NOT NOT1_5447(.VSS(VSS),.VDD(VDD),.Y(g17673),.A(g14723));
  NOT NOT1_5448(.VSS(VSS),.VDD(VDD),.Y(g17847),.A(I18839));
  NOT NOT1_5449(.VSS(VSS),.VDD(VDD),.Y(I26430),.A(g26856));
  NOT NOT1_5450(.VSS(VSS),.VDD(VDD),.Y(g13008),.A(g11855));
  NOT NOT1_5451(.VSS(VSS),.VDD(VDD),.Y(g15656),.A(I17198));
  NOT NOT1_5452(.VSS(VSS),.VDD(VDD),.Y(I21483),.A(g18726));
  NOT NOT1_5453(.VSS(VSS),.VDD(VDD),.Y(g20329),.A(g15277));
  NOT NOT1_5454(.VSS(VSS),.VDD(VDD),.Y(I33267),.A(g34979));
  NOT NOT1_5455(.VSS(VSS),.VDD(VDD),.Y(g8052),.A(g1211));
  NOT NOT1_5456(.VSS(VSS),.VDD(VDD),.Y(I18861),.A(g14307));
  NOT NOT1_5457(.VSS(VSS),.VDD(VDD),.Y(g21293),.A(I21036));
  NOT NOT1_5458(.VSS(VSS),.VDD(VDD),.Y(g20207),.A(g17015));
  NOT NOT1_5459(.VSS(VSS),.VDD(VDD),.Y(g23230),.A(I22327));
  NOT NOT1_5460(.VSS(VSS),.VDD(VDD),.Y(g15680),.A(I17207));
  NOT NOT1_5461(.VSS(VSS),.VDD(VDD),.Y(g20539),.A(g15483));
  NOT NOT1_5462(.VSS(VSS),.VDD(VDD),.Y(g25001),.A(g23666));
  NOT NOT1_5463(.VSS(VSS),.VDD(VDD),.Y(g17062),.A(I18154));
  NOT NOT1_5464(.VSS(VSS),.VDD(VDD),.Y(g20005),.A(g17433));
  NOT NOT1_5465(.VSS(VSS),.VDD(VDD),.Y(g13485),.A(g10476));
  NOT NOT1_5466(.VSS(VSS),.VDD(VDD),.Y(g20328),.A(g15867));
  NOT NOT1_5467(.VSS(VSS),.VDD(VDD),.Y(g32595),.A(g30825));
  NOT NOT1_5468(.VSS(VSS),.VDD(VDD),.Y(g32467),.A(g31194));
  NOT NOT1_5469(.VSS(VSS),.VDD(VDD),.Y(g32494),.A(g30825));
  NOT NOT1_5470(.VSS(VSS),.VDD(VDD),.Y(g19902),.A(g17200));
  NOT NOT1_5471(.VSS(VSS),.VDD(VDD),.Y(g24005),.A(I23149));
  NOT NOT1_5472(.VSS(VSS),.VDD(VDD),.Y(g17509),.A(I18446));
  NOT NOT1_5473(.VSS(VSS),.VDD(VDD),.Y(g14034),.A(g11048));
  NOT NOT1_5474(.VSS(VSS),.VDD(VDD),.Y(g19957),.A(g16540));
  NOT NOT1_5475(.VSS(VSS),.VDD(VDD),.Y(g16816),.A(I18028));
  NOT NOT1_5476(.VSS(VSS),.VDD(VDD),.Y(g20538),.A(g15348));
  NOT NOT1_5477(.VSS(VSS),.VDD(VDD),.Y(g9688),.A(g113));
  NOT NOT1_5478(.VSS(VSS),.VDD(VDD),.Y(g28606),.A(g27762));
  NOT NOT1_5479(.VSS(VSS),.VDD(VDD),.Y(g6847),.A(g2283));
  NOT NOT1_5480(.VSS(VSS),.VDD(VDD),.Y(g13555),.A(g12692));
  NOT NOT1_5481(.VSS(VSS),.VDD(VDD),.Y(g18882),.A(I19674));
  NOT NOT1_5482(.VSS(VSS),.VDD(VDD),.Y(g32623),.A(g30735));
  NOT NOT1_5483(.VSS(VSS),.VDD(VDD),.Y(g18991),.A(g16136));
  NOT NOT1_5484(.VSS(VSS),.VDD(VDD),.Y(I28897),.A(g30155));
  NOT NOT1_5485(.VSS(VSS),.VDD(VDD),.Y(g19739),.A(g16931));
  NOT NOT1_5486(.VSS(VSS),.VDD(VDD),.Y(I25391),.A(g24483));
  NOT NOT1_5487(.VSS(VSS),.VDD(VDD),.Y(g9976),.A(g2537));
  NOT NOT1_5488(.VSS(VSS),.VDD(VDD),.Y(g17508),.A(I18443));
  NOT NOT1_5489(.VSS(VSS),.VDD(VDD),.Y(g29317),.A(I27677));
  NOT NOT1_5490(.VSS(VSS),.VDD(VDD),.Y(g10153),.A(g2417));
  NOT NOT1_5491(.VSS(VSS),.VDD(VDD),.Y(g23841),.A(g19074));
  NOT NOT1_5492(.VSS(VSS),.VDD(VDD),.Y(I22096),.A(g19890));
  NOT NOT1_5493(.VSS(VSS),.VDD(VDD),.Y(g23992),.A(g19210));
  NOT NOT1_5494(.VSS(VSS),.VDD(VDD),.Y(g32782),.A(g30735));
  NOT NOT1_5495(.VSS(VSS),.VDD(VDD),.Y(g23391),.A(g20645));
  NOT NOT1_5496(.VSS(VSS),.VDD(VDD),.Y(g19146),.A(g15574));
  NOT NOT1_5497(.VSS(VSS),.VDD(VDD),.Y(g19738),.A(g15992));
  NOT NOT1_5498(.VSS(VSS),.VDD(VDD),.Y(g33080),.A(I30644));
  NOT NOT1_5499(.VSS(VSS),.VDD(VDD),.Y(g21510),.A(g15647));
  NOT NOT1_5500(.VSS(VSS),.VDD(VDD),.Y(g23510),.A(g18833));
  NOT NOT1_5501(.VSS(VSS),.VDD(VDD),.Y(g10409),.A(g7087));
  NOT NOT1_5502(.VSS(VSS),.VDD(VDD),.Y(g16752),.A(I17976));
  NOT NOT1_5503(.VSS(VSS),.VDD(VDD),.Y(I21757),.A(g21308));
  NOT NOT1_5504(.VSS(VSS),.VDD(VDD),.Y(I33218),.A(g34955));
  NOT NOT1_5505(.VSS(VSS),.VDD(VDD),.Y(I25579),.A(g25297));
  NOT NOT1_5506(.VSS(VSS),.VDD(VDD),.Y(g16954),.A(I18104));
  NOT NOT1_5507(.VSS(VSS),.VDD(VDD),.Y(g29129),.A(g27858));
  NOT NOT1_5508(.VSS(VSS),.VDD(VDD),.Y(g22213),.A(g19147));
  NOT NOT1_5509(.VSS(VSS),.VDD(VDD),.Y(g19699),.A(I20116));
  NOT NOT1_5510(.VSS(VSS),.VDD(VDD),.Y(g8504),.A(g3451));
  NOT NOT1_5511(.VSS(VSS),.VDD(VDD),.Y(g34511),.A(g34419));
  NOT NOT1_5512(.VSS(VSS),.VDD(VDD),.Y(g10136),.A(g6113));
  NOT NOT1_5513(.VSS(VSS),.VDD(VDD),.Y(g16643),.A(I17839));
  NOT NOT1_5514(.VSS(VSS),.VDD(VDD),.Y(g10408),.A(g7049));
  NOT NOT1_5515(.VSS(VSS),.VDD(VDD),.Y(g9000),.A(g632));
  NOT NOT1_5516(.VSS(VSS),.VDD(VDD),.Y(g32822),.A(g30937));
  NOT NOT1_5517(.VSS(VSS),.VDD(VDD),.Y(g13074),.A(I15702));
  NOT NOT1_5518(.VSS(VSS),.VDD(VDD),.Y(I24191),.A(g22360));
  NOT NOT1_5519(.VSS(VSS),.VDD(VDD),.Y(g29128),.A(g27800));
  NOT NOT1_5520(.VSS(VSS),.VDD(VDD),.Y(g14635),.A(I16741));
  NOT NOT1_5521(.VSS(VSS),.VDD(VDD),.Y(I12227),.A(g34));
  NOT NOT1_5522(.VSS(VSS),.VDD(VDD),.Y(g13239),.A(g10632));
  NOT NOT1_5523(.VSS(VSS),.VDD(VDD),.Y(g19698),.A(g16971));
  NOT NOT1_5524(.VSS(VSS),.VDD(VDD),.Y(g9326),.A(g6203));
  NOT NOT1_5525(.VSS(VSS),.VDD(VDD),.Y(I15238),.A(g6351));
  NOT NOT1_5526(.VSS(VSS),.VDD(VDD),.Y(g12951),.A(I15569));
  NOT NOT1_5527(.VSS(VSS),.VDD(VDD),.Y(g25157),.A(g22498));
  NOT NOT1_5528(.VSS(VSS),.VDD(VDD),.Y(g23578),.A(I22725));
  NOT NOT1_5529(.VSS(VSS),.VDD(VDD),.Y(g8070),.A(g3518));
  NOT NOT1_5530(.VSS(VSS),.VDD(VDD),.Y(g13594),.A(g11012));
  NOT NOT1_5531(.VSS(VSS),.VDD(VDD),.Y(I16438),.A(g11165));
  NOT NOT1_5532(.VSS(VSS),.VDD(VDD),.Y(g23014),.A(g20391));
  NOT NOT1_5533(.VSS(VSS),.VDD(VDD),.Y(I25586),.A(g25537));
  NOT NOT1_5534(.VSS(VSS),.VDD(VDD),.Y(g8470),.A(I12605));
  NOT NOT1_5535(.VSS(VSS),.VDD(VDD),.Y(g20100),.A(I20369));
  NOT NOT1_5536(.VSS(VSS),.VDD(VDD),.Y(g7512),.A(g5283));
  NOT NOT1_5537(.VSS(VSS),.VDD(VDD),.Y(g34660),.A(g34473));
  NOT NOT1_5538(.VSS(VSS),.VDD(VDD),.Y(I30983),.A(g32433));
  NOT NOT1_5539(.VSS(VSS),.VDD(VDD),.Y(g9760),.A(g2315));
  NOT NOT1_5540(.VSS(VSS),.VDD(VDD),.Y(g20771),.A(g15171));
  NOT NOT1_5541(.VSS(VSS),.VDD(VDD),.Y(g22311),.A(g18935));
  NOT NOT1_5542(.VSS(VSS),.VDD(VDD),.Y(g24100),.A(g20857));
  NOT NOT1_5543(.VSS(VSS),.VDD(VDD),.Y(g26054),.A(g24804));
  NOT NOT1_5544(.VSS(VSS),.VDD(VDD),.Y(g7490),.A(g2629));
  NOT NOT1_5545(.VSS(VSS),.VDD(VDD),.Y(I15382),.A(g9071));
  NOT NOT1_5546(.VSS(VSS),.VDD(VDD),.Y(I14647),.A(g7717));
  NOT NOT1_5547(.VSS(VSS),.VDD(VDD),.Y(g25231),.A(g22228));
  NOT NOT1_5548(.VSS(VSS),.VDD(VDD),.Y(g7166),.A(g4311));
  NOT NOT1_5549(.VSS(VSS),.VDD(VDD),.Y(g20235),.A(g15277));
  NOT NOT1_5550(.VSS(VSS),.VDD(VDD),.Y(g19427),.A(g16292));
  NOT NOT1_5551(.VSS(VSS),.VDD(VDD),.Y(I26130),.A(g26510));
  NOT NOT1_5552(.VSS(VSS),.VDD(VDD),.Y(g11941),.A(I14761));
  NOT NOT1_5553(.VSS(VSS),.VDD(VDD),.Y(g19366),.A(g15885));
  NOT NOT1_5554(.VSS(VSS),.VDD(VDD),.Y(I17857),.A(g3969));
  NOT NOT1_5555(.VSS(VSS),.VDD(VDD),.Y(g32853),.A(g30673));
  NOT NOT1_5556(.VSS(VSS),.VDD(VDD),.Y(g24683),.A(g23112));
  NOT NOT1_5557(.VSS(VSS),.VDD(VDD),.Y(g33736),.A(I31597));
  NOT NOT1_5558(.VSS(VSS),.VDD(VDD),.Y(g11519),.A(g8481));
  NOT NOT1_5559(.VSS(VSS),.VDD(VDD),.Y(I14999),.A(g10030));
  NOT NOT1_5560(.VSS(VSS),.VDD(VDD),.Y(g16195),.A(g13437));
  NOT NOT1_5561(.VSS(VSS),.VDD(VDD),.Y(g34480),.A(I32535));
  NOT NOT1_5562(.VSS(VSS),.VDD(VDD),.Y(g16489),.A(I17699));
  NOT NOT1_5563(.VSS(VSS),.VDD(VDD),.Y(g34916),.A(I33140));
  NOT NOT1_5564(.VSS(VSS),.VDD(VDD),.Y(g13675),.A(g10556));
  NOT NOT1_5565(.VSS(VSS),.VDD(VDD),.Y(I20861),.A(g16960));
  NOT NOT1_5566(.VSS(VSS),.VDD(VDD),.Y(g32589),.A(g31070));
  NOT NOT1_5567(.VSS(VSS),.VDD(VDD),.Y(g7456),.A(g2495));
  NOT NOT1_5568(.VSS(VSS),.VDD(VDD),.Y(g15224),.A(I17101));
  NOT NOT1_5569(.VSS(VSS),.VDD(VDD),.Y(g7148),.A(I11835));
  NOT NOT1_5570(.VSS(VSS),.VDD(VDD),.Y(g6817),.A(g956));
  NOT NOT1_5571(.VSS(VSS),.VDD(VDD),.Y(g7649),.A(g1345));
  NOT NOT1_5572(.VSS(VSS),.VDD(VDD),.Y(g22592),.A(I21930));
  NOT NOT1_5573(.VSS(VSS),.VDD(VDD),.Y(g22756),.A(g20436));
  NOT NOT1_5574(.VSS(VSS),.VDD(VDD),.Y(g16525),.A(I17723));
  NOT NOT1_5575(.VSS(VSS),.VDD(VDD),.Y(g15571),.A(g13211));
  NOT NOT1_5576(.VSS(VSS),.VDD(VDD),.Y(g26942),.A(I25692));
  NOT NOT1_5577(.VSS(VSS),.VDD(VDD),.Y(g9924),.A(g5644));
  NOT NOT1_5578(.VSS(VSS),.VDD(VDD),.Y(g10474),.A(g8841));
  NOT NOT1_5579(.VSS(VSS),.VDD(VDD),.Y(g32588),.A(g30825));
  NOT NOT1_5580(.VSS(VSS),.VDD(VDD),.Y(g32524),.A(g31070));
  NOT NOT1_5581(.VSS(VSS),.VDD(VDD),.Y(g9220),.A(g843));
  NOT NOT1_5582(.VSS(VSS),.VDD(VDD),.Y(g31843),.A(g29385));
  NOT NOT1_5583(.VSS(VSS),.VDD(VDD),.Y(g32836),.A(g31021));
  NOT NOT1_5584(.VSS(VSS),.VDD(VDD),.Y(g33696),.A(I31535));
  NOT NOT1_5585(.VSS(VSS),.VDD(VDD),.Y(g30076),.A(g29085));
  NOT NOT1_5586(.VSS(VSS),.VDD(VDD),.Y(g30085),.A(g29082));
  NOT NOT1_5587(.VSS(VSS),.VDD(VDD),.Y(g7851),.A(g921));
  NOT NOT1_5588(.VSS(VSS),.VDD(VDD),.Y(I33075),.A(g34843));
  NOT NOT1_5589(.VSS(VSS),.VDD(VDD),.Y(g9779),.A(g5156));
  NOT NOT1_5590(.VSS(VSS),.VDD(VDD),.Y(g26655),.A(g25492));
  NOT NOT1_5591(.VSS(VSS),.VDD(VDD),.Y(g13637),.A(g10556));
  NOT NOT1_5592(.VSS(VSS),.VDD(VDD),.Y(g20515),.A(g15483));
  NOT NOT1_5593(.VSS(VSS),.VDD(VDD),.Y(g34307),.A(g34087));
  NOT NOT1_5594(.VSS(VSS),.VDD(VDD),.Y(g23041),.A(g19882));
  NOT NOT1_5595(.VSS(VSS),.VDD(VDD),.Y(I20388),.A(g17724));
  NOT NOT1_5596(.VSS(VSS),.VDD(VDD),.Y(g32477),.A(g31566));
  NOT NOT1_5597(.VSS(VSS),.VDD(VDD),.Y(I18360),.A(g1426));
  NOT NOT1_5598(.VSS(VSS),.VDD(VDD),.Y(g21275),.A(g15426));
  NOT NOT1_5599(.VSS(VSS),.VDD(VDD),.Y(g24515),.A(g22689));
  NOT NOT1_5600(.VSS(VSS),.VDD(VDD),.Y(I31494),.A(g33283));
  NOT NOT1_5601(.VSS(VSS),.VDD(VDD),.Y(g24991),.A(g22369));
  NOT NOT1_5602(.VSS(VSS),.VDD(VDD),.Y(I12120),.A(g632));
  NOT NOT1_5603(.VSS(VSS),.VDD(VDD),.Y(g10109),.A(g135));
  NOT NOT1_5604(.VSS(VSS),.VDD(VDD),.Y(g30054),.A(g29134));
  NOT NOT1_5605(.VSS(VSS),.VDD(VDD),.Y(g21430),.A(g15608));
  NOT NOT1_5606(.VSS(VSS),.VDD(VDD),.Y(g27163),.A(I25869));
  NOT NOT1_5607(.VSS(VSS),.VDD(VDD),.Y(g34596),.A(I32696));
  NOT NOT1_5608(.VSS(VSS),.VDD(VDD),.Y(g8406),.A(g232));
  NOT NOT1_5609(.VSS(VSS),.VDD(VDD),.Y(g17756),.A(g14858));
  NOT NOT1_5610(.VSS(VSS),.VDD(VDD),.Y(I27738),.A(g28140));
  NOT NOT1_5611(.VSS(VSS),.VDD(VDD),.Y(g23430),.A(I22547));
  NOT NOT1_5612(.VSS(VSS),.VDD(VDD),.Y(g23746),.A(g20902));
  NOT NOT1_5613(.VSS(VSS),.VDD(VDD),.Y(g23493),.A(g21611));
  NOT NOT1_5614(.VSS(VSS),.VDD(VDD),.Y(g7964),.A(g3155));
  NOT NOT1_5615(.VSS(VSS),.VDD(VDD),.Y(g7260),.A(I11908));
  NOT NOT1_5616(.VSS(VSS),.VDD(VDD),.Y(g8635),.A(g2783));
  NOT NOT1_5617(.VSS(VSS),.VDD(VDD),.Y(g24407),.A(g22594));
  NOT NOT1_5618(.VSS(VSS),.VDD(VDD),.Y(g34243),.A(I32228));
  NOT NOT1_5619(.VSS(VSS),.VDD(VDD),.Y(g29697),.A(g28336));
  NOT NOT1_5620(.VSS(VSS),.VDD(VDD),.Y(g9977),.A(g2667));
  NOT NOT1_5621(.VSS(VSS),.VDD(VDD),.Y(g19481),.A(g16349));
  NOT NOT1_5622(.VSS(VSS),.VDD(VDD),.Y(g10108),.A(g120));
  NOT NOT1_5623(.VSS(VSS),.VDD(VDD),.Y(I14932),.A(g9901));
  NOT NOT1_5624(.VSS(VSS),.VDD(VDD),.Y(g29995),.A(g28955));
  NOT NOT1_5625(.VSS(VSS),.VDD(VDD),.Y(I33037),.A(g34770));
  NOT NOT1_5626(.VSS(VSS),.VDD(VDD),.Y(g34431),.A(I32464));
  NOT NOT1_5627(.VSS(VSS),.VDD(VDD),.Y(g12012),.A(g9213));
  NOT NOT1_5628(.VSS(VSS),.VDD(VDD),.Y(g32118),.A(g31008));
  NOT NOT1_5629(.VSS(VSS),.VDD(VDD),.Y(g15816),.A(I17314));
  NOT NOT1_5630(.VSS(VSS),.VDD(VDD),.Y(g8766),.A(g572));
  NOT NOT1_5631(.VSS(VSS),.VDD(VDD),.Y(g18940),.A(I19719));
  NOT NOT1_5632(.VSS(VSS),.VDD(VDD),.Y(g8087),.A(g1157));
  NOT NOT1_5633(.VSS(VSS),.VDD(VDD),.Y(I31782),.A(g33219));
  NOT NOT1_5634(.VSS(VSS),.VDD(VDD),.Y(g32864),.A(g30937));
  NOT NOT1_5635(.VSS(VSS),.VDD(VDD),.Y(g23237),.A(g20924));
  NOT NOT1_5636(.VSS(VSS),.VDD(VDD),.Y(I19734),.A(g17725));
  NOT NOT1_5637(.VSS(VSS),.VDD(VDD),.Y(g7063),.A(g4831));
  NOT NOT1_5638(.VSS(VSS),.VDD(VDD),.Y(g10606),.A(g10233));
  NOT NOT1_5639(.VSS(VSS),.VDD(VDD),.Y(g21340),.A(I21074));
  NOT NOT1_5640(.VSS(VSS),.VDD(VDD),.Y(g32749),.A(g31021));
  NOT NOT1_5641(.VSS(VSS),.VDD(VDD),.Y(g32616),.A(g30735));
  NOT NOT1_5642(.VSS(VSS),.VDD(VDD),.Y(g23340),.A(g21070));
  NOT NOT1_5643(.VSS(VSS),.VDD(VDD),.Y(g23983),.A(g19210));
  NOT NOT1_5644(.VSS(VSS),.VDD(VDD),.Y(I22128),.A(g19968));
  NOT NOT1_5645(.VSS(VSS),.VDD(VDD),.Y(g34773),.A(I32963));
  NOT NOT1_5646(.VSS(VSS),.VDD(VDD),.Y(g9051),.A(g1426));
  NOT NOT1_5647(.VSS(VSS),.VDD(VDD),.Y(g23684),.A(I22819));
  NOT NOT1_5648(.VSS(VSS),.VDD(VDD),.Y(g25480),.A(g22228));
  NOT NOT1_5649(.VSS(VSS),.VDD(VDD),.Y(g34942),.A(g34928));
  NOT NOT1_5650(.VSS(VSS),.VDD(VDD),.Y(g32748),.A(g31710));
  NOT NOT1_5651(.VSS(VSS),.VDD(VDD),.Y(I15577),.A(g10430));
  NOT NOT1_5652(.VSS(VSS),.VDD(VDD),.Y(g8748),.A(g776));
  NOT NOT1_5653(.VSS(VSS),.VDD(VDD),.Y(g11215),.A(g8285));
  NOT NOT1_5654(.VSS(VSS),.VDD(VDD),.Y(g19127),.A(I19775));
  NOT NOT1_5655(.VSS(VSS),.VDD(VDD),.Y(g9451),.A(g5873));
  NOT NOT1_5656(.VSS(VSS),.VDD(VDD),.Y(g28326),.A(g27414));
  NOT NOT1_5657(.VSS(VSS),.VDD(VDD),.Y(I32991),.A(g34759));
  NOT NOT1_5658(.VSS(VSS),.VDD(VDD),.Y(I14505),.A(g10140));
  NOT NOT1_5659(.VSS(VSS),.VDD(VDD),.Y(I33155),.A(g34897));
  NOT NOT1_5660(.VSS(VSS),.VDD(VDD),.Y(g13215),.A(g10909));
  NOT NOT1_5661(.VSS(VSS),.VDD(VDD),.Y(g26131),.A(I25161));
  NOT NOT1_5662(.VSS(VSS),.VDD(VDD),.Y(g34156),.A(g33907));
  NOT NOT1_5663(.VSS(VSS),.VDD(VDD),.Y(g13729),.A(g10951));
  NOT NOT1_5664(.VSS(VSS),.VDD(VDD),.Y(g25550),.A(g22763));
  NOT NOT1_5665(.VSS(VSS),.VDD(VDD),.Y(g20441),.A(g17873));
  NOT NOT1_5666(.VSS(VSS),.VDD(VDD),.Y(g20584),.A(g17873));
  NOT NOT1_5667(.VSS(VSS),.VDD(VDD),.Y(g32704),.A(g31070));
  NOT NOT1_5668(.VSS(VSS),.VDD(VDD),.Y(I21047),.A(g17429));
  NOT NOT1_5669(.VSS(VSS),.VDD(VDD),.Y(g10381),.A(g6957));
  NOT NOT1_5670(.VSS(VSS),.VDD(VDD),.Y(g28040),.A(g26365));
  NOT NOT1_5671(.VSS(VSS),.VDD(VDD),.Y(g33708),.A(I31555));
  NOT NOT1_5672(.VSS(VSS),.VDD(VDD),.Y(I33170),.A(g34890));
  NOT NOT1_5673(.VSS(VSS),.VDD(VDD),.Y(g19490),.A(g16489));
  NOT NOT1_5674(.VSS(VSS),.VDD(VDD),.Y(g25287),.A(g22228));
  NOT NOT1_5675(.VSS(VSS),.VDD(VDD),.Y(g34670),.A(I32794));
  NOT NOT1_5676(.VSS(VSS),.VDD(VDD),.Y(I29939),.A(g31667));
  NOT NOT1_5677(.VSS(VSS),.VDD(VDD),.Y(g9999),.A(g6109));
  NOT NOT1_5678(.VSS(VSS),.VDD(VDD),.Y(I17128),.A(g13835));
  NOT NOT1_5679(.VSS(VSS),.VDD(VDD),.Y(g23517),.A(g21070));
  NOT NOT1_5680(.VSS(VSS),.VDD(VDD),.Y(g33258),.A(g32296));
  NOT NOT1_5681(.VSS(VSS),.VDD(VDD),.Y(g32809),.A(g31327));
  NOT NOT1_5682(.VSS(VSS),.VDD(VDD),.Y(g32900),.A(g30937));
  NOT NOT1_5683(.VSS(VSS),.VDD(VDD),.Y(g25307),.A(g22763));
  NOT NOT1_5684(.VSS(VSS),.VDD(VDD),.Y(g32466),.A(g31070));
  NOT NOT1_5685(.VSS(VSS),.VDD(VDD),.Y(g7118),.A(g832));
  NOT NOT1_5686(.VSS(VSS),.VDD(VDD),.Y(g7619),.A(g1296));
  NOT NOT1_5687(.VSS(VSS),.VDD(VDD),.Y(g16124),.A(g13555));
  NOT NOT1_5688(.VSS(VSS),.VDD(VDD),.Y(I19487),.A(g15125));
  NOT NOT1_5689(.VSS(VSS),.VDD(VDD),.Y(g19376),.A(g17509));
  NOT NOT1_5690(.VSS(VSS),.VDD(VDD),.Y(g19385),.A(g16326));
  NOT NOT1_5691(.VSS(VSS),.VDD(VDD),.Y(I17626),.A(g14582));
  NOT NOT1_5692(.VSS(VSS),.VDD(VDD),.Y(g17413),.A(I18350));
  NOT NOT1_5693(.VSS(VSS),.VDD(VDD),.Y(g9103),.A(g5774));
  NOT NOT1_5694(.VSS(VSS),.VDD(VDD),.Y(g32808),.A(g30937));
  NOT NOT1_5695(.VSS(VSS),.VDD(VDD),.Y(I26952),.A(g27972));
  NOT NOT1_5696(.VSS(VSS),.VDD(VDD),.Y(g24759),.A(g23003));
  NOT NOT1_5697(.VSS(VSS),.VDD(VDD),.Y(I18071),.A(g13680));
  NOT NOT1_5698(.VSS(VSS),.VDD(VDD),.Y(g19980),.A(g17226));
  NOT NOT1_5699(.VSS(VSS),.VDD(VDD),.Y(g25243),.A(g22763));
  NOT NOT1_5700(.VSS(VSS),.VDD(VDD),.Y(g34839),.A(I33053));
  NOT NOT1_5701(.VSS(VSS),.VDD(VDD),.Y(g17691),.A(I18674));
  NOT NOT1_5702(.VSS(VSS),.VDD(VDD),.Y(g20114),.A(I20385));
  NOT NOT1_5703(.VSS(VSS),.VDD(VDD),.Y(g16686),.A(I17892));
  NOT NOT1_5704(.VSS(VSS),.VDD(VDD),.Y(g34930),.A(I33182));
  NOT NOT1_5705(.VSS(VSS),.VDD(VDD),.Y(g11349),.A(I14365));
  NOT NOT1_5706(.VSS(VSS),.VDD(VDD),.Y(g34993),.A(I33279));
  NOT NOT1_5707(.VSS(VSS),.VDD(VDD),.Y(g12946),.A(I15564));
  NOT NOT1_5708(.VSS(VSS),.VDD(VDD),.Y(g15842),.A(g13469));
  NOT NOT1_5709(.VSS(VSS),.VDD(VDD),.Y(g32560),.A(g31070));
  NOT NOT1_5710(.VSS(VSS),.VDD(VDD),.Y(g20435),.A(g15348));
  NOT NOT1_5711(.VSS(VSS),.VDD(VDD),.Y(g8373),.A(g2485));
  NOT NOT1_5712(.VSS(VSS),.VDD(VDD),.Y(I15906),.A(g10430));
  NOT NOT1_5713(.VSS(VSS),.VDD(VDD),.Y(g24114),.A(g20720));
  NOT NOT1_5714(.VSS(VSS),.VDD(VDD),.Y(g8091),.A(g1579));
  NOT NOT1_5715(.VSS(VSS),.VDD(VDD),.Y(I33167),.A(g34890));
  NOT NOT1_5716(.VSS(VSS),.VDD(VDD),.Y(g6772),.A(I11629));
  NOT NOT1_5717(.VSS(VSS),.VDD(VDD),.Y(g29498),.A(I27784));
  NOT NOT1_5718(.VSS(VSS),.VDD(VDD),.Y(g24082),.A(g19890));
  NOT NOT1_5719(.VSS(VSS),.VDD(VDD),.Y(I15284),.A(g6697));
  NOT NOT1_5720(.VSS(VSS),.VDD(VDD),.Y(g16030),.A(g13570));
  NOT NOT1_5721(.VSS(VSS),.VDD(VDD),.Y(g7393),.A(g5320));
  NOT NOT1_5722(.VSS(VSS),.VDD(VDD),.Y(g13906),.A(I16201));
  NOT NOT1_5723(.VSS(VSS),.VDD(VDD),.Y(g10390),.A(g6987));
  NOT NOT1_5724(.VSS(VSS),.VDD(VDD),.Y(g21362),.A(g17873));
  NOT NOT1_5725(.VSS(VSS),.VDD(VDD),.Y(g24107),.A(g20857));
  NOT NOT1_5726(.VSS(VSS),.VDD(VDD),.Y(g32642),.A(g31542));
  NOT NOT1_5727(.VSS(VSS),.VDD(VDD),.Y(g9732),.A(g5481));
  NOT NOT1_5728(.VSS(VSS),.VDD(VDD),.Y(g23362),.A(I22467));
  NOT NOT1_5729(.VSS(VSS),.VDD(VDD),.Y(g34131),.A(I32074));
  NOT NOT1_5730(.VSS(VSS),.VDD(VDD),.Y(g29056),.A(g27800));
  NOT NOT1_5731(.VSS(VSS),.VDD(VDD),.Y(g22928),.A(I22131));
  NOT NOT1_5732(.VSS(VSS),.VDD(VDD),.Y(g9753),.A(g1890));
  NOT NOT1_5733(.VSS(VSS),.VDD(VDD),.Y(I26516),.A(g26824));
  NOT NOT1_5734(.VSS(VSS),.VDD(VDD),.Y(g23523),.A(g21514));
  NOT NOT1_5735(.VSS(VSS),.VDD(VDD),.Y(g31810),.A(g29385));
  NOT NOT1_5736(.VSS(VSS),.VDD(VDD),.Y(g8283),.A(I12493));
  NOT NOT1_5737(.VSS(VSS),.VDD(VDD),.Y(g25773),.A(g24453));
  NOT NOT1_5738(.VSS(VSS),.VDD(VDD),.Y(I27481),.A(g27928));
  NOT NOT1_5739(.VSS(VSS),.VDD(VDD),.Y(g18833),.A(I19661));
  NOT NOT1_5740(.VSS(VSS),.VDD(VDD),.Y(g31657),.A(I29239));
  NOT NOT1_5741(.VSS(VSS),.VDD(VDD),.Y(g7971),.A(g4818));
  NOT NOT1_5742(.VSS(VSS),.VDD(VDD),.Y(g13304),.A(I15872));
  NOT NOT1_5743(.VSS(VSS),.VDD(VDD),.Y(I20447),.A(g16244));
  NOT NOT1_5744(.VSS(VSS),.VDD(VDD),.Y(I28582),.A(g30116));
  NOT NOT1_5745(.VSS(VSS),.VDD(VDD),.Y(I18825),.A(g6019));
  NOT NOT1_5746(.VSS(VSS),.VDD(VDD),.Y(I18370),.A(g14873));
  NOT NOT1_5747(.VSS(VSS),.VDD(VDD),.Y(g24744),.A(g22202));
  NOT NOT1_5748(.VSS(VSS),.VDD(VDD),.Y(I31477),.A(g33391));
  NOT NOT1_5749(.VSS(VSS),.VDD(VDD),.Y(g29080),.A(g27779));
  NOT NOT1_5750(.VSS(VSS),.VDD(VDD),.Y(g7686),.A(g4659));
  NOT NOT1_5751(.VSS(VSS),.VDD(VDD),.Y(g33375),.A(g32377));
  NOT NOT1_5752(.VSS(VSS),.VDD(VDD),.Y(g8407),.A(g1171));
  NOT NOT1_5753(.VSS(VSS),.VDD(VDD),.Y(g17929),.A(I18855));
  NOT NOT1_5754(.VSS(VSS),.VDD(VDD),.Y(g9072),.A(g2994));
  NOT NOT1_5755(.VSS(VSS),.VDD(VDD),.Y(g25156),.A(g22498));
  NOT NOT1_5756(.VSS(VSS),.VDD(VDD),.Y(I29218),.A(g30304));
  NOT NOT1_5757(.VSS(VSS),.VDD(VDD),.Y(g8920),.A(I12899));
  NOT NOT1_5758(.VSS(VSS),.VDD(VDD),.Y(g8059),.A(g3171));
  NOT NOT1_5759(.VSS(VSS),.VDD(VDD),.Y(g32733),.A(g31672));
  NOT NOT1_5760(.VSS(VSS),.VDD(VDD),.Y(I33119),.A(g34852));
  NOT NOT1_5761(.VSS(VSS),.VDD(VDD),.Y(g14192),.A(g11385));
  NOT NOT1_5762(.VSS(VSS),.VDD(VDD),.Y(I18858),.A(g13835));
  NOT NOT1_5763(.VSS(VSS),.VDD(VDD),.Y(g9472),.A(g6555));
  NOT NOT1_5764(.VSS(VSS),.VDD(VDD),.Y(g19931),.A(g17200));
  NOT NOT1_5765(.VSS(VSS),.VDD(VDD),.Y(g25180),.A(g23529));
  NOT NOT1_5766(.VSS(VSS),.VDD(VDD),.Y(g6856),.A(I11682));
  NOT NOT1_5767(.VSS(VSS),.VDD(VDD),.Y(I12572),.A(g51));
  NOT NOT1_5768(.VSS(VSS),.VDD(VDD),.Y(g15830),.A(g13432));
  NOT NOT1_5769(.VSS(VSS),.VDD(VDD),.Y(g17583),.A(g14968));
  NOT NOT1_5770(.VSS(VSS),.VDD(VDD),.Y(g8718),.A(g3333));
  NOT NOT1_5771(.VSS(VSS),.VDD(VDD),.Y(I18151),.A(g13144));
  NOT NOT1_5772(.VSS(VSS),.VDD(VDD),.Y(g34210),.A(I32173));
  NOT NOT1_5773(.VSS(VSS),.VDD(VDD),.Y(g32874),.A(g30673));
  NOT NOT1_5774(.VSS(VSS),.VDD(VDD),.Y(I28925),.A(g29987));
  NOT NOT1_5775(.VSS(VSS),.VDD(VDD),.Y(g9443),.A(g5489));
  NOT NOT1_5776(.VSS(VSS),.VDD(VDD),.Y(g21727),.A(I21300));
  NOT NOT1_5777(.VSS(VSS),.VDD(VDD),.Y(I22512),.A(g19389));
  NOT NOT1_5778(.VSS(VSS),.VDD(VDD),.Y(g20652),.A(I20744));
  NOT NOT1_5779(.VSS(VSS),.VDD(VDD),.Y(g28508),.A(I26989));
  NOT NOT1_5780(.VSS(VSS),.VDD(VDD),.Y(g32630),.A(g30735));
  NOT NOT1_5781(.VSS(VSS),.VDD(VDD),.Y(g7121),.A(I11820));
  NOT NOT1_5782(.VSS(VSS),.VDD(VDD),.Y(g23863),.A(g19210));
  NOT NOT1_5783(.VSS(VSS),.VDD(VDD),.Y(g32693),.A(g31579));
  NOT NOT1_5784(.VSS(VSS),.VDD(VDD),.Y(I31616),.A(g33219));
  NOT NOT1_5785(.VSS(VSS),.VDD(VDD),.Y(g21222),.A(g17430));
  NOT NOT1_5786(.VSS(VSS),.VDD(VDD),.Y(I23396),.A(g23427));
  NOT NOT1_5787(.VSS(VSS),.VDD(VDD),.Y(g7670),.A(g4104));
  NOT NOT1_5788(.VSS(VSS),.VDD(VDD),.Y(g23222),.A(g20785));
  NOT NOT1_5789(.VSS(VSS),.VDD(VDD),.Y(I18367),.A(g13010));
  NOT NOT1_5790(.VSS(VSS),.VDD(VDD),.Y(g26187),.A(I25190));
  NOT NOT1_5791(.VSS(VSS),.VDD(VDD),.Y(g29342),.A(g28188));
  NOT NOT1_5792(.VSS(VSS),.VDD(VDD),.Y(g9316),.A(g5742));
  NOT NOT1_5793(.VSS(VSS),.VDD(VDD),.Y(g25930),.A(I25028));
  NOT NOT1_5794(.VSS(VSS),.VDD(VDD),.Y(g7625),.A(I12109));
  NOT NOT1_5795(.VSS(VSS),.VDD(VDD),.Y(g32665),.A(g31579));
  NOT NOT1_5796(.VSS(VSS),.VDD(VDD),.Y(I31748),.A(g33228));
  NOT NOT1_5797(.VSS(VSS),.VDD(VDD),.Y(I13473),.A(g4157));
  NOT NOT1_5798(.VSS(VSS),.VDD(VDD),.Y(g19520),.A(g16826));
  NOT NOT1_5799(.VSS(VSS),.VDD(VDD),.Y(g6992),.A(g4899));
  NOT NOT1_5800(.VSS(VSS),.VDD(VDD),.Y(g12760),.A(g10272));
  NOT NOT1_5801(.VSS(VSS),.VDD(VDD),.Y(g9434),.A(g5385));
  NOT NOT1_5802(.VSS(VSS),.VDD(VDD),.Y(g13138),.A(I15765));
  NOT NOT1_5803(.VSS(VSS),.VDD(VDD),.Y(g17787),.A(I18795));
  NOT NOT1_5804(.VSS(VSS),.VDD(VDD),.Y(g7232),.A(g4411));
  NOT NOT1_5805(.VSS(VSS),.VDD(VDD),.Y(g10553),.A(g8971));
  NOT NOT1_5806(.VSS(VSS),.VDD(VDD),.Y(g25838),.A(g25250));
  NOT NOT1_5807(.VSS(VSS),.VDD(VDD),.Y(I27784),.A(g29013));
  NOT NOT1_5808(.VSS(VSS),.VDD(VDD),.Y(I15636),.A(g12075));
  NOT NOT1_5809(.VSS(VSS),.VDD(VDD),.Y(I33276),.A(g34985));
  NOT NOT1_5810(.VSS(VSS),.VDD(VDD),.Y(I33285),.A(g34988));
  NOT NOT1_5811(.VSS(VSS),.VDD(VDD),.Y(g18947),.A(g16136));
  NOT NOT1_5812(.VSS(VSS),.VDD(VDD),.Y(I27385),.A(g27438));
  NOT NOT1_5813(.VSS(VSS),.VDD(VDD),.Y(g30039),.A(g29134));
  NOT NOT1_5814(.VSS(VSS),.VDD(VDD),.Y(g30306),.A(g28796));
  NOT NOT1_5815(.VSS(VSS),.VDD(VDD),.Y(g25131),.A(g23699));
  NOT NOT1_5816(.VSS(VSS),.VDD(VDD),.Y(I33053),.A(g34778));
  NOT NOT1_5817(.VSS(VSS),.VDD(VDD),.Y(g15705),.A(g13217));
  NOT NOT1_5818(.VSS(VSS),.VDD(VDD),.Y(g26937),.A(I25683));
  NOT NOT1_5819(.VSS(VSS),.VDD(VDD),.Y(g17302),.A(I18285));
  NOT NOT1_5820(.VSS(VSS),.VDD(VDD),.Y(g32892),.A(g31021));
  NOT NOT1_5821(.VSS(VSS),.VDD(VDD),.Y(g23347),.A(I22444));
  NOT NOT1_5822(.VSS(VSS),.VDD(VDD),.Y(g24135),.A(g20720));
  NOT NOT1_5823(.VSS(VSS),.VDD(VDD),.Y(g32476),.A(g30673));
  NOT NOT1_5824(.VSS(VSS),.VDD(VDD),.Y(g32485),.A(g31376));
  NOT NOT1_5825(.VSS(VSS),.VDD(VDD),.Y(g33459),.A(I30995));
  NOT NOT1_5826(.VSS(VSS),.VDD(VDD),.Y(I31466),.A(g33318));
  NOT NOT1_5827(.VSS(VSS),.VDD(VDD),.Y(g7909),.A(g936));
  NOT NOT1_5828(.VSS(VSS),.VDD(VDD),.Y(g30038),.A(g29097));
  NOT NOT1_5829(.VSS(VSS),.VDD(VDD),.Y(g23253),.A(g21037));
  NOT NOT1_5830(.VSS(VSS),.VDD(VDD),.Y(I12103),.A(g572));
  NOT NOT1_5831(.VSS(VSS),.VDD(VDD),.Y(g11852),.A(I14668));
  NOT NOT1_5832(.VSS(VSS),.VDD(VDD),.Y(g17743),.A(I18734));
  NOT NOT1_5833(.VSS(VSS),.VDD(VDD),.Y(g9681),.A(g5798));
  NOT NOT1_5834(.VSS(VSS),.VDD(VDD),.Y(I22499),.A(g21160));
  NOT NOT1_5835(.VSS(VSS),.VDD(VDD),.Y(g10040),.A(g2652));
  NOT NOT1_5836(.VSS(VSS),.VDD(VDD),.Y(I22316),.A(g19361));
  NOT NOT1_5837(.VSS(VSS),.VDD(VDD),.Y(g32555),.A(g30673));
  NOT NOT1_5838(.VSS(VSS),.VDD(VDD),.Y(I18446),.A(g13028));
  NOT NOT1_5839(.VSS(VSS),.VDD(VDD),.Y(g14536),.A(I16651));
  NOT NOT1_5840(.VSS(VSS),.VDD(VDD),.Y(g19860),.A(g17226));
  NOT NOT1_5841(.VSS(VSS),.VDD(VDD),.Y(g33458),.A(I30992));
  NOT NOT1_5842(.VSS(VSS),.VDD(VDD),.Y(g7519),.A(g1157));
  NOT NOT1_5843(.VSS(VSS),.VDD(VDD),.Y(g24361),.A(g22885));
  NOT NOT1_5844(.VSS(VSS),.VDD(VDD),.Y(g11963),.A(g9153));
  NOT NOT1_5845(.VSS(VSS),.VDD(VDD),.Y(g25557),.A(g22763));
  NOT NOT1_5846(.VSS(VSS),.VDD(VDD),.Y(g32570),.A(g31554));
  NOT NOT1_5847(.VSS(VSS),.VDD(VDD),.Y(g32712),.A(g30614));
  NOT NOT1_5848(.VSS(VSS),.VDD(VDD),.Y(g25210),.A(g23802));
  NOT NOT1_5849(.VSS(VSS),.VDD(VDD),.Y(g32914),.A(g31672));
  NOT NOT1_5850(.VSS(VSS),.VDD(VDD),.Y(I25351),.A(g24466));
  NOT NOT1_5851(.VSS(VSS),.VDD(VDD),.Y(g9914),.A(g2533));
  NOT NOT1_5852(.VSS(VSS),.VDD(VDD),.Y(I20355),.A(g17613));
  NOT NOT1_5853(.VSS(VSS),.VDD(VDD),.Y(g33918),.A(I31782));
  NOT NOT1_5854(.VSS(VSS),.VDD(VDD),.Y(g23236),.A(g20785));
  NOT NOT1_5855(.VSS(VSS),.VDD(VDD),.Y(g20500),.A(g17873));
  NOT NOT1_5856(.VSS(VSS),.VDD(VDD),.Y(g10621),.A(g7567));
  NOT NOT1_5857(.VSS(VSS),.VDD(VDD),.Y(g34677),.A(I32815));
  NOT NOT1_5858(.VSS(VSS),.VDD(VDD),.Y(g29365),.A(g29067));
  NOT NOT1_5859(.VSS(VSS),.VDD(VDD),.Y(g14252),.A(I16438));
  NOT NOT1_5860(.VSS(VSS),.VDD(VDD),.Y(I22989),.A(g21175));
  NOT NOT1_5861(.VSS(VSS),.VDD(VDD),.Y(g13664),.A(g11252));
  NOT NOT1_5862(.VSS(VSS),.VDD(VDD),.Y(g20049),.A(I20318));
  NOT NOT1_5863(.VSS(VSS),.VDD(VDD),.Y(g23952),.A(g19277));
  NOT NOT1_5864(.VSS(VSS),.VDD(VDD),.Y(g23351),.A(g20924));
  NOT NOT1_5865(.VSS(VSS),.VDD(VDD),.Y(g32907),.A(g30937));
  NOT NOT1_5866(.VSS(VSS),.VDD(VDD),.Y(I31642),.A(g33204));
  NOT NOT1_5867(.VSS(VSS),.VDD(VDD),.Y(g33079),.A(I30641));
  NOT NOT1_5868(.VSS(VSS),.VDD(VDD),.Y(g24049),.A(g20014));
  NOT NOT1_5869(.VSS(VSS),.VDD(VDD),.Y(I14896),.A(g9820));
  NOT NOT1_5870(.VSS(VSS),.VDD(VDD),.Y(g29960),.A(g28885));
  NOT NOT1_5871(.VSS(VSS),.VDD(VDD),.Y(g21175),.A(I20951));
  NOT NOT1_5872(.VSS(VSS),.VDD(VDD),.Y(g22881),.A(I22096));
  NOT NOT1_5873(.VSS(VSS),.VDD(VDD),.Y(g23821),.A(g19210));
  NOT NOT1_5874(.VSS(VSS),.VDD(VDD),.Y(g10564),.A(g9462));
  NOT NOT1_5875(.VSS(VSS),.VDD(VDD),.Y(g15938),.A(I17401));
  NOT NOT1_5876(.VSS(VSS),.VDD(VDD),.Y(g16075),.A(g13597));
  NOT NOT1_5877(.VSS(VSS),.VDD(VDD),.Y(g9413),.A(g1744));
  NOT NOT1_5878(.VSS(VSS),.VDD(VDD),.Y(g19659),.A(g17062));
  NOT NOT1_5879(.VSS(VSS),.VDD(VDD),.Y(g14564),.A(I16679));
  NOT NOT1_5880(.VSS(VSS),.VDD(VDD),.Y(g24048),.A(g19968));
  NOT NOT1_5881(.VSS(VSS),.VDD(VDD),.Y(I11682),.A(g2756));
  NOT NOT1_5882(.VSS(VSS),.VDD(VDD),.Y(g11576),.A(g8542));
  NOT NOT1_5883(.VSS(VSS),.VDD(VDD),.Y(I33064),.A(g34784));
  NOT NOT1_5884(.VSS(VSS),.VDD(VDD),.Y(I25790),.A(g26424));
  NOT NOT1_5885(.VSS(VSS),.VDD(VDD),.Y(I17989),.A(g14173));
  NOT NOT1_5886(.VSS(VSS),.VDD(VDD),.Y(g20004),.A(g17249));
  NOT NOT1_5887(.VSS(VSS),.VDD(VDD),.Y(g13484),.A(g10981));
  NOT NOT1_5888(.VSS(VSS),.VDD(VDD),.Y(g32567),.A(g31070));
  NOT NOT1_5889(.VSS(VSS),.VDD(VDD),.Y(g32594),.A(g30735));
  NOT NOT1_5890(.VSS(VSS),.VDD(VDD),.Y(g19658),.A(g16987));
  NOT NOT1_5891(.VSS(VSS),.VDD(VDD),.Y(g23264),.A(g21037));
  NOT NOT1_5892(.VSS(VSS),.VDD(VDD),.Y(g25286),.A(g22228));
  NOT NOT1_5893(.VSS(VSS),.VDD(VDD),.Y(g16623),.A(g14127));
  NOT NOT1_5894(.VSS(VSS),.VDD(VDD),.Y(g10183),.A(g2595));
  NOT NOT1_5895(.VSS(VSS),.VDD(VDD),.Y(I15609),.A(g12013));
  NOT NOT1_5896(.VSS(VSS),.VDD(VDD),.Y(g7586),.A(I12056));
  NOT NOT1_5897(.VSS(VSS),.VDD(VDD),.Y(g23516),.A(g20924));
  NOT NOT1_5898(.VSS(VSS),.VDD(VDD),.Y(g25039),.A(g22498));
  NOT NOT1_5899(.VSS(VSS),.VDD(VDD),.Y(I28548),.A(g28147));
  NOT NOT1_5900(.VSS(VSS),.VDD(VDD),.Y(g10397),.A(g7018));
  NOT NOT1_5901(.VSS(VSS),.VDD(VDD),.Y(g6976),.A(I11750));
  NOT NOT1_5902(.VSS(VSS),.VDD(VDD),.Y(g14183),.A(g12381));
  NOT NOT1_5903(.VSS(VSS),.VDD(VDD),.Y(g14673),.A(I16770));
  NOT NOT1_5904(.VSS(VSS),.VDD(VDD),.Y(g11609),.A(g7660));
  NOT NOT1_5905(.VSS(VSS),.VDD(VDD),.Y(g9820),.A(g99));
  NOT NOT1_5906(.VSS(VSS),.VDD(VDD),.Y(g16782),.A(I18006));
  NOT NOT1_5907(.VSS(VSS),.VDD(VDD),.Y(g12903),.A(g10411));
  NOT NOT1_5908(.VSS(VSS),.VDD(VDD),.Y(g20613),.A(g15224));
  NOT NOT1_5909(.VSS(VSS),.VDD(VDD),.Y(I21787),.A(g19422));
  NOT NOT1_5910(.VSS(VSS),.VDD(VDD),.Y(I22461),.A(g21225));
  NOT NOT1_5911(.VSS(VSS),.VDD(VDD),.Y(g31817),.A(g29385));
  NOT NOT1_5912(.VSS(VSS),.VDD(VDD),.Y(g13312),.A(g11048));
  NOT NOT1_5913(.VSS(VSS),.VDD(VDD),.Y(I18301),.A(g12976));
  NOT NOT1_5914(.VSS(VSS),.VDD(VDD),.Y(g32941),.A(g30735));
  NOT NOT1_5915(.VSS(VSS),.VDD(VDD),.Y(g32382),.A(g31657));
  NOT NOT1_5916(.VSS(VSS),.VDD(VDD),.Y(g11608),.A(g7659));
  NOT NOT1_5917(.VSS(VSS),.VDD(VDD),.Y(g19644),.A(g17953));
  NOT NOT1_5918(.VSS(VSS),.VDD(VDD),.Y(g10509),.A(g10233));
  NOT NOT1_5919(.VSS(VSS),.VDD(VDD),.Y(I18120),.A(g13350));
  NOT NOT1_5920(.VSS(VSS),.VDD(VDD),.Y(g32519),.A(g30673));
  NOT NOT1_5921(.VSS(VSS),.VDD(VDD),.Y(I22031),.A(g21387));
  NOT NOT1_5922(.VSS(VSS),.VDD(VDD),.Y(I27546),.A(g29041));
  NOT NOT1_5923(.VSS(VSS),.VDD(VDD),.Y(g32185),.A(I29717));
  NOT NOT1_5924(.VSS(VSS),.VDD(VDD),.Y(g18421),.A(I19235));
  NOT NOT1_5925(.VSS(VSS),.VDD(VDD),.Y(g14509),.A(I16626));
  NOT NOT1_5926(.VSS(VSS),.VDD(VDD),.Y(I15921),.A(g12381));
  NOT NOT1_5927(.VSS(VSS),.VDD(VDD),.Y(g32675),.A(g31070));
  NOT NOT1_5928(.VSS(VSS),.VDD(VDD),.Y(g8388),.A(g3010));
  NOT NOT1_5929(.VSS(VSS),.VDD(VDD),.Y(I23357),.A(g23359));
  NOT NOT1_5930(.VSS(VSS),.VDD(VDD),.Y(g20273),.A(g17128));
  NOT NOT1_5931(.VSS(VSS),.VDD(VDD),.Y(g20106),.A(g17328));
  NOT NOT1_5932(.VSS(VSS),.VDD(VDD),.Y(g12563),.A(g9864));
  NOT NOT1_5933(.VSS(VSS),.VDD(VDD),.Y(g20605),.A(g17955));
  NOT NOT1_5934(.VSS(VSS),.VDD(VDD),.Y(g21422),.A(g15373));
  NOT NOT1_5935(.VSS(VSS),.VDD(VDD),.Y(I26409),.A(g26187));
  NOT NOT1_5936(.VSS(VSS),.VDD(VDD),.Y(g30217),.A(I28458));
  NOT NOT1_5937(.VSS(VSS),.VDD(VDD),.Y(g8216),.A(g3092));
  NOT NOT1_5938(.VSS(VSS),.VDD(VDD),.Y(g10851),.A(I14069));
  NOT NOT1_5939(.VSS(VSS),.VDD(VDD),.Y(I12089),.A(g744));
  NOT NOT1_5940(.VSS(VSS),.VDD(VDD),.Y(g10872),.A(g7567));
  NOT NOT1_5941(.VSS(VSS),.VDD(VDD),.Y(g9601),.A(g4005));
  NOT NOT1_5942(.VSS(VSS),.VDD(VDD),.Y(g23422),.A(g21611));
  NOT NOT1_5943(.VSS(VSS),.VDD(VDD),.Y(g32518),.A(g30614));
  NOT NOT1_5944(.VSS(VSS),.VDD(VDD),.Y(I16328),.A(g878));
  NOT NOT1_5945(.VSS(VSS),.VDD(VDD),.Y(g24106),.A(g19984));
  NOT NOT1_5946(.VSS(VSS),.VDD(VDD),.Y(g24605),.A(g23139));
  NOT NOT1_5947(.VSS(VSS),.VDD(VDD),.Y(I14050),.A(g9963));
  NOT NOT1_5948(.VSS(VSS),.VDD(VDD),.Y(g29043),.A(I27391));
  NOT NOT1_5949(.VSS(VSS),.VDD(VDD),.Y(I16538),.A(g10417));
  NOT NOT1_5950(.VSS(VSS),.VDD(VDD),.Y(g13745),.A(I16102));
  NOT NOT1_5951(.VSS(VSS),.VDD(VDD),.Y(g32637),.A(g30735));
  NOT NOT1_5952(.VSS(VSS),.VDD(VDD),.Y(g31656),.A(I29236));
  NOT NOT1_5953(.VSS(VSS),.VDD(VDD),.Y(I20318),.A(g16920));
  NOT NOT1_5954(.VSS(VSS),.VDD(VDD),.Y(g17249),.A(I18265));
  NOT NOT1_5955(.VSS(VSS),.VDD(VDD),.Y(I28002),.A(g28153));
  NOT NOT1_5956(.VSS(VSS),.VDD(VDD),.Y(g32935),.A(g31672));
  NOT NOT1_5957(.VSS(VSS),.VDD(VDD),.Y(g24463),.A(g23578));
  NOT NOT1_5958(.VSS(VSS),.VDD(VDD),.Y(I21769),.A(g19402));
  NOT NOT1_5959(.VSS(VSS),.VDD(VDD),.Y(I17650),.A(g13271));
  NOT NOT1_5960(.VSS(VSS),.VDD(VDD),.Y(I28128),.A(g28314));
  NOT NOT1_5961(.VSS(VSS),.VDD(VDD),.Y(g20033),.A(g16579));
  NOT NOT1_5962(.VSS(VSS),.VDD(VDD),.Y(g31823),.A(g29385));
  NOT NOT1_5963(.VSS(VSS),.VDD(VDD),.Y(I32613),.A(g34329));
  NOT NOT1_5964(.VSS(VSS),.VDD(VDD),.Y(g32883),.A(g30735));
  NOT NOT1_5965(.VSS(VSS),.VDD(VDD),.Y(g17248),.A(I18262));
  NOT NOT1_5966(.VSS(VSS),.VDD(VDD),.Y(I30641),.A(g32024));
  NOT NOT1_5967(.VSS(VSS),.VDD(VDD),.Y(I31555),.A(g33212));
  NOT NOT1_5968(.VSS(VSS),.VDD(VDD),.Y(I14742),.A(g9534));
  NOT NOT1_5969(.VSS(VSS),.VDD(VDD),.Y(g19411),.A(g16489));
  NOT NOT1_5970(.VSS(VSS),.VDD(VDD),.Y(g19527),.A(g16349));
  NOT NOT1_5971(.VSS(VSS),.VDD(VDD),.Y(g17710),.A(g14764));
  NOT NOT1_5972(.VSS(VSS),.VDD(VDD),.Y(g24033),.A(g19919));
  NOT NOT1_5973(.VSS(VSS),.VDD(VDD),.Y(I17198),.A(g13809));
  NOT NOT1_5974(.VSS(VSS),.VDD(VDD),.Y(g12845),.A(g10358));
  NOT NOT1_5975(.VSS(VSS),.VDD(VDD),.Y(g27990),.A(g26770));
  NOT NOT1_5976(.VSS(VSS),.VDD(VDD),.Y(g16853),.A(g13584));
  NOT NOT1_5977(.VSS(VSS),.VDD(VDD),.Y(I12497),.A(g49));
  NOT NOT1_5978(.VSS(VSS),.VDD(VDD),.Y(g23542),.A(g21514));
  NOT NOT1_5979(.VSS(VSS),.VDD(VDD),.Y(g9581),.A(g91));
  NOT NOT1_5980(.VSS(VSS),.VDD(VDD),.Y(g23021),.A(g20283));
  NOT NOT1_5981(.VSS(VSS),.VDD(VDD),.Y(g23453),.A(I22576));
  NOT NOT1_5982(.VSS(VSS),.VDD(VDD),.Y(g10213),.A(g6732));
  NOT NOT1_5983(.VSS(VSS),.VDD(VDD),.Y(I32947),.A(g34659));
  NOT NOT1_5984(.VSS(VSS),.VDD(VDD),.Y(g12899),.A(g10407));
  NOT NOT1_5985(.VSS(VSS),.VDD(VDD),.Y(g21726),.A(I21297));
  NOT NOT1_5986(.VSS(VSS),.VDD(VDD),.Y(g16589),.A(g14082));
  NOT NOT1_5987(.VSS(VSS),.VDD(VDD),.Y(g25169),.A(g22763));
  NOT NOT1_5988(.VSS(VSS),.VDD(VDD),.Y(g29955),.A(g28950));
  NOT NOT1_5989(.VSS(VSS),.VDD(VDD),.Y(g9060),.A(g3355));
  NOT NOT1_5990(.VSS(VSS),.VDD(VDD),.Y(I32106),.A(g33653));
  NOT NOT1_5991(.VSS(VSS),.VDD(VDD),.Y(g23913),.A(g19147));
  NOT NOT1_5992(.VSS(VSS),.VDD(VDD),.Y(g15915),.A(I17392));
  NOT NOT1_5993(.VSS(VSS),.VDD(VDD),.Y(g9460),.A(g6154));
  NOT NOT1_5994(.VSS(VSS),.VDD(VDD),.Y(g24795),.A(g23342));
  NOT NOT1_5995(.VSS(VSS),.VDD(VDD),.Y(g29970),.A(I28199));
  NOT NOT1_5996(.VSS(VSS),.VDD(VDD),.Y(g7659),.A(I12141));
  NOT NOT1_5997(.VSS(VSS),.VDD(VDD),.Y(g12898),.A(g10405));
  NOT NOT1_5998(.VSS(VSS),.VDD(VDD),.Y(g22647),.A(I21959));
  NOT NOT1_5999(.VSS(VSS),.VDD(VDD),.Y(g17778),.A(I18778));
  NOT NOT1_6000(.VSS(VSS),.VDD(VDD),.Y(g16588),.A(g13929));
  NOT NOT1_6001(.VSS(VSS),.VDD(VDD),.Y(g25168),.A(I24334));
  NOT NOT1_6002(.VSS(VSS),.VDD(VDD),.Y(g23614),.A(g20248));
  NOT NOT1_6003(.VSS(VSS),.VDD(VDD),.Y(g25410),.A(g22228));
  NOT NOT1_6004(.VSS(VSS),.VDD(VDD),.Y(g18829),.A(g15171));
  NOT NOT1_6005(.VSS(VSS),.VDD(VDD),.Y(I12987),.A(g12));
  NOT NOT1_6006(.VSS(VSS),.VDD(VDD),.Y(I15732),.A(g6692));
  NOT NOT1_6007(.VSS(VSS),.VDD(VDD),.Y(g8741),.A(g4821));
  NOT NOT1_6008(.VSS(VSS),.VDD(VDD),.Y(g10047),.A(g5421));
  NOT NOT1_6009(.VSS(VSS),.VDD(VDD),.Y(I32812),.A(g34588));
  NOT NOT1_6010(.VSS(VSS),.VDD(VDD),.Y(g19503),.A(g16349));
  NOT NOT1_6011(.VSS(VSS),.VDD(VDD),.Y(g29878),.A(g28421));
  NOT NOT1_6012(.VSS(VSS),.VDD(VDD),.Y(g15277),.A(I17104));
  NOT NOT1_6013(.VSS(VSS),.VDD(VDD),.Y(g21607),.A(g17873));
  NOT NOT1_6014(.VSS(VSS),.VDD(VDD),.Y(g22999),.A(g20453));
  NOT NOT1_6015(.VSS(VSS),.VDD(VDD),.Y(g23607),.A(g21611));
  NOT NOT1_6016(.VSS(VSS),.VDD(VDD),.Y(g21905),.A(I21486));
  NOT NOT1_6017(.VSS(VSS),.VDD(VDD),.Y(g14205),.A(g12381));
  NOT NOT1_6018(.VSS(VSS),.VDD(VDD),.Y(g26654),.A(g25275));
  NOT NOT1_6019(.VSS(VSS),.VDD(VDD),.Y(g20514),.A(g15348));
  NOT NOT1_6020(.VSS(VSS),.VDD(VDD),.Y(I25530),.A(g25222));
  NOT NOT1_6021(.VSS(VSS),.VDD(VDD),.Y(g32501),.A(g30825));
  NOT NOT1_6022(.VSS(VSS),.VDD(VDD),.Y(g32729),.A(g30937));
  NOT NOT1_6023(.VSS(VSS),.VDD(VDD),.Y(g18828),.A(g17955));
  NOT NOT1_6024(.VSS(VSS),.VDD(VDD),.Y(g31631),.A(I29221));
  NOT NOT1_6025(.VSS(VSS),.VDD(VDD),.Y(g10311),.A(g4633));
  NOT NOT1_6026(.VSS(VSS),.VDD(VDD),.Y(g23320),.A(I22419));
  NOT NOT1_6027(.VSS(VSS),.VDD(VDD),.Y(g23905),.A(g21514));
  NOT NOT1_6028(.VSS(VSS),.VDD(VDD),.Y(g9739),.A(g5752));
  NOT NOT1_6029(.VSS(VSS),.VDD(VDD),.Y(g32577),.A(g31554));
  NOT NOT1_6030(.VSS(VSS),.VDD(VDD),.Y(g33631),.A(I31459));
  NOT NOT1_6031(.VSS(VSS),.VDD(VDD),.Y(I14730),.A(g7717));
  NOT NOT1_6032(.VSS(VSS),.VDD(VDD),.Y(g18946),.A(g16100));
  NOT NOT1_6033(.VSS(VSS),.VDD(VDD),.Y(g29171),.A(g27937));
  NOT NOT1_6034(.VSS(VSS),.VDD(VDD),.Y(g21274),.A(g15373));
  NOT NOT1_6035(.VSS(VSS),.VDD(VDD),.Y(g14912),.A(I16917));
  NOT NOT1_6036(.VSS(VSS),.VDD(VDD),.Y(g30321),.A(I28572));
  NOT NOT1_6037(.VSS(VSS),.VDD(VDD),.Y(g23274),.A(g21070));
  NOT NOT1_6038(.VSS(VSS),.VDD(VDD),.Y(g20507),.A(g15509));
  NOT NOT1_6039(.VSS(VSS),.VDD(VDD),.Y(g23530),.A(g20248));
  NOT NOT1_6040(.VSS(VSS),.VDD(VDD),.Y(g22998),.A(g20391));
  NOT NOT1_6041(.VSS(VSS),.VDD(VDD),.Y(g27832),.A(I26409));
  NOT NOT1_6042(.VSS(VSS),.VDD(VDD),.Y(I32234),.A(g34126));
  NOT NOT1_6043(.VSS(VSS),.VDD(VDD),.Y(g34922),.A(I33158));
  NOT NOT1_6044(.VSS(VSS),.VDD(VDD),.Y(I24281),.A(g23440));
  NOT NOT1_6045(.VSS(VSS),.VDD(VDD),.Y(g26936),.A(I25680));
  NOT NOT1_6046(.VSS(VSS),.VDD(VDD),.Y(g15595),.A(I17173));
  NOT NOT1_6047(.VSS(VSS),.VDD(VDD),.Y(g32728),.A(g31021));
  NOT NOT1_6048(.VSS(VSS),.VDD(VDD),.Y(g21346),.A(g17821));
  NOT NOT1_6049(.VSS(VSS),.VDD(VDD),.Y(g25015),.A(g23662));
  NOT NOT1_6050(.VSS(VSS),.VDD(VDD),.Y(g6977),.A(I11753));
  NOT NOT1_6051(.VSS(VSS),.VDD(VDD),.Y(I20957),.A(g16228));
  NOT NOT1_6052(.VSS(VSS),.VDD(VDD),.Y(g19714),.A(g16821));
  NOT NOT1_6053(.VSS(VSS),.VDD(VDD),.Y(I13240),.A(g5794));
  NOT NOT1_6054(.VSS(VSS),.VDD(VDD),.Y(g7275),.A(g1728));
  NOT NOT1_6055(.VSS(VSS),.VDD(VDD),.Y(g22182),.A(I21766));
  NOT NOT1_6056(.VSS(VSS),.VDD(VDD),.Y(g29967),.A(g28946));
  NOT NOT1_6057(.VSS(VSS),.VDD(VDD),.Y(g29994),.A(g29049));
  NOT NOT1_6058(.VSS(VSS),.VDD(VDD),.Y(g34531),.A(I32594));
  NOT NOT1_6059(.VSS(VSS),.VDD(VDD),.Y(g9995),.A(g6035));
  NOT NOT1_6060(.VSS(VSS),.VDD(VDD),.Y(I12644),.A(g3689));
  NOT NOT1_6061(.VSS(VSS),.VDD(VDD),.Y(I11903),.A(g4414));
  NOT NOT1_6062(.VSS(VSS),.VDD(VDD),.Y(g23565),.A(g21562));
  NOT NOT1_6063(.VSS(VSS),.VDD(VDD),.Y(g10072),.A(g9));
  NOT NOT1_6064(.VSS(VSS),.VDD(VDD),.Y(g32438),.A(g30991));
  NOT NOT1_6065(.VSS(VSS),.VDD(VDD),.Y(I14690),.A(g9340));
  NOT NOT1_6066(.VSS(VSS),.VDD(VDD),.Y(g8883),.A(g4709));
  NOT NOT1_6067(.VSS(VSS),.VDD(VDD),.Y(g7615),.A(I12083));
  NOT NOT1_6068(.VSS(VSS),.VDD(VDD),.Y(g12440),.A(g9985));
  NOT NOT1_6069(.VSS(VSS),.VDD(VDD),.Y(g27573),.A(g26667));
  NOT NOT1_6070(.VSS(VSS),.VDD(VDD),.Y(I20562),.A(g16525));
  NOT NOT1_6071(.VSS(VSS),.VDD(VDD),.Y(g25556),.A(g22763));
  NOT NOT1_6072(.VSS(VSS),.VDD(VDD),.Y(g24163),.A(I23333));
  NOT NOT1_6073(.VSS(VSS),.VDD(VDD),.Y(I33176),.A(g34887));
  NOT NOT1_6074(.VSS(VSS),.VDD(VDD),.Y(g7174),.A(g6052));
  NOT NOT1_6075(.VSS(VSS),.VDD(VDD),.Y(g19979),.A(g17226));
  NOT NOT1_6076(.VSS(VSS),.VDD(VDD),.Y(g16748),.A(I17970));
  NOT NOT1_6077(.VSS(VSS),.VDD(VDD),.Y(g7374),.A(g2227));
  NOT NOT1_6078(.VSS(VSS),.VDD(VDD),.Y(g12861),.A(g10367));
  NOT NOT1_6079(.VSS(VSS),.VDD(VDD),.Y(g17651),.A(g14868));
  NOT NOT1_6080(.VSS(VSS),.VDD(VDD),.Y(g17672),.A(g14720));
  NOT NOT1_6081(.VSS(VSS),.VDD(VDD),.Y(g34676),.A(I32812));
  NOT NOT1_6082(.VSS(VSS),.VDD(VDD),.Y(g8217),.A(g3143));
  NOT NOT1_6083(.VSS(VSS),.VDD(VDD),.Y(I16515),.A(g12477));
  NOT NOT1_6084(.VSS(VSS),.VDD(VDD),.Y(I17471),.A(g13394));
  NOT NOT1_6085(.VSS(VSS),.VDD(VDD),.Y(g9390),.A(g5808));
  NOT NOT1_6086(.VSS(VSS),.VDD(VDD),.Y(g21292),.A(I21033));
  NOT NOT1_6087(.VSS(VSS),.VDD(VDD),.Y(g11214),.A(g9602));
  NOT NOT1_6088(.VSS(VSS),.VDD(VDD),.Y(g32906),.A(g31021));
  NOT NOT1_6089(.VSS(VSS),.VDD(VDD),.Y(g7985),.A(g3506));
  NOT NOT1_6090(.VSS(VSS),.VDD(VDD),.Y(g16285),.A(I17612));
  NOT NOT1_6091(.VSS(VSS),.VDD(VDD),.Y(g8466),.A(g1514));
  NOT NOT1_6092(.VSS(VSS),.VDD(VDD),.Y(I19762),.A(g15732));
  NOT NOT1_6093(.VSS(VSS),.VDD(VDD),.Y(g22449),.A(g19597));
  NOT NOT1_6094(.VSS(VSS),.VDD(VDD),.Y(g34654),.A(I32766));
  NOT NOT1_6095(.VSS(VSS),.VDD(VDD),.Y(g20541),.A(g17821));
  NOT NOT1_6096(.VSS(VSS),.VDD(VDD),.Y(I12855),.A(g4311));
  NOT NOT1_6097(.VSS(VSS),.VDD(VDD),.Y(g16305),.A(g13346));
  NOT NOT1_6098(.VSS(VSS),.VDD(VDD),.Y(g10350),.A(g6800));
  NOT NOT1_6099(.VSS(VSS),.VDD(VDD),.Y(g13329),.A(I15893));
  NOT NOT1_6100(.VSS(VSS),.VDD(VDD),.Y(g16053),.A(I17442));
  NOT NOT1_6101(.VSS(VSS),.VDD(VDD),.Y(g9501),.A(g5731));
  NOT NOT1_6102(.VSS(VSS),.VDD(VDD),.Y(g6999),.A(g86));
  NOT NOT1_6103(.VSS(VSS),.VDD(VDD),.Y(g16809),.A(g14387));
  NOT NOT1_6104(.VSS(VSS),.VDD(VDD),.Y(g21409),.A(g18008));
  NOT NOT1_6105(.VSS(VSS),.VDD(VDD),.Y(g22897),.A(g21024));
  NOT NOT1_6106(.VSS(VSS),.VDD(VDD),.Y(g7239),.A(g5033));
  NOT NOT1_6107(.VSS(VSS),.VDD(VDD),.Y(I12411),.A(g4809));
  NOT NOT1_6108(.VSS(VSS),.VDD(VDD),.Y(g23409),.A(g21514));
  NOT NOT1_6109(.VSS(VSS),.VDD(VDD),.Y(g8165),.A(g3530));
  NOT NOT1_6110(.VSS(VSS),.VDD(VDD),.Y(g32622),.A(g31376));
  NOT NOT1_6111(.VSS(VSS),.VDD(VDD),.Y(g8571),.A(g57));
  NOT NOT1_6112(.VSS(VSS),.VDD(VDD),.Y(g8365),.A(g2060));
  NOT NOT1_6113(.VSS(VSS),.VDD(VDD),.Y(I26381),.A(g26851));
  NOT NOT1_6114(.VSS(VSS),.VDD(VDD),.Y(g24789),.A(g23309));
  NOT NOT1_6115(.VSS(VSS),.VDD(VDD),.Y(g32566),.A(g30825));
  NOT NOT1_6116(.VSS(VSS),.VDD(VDD),.Y(g19741),.A(g16987));
  NOT NOT1_6117(.VSS(VSS),.VDD(VDD),.Y(I30537),.A(g32027));
  NOT NOT1_6118(.VSS(VSS),.VDD(VDD),.Y(g29079),.A(g27742));
  NOT NOT1_6119(.VSS(VSS),.VDD(VDD),.Y(g7380),.A(g2331));
  NOT NOT1_6120(.VSS(VSS),.VDD(VDD),.Y(g21408),.A(g15373));
  NOT NOT1_6121(.VSS(VSS),.VDD(VDD),.Y(g10152),.A(g2122));
  NOT NOT1_6122(.VSS(VSS),.VDD(VDD),.Y(g7591),.A(g6668));
  NOT NOT1_6123(.VSS(VSS),.VDD(VDD),.Y(g23408),.A(g21468));
  NOT NOT1_6124(.VSS(VSS),.VDD(VDD),.Y(g8055),.A(g1236));
  NOT NOT1_6125(.VSS(VSS),.VDD(VDD),.Y(g10396),.A(g6997));
  NOT NOT1_6126(.VSS(VSS),.VDD(VDD),.Y(g20325),.A(g15171));
  NOT NOT1_6127(.VSS(VSS),.VDD(VDD),.Y(g24359),.A(g22550));
  NOT NOT1_6128(.VSS(VSS),.VDD(VDD),.Y(g19067),.A(g15979));
  NOT NOT1_6129(.VSS(VSS),.VDD(VDD),.Y(g20920),.A(g15426));
  NOT NOT1_6130(.VSS(VSS),.VDD(VDD),.Y(g20535),.A(g17847));
  NOT NOT1_6131(.VSS(VSS),.VDD(VDD),.Y(I13990),.A(g7636));
  NOT NOT1_6132(.VSS(VSS),.VDD(VDD),.Y(g20434),.A(g18065));
  NOT NOT1_6133(.VSS(VSS),.VDD(VDD),.Y(g9704),.A(g2575));
  NOT NOT1_6134(.VSS(VSS),.VDD(VDD),.Y(g31816),.A(g29385));
  NOT NOT1_6135(.VSS(VSS),.VDD(VDD),.Y(g8133),.A(g4809));
  NOT NOT1_6136(.VSS(VSS),.VDD(VDD),.Y(g24920),.A(I24089));
  NOT NOT1_6137(.VSS(VSS),.VDD(VDD),.Y(g24535),.A(g22942));
  NOT NOT1_6138(.VSS(VSS),.VDD(VDD),.Y(I18376),.A(g14332));
  NOT NOT1_6139(.VSS(VSS),.VDD(VDD),.Y(g24358),.A(g22550));
  NOT NOT1_6140(.VSS(VSS),.VDD(VDD),.Y(I18297),.A(g1418));
  NOT NOT1_6141(.VSS(VSS),.VDD(VDD),.Y(I12503),.A(g215));
  NOT NOT1_6142(.VSS(VSS),.VDD(VDD),.Y(g17505),.A(g14899));
  NOT NOT1_6143(.VSS(VSS),.VDD(VDD),.Y(g17404),.A(I18337));
  NOT NOT1_6144(.VSS(VSS),.VDD(VDD),.Y(g10413),.A(g7110));
  NOT NOT1_6145(.VSS(VSS),.VDD(VDD),.Y(g8774),.A(g781));
  NOT NOT1_6146(.VSS(VSS),.VDD(VDD),.Y(g32653),.A(g30825));
  NOT NOT1_6147(.VSS(VSS),.VDD(VDD),.Y(g19801),.A(I20216));
  NOT NOT1_6148(.VSS(VSS),.VDD(VDD),.Y(I32473),.A(g34248));
  NOT NOT1_6149(.VSS(VSS),.VDD(VDD),.Y(g17717),.A(g14937));
  NOT NOT1_6150(.VSS(VSS),.VDD(VDD),.Y(I17879),.A(g14386));
  NOT NOT1_6151(.VSS(VSS),.VDD(VDD),.Y(g34423),.A(g34222));
  NOT NOT1_6152(.VSS(VSS),.VDD(VDD),.Y(g15588),.A(I17166));
  NOT NOT1_6153(.VSS(VSS),.VDD(VDD),.Y(I22886),.A(g18926));
  NOT NOT1_6154(.VSS(VSS),.VDD(VDD),.Y(g32138),.A(g31233));
  NOT NOT1_6155(.VSS(VSS),.VDD(VDD),.Y(I17970),.A(g4027));
  NOT NOT1_6156(.VSS(VSS),.VDD(VDD),.Y(I20895),.A(g16954));
  NOT NOT1_6157(.VSS(VSS),.VDD(VDD),.Y(g24121),.A(g20720));
  NOT NOT1_6158(.VSS(VSS),.VDD(VDD),.Y(I18888),.A(g16644));
  NOT NOT1_6159(.VSS(VSS),.VDD(VDD),.Y(g8396),.A(g3401));
  NOT NOT1_6160(.VSS(VSS),.VDD(VDD),.Y(g9250),.A(g1600));
  NOT NOT1_6161(.VSS(VSS),.VDD(VDD),.Y(g34587),.A(I32671));
  NOT NOT1_6162(.VSS(VSS),.VDD(VDD),.Y(I13718),.A(g890));
  NOT NOT1_6163(.VSS(VSS),.VDD(VDD),.Y(g12997),.A(g11826));
  NOT NOT1_6164(.VSS(VSS),.VDD(VDD),.Y(g10405),.A(g7064));
  NOT NOT1_6165(.VSS(VSS),.VDD(VDD),.Y(g32636),.A(g31376));
  NOT NOT1_6166(.VSS(VSS),.VDD(VDD),.Y(I23998),.A(g22182));
  NOT NOT1_6167(.VSS(VSS),.VDD(VDD),.Y(I32788),.A(g34577));
  NOT NOT1_6168(.VSS(VSS),.VDD(VDD),.Y(g32415),.A(g31591));
  NOT NOT1_6169(.VSS(VSS),.VDD(VDD),.Y(g14405),.A(g12170));
  NOT NOT1_6170(.VSS(VSS),.VDD(VDD),.Y(g19695),.A(g17015));
  NOT NOT1_6171(.VSS(VSS),.VDD(VDD),.Y(g8538),.A(g3412));
  NOT NOT1_6172(.VSS(VSS),.VDD(VDD),.Y(I12819),.A(g4277));
  NOT NOT1_6173(.VSS(VSS),.VDD(VDD),.Y(g29977),.A(g28920));
  NOT NOT1_6174(.VSS(VSS),.VDD(VDD),.Y(I12910),.A(g4340));
  NOT NOT1_6175(.VSS(VSS),.VDD(VDD),.Y(g16874),.A(I18066));
  NOT NOT1_6176(.VSS(VSS),.VDD(VDD),.Y(g32852),.A(g30614));
  NOT NOT1_6177(.VSS(VSS),.VDD(VDD),.Y(g11235),.A(I14301));
  NOT NOT1_6178(.VSS(VSS),.VDD(VDD),.Y(I32535),.A(g34296));
  NOT NOT1_6179(.VSS(VSS),.VDD(VDD),.Y(I25327),.A(g24641));
  NOT NOT1_6180(.VSS(VSS),.VDD(VDD),.Y(g8509),.A(g4141));
  NOT NOT1_6181(.VSS(VSS),.VDD(VDD),.Y(g35002),.A(I33300));
  NOT NOT1_6182(.VSS(VSS),.VDD(VDD),.Y(g19526),.A(g16349));
  NOT NOT1_6183(.VSS(VSS),.VDD(VDD),.Y(g16630),.A(g14142));
  NOT NOT1_6184(.VSS(VSS),.VDD(VDD),.Y(g16693),.A(I17901));
  NOT NOT1_6185(.VSS(VSS),.VDD(VDD),.Y(g26814),.A(g25221));
  NOT NOT1_6186(.VSS(VSS),.VDD(VDD),.Y(g34543),.A(g34359));
  NOT NOT1_6187(.VSS(VSS),.VDD(VDD),.Y(I22425),.A(g19379));
  NOT NOT1_6188(.VSS(VSS),.VDD(VDD),.Y(g24173),.A(I23363));
  NOT NOT1_6189(.VSS(VSS),.VDD(VDD),.Y(g32963),.A(g30825));
  NOT NOT1_6190(.VSS(VSS),.VDD(VDD),.Y(g22148),.A(g19074));
  NOT NOT1_6191(.VSS(VSS),.VDD(VDD),.Y(g7515),.A(I12000));
  NOT NOT1_6192(.VSS(VSS),.VDD(VDD),.Y(g12871),.A(g10378));
  NOT NOT1_6193(.VSS(VSS),.VDD(VDD),.Y(g29353),.A(I27713));
  NOT NOT1_6194(.VSS(VSS),.VDD(VDD),.Y(I12070),.A(g785));
  NOT NOT1_6195(.VSS(VSS),.VDD(VDD),.Y(I22458),.A(g18954));
  NOT NOT1_6196(.VSS(VSS),.VDD(VDD),.Y(g23537),.A(g20785));
  NOT NOT1_6197(.VSS(VSS),.VDD(VDD),.Y(g9568),.A(g6181));
  NOT NOT1_6198(.VSS(VSS),.VDD(VDD),.Y(g31842),.A(g29385));
  NOT NOT1_6199(.VSS(VSS),.VDD(VDD),.Y(g32664),.A(g31528));
  NOT NOT1_6200(.VSS(VSS),.VDD(VDD),.Y(g30569),.A(I28838));
  NOT NOT1_6201(.VSS(VSS),.VDD(VDD),.Y(I16345),.A(g881));
  NOT NOT1_6202(.VSS(VSS),.VDD(VDD),.Y(g8418),.A(g2619));
  NOT NOT1_6203(.VSS(VSS),.VDD(VDD),.Y(I19772),.A(g17818));
  NOT NOT1_6204(.VSS(VSS),.VDD(VDD),.Y(g34569),.A(I32639));
  NOT NOT1_6205(.VSS(VSS),.VDD(VDD),.Y(g22646),.A(g19389));
  NOT NOT1_6206(.VSS(VSS),.VDD(VDD),.Y(I22918),.A(g21451));
  NOT NOT1_6207(.VSS(VSS),.VDD(VDD),.Y(g17433),.A(I18382));
  NOT NOT1_6208(.VSS(VSS),.VDD(VDD),.Y(I25606),.A(g25465));
  NOT NOT1_6209(.VSS(VSS),.VDD(VDD),.Y(g8290),.A(g218));
  NOT NOT1_6210(.VSS(VSS),.VDD(VDD),.Y(I17425),.A(g13416));
  NOT NOT1_6211(.VSS(VSS),.VDD(VDD),.Y(g18903),.A(g15758));
  NOT NOT1_6212(.VSS(VSS),.VDD(VDD),.Y(g30568),.A(g29339));
  NOT NOT1_6213(.VSS(VSS),.VDD(VDD),.Y(g23283),.A(g20785));
  NOT NOT1_6214(.VSS(VSS),.VDD(VDD),.Y(g19866),.A(g16540));
  NOT NOT1_6215(.VSS(VSS),.VDD(VDD),.Y(g11991),.A(g9485));
  NOT NOT1_6216(.VSS(VSS),.VDD(VDD),.Y(I17919),.A(g14609));
  NOT NOT1_6217(.VSS(VSS),.VDD(VDD),.Y(g13414),.A(g11048));
  NOT NOT1_6218(.VSS(VSS),.VDD(VDD),.Y(I22444),.A(g19626));
  NOT NOT1_6219(.VSS(VSS),.VDD(VDD),.Y(g23492),.A(g21562));
  NOT NOT1_6220(.VSS(VSS),.VDD(VDD),.Y(g25423),.A(I24558));
  NOT NOT1_6221(.VSS(VSS),.VDD(VDD),.Y(g23303),.A(g20785));
  NOT NOT1_6222(.VSS(VSS),.VDD(VDD),.Y(I31622),.A(g33204));
  NOT NOT1_6223(.VSS(VSS),.VDD(VDD),.Y(g32576),.A(g30614));
  NOT NOT1_6224(.VSS(VSS),.VDD(VDD),.Y(g24134),.A(g19984));
  NOT NOT1_6225(.VSS(VSS),.VDD(VDD),.Y(g8093),.A(g1624));
  NOT NOT1_6226(.VSS(VSS),.VDD(VDD),.Y(g32484),.A(g31566));
  NOT NOT1_6227(.VSS(VSS),.VDD(VDD),.Y(g34242),.A(I32225));
  NOT NOT1_6228(.VSS(VSS),.VDD(VDD),.Y(g24029),.A(g20982));
  NOT NOT1_6229(.VSS(VSS),.VDD(VDD),.Y(g33424),.A(g32415));
  NOT NOT1_6230(.VSS(VSS),.VDD(VDD),.Y(I11701),.A(g4164));
  NOT NOT1_6231(.VSS(VSS),.VDD(VDD),.Y(g10113),.A(g2084));
  NOT NOT1_6232(.VSS(VSS),.VDD(VDD),.Y(g17811),.A(g12925));
  NOT NOT1_6233(.VSS(VSS),.VDD(VDD),.Y(g17646),.A(I18609));
  NOT NOT1_6234(.VSS(VSS),.VDD(VDD),.Y(I11777),.A(g5357));
  NOT NOT1_6235(.VSS(VSS),.VDD(VDD),.Y(g20506),.A(g15426));
  NOT NOT1_6236(.VSS(VSS),.VDD(VDD),.Y(I28199),.A(g28803));
  NOT NOT1_6237(.VSS(VSS),.VDD(VDD),.Y(I25750),.A(g26823));
  NOT NOT1_6238(.VSS(VSS),.VDD(VDD),.Y(g20028),.A(g15371));
  NOT NOT1_6239(.VSS(VSS),.VDD(VDD),.Y(I12067),.A(g739));
  NOT NOT1_6240(.VSS(VSS),.VDD(VDD),.Y(I32173),.A(g33645));
  NOT NOT1_6241(.VSS(VSS),.VDD(VDD),.Y(g32554),.A(g30614));
  NOT NOT1_6242(.VSS(VSS),.VDD(VDD),.Y(I18089),.A(g13144));
  NOT NOT1_6243(.VSS(VSS),.VDD(VDD),.Y(g24506),.A(I23711));
  NOT NOT1_6244(.VSS(VSS),.VDD(VDD),.Y(I20385),.A(g16194));
  NOT NOT1_6245(.VSS(VSS),.VDD(VDD),.Y(g7750),.A(g1070));
  NOT NOT1_6246(.VSS(VSS),.VDD(VDD),.Y(g24028),.A(g20841));
  NOT NOT1_6247(.VSS(VSS),.VDD(VDD),.Y(I24784),.A(g24265));
  NOT NOT1_6248(.VSS(VSS),.VDD(VDD),.Y(g34123),.A(I32062));
  NOT NOT1_6249(.VSS(VSS),.VDD(VDD),.Y(g16712),.A(g13223));
  NOT NOT1_6250(.VSS(VSS),.VDD(VDD),.Y(g26841),.A(g24893));
  NOT NOT1_6251(.VSS(VSS),.VDD(VDD),.Y(g32609),.A(g30735));
  NOT NOT1_6252(.VSS(VSS),.VDD(VDD),.Y(g21381),.A(g18008));
  NOT NOT1_6253(.VSS(VSS),.VDD(VDD),.Y(I27735),.A(g28779));
  NOT NOT1_6254(.VSS(VSS),.VDD(VDD),.Y(I29239),.A(g29498));
  NOT NOT1_6255(.VSS(VSS),.VDD(VDD),.Y(g31830),.A(g29385));
  NOT NOT1_6256(.VSS(VSS),.VDD(VDD),.Y(g23982),.A(g19147));
  NOT NOT1_6257(.VSS(VSS),.VDD(VDD),.Y(g10357),.A(g6825));
  NOT NOT1_6258(.VSS(VSS),.VDD(VDD),.Y(g26510),.A(I25369));
  NOT NOT1_6259(.VSS(VSS),.VDD(VDD),.Y(g14357),.A(g12181));
  NOT NOT1_6260(.VSS(VSS),.VDD(VDD),.Y(g34772),.A(I32960));
  NOT NOT1_6261(.VSS(VSS),.VDD(VDD),.Y(I12735),.A(g4572));
  NOT NOT1_6262(.VSS(VSS),.VDD(VDD),.Y(g8181),.A(g424));
  NOT NOT1_6263(.VSS(VSS),.VDD(VDD),.Y(g28779),.A(I27253));
  NOT NOT1_6264(.VSS(VSS),.VDD(VDD),.Y(g32608),.A(g31376));
  NOT NOT1_6265(.VSS(VSS),.VDD(VDD),.Y(g8381),.A(g2610));
  NOT NOT1_6266(.VSS(VSS),.VDD(VDD),.Y(g19689),.A(g16795));
  NOT NOT1_6267(.VSS(VSS),.VDD(VDD),.Y(g7040),.A(g4821));
  NOT NOT1_6268(.VSS(VSS),.VDD(VDD),.Y(g25117),.A(g22417));
  NOT NOT1_6269(.VSS(VSS),.VDD(VDD),.Y(I16135),.A(g10430));
  NOT NOT1_6270(.VSS(VSS),.VDD(VDD),.Y(g25000),.A(g23630));
  NOT NOT1_6271(.VSS(VSS),.VDD(VDD),.Y(g8685),.A(g1430));
  NOT NOT1_6272(.VSS(VSS),.VDD(VDD),.Y(g7440),.A(g329));
  NOT NOT1_6273(.VSS(VSS),.VDD(VDD),.Y(g8700),.A(g4054));
  NOT NOT1_6274(.VSS(VSS),.VDD(VDD),.Y(g28081),.A(I26584));
  NOT NOT1_6275(.VSS(VSS),.VDD(VDD),.Y(g32921),.A(g31672));
  NOT NOT1_6276(.VSS(VSS),.VDD(VDD),.Y(g33713),.A(I31564));
  NOT NOT1_6277(.VSS(VSS),.VDD(VDD),.Y(g8397),.A(g3470));
  NOT NOT1_6278(.VSS(VSS),.VDD(VDD),.Y(g19688),.A(g16777));
  NOT NOT1_6279(.VSS(VSS),.VDD(VDD),.Y(g9626),.A(g6466));
  NOT NOT1_6280(.VSS(VSS),.VDD(VDD),.Y(g8021),.A(g3512));
  NOT NOT1_6281(.VSS(VSS),.VDD(VDD),.Y(g16594),.A(I17772));
  NOT NOT1_6282(.VSS(VSS),.VDD(VDD),.Y(g26835),.A(I25555));
  NOT NOT1_6283(.VSS(VSS),.VDD(VDD),.Y(g13584),.A(g12735));
  NOT NOT1_6284(.VSS(VSS),.VDD(VDD),.Y(g18990),.A(g16136));
  NOT NOT1_6285(.VSS(VSS),.VDD(VDD),.Y(g32745),.A(g31376));
  NOT NOT1_6286(.VSS(VSS),.VDD(VDD),.Y(I29185),.A(g30012));
  NOT NOT1_6287(.VSS(VSS),.VDD(VDD),.Y(g22896),.A(g21012));
  NOT NOT1_6288(.VSS(VSS),.VDD(VDD),.Y(I18700),.A(g6027));
  NOT NOT1_6289(.VSS(VSS),.VDD(VDD),.Y(g23840),.A(g19074));
  NOT NOT1_6290(.VSS(VSS),.VDD(VDD),.Y(g15733),.A(I17249));
  NOT NOT1_6291(.VSS(VSS),.VDD(VDD),.Y(g32799),.A(g31710));
  NOT NOT1_6292(.VSS(VSS),.VDD(VDD),.Y(g18898),.A(g15566));
  NOT NOT1_6293(.VSS(VSS),.VDD(VDD),.Y(g23390),.A(g21468));
  NOT NOT1_6294(.VSS(VSS),.VDD(VDD),.Y(g32813),.A(g31710));
  NOT NOT1_6295(.VSS(VSS),.VDD(VDD),.Y(g22228),.A(I21810));
  NOT NOT1_6296(.VSS(VSS),.VDD(VDD),.Y(g6820),.A(g1070));
  NOT NOT1_6297(.VSS(VSS),.VDD(VDD),.Y(g33705),.A(I31550));
  NOT NOT1_6298(.VSS(VSS),.VDD(VDD),.Y(g25242),.A(g23684));
  NOT NOT1_6299(.VSS(VSS),.VDD(VDD),.Y(g7666),.A(g4076));
  NOT NOT1_6300(.VSS(VSS),.VDD(VDD),.Y(I17159),.A(g13350));
  NOT NOT1_6301(.VSS(VSS),.VDD(VDD),.Y(g20649),.A(g18065));
  NOT NOT1_6302(.VSS(VSS),.VDD(VDD),.Y(I17125),.A(g13809));
  NOT NOT1_6303(.VSS(VSS),.VDD(VDD),.Y(I22561),.A(g20841));
  NOT NOT1_6304(.VSS(VSS),.VDD(VDD),.Y(I23149),.A(g19061));
  NOT NOT1_6305(.VSS(VSS),.VDD(VDD),.Y(g31189),.A(I29002));
  NOT NOT1_6306(.VSS(VSS),.VDD(VDD),.Y(g34992),.A(I33276));
  NOT NOT1_6307(.VSS(VSS),.VDD(VDD),.Y(I17901),.A(g3976));
  NOT NOT1_6308(.VSS(VSS),.VDD(VDD),.Y(g34391),.A(g34200));
  NOT NOT1_6309(.VSS(VSS),.VDD(VDD),.Y(g32798),.A(g31672));
  NOT NOT1_6310(.VSS(VSS),.VDD(VDD),.Y(I22353),.A(g19375));
  NOT NOT1_6311(.VSS(VSS),.VDD(VDD),.Y(g28380),.A(g27064));
  NOT NOT1_6312(.VSS(VSS),.VDD(VDD),.Y(g20240),.A(g17847));
  NOT NOT1_6313(.VSS(VSS),.VDD(VDD),.Y(I23387),.A(g23394));
  NOT NOT1_6314(.VSS(VSS),.VDD(VDD),.Y(g32973),.A(g31021));
  NOT NOT1_6315(.VSS(VSS),.VDD(VDD),.Y(I30904),.A(g32424));
  NOT NOT1_6316(.VSS(VSS),.VDD(VDD),.Y(g34510),.A(g34418));
  NOT NOT1_6317(.VSS(VSS),.VDD(VDD),.Y(g22716),.A(g19795));
  NOT NOT1_6318(.VSS(VSS),.VDD(VDD),.Y(g23192),.A(g20248));
  NOT NOT1_6319(.VSS(VSS),.VDD(VDD),.Y(g16675),.A(I17873));
  NOT NOT1_6320(.VSS(VSS),.VDD(VDD),.Y(g20648),.A(g15615));
  NOT NOT1_6321(.VSS(VSS),.VDD(VDD),.Y(g10881),.A(g7567));
  NOT NOT1_6322(.VSS(VSS),.VDD(VDD),.Y(I17783),.A(g13304));
  NOT NOT1_6323(.VSS(VSS),.VDD(VDD),.Y(g20903),.A(g17249));
  NOT NOT1_6324(.VSS(VSS),.VDD(VDD),.Y(g32805),.A(g31672));
  NOT NOT1_6325(.VSS(VSS),.VDD(VDD),.Y(g13082),.A(g10981));
  NOT NOT1_6326(.VSS(VSS),.VDD(VDD),.Y(g32674),.A(g30735));
  NOT NOT1_6327(.VSS(VSS),.VDD(VDD),.Y(g24648),.A(g23148));
  NOT NOT1_6328(.VSS(VSS),.VDD(VDD),.Y(g7528),.A(g930));
  NOT NOT1_6329(.VSS(VSS),.VDD(VDD),.Y(g12859),.A(g10366));
  NOT NOT1_6330(.VSS(VSS),.VDD(VDD),.Y(g13107),.A(g10476));
  NOT NOT1_6331(.VSS(VSS),.VDD(VDD),.Y(g34579),.A(I32659));
  NOT NOT1_6332(.VSS(VSS),.VDD(VDD),.Y(g7648),.A(I12135));
  NOT NOT1_6333(.VSS(VSS),.VDD(VDD),.Y(g26615),.A(g25432));
  NOT NOT1_6334(.VSS(VSS),.VDD(VDD),.Y(g12950),.A(g12708));
  NOT NOT1_6335(.VSS(VSS),.VDD(VDD),.Y(g20604),.A(g17873));
  NOT NOT1_6336(.VSS(VSS),.VDD(VDD),.Y(g9683),.A(g6140));
  NOT NOT1_6337(.VSS(VSS),.VDD(VDD),.Y(g23522),.A(g21514));
  NOT NOT1_6338(.VSS(VSS),.VDD(VDD),.Y(g18832),.A(g15634));
  NOT NOT1_6339(.VSS(VSS),.VDD(VDD),.Y(I13360),.A(g5343));
  NOT NOT1_6340(.VSS(VSS),.VDD(VDD),.Y(g24604),.A(g23112));
  NOT NOT1_6341(.VSS(VSS),.VDD(VDD),.Y(g30578),.A(g29956));
  NOT NOT1_6342(.VSS(VSS),.VDD(VDD),.Y(g33460),.A(I30998));
  NOT NOT1_6343(.VSS(VSS),.VDD(VDD),.Y(g33686),.A(g33187));
  NOT NOT1_6344(.VSS(VSS),.VDD(VDD),.Y(g19885),.A(g17249));
  NOT NOT1_6345(.VSS(VSS),.VDD(VDD),.Y(g26720),.A(g25275));
  NOT NOT1_6346(.VSS(VSS),.VDD(VDD),.Y(g7655),.A(g4332));
  NOT NOT1_6347(.VSS(VSS),.VDD(VDD),.Y(g11744),.A(I14602));
  NOT NOT1_6348(.VSS(VSS),.VDD(VDD),.Y(g20770),.A(g17955));
  NOT NOT1_6349(.VSS(VSS),.VDD(VDD),.Y(I26508),.A(g26814));
  NOT NOT1_6350(.VSS(VSS),.VDD(VDD),.Y(g9778),.A(g5069));
  NOT NOT1_6351(.VSS(VSS),.VDD(VDD),.Y(I14271),.A(g8456));
  NOT NOT1_6352(.VSS(VSS),.VDD(VDD),.Y(g20563),.A(g15171));
  NOT NOT1_6353(.VSS(VSS),.VDD(VDD),.Y(g27996),.A(I26508));
  NOT NOT1_6354(.VSS(VSS),.VDD(VDD),.Y(g32732),.A(g30825));
  NOT NOT1_6355(.VSS(VSS),.VDD(VDD),.Y(g24770),.A(g22763));
  NOT NOT1_6356(.VSS(VSS),.VDD(VDD),.Y(g8631),.A(g283));
  NOT NOT1_6357(.VSS(VSS),.VDD(VDD),.Y(g25230),.A(g23314));
  NOT NOT1_6358(.VSS(VSS),.VDD(VDD),.Y(g32934),.A(g30735));
  NOT NOT1_6359(.VSS(VSS),.VDD(VDD),.Y(g24981),.A(g22763));
  NOT NOT1_6360(.VSS(VSS),.VDD(VDD),.Y(I24089),.A(g22409));
  NOT NOT1_6361(.VSS(VSS),.VDD(VDD),.Y(g11849),.A(g7601));
  NOT NOT1_6362(.VSS(VSS),.VDD(VDD),.Y(I16613),.A(g10430));
  NOT NOT1_6363(.VSS(VSS),.VDD(VDD),.Y(g17582),.A(g14768));
  NOT NOT1_6364(.VSS(VSS),.VDD(VDD),.Y(g12996),.A(g11823));
  NOT NOT1_6365(.VSS(VSS),.VDD(VDD),.Y(g10027),.A(g6523));
  NOT NOT1_6366(.VSS(VSS),.VDD(VDD),.Y(g23483),.A(g18833));
  NOT NOT1_6367(.VSS(VSS),.VDD(VDD),.Y(I18060),.A(g14198));
  NOT NOT1_6368(.VSS(VSS),.VDD(VDD),.Y(I23369),.A(g23347));
  NOT NOT1_6369(.VSS(VSS),.VDD(VDD),.Y(g14662),.A(I16762));
  NOT NOT1_6370(.VSS(VSS),.VDD(VDD),.Y(g8301),.A(g1399));
  NOT NOT1_6371(.VSS(VSS),.VDD(VDD),.Y(g19763),.A(g16431));
  NOT NOT1_6372(.VSS(VSS),.VDD(VDD),.Y(g25265),.A(I24455));
  NOT NOT1_6373(.VSS(VSS),.VDD(VDD),.Y(I32240),.A(g34131));
  NOT NOT1_6374(.VSS(VSS),.VDD(VDD),.Y(g29976),.A(g29018));
  NOT NOT1_6375(.VSS(VSS),.VDD(VDD),.Y(g12844),.A(g10360));
  NOT NOT1_6376(.VSS(VSS),.VDD(VDD),.Y(g7410),.A(g2008));
  NOT NOT1_6377(.VSS(VSS),.VDD(VDD),.Y(g11398),.A(I14409));
  NOT NOT1_6378(.VSS(VSS),.VDD(VDD),.Y(g23862),.A(g19147));
  NOT NOT1_6379(.VSS(VSS),.VDD(VDD),.Y(g12367),.A(I15205));
  NOT NOT1_6380(.VSS(VSS),.VDD(VDD),.Y(g32692),.A(g31528));
  NOT NOT1_6381(.VSS(VSS),.VDD(VDD),.Y(g32761),.A(g30825));
  NOT NOT1_6382(.VSS(VSS),.VDD(VDD),.Y(I32648),.A(g34371));
  NOT NOT1_6383(.VSS(VSS),.VDD(VDD),.Y(g18926),.A(I19707));
  NOT NOT1_6384(.VSS(VSS),.VDD(VDD),.Y(I18855),.A(g13745));
  NOT NOT1_6385(.VSS(VSS),.VDD(VDD),.Y(I11629),.A(g19));
  NOT NOT1_6386(.VSS(VSS),.VDD(VDD),.Y(g11652),.A(g7674));
  NOT NOT1_6387(.VSS(VSS),.VDD(VDD),.Y(g9661),.A(g3661));
  NOT NOT1_6388(.VSS(VSS),.VDD(VDD),.Y(g13141),.A(g11374));
  NOT NOT1_6389(.VSS(VSS),.VDD(VDD),.Y(g29374),.A(I27742));
  NOT NOT1_6390(.VSS(VSS),.VDD(VDD),.Y(g20767),.A(g17873));
  NOT NOT1_6391(.VSS(VSS),.VDD(VDD),.Y(g26340),.A(g24953));
  NOT NOT1_6392(.VSS(VSS),.VDD(VDD),.Y(g21326),.A(I21058));
  NOT NOT1_6393(.VSS(VSS),.VDD(VDD),.Y(g18099),.A(I18903));
  NOT NOT1_6394(.VSS(VSS),.VDD(VDD),.Y(I18411),.A(g13018));
  NOT NOT1_6395(.VSS(VSS),.VDD(VDD),.Y(g30116),.A(I28349));
  NOT NOT1_6396(.VSS(VSS),.VDD(VDD),.Y(I14650),.A(g9340));
  NOT NOT1_6397(.VSS(VSS),.VDD(VDD),.Y(g33875),.A(I31727));
  NOT NOT1_6398(.VSS(VSS),.VDD(VDD),.Y(I24497),.A(g22592));
  NOT NOT1_6399(.VSS(VSS),.VDD(VDD),.Y(g10710),.A(I14006));
  NOT NOT1_6400(.VSS(VSS),.VDD(VDD),.Y(g20899),.A(I20861));
  NOT NOT1_6401(.VSS(VSS),.VDD(VDD),.Y(I12300),.A(g1157));
  NOT NOT1_6402(.VSS(VSS),.VDD(VDD),.Y(g10003),.A(I13539));
  NOT NOT1_6403(.VSS(VSS),.VDD(VDD),.Y(g23948),.A(g21012));
  NOT NOT1_6404(.VSS(VSS),.VDD(VDD),.Y(I32770),.A(g34505));
  NOT NOT1_6405(.VSS(VSS),.VDD(VDD),.Y(g18098),.A(I18900));
  NOT NOT1_6406(.VSS(VSS),.VDD(VDD),.Y(g10204),.A(g2685));
  NOT NOT1_6407(.VSS(VSS),.VDD(VDD),.Y(I29438),.A(g30610));
  NOT NOT1_6408(.VSS(VSS),.VDD(VDD),.Y(g21904),.A(I21483));
  NOT NOT1_6409(.VSS(VSS),.VDD(VDD),.Y(g14204),.A(g12155));
  NOT NOT1_6410(.VSS(VSS),.VDD(VDD),.Y(g16577),.A(I17747));
  NOT NOT1_6411(.VSS(VSS),.VDD(VDD),.Y(g20633),.A(g15171));
  NOT NOT1_6412(.VSS(VSS),.VDD(VDD),.Y(g23904),.A(g18997));
  NOT NOT1_6413(.VSS(VSS),.VDD(VDD),.Y(I16371),.A(g887));
  NOT NOT1_6414(.VSS(VSS),.VDD(VDD),.Y(g31837),.A(g29385));
  NOT NOT1_6415(.VSS(VSS),.VDD(VDD),.Y(g14779),.A(I16847));
  NOT NOT1_6416(.VSS(VSS),.VDD(VDD),.Y(g21252),.A(g15656));
  NOT NOT1_6417(.VSS(VSS),.VDD(VDD),.Y(I22289),.A(g19446));
  NOT NOT1_6418(.VSS(VSS),.VDD(VDD),.Y(g32329),.A(g31522));
  NOT NOT1_6419(.VSS(VSS),.VDD(VDD),.Y(g29669),.A(I27941));
  NOT NOT1_6420(.VSS(VSS),.VDD(VDD),.Y(g34275),.A(g34047));
  NOT NOT1_6421(.VSS(VSS),.VDD(VDD),.Y(g19480),.A(g16349));
  NOT NOT1_6422(.VSS(VSS),.VDD(VDD),.Y(g23252),.A(I22353));
  NOT NOT1_6423(.VSS(VSS),.VDD(VDD),.Y(g17603),.A(g14993));
  NOT NOT1_6424(.VSS(VSS),.VDD(VDD),.Y(g20191),.A(g17821));
  NOT NOT1_6425(.VSS(VSS),.VDD(VDD),.Y(g34430),.A(I32461));
  NOT NOT1_6426(.VSS(VSS),.VDD(VDD),.Y(g17742),.A(g14971));
  NOT NOT1_6427(.VSS(VSS),.VDD(VDD),.Y(g32539),.A(g31170));
  NOT NOT1_6428(.VSS(VSS),.VDD(VDD),.Y(g10081),.A(g2279));
  NOT NOT1_6429(.VSS(VSS),.VDD(VDD),.Y(g17096),.A(I18168));
  NOT NOT1_6430(.VSS(VSS),.VDD(VDD),.Y(I18894),.A(g16708));
  NOT NOT1_6431(.VSS(VSS),.VDD(VDD),.Y(g6995),.A(g4944));
  NOT NOT1_6432(.VSS(VSS),.VDD(VDD),.Y(g7618),.A(I12092));
  NOT NOT1_6433(.VSS(VSS),.VDD(VDD),.Y(g8441),.A(g3361));
  NOT NOT1_6434(.VSS(VSS),.VDD(VDD),.Y(g22857),.A(g20739));
  NOT NOT1_6435(.VSS(VSS),.VDD(VDD),.Y(I22571),.A(g20097));
  NOT NOT1_6436(.VSS(VSS),.VDD(VDD),.Y(I11785),.A(g5703));
  NOT NOT1_6437(.VSS(VSS),.VDD(VDD),.Y(g7235),.A(g4521));
  NOT NOT1_6438(.VSS(VSS),.VDD(VDD),.Y(g7343),.A(g5290));
  NOT NOT1_6439(.VSS(VSS),.VDD(VDD),.Y(I14365),.A(g3303));
  NOT NOT1_6440(.VSS(VSS),.VDD(VDD),.Y(g30237),.A(I28480));
  NOT NOT1_6441(.VSS(VSS),.VDD(VDD),.Y(I16795),.A(g5637));
  NOT NOT1_6442(.VSS(VSS),.VDD(VDD),.Y(g25007),.A(g22457));
  NOT NOT1_6443(.VSS(VSS),.VDD(VDD),.Y(g32538),.A(g31070));
  NOT NOT1_6444(.VSS(VSS),.VDD(VDD),.Y(g24718),.A(g22182));
  NOT NOT1_6445(.VSS(VSS),.VDD(VDD),.Y(I32794),.A(g34580));
  NOT NOT1_6446(.VSS(VSS),.VDD(VDD),.Y(g14786),.A(g12471));
  NOT NOT1_6447(.VSS(VSS),.VDD(VDD),.Y(g29195),.A(I27495));
  NOT NOT1_6448(.VSS(VSS),.VDD(VDD),.Y(g9484),.A(g1612));
  NOT NOT1_6449(.VSS(VSS),.VDD(VDD),.Y(g30983),.A(g29657));
  NOT NOT1_6450(.VSS(VSS),.VDD(VDD),.Y(g9439),.A(g5428));
  NOT NOT1_6451(.VSS(VSS),.VDD(VDD),.Y(g17681),.A(g14735));
  NOT NOT1_6452(.VSS(VSS),.VDD(VDD),.Y(g7566),.A(I12049));
  NOT NOT1_6453(.VSS(VSS),.VDD(VDD),.Y(g6840),.A(g1992));
  NOT NOT1_6454(.VSS(VSS),.VDD(VDD),.Y(g8673),.A(g4737));
  NOT NOT1_6455(.VSS(VSS),.VDD(VDD),.Y(g16349),.A(I17661));
  NOT NOT1_6456(.VSS(VSS),.VDD(VDD),.Y(g34983),.A(I33249));
  NOT NOT1_6457(.VSS(VSS),.VDD(VDD),.Y(g18997),.A(I19756));
  NOT NOT1_6458(.VSS(VSS),.VDD(VDD),.Y(g10356),.A(g6819));
  NOT NOT1_6459(.VSS(VSS),.VDD(VDD),.Y(g33455),.A(I30983));
  NOT NOT1_6460(.VSS(VSS),.VDD(VDD),.Y(g21183),.A(g15509));
  NOT NOT1_6461(.VSS(VSS),.VDD(VDD),.Y(g21673),.A(I21234));
  NOT NOT1_6462(.VSS(VSS),.VDD(VDD),.Y(g7693),.A(g4849));
  NOT NOT1_6463(.VSS(VSS),.VDD(VDD),.Y(g11833),.A(g8026));
  NOT NOT1_6464(.VSS(VSS),.VDD(VDD),.Y(g17429),.A(I18370));
  NOT NOT1_6465(.VSS(VSS),.VDD(VDD),.Y(g7134),.A(g5029));
  NOT NOT1_6466(.VSS(VSS),.VDD(VDD),.Y(g21397),.A(g15171));
  NOT NOT1_6467(.VSS(VSS),.VDD(VDD),.Y(g23847),.A(g19210));
  NOT NOT1_6468(.VSS(VSS),.VDD(VDD),.Y(g13049),.A(I15677));
  NOT NOT1_6469(.VSS(VSS),.VDD(VDD),.Y(g10380),.A(g6960));
  NOT NOT1_6470(.VSS(VSS),.VDD(VDD),.Y(g30142),.A(g28754));
  NOT NOT1_6471(.VSS(VSS),.VDD(VDD),.Y(g18061),.A(g14800));
  NOT NOT1_6472(.VSS(VSS),.VDD(VDD),.Y(g16284),.A(I17609));
  NOT NOT1_6473(.VSS(VSS),.VDD(VDD),.Y(g19431),.A(g16249));
  NOT NOT1_6474(.VSS(VSS),.VDD(VDD),.Y(g34142),.A(I32089));
  NOT NOT1_6475(.VSS(VSS),.VDD(VDD),.Y(g25116),.A(g22369));
  NOT NOT1_6476(.VSS(VSS),.VDD(VDD),.Y(g17428),.A(I18367));
  NOT NOT1_6477(.VSS(VSS),.VDD(VDD),.Y(I22816),.A(g19862));
  NOT NOT1_6478(.VSS(VSS),.VDD(VDD),.Y(g7548),.A(g1036));
  NOT NOT1_6479(.VSS(VSS),.VDD(VDD),.Y(g11048),.A(I14158));
  NOT NOT1_6480(.VSS(VSS),.VDD(VDD),.Y(g8669),.A(g3767));
  NOT NOT1_6481(.VSS(VSS),.VDD(VDD),.Y(g10090),.A(g5348));
  NOT NOT1_6482(.VSS(VSS),.VDD(VDD),.Y(g20573),.A(g17384));
  NOT NOT1_6483(.VSS(VSS),.VDD(VDD),.Y(g10233),.A(I13699));
  NOT NOT1_6484(.VSS(VSS),.VDD(VDD),.Y(g20247),.A(g17015));
  NOT NOT1_6485(.VSS(VSS),.VDD(VDD),.Y(g29893),.A(g28755));
  NOT NOT1_6486(.VSS(VSS),.VDD(VDD),.Y(I24060),.A(g22202));
  NOT NOT1_6487(.VSS(VSS),.VDD(VDD),.Y(g16622),.A(g14104));
  NOT NOT1_6488(.VSS(VSS),.VDD(VDD),.Y(g23509),.A(g21611));
  NOT NOT1_6489(.VSS(VSS),.VDD(VDD),.Y(g10182),.A(g2681));
  NOT NOT1_6490(.VSS(VSS),.VDD(VDD),.Y(g28620),.A(g27679));
  NOT NOT1_6491(.VSS(VSS),.VDD(VDD),.Y(I21959),.A(g20242));
  NOT NOT1_6492(.VSS(VSS),.VDD(VDD),.Y(g20389),.A(g15277));
  NOT NOT1_6493(.VSS(VSS),.VDD(VDD),.Y(g8058),.A(g3115));
  NOT NOT1_6494(.VSS(VSS),.VDD(VDD),.Y(I14708),.A(g9417));
  NOT NOT1_6495(.VSS(VSS),.VDD(VDD),.Y(I28458),.A(g28443));
  NOT NOT1_6496(.VSS(VSS),.VDD(VDD),.Y(I29139),.A(g29382));
  NOT NOT1_6497(.VSS(VSS),.VDD(VDD),.Y(g8531),.A(g3288));
  NOT NOT1_6498(.VSS(VSS),.VDD(VDD),.Y(g19773),.A(g17615));
  NOT NOT1_6499(.VSS(VSS),.VDD(VDD),.Y(g24389),.A(g22908));
  NOT NOT1_6500(.VSS(VSS),.VDD(VDD),.Y(g8458),.A(g294));
  NOT NOT1_6501(.VSS(VSS),.VDD(VDD),.Y(g24045),.A(g21193));
  NOT NOT1_6502(.VSS(VSS),.VDD(VDD),.Y(g12902),.A(g10409));
  NOT NOT1_6503(.VSS(VSS),.VDD(VDD),.Y(g20612),.A(g18008));
  NOT NOT1_6504(.VSS(VSS),.VDD(VDD),.Y(g23508),.A(g21562));
  NOT NOT1_6505(.VSS(VSS),.VDD(VDD),.Y(I16163),.A(g11930));
  NOT NOT1_6506(.VSS(VSS),.VDD(VDD),.Y(I20870),.A(g16216));
  NOT NOT1_6507(.VSS(VSS),.VDD(VDD),.Y(g32771),.A(g31021));
  NOT NOT1_6508(.VSS(VSS),.VDD(VDD),.Y(g8743),.A(g550));
  NOT NOT1_6509(.VSS(VSS),.VDD(VDD),.Y(g20388),.A(g17297));
  NOT NOT1_6510(.VSS(VSS),.VDD(VDD),.Y(g20324),.A(g17955));
  NOT NOT1_6511(.VSS(VSS),.VDD(VDD),.Y(g8890),.A(g376));
  NOT NOT1_6512(.VSS(VSS),.VDD(VDD),.Y(I23378),.A(g23426));
  NOT NOT1_6513(.VSS(VSS),.VDD(VDD),.Y(g29713),.A(I27970));
  NOT NOT1_6514(.VSS(VSS),.VDD(VDD),.Y(g24099),.A(g20720));
  NOT NOT1_6515(.VSS(VSS),.VDD(VDD),.Y(g24388),.A(g22885));
  NOT NOT1_6516(.VSS(VSS),.VDD(VDD),.Y(g20701),.A(g17955));
  NOT NOT1_6517(.VSS(VSS),.VDD(VDD),.Y(g20777),.A(g15224));
  NOT NOT1_6518(.VSS(VSS),.VDD(VDD),.Y(g20534),.A(g17183));
  NOT NOT1_6519(.VSS(VSS),.VDD(VDD),.Y(g22317),.A(g19801));
  NOT NOT1_6520(.VSS(VSS),.VDD(VDD),.Y(g31623),.A(g29669));
  NOT NOT1_6521(.VSS(VSS),.VDD(VDD),.Y(g32683),.A(g30614));
  NOT NOT1_6522(.VSS(VSS),.VDD(VDD),.Y(I17976),.A(g13638));
  NOT NOT1_6523(.VSS(VSS),.VDD(VDD),.Y(g25465),.A(g23824));
  NOT NOT1_6524(.VSS(VSS),.VDD(VDD),.Y(g19670),.A(g16897));
  NOT NOT1_6525(.VSS(VSS),.VDD(VDD),.Y(g24534),.A(g22670));
  NOT NOT1_6526(.VSS(VSS),.VDD(VDD),.Y(g8505),.A(g3480));
  NOT NOT1_6527(.VSS(VSS),.VDD(VDD),.Y(g20272),.A(g17239));
  NOT NOT1_6528(.VSS(VSS),.VDD(VDD),.Y(g34130),.A(I32071));
  NOT NOT1_6529(.VSS(VSS),.VDD(VDD),.Y(g24098),.A(g19984));
  NOT NOT1_6530(.VSS(VSS),.VDD(VDD),.Y(g14331),.A(I16489));
  NOT NOT1_6531(.VSS(VSS),.VDD(VDD),.Y(g12738),.A(g9374));
  NOT NOT1_6532(.VSS(VSS),.VDD(VDD),.Y(I19863),.A(g16675));
  NOT NOT1_6533(.VSS(VSS),.VDD(VDD),.Y(g9616),.A(g5452));
  NOT NOT1_6534(.VSS(VSS),.VDD(VDD),.Y(g17504),.A(g15021));
  NOT NOT1_6535(.VSS(VSS),.VDD(VDD),.Y(I16541),.A(g11929));
  NOT NOT1_6536(.VSS(VSS),.VDD(VDD),.Y(g8011),.A(g3167));
  NOT NOT1_6537(.VSS(VSS),.VDD(VDD),.Y(g25340),.A(g22763));
  NOT NOT1_6538(.VSS(VSS),.VDD(VDD),.Y(g25035),.A(g23699));
  NOT NOT1_6539(.VSS(VSS),.VDD(VDD),.Y(I17374),.A(g13638));
  NOT NOT1_6540(.VSS(VSS),.VDD(VDD),.Y(g8411),.A(I12577));
  NOT NOT1_6541(.VSS(VSS),.VDD(VDD),.Y(g8734),.A(g4045));
  NOT NOT1_6542(.VSS(VSS),.VDD(VDD),.Y(g19734),.A(g16861));
  NOT NOT1_6543(.VSS(VSS),.VDD(VDD),.Y(g13106),.A(g10981));
  NOT NOT1_6544(.VSS(VSS),.VDD(VDD),.Y(g27698),.A(g26648));
  NOT NOT1_6545(.VSS(VSS),.VDD(VDD),.Y(g29042),.A(I27388));
  NOT NOT1_6546(.VSS(VSS),.VDD(VDD),.Y(g13605),.A(I16040));
  NOT NOT1_6547(.VSS(VSS),.VDD(VDD),.Y(g10897),.A(g7601));
  NOT NOT1_6548(.VSS(VSS),.VDD(VDD),.Y(I33214),.A(g34954));
  NOT NOT1_6549(.VSS(VSS),.VDD(VDD),.Y(I20867),.A(g16216));
  NOT NOT1_6550(.VSS(VSS),.VDD(VDD),.Y(I27314),.A(g28009));
  NOT NOT1_6551(.VSS(VSS),.VDD(VDD),.Y(g6954),.A(g4138));
  NOT NOT1_6552(.VSS(VSS),.VDD(VDD),.Y(g19930),.A(g17200));
  NOT NOT1_6553(.VSS(VSS),.VDD(VDD),.Y(g6810),.A(g723));
  NOT NOT1_6554(.VSS(VSS),.VDD(VDD),.Y(g9527),.A(g6500));
  NOT NOT1_6555(.VSS(VSS),.VDD(VDD),.Y(I14069),.A(g9104));
  NOT NOT1_6556(.VSS(VSS),.VDD(VDD),.Y(g11812),.A(g7567));
  NOT NOT1_6557(.VSS(VSS),.VDD(VDD),.Y(g7202),.A(g4639));
  NOT NOT1_6558(.VSS(VSS),.VDD(VDD),.Y(I16724),.A(g12108));
  NOT NOT1_6559(.VSS(VSS),.VDD(VDD),.Y(g10404),.A(g7026));
  NOT NOT1_6560(.VSS(VSS),.VDD(VDD),.Y(I12314),.A(g1500));
  NOT NOT1_6561(.VSS(VSS),.VDD(VDD),.Y(g13463),.A(g10476));
  NOT NOT1_6562(.VSS(VSS),.VDD(VDD),.Y(g31822),.A(g29385));
  NOT NOT1_6563(.VSS(VSS),.VDD(VDD),.Y(g32515),.A(g30825));
  NOT NOT1_6564(.VSS(VSS),.VDD(VDD),.Y(I31539),.A(g33212));
  NOT NOT1_6565(.VSS(VSS),.VDD(VDD),.Y(g32882),.A(g31376));
  NOT NOT1_6566(.VSS(VSS),.VDD(VDD),.Y(I14602),.A(g9340));
  NOT NOT1_6567(.VSS(VSS),.VDD(VDD),.Y(I15033),.A(g10273));
  NOT NOT1_6568(.VSS(VSS),.VDD(VDD),.Y(g19694),.A(g16429));
  NOT NOT1_6569(.VSS(VSS),.VDD(VDD),.Y(g7908),.A(g4157));
  NOT NOT1_6570(.VSS(VSS),.VDD(VDD),.Y(I32388),.A(g34153));
  NOT NOT1_6571(.VSS(VSS),.VDD(VDD),.Y(g24032),.A(g21256));
  NOT NOT1_6572(.VSS(VSS),.VDD(VDD),.Y(g22626),.A(I21941));
  NOT NOT1_6573(.VSS(VSS),.VDD(VDD),.Y(I21802),.A(g21308));
  NOT NOT1_6574(.VSS(VSS),.VDD(VDD),.Y(I16829),.A(g6715));
  NOT NOT1_6575(.VSS(VSS),.VDD(VDD),.Y(g25517),.A(g22228));
  NOT NOT1_6576(.VSS(VSS),.VDD(VDD),.Y(g11033),.A(g8500));
  NOT NOT1_6577(.VSS(VSS),.VDD(VDD),.Y(g11371),.A(g7565));
  NOT NOT1_6578(.VSS(VSS),.VDD(VDD),.Y(I16535),.A(g11235));
  NOT NOT1_6579(.VSS(VSS),.VDD(VDD),.Y(g18911),.A(g15169));
  NOT NOT1_6580(.VSS(VSS),.VDD(VDD),.Y(g23452),.A(g21468));
  NOT NOT1_6581(.VSS(VSS),.VDD(VDD),.Y(g10026),.A(g6494));
  NOT NOT1_6582(.VSS(VSS),.VDD(VDD),.Y(g32407),.A(I29939));
  NOT NOT1_6583(.VSS(VSS),.VDD(VDD),.Y(g9546),.A(g2437));
  NOT NOT1_6584(.VSS(VSS),.VDD(VDD),.Y(g13033),.A(g11917));
  NOT NOT1_6585(.VSS(VSS),.VDD(VDD),.Y(g21205),.A(g15656));
  NOT NOT1_6586(.VSS(VSS),.VDD(VDD),.Y(g11234),.A(g8355));
  NOT NOT1_6587(.VSS(VSS),.VDD(VDD),.Y(g10212),.A(g6390));
  NOT NOT1_6588(.VSS(VSS),.VDD(VDD),.Y(I14970),.A(g9965));
  NOT NOT1_6589(.VSS(VSS),.VDD(VDD),.Y(g29939),.A(g28857));
  NOT NOT1_6590(.VSS(VSS),.VDD(VDD),.Y(g17128),.A(I18180));
  NOT NOT1_6591(.VSS(VSS),.VDD(VDD),.Y(g7518),.A(g1024));
  NOT NOT1_6592(.VSS(VSS),.VDD(VDD),.Y(I17668),.A(g13279));
  NOT NOT1_6593(.VSS(VSS),.VDD(VDD),.Y(I20819),.A(g17088));
  NOT NOT1_6594(.VSS(VSS),.VDD(VDD),.Y(I22525),.A(g19345));
  NOT NOT1_6595(.VSS(VSS),.VDD(VDD),.Y(I22488),.A(g18984));
  NOT NOT1_6596(.VSS(VSS),.VDD(VDD),.Y(I17842),.A(g13051));
  NOT NOT1_6597(.VSS(VSS),.VDD(VDD),.Y(I20910),.A(g17197));
  NOT NOT1_6598(.VSS(VSS),.VDD(VDD),.Y(g16963),.A(I18117));
  NOT NOT1_6599(.VSS(VSS),.VDD(VDD),.Y(g23912),.A(g19147));
  NOT NOT1_6600(.VSS(VSS),.VDD(VDD),.Y(I17392),.A(g13680));
  NOT NOT1_6601(.VSS(VSS),.VDD(VDD),.Y(g34222),.A(I32195));
  NOT NOT1_6602(.VSS(VSS),.VDD(VDD),.Y(g9970),.A(g1714));
  NOT NOT1_6603(.VSS(VSS),.VDD(VDD),.Y(g24061),.A(g19919));
  NOT NOT1_6604(.VSS(VSS),.VDD(VDD),.Y(I29585),.A(g31655));
  NOT NOT1_6605(.VSS(VSS),.VDD(VDD),.Y(g29093),.A(g27858));
  NOT NOT1_6606(.VSS(VSS),.VDD(VDD),.Y(g34437),.A(I32482));
  NOT NOT1_6607(.VSS(VSS),.VDD(VDD),.Y(g20766),.A(g17433));
  NOT NOT1_6608(.VSS(VSS),.VDD(VDD),.Y(I26929),.A(g27980));
  NOT NOT1_6609(.VSS(VSS),.VDD(VDD),.Y(g8080),.A(g3863));
  NOT NOT1_6610(.VSS(VSS),.VDD(VDD),.Y(I18526),.A(g13055));
  NOT NOT1_6611(.VSS(VSS),.VDD(VDD),.Y(g31853),.A(g29385));
  NOT NOT1_6612(.VSS(VSS),.VDD(VDD),.Y(g19502),.A(g15674));
  NOT NOT1_6613(.VSS(VSS),.VDD(VDD),.Y(g8480),.A(g3147));
  NOT NOT1_6614(.VSS(VSS),.VDD(VDD),.Y(g19210),.A(I19796));
  NOT NOT1_6615(.VSS(VSS),.VDD(VDD),.Y(g17533),.A(I18482));
  NOT NOT1_6616(.VSS(VSS),.VDD(VDD),.Y(g25193),.A(g22763));
  NOT NOT1_6617(.VSS(VSS),.VDD(VDD),.Y(g8713),.A(g4826));
  NOT NOT1_6618(.VSS(VSS),.VDD(VDD),.Y(g21051),.A(g15171));
  NOT NOT1_6619(.VSS(VSS),.VDD(VDD),.Y(g7593),.A(I12061));
  NOT NOT1_6620(.VSS(VSS),.VDD(VDD),.Y(I17488),.A(g13394));
  NOT NOT1_6621(.VSS(VSS),.VDD(VDD),.Y(g15348),.A(I17111));
  NOT NOT1_6622(.VSS(VSS),.VDD(VDD),.Y(g19618),.A(g16349));
  NOT NOT1_6623(.VSS(VSS),.VDD(VDD),.Y(g19443),.A(g16449));
  NOT NOT1_6624(.VSS(VSS),.VDD(VDD),.Y(I14967),.A(g9964));
  NOT NOT1_6625(.VSS(VSS),.VDD(VDD),.Y(g12895),.A(g10403));
  NOT NOT1_6626(.VSS(VSS),.VDD(VDD),.Y(I12773),.A(g4204));
  NOT NOT1_6627(.VSS(VSS),.VDD(VDD),.Y(g16585),.A(g14075));
  NOT NOT1_6628(.VSS(VSS),.VDD(VDD),.Y(g13514),.A(I15987));
  NOT NOT1_6629(.VSS(VSS),.VDD(VDD),.Y(g25523),.A(g22550));
  NOT NOT1_6630(.VSS(VSS),.VDD(VDD),.Y(g31836),.A(g29385));
  NOT NOT1_6631(.VSS(VSS),.VDD(VDD),.Y(g32441),.A(I29969));
  NOT NOT1_6632(.VSS(VSS),.VDD(VDD),.Y(g32584),.A(g30673));
  NOT NOT1_6633(.VSS(VSS),.VDD(VDD),.Y(I32997),.A(g34760));
  NOT NOT1_6634(.VSS(VSS),.VDD(VDD),.Y(g24360),.A(g22228));
  NOT NOT1_6635(.VSS(VSS),.VDD(VDD),.Y(g29219),.A(I27573));
  NOT NOT1_6636(.VSS(VSS),.VDD(VDD),.Y(g15566),.A(I17143));
  NOT NOT1_6637(.VSS(VSS),.VDD(VDD),.Y(g20447),.A(g15426));
  NOT NOT1_6638(.VSS(VSS),.VDD(VDD),.Y(g14149),.A(g12381));
  NOT NOT1_6639(.VSS(VSS),.VDD(VDD),.Y(g10387),.A(g6996));
  NOT NOT1_6640(.VSS(VSS),.VDD(VDD),.Y(g16609),.A(g14454));
  NOT NOT1_6641(.VSS(VSS),.VDD(VDD),.Y(g19469),.A(g16326));
  NOT NOT1_6642(.VSS(VSS),.VDD(VDD),.Y(I28336),.A(g29147));
  NOT NOT1_6643(.VSS(VSS),.VDD(VDD),.Y(g10620),.A(g10233));
  NOT NOT1_6644(.VSS(VSS),.VDD(VDD),.Y(g17737),.A(g14810));
  NOT NOT1_6645(.VSS(VSS),.VDD(VDD),.Y(g22856),.A(g20453));
  NOT NOT1_6646(.VSS(VSS),.VDD(VDD),.Y(g29218),.A(I27570));
  NOT NOT1_6647(.VSS(VSS),.VDD(VDD),.Y(g22995),.A(g20330));
  NOT NOT1_6648(.VSS(VSS),.VDD(VDD),.Y(g32759),.A(g31376));
  NOT NOT1_6649(.VSS(VSS),.VDD(VDD),.Y(g16200),.A(g13584));
  NOT NOT1_6650(.VSS(VSS),.VDD(VDD),.Y(I33235),.A(g34957));
  NOT NOT1_6651(.VSS(VSS),.VDD(VDD),.Y(g23350),.A(g20785));
  NOT NOT1_6652(.VSS(VSS),.VDD(VDD),.Y(g25006),.A(g22417));
  NOT NOT1_6653(.VSS(VSS),.VDD(VDD),.Y(g32725),.A(g30825));
  NOT NOT1_6654(.VSS(VSS),.VDD(VDD),.Y(g24162),.A(I23330));
  NOT NOT1_6655(.VSS(VSS),.VDD(VDD),.Y(I32766),.A(g34522));
  NOT NOT1_6656(.VSS(VSS),.VDD(VDD),.Y(g7933),.A(g907));
  NOT NOT1_6657(.VSS(VSS),.VDD(VDD),.Y(g16608),.A(g14116));
  NOT NOT1_6658(.VSS(VSS),.VDD(VDD),.Y(g19468),.A(g15938));
  NOT NOT1_6659(.VSS(VSS),.VDD(VDD),.Y(g9617),.A(I13240));
  NOT NOT1_6660(.VSS(VSS),.VDD(VDD),.Y(g23820),.A(g19147));
  NOT NOT1_6661(.VSS(VSS),.VDD(VDD),.Y(g34952),.A(g34942));
  NOT NOT1_6662(.VSS(VSS),.VDD(VDD),.Y(g34351),.A(g34174));
  NOT NOT1_6663(.VSS(VSS),.VDD(VDD),.Y(g13012),.A(I15626));
  NOT NOT1_6664(.VSS(VSS),.VDD(VDD),.Y(g32758),.A(g31327));
  NOT NOT1_6665(.VSS(VSS),.VDD(VDD),.Y(g7521),.A(g5630));
  NOT NOT1_6666(.VSS(VSS),.VDD(VDD),.Y(I32871),.A(g34521));
  NOT NOT1_6667(.VSS(VSS),.VDD(VDD),.Y(g25222),.A(I24400));
  NOT NOT1_6668(.VSS(VSS),.VDD(VDD),.Y(g7050),.A(g5845));
  NOT NOT1_6669(.VSS(VSS),.VDD(VDD),.Y(g20629),.A(g17955));
  NOT NOT1_6670(.VSS(VSS),.VDD(VDD),.Y(g23152),.A(g20283));
  NOT NOT1_6671(.VSS(VSS),.VDD(VDD),.Y(I12930),.A(g4349));
  NOT NOT1_6672(.VSS(VSS),.VDD(VDD),.Y(I13699),.A(g4581));
  NOT NOT1_6673(.VSS(VSS),.VDD(VDD),.Y(g9516),.A(g6116));
  NOT NOT1_6674(.VSS(VSS),.VDD(VDD),.Y(I21002),.A(g16709));
  NOT NOT1_6675(.VSS(VSS),.VDD(VDD),.Y(g20451),.A(g15277));
  NOT NOT1_6676(.VSS(VSS),.VDD(VDD),.Y(g21396),.A(g17955));
  NOT NOT1_6677(.VSS(VSS),.VDD(VDD),.Y(g31616),.A(I29214));
  NOT NOT1_6678(.VSS(VSS),.VDD(VDD),.Y(I14079),.A(g7231));
  NOT NOT1_6679(.VSS(VSS),.VDD(VDD),.Y(g30063),.A(g29015));
  NOT NOT1_6680(.VSS(VSS),.VDD(VDD),.Y(I22124),.A(g21300));
  NOT NOT1_6681(.VSS(VSS),.VDD(VDD),.Y(g9771),.A(g3969));
  NOT NOT1_6682(.VSS(VSS),.VDD(VDD),.Y(I29973),.A(g31213));
  NOT NOT1_6683(.VSS(VSS),.VDD(VDD),.Y(g26834),.A(I25552));
  NOT NOT1_6684(.VSS(VSS),.VDD(VDD),.Y(g20911),.A(g15171));
  NOT NOT1_6685(.VSS(VSS),.VDD(VDD),.Y(I16028),.A(g12381));
  NOT NOT1_6686(.VSS(VSS),.VDD(VDD),.Y(g10369),.A(g6873));
  NOT NOT1_6687(.VSS(VSS),.VDD(VDD),.Y(g32744),.A(g31327));
  NOT NOT1_6688(.VSS(VSS),.VDD(VDD),.Y(I31515),.A(g33187));
  NOT NOT1_6689(.VSS(VSS),.VDD(VDD),.Y(g24911),.A(I24078));
  NOT NOT1_6690(.VSS(VSS),.VDD(VDD),.Y(g19677),.A(g17096));
  NOT NOT1_6691(.VSS(VSS),.VDD(VDD),.Y(I18280),.A(g12951));
  NOT NOT1_6692(.VSS(VSS),.VDD(VDD),.Y(g12490),.A(I15316));
  NOT NOT1_6693(.VSS(VSS),.VDD(VDD),.Y(g17512),.A(g12983));
  NOT NOT1_6694(.VSS(VSS),.VDD(VDD),.Y(I17679),.A(g13416));
  NOT NOT1_6695(.VSS(VSS),.VDD(VDD),.Y(g21413),.A(g15585));
  NOT NOT1_6696(.VSS(VSS),.VDD(VDD),.Y(g9299),.A(g5124));
  NOT NOT1_6697(.VSS(VSS),.VDD(VDD),.Y(I15788),.A(g10430));
  NOT NOT1_6698(.VSS(VSS),.VDD(VDD),.Y(g23413),.A(g21012));
  NOT NOT1_6699(.VSS(VSS),.VDD(VDD),.Y(g27956),.A(I26466));
  NOT NOT1_6700(.VSS(VSS),.VDD(VDD),.Y(g32849),.A(g31021));
  NOT NOT1_6701(.VSS(VSS),.VDD(VDD),.Y(g9547),.A(g2735));
  NOT NOT1_6702(.VSS(VSS),.VDD(VDD),.Y(g10368),.A(g6887));
  NOT NOT1_6703(.VSS(VSS),.VDD(VDD),.Y(g32940),.A(g31376));
  NOT NOT1_6704(.VSS(VSS),.VDD(VDD),.Y(g7379),.A(g2299));
  NOT NOT1_6705(.VSS(VSS),.VDD(VDD),.Y(g8400),.A(g4836));
  NOT NOT1_6706(.VSS(VSS),.VDD(VDD),.Y(g11724),.A(I14593));
  NOT NOT1_6707(.VSS(VSS),.VDD(VDD),.Y(I17188),.A(g13782));
  NOT NOT1_6708(.VSS(VSS),.VDD(VDD),.Y(g31809),.A(g29385));
  NOT NOT1_6709(.VSS(VSS),.VDD(VDD),.Y(I12487),.A(g3443));
  NOT NOT1_6710(.VSS(VSS),.VDD(VDD),.Y(g11325),.A(g7543));
  NOT NOT1_6711(.VSS(VSS),.VDD(VDD),.Y(g20071),.A(g16826));
  NOT NOT1_6712(.VSS(VSS),.VDD(VDD),.Y(g32848),.A(g30825));
  NOT NOT1_6713(.VSS(VSS),.VDD(VDD),.Y(g9892),.A(g6428));
  NOT NOT1_6714(.VSS(VSS),.VDD(VDD),.Y(g24071),.A(g20841));
  NOT NOT1_6715(.VSS(VSS),.VDD(VDD),.Y(g11829),.A(I14653));
  NOT NOT1_6716(.VSS(VSS),.VDD(VDD),.Y(g12889),.A(g10396));
  NOT NOT1_6717(.VSS(VSS),.VDD(VDD),.Y(g11920),.A(I14730));
  NOT NOT1_6718(.VSS(VSS),.VDD(VDD),.Y(I11632),.A(g16));
  NOT NOT1_6719(.VSS(VSS),.VDD(VDD),.Y(g20591),.A(g15509));
  NOT NOT1_6720(.VSS(VSS),.VDD(VDD),.Y(g25781),.A(g24510));
  NOT NOT1_6721(.VSS(VSS),.VDD(VDD),.Y(g10412),.A(g7072));
  NOT NOT1_6722(.VSS(VSS),.VDD(VDD),.Y(g20776),.A(g18008));
  NOT NOT1_6723(.VSS(VSS),.VDD(VDD),.Y(g20785),.A(I20846));
  NOT NOT1_6724(.VSS(VSS),.VDD(VDD),.Y(g31808),.A(g29385));
  NOT NOT1_6725(.VSS(VSS),.VDD(VDD),.Y(g32652),.A(g30735));
  NOT NOT1_6726(.VSS(VSS),.VDD(VDD),.Y(g32804),.A(g30735));
  NOT NOT1_6727(.VSS(VSS),.VDD(VDD),.Y(g14412),.A(I16564));
  NOT NOT1_6728(.VSS(VSS),.VDD(VDD),.Y(g7289),.A(g4382));
  NOT NOT1_6729(.VSS(VSS),.VDD(VDD),.Y(I12618),.A(g3338));
  NOT NOT1_6730(.VSS(VSS),.VDD(VDD),.Y(g12888),.A(g10395));
  NOT NOT1_6731(.VSS(VSS),.VDD(VDD),.Y(g26614),.A(g25426));
  NOT NOT1_6732(.VSS(VSS),.VDD(VDD),.Y(g10133),.A(g6049));
  NOT NOT1_6733(.VSS(VSS),.VDD(VDD),.Y(g20147),.A(g17328));
  NOT NOT1_6734(.VSS(VSS),.VDD(VDD),.Y(I17938),.A(g3676));
  NOT NOT1_6735(.VSS(VSS),.VDD(VDD),.Y(g34209),.A(I32170));
  NOT NOT1_6736(.VSS(VSS),.VDD(VDD),.Y(g7835),.A(g4125));
  NOT NOT1_6737(.VSS(VSS),.VDD(VDD),.Y(g24147),.A(g19402));
  NOT NOT1_6738(.VSS(VSS),.VDD(VDD),.Y(g10229),.A(g6736));
  NOT NOT1_6739(.VSS(VSS),.VDD(VDD),.Y(I18066),.A(g3317));
  NOT NOT1_6740(.VSS(VSS),.VDD(VDD),.Y(g12181),.A(g9478));
  NOT NOT1_6741(.VSS(VSS),.VDD(VDD),.Y(g26607),.A(g25382));
  NOT NOT1_6742(.VSS(VSS),.VDD(VDD),.Y(g17499),.A(g14885));
  NOT NOT1_6743(.VSS(VSS),.VDD(VDD),.Y(g22989),.A(g20453));
  NOT NOT1_6744(.VSS(VSS),.VDD(VDD),.Y(g23929),.A(g19147));
  NOT NOT1_6745(.VSS(VSS),.VDD(VDD),.Y(g17316),.A(I18293));
  NOT NOT1_6746(.VSS(VSS),.VDD(VDD),.Y(g11344),.A(g9015));
  NOT NOT1_6747(.VSS(VSS),.VDD(VDD),.Y(g34208),.A(g33838));
  NOT NOT1_6748(.VSS(VSS),.VDD(VDD),.Y(I14158),.A(g8806));
  NOT NOT1_6749(.VSS(VSS),.VDD(VDD),.Y(g19410),.A(g16449));
  NOT NOT1_6750(.VSS(VSS),.VDD(VDD),.Y(g24825),.A(g23204));
  NOT NOT1_6751(.VSS(VSS),.VDD(VDD),.Y(g22722),.A(I22031));
  NOT NOT1_6752(.VSS(VSS),.VDD(VDD),.Y(g17498),.A(g14688));
  NOT NOT1_6753(.VSS(VSS),.VDD(VDD),.Y(g22988),.A(g20391));
  NOT NOT1_6754(.VSS(VSS),.VDD(VDD),.Y(g8183),.A(g482));
  NOT NOT1_6755(.VSS(VSS),.VDD(VDD),.Y(g23020),.A(g19869));
  NOT NOT1_6756(.VSS(VSS),.VDD(VDD),.Y(I15682),.A(g12182));
  NOT NOT1_6757(.VSS(VSS),.VDD(VDD),.Y(g23928),.A(g21562));
  NOT NOT1_6758(.VSS(VSS),.VDD(VDD),.Y(g8608),.A(g278));
  NOT NOT1_6759(.VSS(VSS),.VDD(VDD),.Y(I18885),.A(g16643));
  NOT NOT1_6760(.VSS(VSS),.VDD(VDD),.Y(g30021),.A(g28994));
  NOT NOT1_6761(.VSS(VSS),.VDD(VDD),.Y(I32071),.A(g33665));
  NOT NOT1_6762(.VSS(VSS),.VDD(VDD),.Y(g19479),.A(g16449));
  NOT NOT1_6763(.VSS(VSS),.VDD(VDD),.Y(g19666),.A(g17188));
  NOT NOT1_6764(.VSS(VSS),.VDD(VDD),.Y(g6782),.A(I11632));
  NOT NOT1_6765(.VSS(VSS),.VDD(VDD),.Y(g25264),.A(g23828));
  NOT NOT1_6766(.VSS(VSS),.VDD(VDD),.Y(g16692),.A(g14170));
  NOT NOT1_6767(.VSS(VSS),.VDD(VDD),.Y(g25790),.A(g25027));
  NOT NOT1_6768(.VSS(VSS),.VDD(VDD),.Y(I29013),.A(g29705));
  NOT NOT1_6769(.VSS(VSS),.VDD(VDD),.Y(g25137),.A(g22432));
  NOT NOT1_6770(.VSS(VSS),.VDD(VDD),.Y(g9340),.A(I13094));
  NOT NOT1_6771(.VSS(VSS),.VDD(VDD),.Y(I13715),.A(g71));
  NOT NOT1_6772(.VSS(VSS),.VDD(VDD),.Y(g17056),.A(g13437));
  NOT NOT1_6773(.VSS(VSS),.VDD(VDD),.Y(I29214),.A(g30300));
  NOT NOT1_6774(.VSS(VSS),.VDD(VDD),.Y(g11291),.A(g7526));
  NOT NOT1_6775(.VSS(VSS),.VDD(VDD),.Y(I32591),.A(g34287));
  NOT NOT1_6776(.VSS(VSS),.VDD(VDD),.Y(g24172),.A(I23360));
  NOT NOT1_6777(.VSS(VSS),.VDD(VDD),.Y(g23046),.A(g20283));
  NOT NOT1_6778(.VSS(VSS),.VDD(VDD),.Y(g32962),.A(g30735));
  NOT NOT1_6779(.VSS(VSS),.VDD(VDD),.Y(g9478),.A(I13152));
  NOT NOT1_6780(.VSS(VSS),.VDD(VDD),.Y(I14823),.A(g8056));
  NOT NOT1_6781(.VSS(VSS),.VDD(VDD),.Y(g19478),.A(g16000));
  NOT NOT1_6782(.VSS(VSS),.VDD(VDD),.Y(g24996),.A(g22763));
  NOT NOT1_6783(.VSS(VSS),.VDD(VDD),.Y(g17611),.A(g14822));
  NOT NOT1_6784(.VSS(VSS),.VDD(VDD),.Y(g17722),.A(I18709));
  NOT NOT1_6785(.VSS(VSS),.VDD(VDD),.Y(g9907),.A(g1959));
  NOT NOT1_6786(.VSS(VSS),.VDD(VDD),.Y(g13173),.A(g10632));
  NOT NOT1_6787(.VSS(VSS),.VDD(VDD),.Y(g34913),.A(I33131));
  NOT NOT1_6788(.VSS(VSS),.VDD(VDD),.Y(g10582),.A(g7116));
  NOT NOT1_6789(.VSS(VSS),.VDD(VDD),.Y(I16755),.A(g12377));
  NOT NOT1_6790(.VSS(VSS),.VDD(VDD),.Y(I29207),.A(g30293));
  NOT NOT1_6791(.VSS(VSS),.VDD(VDD),.Y(g14582),.A(I16698));
  NOT NOT1_6792(.VSS(VSS),.VDD(VDD),.Y(g33874),.A(I31724));
  NOT NOT1_6793(.VSS(VSS),.VDD(VDD),.Y(g9959),.A(g6177));
  NOT NOT1_6794(.VSS(VSS),.VDD(VDD),.Y(g7674),.A(I12151));
  NOT NOT1_6795(.VSS(VSS),.VDD(VDD),.Y(g8977),.A(g4349));
  NOT NOT1_6796(.VSS(VSS),.VDD(VDD),.Y(g24367),.A(g22550));
  NOT NOT1_6797(.VSS(VSS),.VDD(VDD),.Y(g24394),.A(g22228));
  NOT NOT1_6798(.VSS(VSS),.VDD(VDD),.Y(I16770),.A(g6023));
  NOT NOT1_6799(.VSS(VSS),.VDD(VDD),.Y(g32500),.A(g30735));
  NOT NOT1_6800(.VSS(VSS),.VDD(VDD),.Y(g34436),.A(I32479));
  NOT NOT1_6801(.VSS(VSS),.VDD(VDD),.Y(g9517),.A(g6163));
  NOT NOT1_6802(.VSS(VSS),.VDD(VDD),.Y(g9690),.A(g732));
  NOT NOT1_6803(.VSS(VSS),.VDD(VDD),.Y(g17432),.A(I18379));
  NOT NOT1_6804(.VSS(VSS),.VDD(VDD),.Y(g23787),.A(g18997));
  NOT NOT1_6805(.VSS(VSS),.VDD(VDD),.Y(I27677),.A(g28156));
  NOT NOT1_6806(.VSS(VSS),.VDD(VDD),.Y(g29170),.A(g27907));
  NOT NOT1_6807(.VSS(VSS),.VDD(VDD),.Y(g32833),.A(g30825));
  NOT NOT1_6808(.VSS(VSS),.VDD(VDD),.Y(g18957),.A(I19734));
  NOT NOT1_6809(.VSS(VSS),.VDD(VDD),.Y(g21282),.A(I21019));
  NOT NOT1_6810(.VSS(VSS),.VDD(VDD),.Y(g16214),.A(g13437));
  NOT NOT1_6811(.VSS(VSS),.VDD(VDD),.Y(g17271),.A(I18270));
  NOT NOT1_6812(.VSS(VSS),.VDD(VDD),.Y(I32950),.A(g34713));
  NOT NOT1_6813(.VSS(VSS),.VDD(VDD),.Y(g23282),.A(g20330));
  NOT NOT1_6814(.VSS(VSS),.VDD(VDD),.Y(I26710),.A(g27511));
  NOT NOT1_6815(.VSS(VSS),.VDD(VDD),.Y(g7541),.A(g344));
  NOT NOT1_6816(.VSS(VSS),.VDD(VDD),.Y(g10627),.A(I13968));
  NOT NOT1_6817(.VSS(VSS),.VDD(VDD),.Y(I25105),.A(g25284));
  NOT NOT1_6818(.VSS(VSS),.VDD(VDD),.Y(g34320),.A(g34119));
  NOT NOT1_6819(.VSS(VSS),.VDD(VDD),.Y(g27089),.A(g26703));
  NOT NOT1_6820(.VSS(VSS),.VDD(VDD),.Y(g10379),.A(g6953));
  NOT NOT1_6821(.VSS(VSS),.VDD(VDD),.Y(g23302),.A(g20330));
  NOT NOT1_6822(.VSS(VSS),.VDD(VDD),.Y(I25743),.A(g25903));
  NOT NOT1_6823(.VSS(VSS),.VDD(VDD),.Y(g31665),.A(I29245));
  NOT NOT1_6824(.VSS(VSS),.VDD(VDD),.Y(g25209),.A(g22763));
  NOT NOT1_6825(.VSS(VSS),.VDD(VDD),.Y(g19580),.A(g16164));
  NOT NOT1_6826(.VSS(VSS),.VDD(VDD),.Y(g30593),.A(g29970));
  NOT NOT1_6827(.VSS(VSS),.VDD(VDD),.Y(g33665),.A(I31500));
  NOT NOT1_6828(.VSS(VSS),.VDD(VDD),.Y(g6998),.A(g4932));
  NOT NOT1_6829(.VSS(VSS),.VDD(VDD),.Y(g22199),.A(g19210));
  NOT NOT1_6830(.VSS(VSS),.VDD(VDD),.Y(g34530),.A(I32591));
  NOT NOT1_6831(.VSS(VSS),.VDD(VDD),.Y(g10112),.A(g1988));
  NOT NOT1_6832(.VSS(VSS),.VDD(VDD),.Y(g34593),.A(I32687));
  NOT NOT1_6833(.VSS(VSS),.VDD(VDD),.Y(g7132),.A(g4558));
  NOT NOT1_6834(.VSS(VSS),.VDD(VDD),.Y(g12546),.A(g8740));
  NOT NOT1_6835(.VSS(VSS),.VDD(VDD),.Y(I22470),.A(g21326));
  NOT NOT1_6836(.VSS(VSS),.VDD(VDD),.Y(g10050),.A(g6336));
  NOT NOT1_6837(.VSS(VSS),.VDD(VDD),.Y(g27088),.A(g26694));
  NOT NOT1_6838(.VSS(VSS),.VDD(VDD),.Y(g18562),.A(I19384));
  NOT NOT1_6839(.VSS(VSS),.VDD(VDD),.Y(g34346),.A(g34162));
  NOT NOT1_6840(.VSS(VSS),.VDD(VDD),.Y(g10378),.A(g6926));
  NOT NOT1_6841(.VSS(VSS),.VDD(VDD),.Y(g25208),.A(g22763));
  NOT NOT1_6842(.VSS(VSS),.VDD(VDD),.Y(g30565),.A(I28832));
  NOT NOT1_6843(.VSS(VSS),.VDD(VDD),.Y(g7153),.A(g5373));
  NOT NOT1_6844(.VSS(VSS),.VDD(VDD),.Y(g7680),.A(g4108));
  NOT NOT1_6845(.VSS(VSS),.VDD(VDD),.Y(g8451),.A(g4057));
  NOT NOT1_6846(.VSS(VSS),.VDD(VDD),.Y(g22198),.A(g19147));
  NOT NOT1_6847(.VSS(VSS),.VDD(VDD),.Y(g22529),.A(g19549));
  NOT NOT1_6848(.VSS(VSS),.VDD(VDD),.Y(g34122),.A(I32059));
  NOT NOT1_6849(.VSS(VSS),.VDD(VDD),.Y(g15799),.A(g13110));
  NOT NOT1_6850(.VSS(VSS),.VDD(VDD),.Y(I21831),.A(g19127));
  NOT NOT1_6851(.VSS(VSS),.VDD(VDD),.Y(g13506),.A(g10808));
  NOT NOT1_6852(.VSS(VSS),.VDD(VDD),.Y(g12088),.A(g7701));
  NOT NOT1_6853(.VSS(VSS),.VDD(VDD),.Y(g13028),.A(I15650));
  NOT NOT1_6854(.VSS(VSS),.VDD(VDD),.Y(g20446),.A(g15224));
  NOT NOT1_6855(.VSS(VSS),.VDD(VDD),.Y(g10386),.A(g6982));
  NOT NOT1_6856(.VSS(VSS),.VDD(VDD),.Y(g29194),.A(I27492));
  NOT NOT1_6857(.VSS(VSS),.VDD(VDD),.Y(g9915),.A(g2583));
  NOT NOT1_6858(.VSS(VSS),.VDD(VDD),.Y(g12860),.A(g10368));
  NOT NOT1_6859(.VSS(VSS),.VDD(VDD),.Y(g22528),.A(g19801));
  NOT NOT1_6860(.VSS(VSS),.VDD(VDD),.Y(g6850),.A(g2704));
  NOT NOT1_6861(.VSS(VSS),.VDD(VDD),.Y(g14386),.A(I16544));
  NOT NOT1_6862(.VSS(VSS),.VDD(VDD),.Y(g23769),.A(g19074));
  NOT NOT1_6863(.VSS(VSS),.VDD(VDD),.Y(I11980),.A(g66));
  NOT NOT1_6864(.VSS(VSS),.VDD(VDD),.Y(g22330),.A(g19801));
  NOT NOT1_6865(.VSS(VSS),.VDD(VDD),.Y(I13889),.A(g7598));
  NOT NOT1_6866(.VSS(VSS),.VDD(VDD),.Y(g25542),.A(g22763));
  NOT NOT1_6867(.VSS(VSS),.VDD(VDD),.Y(g7802),.A(g324));
  NOT NOT1_6868(.VSS(VSS),.VDD(VDD),.Y(g20059),.A(g17302));
  NOT NOT1_6869(.VSS(VSS),.VDD(VDD),.Y(g32613),.A(g30673));
  NOT NOT1_6870(.VSS(VSS),.VDD(VDD),.Y(g8146),.A(g1760));
  NOT NOT1_6871(.VSS(VSS),.VDD(VDD),.Y(g10096),.A(g5767));
  NOT NOT1_6872(.VSS(VSS),.VDD(VDD),.Y(g20025),.A(g17271));
  NOT NOT1_6873(.VSS(VSS),.VDD(VDD),.Y(g8346),.A(g3845));
  NOT NOT1_6874(.VSS(VSS),.VDD(VDD),.Y(g24059),.A(g21193));
  NOT NOT1_6875(.VSS(VSS),.VDD(VDD),.Y(g33454),.A(I30980));
  NOT NOT1_6876(.VSS(VSS),.VDD(VDD),.Y(g14096),.A(I16328));
  NOT NOT1_6877(.VSS(VSS),.VDD(VDD),.Y(g24025),.A(g21256));
  NOT NOT1_6878(.VSS(VSS),.VDD(VDD),.Y(g9214),.A(g617));
  NOT NOT1_6879(.VSS(VSS),.VDD(VDD),.Y(g17529),.A(g15039));
  NOT NOT1_6880(.VSS(VSS),.VDD(VDD),.Y(g20540),.A(g16646));
  NOT NOT1_6881(.VSS(VSS),.VDD(VDD),.Y(g12497),.A(g9780));
  NOT NOT1_6882(.VSS(VSS),.VDD(VDD),.Y(g30292),.A(g28736));
  NOT NOT1_6883(.VSS(VSS),.VDD(VDD),.Y(I16898),.A(g10615));
  NOT NOT1_6884(.VSS(VSS),.VDD(VDD),.Y(g23768),.A(g18997));
  NOT NOT1_6885(.VSS(VSS),.VDD(VDD),.Y(I12884),.A(g4213));
  NOT NOT1_6886(.VSS(VSS),.VDD(VDD),.Y(I22467),.A(g19662));
  NOT NOT1_6887(.VSS(VSS),.VDD(VDD),.Y(g20058),.A(g16782));
  NOT NOT1_6888(.VSS(VSS),.VDD(VDD),.Y(g24540),.A(g22942));
  NOT NOT1_6889(.VSS(VSS),.VDD(VDD),.Y(g33712),.A(I31561));
  NOT NOT1_6890(.VSS(VSS),.VDD(VDD),.Y(I26356),.A(g26843));
  NOT NOT1_6891(.VSS(VSS),.VDD(VDD),.Y(I18307),.A(g12977));
  NOT NOT1_6892(.VSS(VSS),.VDD(VDD),.Y(g32947),.A(g31376));
  NOT NOT1_6893(.VSS(VSS),.VDD(VDD),.Y(g19531),.A(g16816));
  NOT NOT1_6894(.VSS(VSS),.VDD(VDD),.Y(g24058),.A(g20982));
  NOT NOT1_6895(.VSS(VSS),.VDD(VDD),.Y(g22869),.A(g20875));
  NOT NOT1_6896(.VSS(VSS),.VDD(VDD),.Y(g17528),.A(g14940));
  NOT NOT1_6897(.VSS(VSS),.VDD(VDD),.Y(g7558),.A(I12041));
  NOT NOT1_6898(.VSS(VSS),.VDD(VDD),.Y(g32605),.A(g30614));
  NOT NOT1_6899(.VSS(VSS),.VDD(VDD),.Y(g8696),.A(g3347));
  NOT NOT1_6900(.VSS(VSS),.VDD(VDD),.Y(g34409),.A(g34145));
  NOT NOT1_6901(.VSS(VSS),.VDD(VDD),.Y(I21722),.A(g19264));
  NOT NOT1_6902(.VSS(VSS),.VDD(VDD),.Y(g22868),.A(g20453));
  NOT NOT1_6903(.VSS(VSS),.VDD(VDD),.Y(I16521),.A(g10430));
  NOT NOT1_6904(.VSS(VSS),.VDD(VDD),.Y(g17764),.A(I18758));
  NOT NOT1_6905(.VSS(VSS),.VDD(VDD),.Y(I12666),.A(g4040));
  NOT NOT1_6906(.VSS(VSS),.VDD(VDD),.Y(g10429),.A(g7148));
  NOT NOT1_6907(.VSS(VSS),.VDD(VDD),.Y(g11927),.A(g10207));
  NOT NOT1_6908(.VSS(VSS),.VDD(VDD),.Y(g23881),.A(g19277));
  NOT NOT1_6909(.VSS(VSS),.VDD(VDD),.Y(g10857),.A(g8712));
  NOT NOT1_6910(.VSS(VSS),.VDD(VDD),.Y(g32812),.A(g30825));
  NOT NOT1_6911(.VSS(VSS),.VDD(VDD),.Y(g25073),.A(I24237));
  NOT NOT1_6912(.VSS(VSS),.VDD(VDD),.Y(g32463),.A(g31566));
  NOT NOT1_6913(.VSS(VSS),.VDD(VDD),.Y(g16100),.A(I17471));
  NOT NOT1_6914(.VSS(VSS),.VDD(VDD),.Y(I32446),.A(g34127));
  NOT NOT1_6915(.VSS(VSS),.VDD(VDD),.Y(g19676),.A(g17062));
  NOT NOT1_6916(.VSS(VSS),.VDD(VDD),.Y(g19685),.A(g16987));
  NOT NOT1_6917(.VSS(VSS),.VDD(VDD),.Y(g31239),.A(g29916));
  NOT NOT1_6918(.VSS(VSS),.VDD(VDD),.Y(g25274),.A(g22763));
  NOT NOT1_6919(.VSS(VSS),.VDD(VDD),.Y(g24044),.A(g21127));
  NOT NOT1_6920(.VSS(VSS),.VDD(VDD),.Y(g16771),.A(g14018));
  NOT NOT1_6921(.VSS(VSS),.VDD(VDD),.Y(g34408),.A(g34144));
  NOT NOT1_6922(.VSS(VSS),.VDD(VDD),.Y(I22419),.A(g19638));
  NOT NOT1_6923(.VSS(VSS),.VDD(VDD),.Y(g19373),.A(g16449));
  NOT NOT1_6924(.VSS(VSS),.VDD(VDD),.Y(g26575),.A(g25268));
  NOT NOT1_6925(.VSS(VSS),.VDD(VDD),.Y(g10428),.A(g9631));
  NOT NOT1_6926(.VSS(VSS),.VDD(VDD),.Y(g32951),.A(g31021));
  NOT NOT1_6927(.VSS(VSS),.VDD(VDD),.Y(g32972),.A(g31710));
  NOT NOT1_6928(.VSS(VSS),.VDD(VDD),.Y(g16235),.A(g13437));
  NOT NOT1_6929(.VSS(VSS),.VDD(VDD),.Y(g32033),.A(g30929));
  NOT NOT1_6930(.VSS(VSS),.VDD(VDD),.Y(I32059),.A(g33648));
  NOT NOT1_6931(.VSS(VSS),.VDD(VDD),.Y(g8508),.A(g3827));
  NOT NOT1_6932(.VSS(VSS),.VDD(VDD),.Y(g19654),.A(g16931));
  NOT NOT1_6933(.VSS(VSS),.VDD(VDD),.Y(I31361),.A(g33120));
  NOT NOT1_6934(.VSS(VSS),.VDD(VDD),.Y(g9402),.A(g6209));
  NOT NOT1_6935(.VSS(VSS),.VDD(VDD),.Y(g9824),.A(g1825));
  NOT NOT1_6936(.VSS(VSS),.VDD(VDD),.Y(g8944),.A(g370));
  NOT NOT1_6937(.VSS(VSS),.VDD(VDD),.Y(g8240),.A(g1333));
  NOT NOT1_6938(.VSS(VSS),.VDD(VDD),.Y(g18661),.A(I19487));
  NOT NOT1_6939(.VSS(VSS),.VDD(VDD),.Y(g20902),.A(I20870));
  NOT NOT1_6940(.VSS(VSS),.VDD(VDD),.Y(g18895),.A(g16000));
  NOT NOT1_6941(.VSS(VSS),.VDD(VDD),.Y(g19800),.A(g17096));
  NOT NOT1_6942(.VSS(VSS),.VDD(VDD),.Y(I18341),.A(g14308));
  NOT NOT1_6943(.VSS(VSS),.VDD(VDD),.Y(g19417),.A(g17178));
  NOT NOT1_6944(.VSS(VSS),.VDD(VDD),.Y(g21662),.A(g16540));
  NOT NOT1_6945(.VSS(VSS),.VDD(VDD),.Y(g24377),.A(g22594));
  NOT NOT1_6946(.VSS(VSS),.VDD(VDD),.Y(g7092),.A(g6483));
  NOT NOT1_6947(.VSS(VSS),.VDD(VDD),.Y(I31500),.A(g33176));
  NOT NOT1_6948(.VSS(VSS),.VDD(VDD),.Y(g24120),.A(g19984));
  NOT NOT1_6949(.VSS(VSS),.VDD(VDD),.Y(g23027),.A(g20391));
  NOT NOT1_6950(.VSS(VSS),.VDD(VDD),.Y(g32795),.A(g31327));
  NOT NOT1_6951(.VSS(VSS),.VDD(VDD),.Y(g25034),.A(g23695));
  NOT NOT1_6952(.VSS(VSS),.VDD(VDD),.Y(I23342),.A(g23299));
  NOT NOT1_6953(.VSS(VSS),.VDD(VDD),.Y(g17709),.A(g14761));
  NOT NOT1_6954(.VSS(VSS),.VDD(VDD),.Y(g33382),.A(g32033));
  NOT NOT1_6955(.VSS(VSS),.VDD(VDD),.Y(I12580),.A(g1239));
  NOT NOT1_6956(.VSS(VSS),.VDD(VDD),.Y(g8443),.A(g3736));
  NOT NOT1_6957(.VSS(VSS),.VDD(VDD),.Y(g19334),.A(I19818));
  NOT NOT1_6958(.VSS(VSS),.VDD(VDD),.Y(g20146),.A(g17533));
  NOT NOT1_6959(.VSS(VSS),.VDD(VDD),.Y(g20738),.A(g15483));
  NOT NOT1_6960(.VSS(VSS),.VDD(VDD),.Y(I18180),.A(g13605));
  NOT NOT1_6961(.VSS(VSS),.VDD(VDD),.Y(g25641),.A(I24784));
  NOT NOT1_6962(.VSS(VSS),.VDD(VDD),.Y(g20562),.A(g17955));
  NOT NOT1_6963(.VSS(VSS),.VDD(VDD),.Y(g9590),.A(g1882));
  NOT NOT1_6964(.VSS(VSS),.VDD(VDD),.Y(g21249),.A(g15509));
  NOT NOT1_6965(.VSS(VSS),.VDD(VDD),.Y(I15981),.A(g11290));
  NOT NOT1_6966(.VSS(VSS),.VDD(VDD),.Y(g24146),.A(g19422));
  NOT NOT1_6967(.VSS(VSS),.VDD(VDD),.Y(g6986),.A(g4743));
  NOT NOT1_6968(.VSS(VSS),.VDD(VDD),.Y(g23249),.A(g21070));
  NOT NOT1_6969(.VSS(VSS),.VDD(VDD),.Y(I14687),.A(g7753));
  NOT NOT1_6970(.VSS(VSS),.VDD(VDD),.Y(g11770),.A(I14619));
  NOT NOT1_6971(.VSS(VSS),.VDD(VDD),.Y(I21199),.A(g17501));
  NOT NOT1_6972(.VSS(VSS),.VDD(VDD),.Y(I30998),.A(g32453));
  NOT NOT1_6973(.VSS(VSS),.VDD(VDD),.Y(g20699),.A(g17873));
  NOT NOT1_6974(.VSS(VSS),.VDD(VDD),.Y(g16515),.A(g13486));
  NOT NOT1_6975(.VSS(VSS),.VDD(VDD),.Y(g10504),.A(g8763));
  NOT NOT1_6976(.VSS(VSS),.VDD(VDD),.Y(g11981),.A(I14823));
  NOT NOT1_6977(.VSS(VSS),.VDD(VDD),.Y(g9657),.A(g2763));
  NOT NOT1_6978(.VSS(VSS),.VDD(VDD),.Y(g12968),.A(g11793));
  NOT NOT1_6979(.VSS(VSS),.VDD(VDD),.Y(g17471),.A(g14454));
  NOT NOT1_6980(.VSS(VSS),.VDD(VDD),.Y(g25153),.A(g23733));
  NOT NOT1_6981(.VSS(VSS),.VDD(VDD),.Y(I26448),.A(g26860));
  NOT NOT1_6982(.VSS(VSS),.VDD(VDD),.Y(g8316),.A(g2351));
  NOT NOT1_6983(.VSS(VSS),.VDD(VDD),.Y(g17087),.A(g14321));
  NOT NOT1_6984(.VSS(VSS),.VDD(VDD),.Y(g23482),.A(g18833));
  NOT NOT1_6985(.VSS(VSS),.VDD(VDD),.Y(I25552),.A(g25240));
  NOT NOT1_6986(.VSS(VSS),.VDD(VDD),.Y(g32514),.A(g30735));
  NOT NOT1_6987(.VSS(VSS),.VDD(VDD),.Y(I18734),.A(g6373));
  NOT NOT1_6988(.VSS(VSS),.VDD(VDD),.Y(g24699),.A(g23047));
  NOT NOT1_6989(.VSS(VSS),.VDD(VDD),.Y(g21248),.A(g15224));
  NOT NOT1_6990(.VSS(VSS),.VDD(VDD),.Y(g14504),.A(g12361));
  NOT NOT1_6991(.VSS(VSS),.VDD(VDD),.Y(g19762),.A(g16326));
  NOT NOT1_6992(.VSS(VSS),.VDD(VDD),.Y(g23248),.A(g20924));
  NOT NOT1_6993(.VSS(VSS),.VDD(VDD),.Y(g19964),.A(g17200));
  NOT NOT1_6994(.VSS(VSS),.VDD(VDD),.Y(I22589),.A(g21340));
  NOT NOT1_6995(.VSS(VSS),.VDD(VDD),.Y(g20698),.A(g17873));
  NOT NOT1_6996(.VSS(VSS),.VDD(VDD),.Y(g27527),.A(I26195));
  NOT NOT1_6997(.VSS(VSS),.VDD(VDD),.Y(g25409),.A(g22228));
  NOT NOT1_6998(.VSS(VSS),.VDD(VDD),.Y(g34575),.A(I32651));
  NOT NOT1_6999(.VSS(VSS),.VDD(VDD),.Y(I25779),.A(g26424));
  NOT NOT1_7000(.VSS(VSS),.VDD(VDD),.Y(g32507),.A(g30735));
  NOT NOT1_7001(.VSS(VSS),.VDD(VDD),.Y(g9556),.A(g5448));
  NOT NOT1_7002(.VSS(VSS),.VDD(VDD),.Y(I18839),.A(g13716));
  NOT NOT1_7003(.VSS(VSS),.VDD(VDD),.Y(g23003),.A(I22180));
  NOT NOT1_7004(.VSS(VSS),.VDD(VDD),.Y(g8565),.A(g3802));
  NOT NOT1_7005(.VSS(VSS),.VDD(VDD),.Y(g21204),.A(g15656));
  NOT NOT1_7006(.VSS(VSS),.VDD(VDD),.Y(g33637),.A(I31466));
  NOT NOT1_7007(.VSS(VSS),.VDD(VDD),.Y(g29177),.A(g27937));
  NOT NOT1_7008(.VSS(VSS),.VDD(VDD),.Y(g30327),.A(I28582));
  NOT NOT1_7009(.VSS(VSS),.VDD(VDD),.Y(g33935),.A(I31817));
  NOT NOT1_7010(.VSS(VSS),.VDD(VDD),.Y(g34711),.A(g34559));
  NOT NOT1_7011(.VSS(VSS),.VDD(VDD),.Y(g12870),.A(g10374));
  NOT NOT1_7012(.VSS(VSS),.VDD(VDD),.Y(I11860),.A(g43));
  NOT NOT1_7013(.VSS(VSS),.VDD(VDD),.Y(g25136),.A(g22457));
  NOT NOT1_7014(.VSS(VSS),.VDD(VDD),.Y(g34327),.A(g34108));
  NOT NOT1_7015(.VSS(VSS),.VDD(VDD),.Y(I18667),.A(g6661));
  NOT NOT1_7016(.VSS(VSS),.VDD(VDD),.Y(I18694),.A(g5666));
  NOT NOT1_7017(.VSS(VSS),.VDD(VDD),.Y(g32421),.A(g31213));
  NOT NOT1_7018(.VSS(VSS),.VDD(VDD),.Y(I23330),.A(g22658));
  NOT NOT1_7019(.VSS(VSS),.VDD(VDD),.Y(I23393),.A(g23414));
  NOT NOT1_7020(.VSS(VSS),.VDD(VDD),.Y(g10129),.A(g5352));
  NOT NOT1_7021(.VSS(VSS),.VDD(VDD),.Y(I29441),.A(g30917));
  NOT NOT1_7022(.VSS(VSS),.VDD(VDD),.Y(g11845),.A(I14663));
  NOT NOT1_7023(.VSS(VSS),.VDD(VDD),.Y(g9064),.A(g4983));
  NOT NOT1_7024(.VSS(VSS),.VDD(VDD),.Y(I18131),.A(g13350));
  NOT NOT1_7025(.VSS(VSS),.VDD(VDD),.Y(g8681),.A(g763));
  NOT NOT1_7026(.VSS(VSS),.VDD(VDD),.Y(g10002),.A(g6195));
  NOT NOT1_7027(.VSS(VSS),.VDD(VDD),.Y(I25786),.A(g26424));
  NOT NOT1_7028(.VSS(VSS),.VDD(VDD),.Y(g10057),.A(g6455));
  NOT NOT1_7029(.VSS(VSS),.VDD(VDD),.Y(g9899),.A(g6513));
  NOT NOT1_7030(.VSS(VSS),.VDD(VDD),.Y(I32645),.A(g34367));
  NOT NOT1_7031(.VSS(VSS),.VDD(VDD),.Y(g7262),.A(g5723));
  NOT NOT1_7032(.VSS(VSS),.VDD(VDD),.Y(g24366),.A(g22594));
  NOT NOT1_7033(.VSS(VSS),.VDD(VDD),.Y(g20632),.A(g15171));
  NOT NOT1_7034(.VSS(VSS),.VDD(VDD),.Y(I15633),.A(g12074));
  NOT NOT1_7035(.VSS(VSS),.VDD(VDD),.Y(I32699),.A(g34569));
  NOT NOT1_7036(.VSS(VSS),.VDD(VDD),.Y(I33273),.A(g34984));
  NOT NOT1_7037(.VSS(VSS),.VDD(VDD),.Y(g30606),.A(I28866));
  NOT NOT1_7038(.VSS(VSS),.VDD(VDD),.Y(g8697),.A(g3694));
  NOT NOT1_7039(.VSS(VSS),.VDD(VDD),.Y(I33106),.A(g34855));
  NOT NOT1_7040(.VSS(VSS),.VDD(VDD),.Y(I14668),.A(g7753));
  NOT NOT1_7041(.VSS(VSS),.VDD(VDD),.Y(I25356),.A(g24374));
  NOT NOT1_7042(.VSS(VSS),.VDD(VDD),.Y(g19543),.A(g16349));
  NOT NOT1_7043(.VSS(VSS),.VDD(VDD),.Y(g30303),.A(g28786));
  NOT NOT1_7044(.VSS(VSS),.VDD(VDD),.Y(g8914),.A(g4264));
  NOT NOT1_7045(.VSS(VSS),.VDD(VDD),.Y(I19796),.A(g17870));
  NOT NOT1_7046(.VSS(VSS),.VDD(VDD),.Y(g17602),.A(g14962));
  NOT NOT1_7047(.VSS(VSS),.VDD(VDD),.Y(g12867),.A(g10375));
  NOT NOT1_7048(.VSS(VSS),.VDD(VDD),.Y(g12894),.A(g10401));
  NOT NOT1_7049(.VSS(VSS),.VDD(VDD),.Y(I17401),.A(g13394));
  NOT NOT1_7050(.VSS(VSS),.VDD(VDD),.Y(g16584),.A(g13920));
  NOT NOT1_7051(.VSS(VSS),.VDD(VDD),.Y(g17774),.A(g14902));
  NOT NOT1_7052(.VSS(VSS),.VDD(VDD),.Y(g23647),.A(g18833));
  NOT NOT1_7053(.VSS(VSS),.VDD(VDD),.Y(g18889),.A(g15509));
  NOT NOT1_7054(.VSS(VSS),.VDD(VDD),.Y(g17955),.A(I18865));
  NOT NOT1_7055(.VSS(VSS),.VDD(VDD),.Y(g18980),.A(g16136));
  NOT NOT1_7056(.VSS(VSS),.VDD(VDD),.Y(g32541),.A(g30673));
  NOT NOT1_7057(.VSS(VSS),.VDD(VDD),.Y(g7623),.A(I12103));
  NOT NOT1_7058(.VSS(VSS),.VDD(VDD),.Y(g10323),.A(I13744));
  NOT NOT1_7059(.VSS(VSS),.VDD(VDD),.Y(g23945),.A(g21611));
  NOT NOT1_7060(.VSS(VSS),.VDD(VDD),.Y(g16206),.A(g13437));
  NOT NOT1_7061(.VSS(VSS),.VDD(VDD),.Y(I25380),.A(g24481));
  NOT NOT1_7062(.VSS(VSS),.VDD(VDD),.Y(g18095),.A(I18891));
  NOT NOT1_7063(.VSS(VSS),.VDD(VDD),.Y(g23356),.A(g21070));
  NOT NOT1_7064(.VSS(VSS),.VDD(VDD),.Y(g32473),.A(g31070));
  NOT NOT1_7065(.VSS(VSS),.VDD(VDD),.Y(I31463),.A(g33318));
  NOT NOT1_7066(.VSS(VSS),.VDD(VDD),.Y(g19908),.A(g16540));
  NOT NOT1_7067(.VSS(VSS),.VDD(VDD),.Y(g22171),.A(g18882));
  NOT NOT1_7068(.VSS(VSS),.VDD(VDD),.Y(g13191),.A(I15788));
  NOT NOT1_7069(.VSS(VSS),.VDD(VDD),.Y(g26840),.A(I25562));
  NOT NOT1_7070(.VSS(VSS),.VDD(VDD),.Y(g20661),.A(g15171));
  NOT NOT1_7071(.VSS(VSS),.VDD(VDD),.Y(I12654),.A(g1585));
  NOT NOT1_7072(.VSS(VSS),.VDD(VDD),.Y(g21380),.A(g17955));
  NOT NOT1_7073(.VSS(VSS),.VDD(VDD),.Y(g10533),.A(g8795));
  NOT NOT1_7074(.VSS(VSS),.VDD(VDD),.Y(g20547),.A(g15224));
  NOT NOT1_7075(.VSS(VSS),.VDD(VDD),.Y(g23999),.A(g21468));
  NOT NOT1_7076(.VSS(VSS),.VDD(VDD),.Y(g32789),.A(g30735));
  NOT NOT1_7077(.VSS(VSS),.VDD(VDD),.Y(g18888),.A(g15426));
  NOT NOT1_7078(.VSS(VSS),.VDD(VDD),.Y(g23380),.A(g20619));
  NOT NOT1_7079(.VSS(VSS),.VDD(VDD),.Y(g33729),.A(I31586));
  NOT NOT1_7080(.VSS(VSS),.VDD(VDD),.Y(I18443),.A(g13027));
  NOT NOT1_7081(.VSS(VSS),.VDD(VDD),.Y(g19569),.A(g16349));
  NOT NOT1_7082(.VSS(VSS),.VDD(VDD),.Y(I14424),.A(g4005));
  NOT NOT1_7083(.VSS(VSS),.VDD(VDD),.Y(I14016),.A(g9104));
  NOT NOT1_7084(.VSS(VSS),.VDD(VDD),.Y(I17118),.A(g14363));
  NOT NOT1_7085(.VSS(VSS),.VDD(VDD),.Y(g16725),.A(g13963));
  NOT NOT1_7086(.VSS(VSS),.VDD(VDD),.Y(I22748),.A(g19458));
  NOT NOT1_7087(.VSS(VSS),.VDD(VDD),.Y(g13521),.A(g11357));
  NOT NOT1_7088(.VSS(VSS),.VDD(VDD),.Y(g22994),.A(g20436));
  NOT NOT1_7089(.VSS(VSS),.VDD(VDD),.Y(g34982),.A(I33246));
  NOT NOT1_7090(.VSS(VSS),.VDD(VDD),.Y(g32788),.A(g31327));
  NOT NOT1_7091(.VSS(VSS),.VDD(VDD),.Y(g32724),.A(g30735));
  NOT NOT1_7092(.VSS(VSS),.VDD(VDD),.Y(g19747),.A(g17015));
  NOT NOT1_7093(.VSS(VSS),.VDD(VDD),.Y(g23233),.A(g21037));
  NOT NOT1_7094(.VSS(VSS),.VDD(VDD),.Y(g21182),.A(g15509));
  NOT NOT1_7095(.VSS(VSS),.VDD(VDD),.Y(g6789),.A(I11635));
  NOT NOT1_7096(.VSS(VSS),.VDD(VDD),.Y(g11832),.A(g8011));
  NOT NOT1_7097(.VSS(VSS),.VDD(VDD),.Y(g23182),.A(g21389));
  NOT NOT1_7098(.VSS(VSS),.VDD(VDD),.Y(g20715),.A(g15277));
  NOT NOT1_7099(.VSS(VSS),.VDD(VDD),.Y(g23651),.A(g20655));
  NOT NOT1_7100(.VSS(VSS),.VDD(VDD),.Y(g32829),.A(g30937));
  NOT NOT1_7101(.VSS(VSS),.VDD(VDD),.Y(g28080),.A(I26581));
  NOT NOT1_7102(.VSS(VSS),.VDD(VDD),.Y(g32920),.A(g30825));
  NOT NOT1_7103(.VSS(VSS),.VDD(VDD),.Y(I18469),.A(g13809));
  NOT NOT1_7104(.VSS(VSS),.VDD(VDD),.Y(g32535),.A(g31554));
  NOT NOT1_7105(.VSS(VSS),.VDD(VDD),.Y(g25327),.A(g22161));
  NOT NOT1_7106(.VSS(VSS),.VDD(VDD),.Y(g32434),.A(g31189));
  NOT NOT1_7107(.VSS(VSS),.VDD(VDD),.Y(I14830),.A(g10141));
  NOT NOT1_7108(.VSS(VSS),.VDD(VDD),.Y(I21258),.A(g16540));
  NOT NOT1_7109(.VSS(VSS),.VDD(VDD),.Y(g24481),.A(I23684));
  NOT NOT1_7110(.VSS(VSS),.VDD(VDD),.Y(I14893),.A(g9819));
  NOT NOT1_7111(.VSS(VSS),.VDD(VDD),.Y(g25109),.A(g23666));
  NOT NOT1_7112(.VSS(VSS),.VDD(VDD),.Y(g12818),.A(g8792));
  NOT NOT1_7113(.VSS(VSS),.VDD(VDD),.Y(g20551),.A(g17302));
  NOT NOT1_7114(.VSS(VSS),.VDD(VDD),.Y(g20572),.A(g15833));
  NOT NOT1_7115(.VSS(VSS),.VDD(VDD),.Y(g9194),.A(g827));
  NOT NOT1_7116(.VSS(VSS),.VDD(VDD),.Y(g32828),.A(g31710));
  NOT NOT1_7117(.VSS(VSS),.VDD(VDD),.Y(g18931),.A(g16031));
  NOT NOT1_7118(.VSS(VSS),.VDD(VDD),.Y(g6987),.A(g4754));
  NOT NOT1_7119(.VSS(VSS),.VDD(VDD),.Y(g32946),.A(g31327));
  NOT NOT1_7120(.VSS(VSS),.VDD(VDD),.Y(g10232),.A(g4527));
  NOT NOT1_7121(.VSS(VSS),.VDD(VDD),.Y(I17276),.A(g13605));
  NOT NOT1_7122(.VSS(VSS),.VDD(VDD),.Y(g7285),.A(g4643));
  NOT NOT1_7123(.VSS(VSS),.VDD(VDD),.Y(g11861),.A(g8070));
  NOT NOT1_7124(.VSS(VSS),.VDD(VDD),.Y(g22919),.A(g21163));
  NOT NOT1_7125(.VSS(VSS),.VDD(VDD),.Y(g16744),.A(I17964));
  NOT NOT1_7126(.VSS(VSS),.VDD(VDD),.Y(I17704),.A(g13144));
  NOT NOT1_7127(.VSS(VSS),.VDD(VDD),.Y(g12978),.A(I15593));
  NOT NOT1_7128(.VSS(VSS),.VDD(VDD),.Y(g14232),.A(g11083));
  NOT NOT1_7129(.VSS(VSS),.VDD(VDD),.Y(g9731),.A(g5366));
  NOT NOT1_7130(.VSS(VSS),.VDD(VDD),.Y(g23331),.A(g20905));
  NOT NOT1_7131(.VSS(VSS),.VDD(VDD),.Y(I13968),.A(g7697));
  NOT NOT1_7132(.VSS(VSS),.VDD(VDD),.Y(I32547),.A(g34397));
  NOT NOT1_7133(.VSS(VSS),.VDD(VDD),.Y(g19751),.A(g16044));
  NOT NOT1_7134(.VSS(VSS),.VDD(VDD),.Y(I24839),.A(g24298));
  NOT NOT1_7135(.VSS(VSS),.VDD(VDD),.Y(g9489),.A(g2303));
  NOT NOT1_7136(.VSS(VSS),.VDD(VDD),.Y(g19772),.A(g17183));
  NOT NOT1_7137(.VSS(VSS),.VDD(VDD),.Y(g25283),.A(g22763));
  NOT NOT1_7138(.VSS(VSS),.VDD(VDD),.Y(g34840),.A(I33056));
  NOT NOT1_7139(.VSS(VSS),.VDD(VDD),.Y(g20127),.A(I20388));
  NOT NOT1_7140(.VSS(VSS),.VDD(VDD),.Y(I22177),.A(g21366));
  NOT NOT1_7141(.VSS(VSS),.VDD(VDD),.Y(g23449),.A(g18833));
  NOT NOT1_7142(.VSS(VSS),.VDD(VDD),.Y(g26483),.A(I25359));
  NOT NOT1_7143(.VSS(VSS),.VDD(VDD),.Y(g28753),.A(I27235));
  NOT NOT1_7144(.VSS(VSS),.VDD(VDD),.Y(g9557),.A(g5499));
  NOT NOT1_7145(.VSS(VSS),.VDD(VDD),.Y(g13926),.A(I16217));
  NOT NOT1_7146(.VSS(VSS),.VDD(VDD),.Y(g24127),.A(g19984));
  NOT NOT1_7147(.VSS(VSS),.VDD(VDD),.Y(g13045),.A(g11941));
  NOT NOT1_7148(.VSS(VSS),.VDD(VDD),.Y(g10261),.A(g4555));
  NOT NOT1_7149(.VSS(VSS),.VDD(VDD),.Y(I17808),.A(g13311));
  NOT NOT1_7150(.VSS(VSS),.VDD(VDD),.Y(g9071),.A(g2831));
  NOT NOT1_7151(.VSS(VSS),.VDD(VDD),.Y(g26862),.A(I25598));
  NOT NOT1_7152(.VSS(VSS),.VDD(VDD),.Y(g11388),.A(I14395));
  NOT NOT1_7153(.VSS(VSS),.VDD(VDD),.Y(g23897),.A(g19210));
  NOT NOT1_7154(.VSS(VSS),.VDD(VDD),.Y(g13099),.A(I15732));
  NOT NOT1_7155(.VSS(VSS),.VDD(VDD),.Y(g11324),.A(g7542));
  NOT NOT1_7156(.VSS(VSS),.VDD(VDD),.Y(g23448),.A(g21611));
  NOT NOT1_7157(.VSS(VSS),.VDD(VDD),.Y(g23961),.A(g19074));
  NOT NOT1_7158(.VSS(VSS),.VDD(VDD),.Y(g32682),.A(g30825));
  NOT NOT1_7159(.VSS(VSS),.VDD(VDD),.Y(g24490),.A(g22594));
  NOT NOT1_7160(.VSS(VSS),.VDD(VDD),.Y(I14705),.A(g7717));
  NOT NOT1_7161(.VSS(VSS),.VDD(VDD),.Y(g19638),.A(g17324));
  NOT NOT1_7162(.VSS(VSS),.VDD(VDD),.Y(I17101),.A(g14338));
  NOT NOT1_7163(.VSS(VSS),.VDD(VDD),.Y(g34192),.A(g33921));
  NOT NOT1_7164(.VSS(VSS),.VDD(VDD),.Y(I21810),.A(g20596));
  NOT NOT1_7165(.VSS(VSS),.VDD(VDD),.Y(I16629),.A(g11987));
  NOT NOT1_7166(.VSS(VSS),.VDD(VDD),.Y(g16652),.A(g13892));
  NOT NOT1_7167(.VSS(VSS),.VDD(VDD),.Y(g17010),.A(I18138));
  NOT NOT1_7168(.VSS(VSS),.VDD(VDD),.Y(g23505),.A(g21514));
  NOT NOT1_7169(.VSS(VSS),.VDD(VDD),.Y(I27543),.A(g28187));
  NOT NOT1_7170(.VSS(VSS),.VDD(VDD),.Y(g26326),.A(g24872));
  NOT NOT1_7171(.VSS(VSS),.VDD(VDD),.Y(g8922),.A(I12907));
  NOT NOT1_7172(.VSS(VSS),.VDD(VDD),.Y(g20385),.A(g18008));
  NOT NOT1_7173(.VSS(VSS),.VDD(VDD),.Y(I14679),.A(g9332));
  NOT NOT1_7174(.VSS(VSS),.VDD(VDD),.Y(g13251),.A(I15814));
  NOT NOT1_7175(.VSS(VSS),.VDD(VDD),.Y(I23375),.A(g23403));
  NOT NOT1_7176(.VSS(VSS),.VDD(VDD),.Y(g13272),.A(I15837));
  NOT NOT1_7177(.VSS(VSS),.VDD(VDD),.Y(g19416),.A(g15885));
  NOT NOT1_7178(.VSS(VSS),.VDD(VDD),.Y(g20103),.A(g17433));
  NOT NOT1_7179(.VSS(VSS),.VDD(VDD),.Y(g7424),.A(g2465));
  NOT NOT1_7180(.VSS(VSS),.VDD(VDD),.Y(g24376),.A(g22722));
  NOT NOT1_7181(.VSS(VSS),.VDD(VDD),.Y(g24385),.A(g22908));
  NOT NOT1_7182(.VSS(VSS),.VDD(VDD),.Y(g34522),.A(g34271));
  NOT NOT1_7183(.VSS(VSS),.VDD(VDD),.Y(g7809),.A(g4864));
  NOT NOT1_7184(.VSS(VSS),.VDD(VDD),.Y(I18143),.A(g13350));
  NOT NOT1_7185(.VSS(VSS),.VDD(VDD),.Y(g24103),.A(g21209));
  NOT NOT1_7186(.VSS(VSS),.VDD(VDD),.Y(g23026),.A(g20391));
  NOT NOT1_7187(.VSS(VSS),.VDD(VDD),.Y(g18088),.A(g13267));
  NOT NOT1_7188(.VSS(VSS),.VDD(VDD),.Y(g24980),.A(g22384));
  NOT NOT1_7189(.VSS(VSS),.VDD(VDD),.Y(I16246),.A(g3983));
  NOT NOT1_7190(.VSS(VSS),.VDD(VDD),.Y(I30971),.A(g32015));
  NOT NOT1_7191(.VSS(VSS),.VDD(VDD),.Y(I12117),.A(g586));
  NOT NOT1_7192(.VSS(VSS),.VDD(VDD),.Y(g24095),.A(g21209));
  NOT NOT1_7193(.VSS(VSS),.VDD(VDD),.Y(g26702),.A(g25309));
  NOT NOT1_7194(.VSS(VSS),.VDD(VDD),.Y(g17599),.A(g14794));
  NOT NOT1_7195(.VSS(VSS),.VDD(VDD),.Y(I12000),.A(g582));
  NOT NOT1_7196(.VSS(VSS),.VDD(VDD),.Y(g25174),.A(g23890));
  NOT NOT1_7197(.VSS(VSS),.VDD(VDD),.Y(g28696),.A(g27858));
  NOT NOT1_7198(.VSS(VSS),.VDD(VDD),.Y(g31653),.A(g29713));
  NOT NOT1_7199(.VSS(VSS),.VDD(VDD),.Y(g6991),.A(g4888));
  NOT NOT1_7200(.VSS(VSS),.VDD(VDD),.Y(g33653),.A(I31486));
  NOT NOT1_7201(.VSS(VSS),.VDD(VDD),.Y(I14939),.A(g10216));
  NOT NOT1_7202(.VSS(VSS),.VDD(VDD),.Y(g7231),.A(g5));
  NOT NOT1_7203(.VSS(VSS),.VDD(VDD),.Y(g20671),.A(g15509));
  NOT NOT1_7204(.VSS(VSS),.VDD(VDD),.Y(I17733),.A(g14844));
  NOT NOT1_7205(.VSS(VSS),.VDD(VDD),.Y(g27018),.A(I25750));
  NOT NOT1_7206(.VSS(VSS),.VDD(VDD),.Y(g31138),.A(g29778));
  NOT NOT1_7207(.VSS(VSS),.VDD(VDD),.Y(g32760),.A(g30735));
  NOT NOT1_7208(.VSS(VSS),.VDD(VDD),.Y(g17086),.A(g14297));
  NOT NOT1_7209(.VSS(VSS),.VDD(VDD),.Y(g24181),.A(I23387));
  NOT NOT1_7210(.VSS(VSS),.VDD(VDD),.Y(g7523),.A(g305));
  NOT NOT1_7211(.VSS(VSS),.VDD(VDD),.Y(g19579),.A(g16000));
  NOT NOT1_7212(.VSS(VSS),.VDD(VDD),.Y(g22159),.A(I21744));
  NOT NOT1_7213(.VSS(VSS),.VDD(VDD),.Y(g29941),.A(g28900));
  NOT NOT1_7214(.VSS(VSS),.VDD(VDD),.Y(g13140),.A(g10632));
  NOT NOT1_7215(.VSS(VSS),.VDD(VDD),.Y(g7643),.A(g4322));
  NOT NOT1_7216(.VSS(VSS),.VDD(VDD),.Y(I21792),.A(g21308));
  NOT NOT1_7217(.VSS(VSS),.VDD(VDD),.Y(I12568),.A(g5005));
  NOT NOT1_7218(.VSS(VSS),.VDD(VDD),.Y(g12018),.A(g9538));
  NOT NOT1_7219(.VSS(VSS),.VDD(VDD),.Y(I22009),.A(g21269));
  NOT NOT1_7220(.VSS(VSS),.VDD(VDD),.Y(g34553),.A(I32621));
  NOT NOT1_7221(.VSS(VSS),.VDD(VDD),.Y(g10499),.A(I13872));
  NOT NOT1_7222(.VSS(VSS),.VDD(VDD),.Y(I22665),.A(g21308));
  NOT NOT1_7223(.VSS(VSS),.VDD(VDD),.Y(I13581),.A(g6727));
  NOT NOT1_7224(.VSS(VSS),.VDD(VDD),.Y(I18168),.A(g13191));
  NOT NOT1_7225(.VSS(VSS),.VDD(VDD),.Y(I24278),.A(g23440));
  NOT NOT1_7226(.VSS(VSS),.VDD(VDD),.Y(I14267),.A(g7835));
  NOT NOT1_7227(.VSS(VSS),.VDD(VDD),.Y(g32506),.A(g31376));
  NOT NOT1_7228(.VSS(VSS),.VDD(VDD),.Y(g8784),.A(I12764));
  NOT NOT1_7229(.VSS(VSS),.VDD(VDD),.Y(I31724),.A(g33076));
  NOT NOT1_7230(.VSS(VSS),.VDD(VDD),.Y(g33636),.A(I31463));
  NOT NOT1_7231(.VSS(VSS),.VDD(VDD),.Y(g29185),.A(I27481));
  NOT NOT1_7232(.VSS(VSS),.VDD(VDD),.Y(I32956),.A(g34654));
  NOT NOT1_7233(.VSS(VSS),.VDD(VDD),.Y(g30326),.A(I28579));
  NOT NOT1_7234(.VSS(VSS),.VDD(VDD),.Y(g21723),.A(I21288));
  NOT NOT1_7235(.VSS(VSS),.VDD(VDD),.Y(g29092),.A(g27800));
  NOT NOT1_7236(.VSS(VSS),.VDD(VDD),.Y(I32297),.A(g34059));
  NOT NOT1_7237(.VSS(VSS),.VDD(VDD),.Y(g34949),.A(g34939));
  NOT NOT1_7238(.VSS(VSS),.VDD(VDD),.Y(g10498),.A(g7161));
  NOT NOT1_7239(.VSS(VSS),.VDD(VDD),.Y(I32103),.A(g33661));
  NOT NOT1_7240(.VSS(VSS),.VDD(VDD),.Y(g34326),.A(g34091));
  NOT NOT1_7241(.VSS(VSS),.VDD(VDD),.Y(g13061),.A(g10981));
  NOT NOT1_7242(.VSS(VSS),.VDD(VDD),.Y(I31829),.A(g33454));
  NOT NOT1_7243(.VSS(VSS),.VDD(VDD),.Y(I18479),.A(g13041));
  NOT NOT1_7244(.VSS(VSS),.VDD(VDD),.Y(g31852),.A(g29385));
  NOT NOT1_7245(.VSS(VSS),.VDD(VDD),.Y(g6959),.A(g4420));
  NOT NOT1_7246(.VSS(VSS),.VDD(VDD),.Y(I31535),.A(g33377));
  NOT NOT1_7247(.VSS(VSS),.VDD(VDD),.Y(g30040),.A(g29025));
  NOT NOT1_7248(.VSS(VSS),.VDD(VDD),.Y(I13202),.A(g5105));
  NOT NOT1_7249(.VSS(VSS),.VDD(VDD),.Y(g19586),.A(g16349));
  NOT NOT1_7250(.VSS(VSS),.VDD(VDD),.Y(I12123),.A(g758));
  NOT NOT1_7251(.VSS(VSS),.VDD(VDD),.Y(g17125),.A(I18177));
  NOT NOT1_7252(.VSS(VSS),.VDD(VDD),.Y(g17532),.A(I18479));
  NOT NOT1_7253(.VSS(VSS),.VDD(VDD),.Y(g27402),.A(I26100));
  NOT NOT1_7254(.VSS(VSS),.VDD(VDD),.Y(g34536),.A(I32601));
  NOT NOT1_7255(.VSS(VSS),.VDD(VDD),.Y(I17166),.A(g14536));
  NOT NOT1_7256(.VSS(VSS),.VDD(VDD),.Y(g28161),.A(I26676));
  NOT NOT1_7257(.VSS(VSS),.VDD(VDD),.Y(g7634),.A(I12123));
  NOT NOT1_7258(.VSS(VSS),.VDD(VDD),.Y(g15758),.A(I17276));
  NOT NOT1_7259(.VSS(VSS),.VDD(VDD),.Y(g21387),.A(I21115));
  NOT NOT1_7260(.VSS(VSS),.VDD(VDD),.Y(I22485),.A(g21308));
  NOT NOT1_7261(.VSS(VSS),.VDD(VDD),.Y(I29221),.A(g30307));
  NOT NOT1_7262(.VSS(VSS),.VDD(VDD),.Y(g23433),.A(g21562));
  NOT NOT1_7263(.VSS(VSS),.VDD(VDD),.Y(I28419),.A(g29195));
  NOT NOT1_7264(.VSS(VSS),.VDD(VDD),.Y(I13979),.A(g7733));
  NOT NOT1_7265(.VSS(VSS),.VDD(VDD),.Y(I32824),.A(g34475));
  NOT NOT1_7266(.VSS(VSS),.VDD(VDD),.Y(g24426),.A(g22722));
  NOT NOT1_7267(.VSS(VSS),.VDD(VDD),.Y(g8479),.A(g3057));
  NOT NOT1_7268(.VSS(VSS),.VDD(VDD),.Y(g20190),.A(g16971));
  NOT NOT1_7269(.VSS(VSS),.VDD(VDD),.Y(g22144),.A(g18997));
  NOT NOT1_7270(.VSS(VSS),.VDD(VDD),.Y(I24038),.A(g22202));
  NOT NOT1_7271(.VSS(VSS),.VDD(VDD),.Y(g23620),.A(I22769));
  NOT NOT1_7272(.VSS(VSS),.VDD(VDD),.Y(g28709),.A(I27192));
  NOT NOT1_7273(.VSS(VSS),.VDD(VDD),.Y(g10080),.A(g1982));
  NOT NOT1_7274(.VSS(VSS),.VDD(VDD),.Y(I17008),.A(g12857));
  NOT NOT1_7275(.VSS(VSS),.VDD(VDD),.Y(I32671),.A(g34388));
  NOT NOT1_7276(.VSS(VSS),.VDD(VDD),.Y(g8840),.A(g4277));
  NOT NOT1_7277(.VSS(VSS),.VDD(VDD),.Y(g9212),.A(g6466));
  NOT NOT1_7278(.VSS(VSS),.VDD(VDD),.Y(g12866),.A(g10369));
  NOT NOT1_7279(.VSS(VSS),.VDD(VDD),.Y(I21918),.A(g21290));
  NOT NOT1_7280(.VSS(VSS),.VDD(VDD),.Y(I17892),.A(g3325));
  NOT NOT1_7281(.VSS(VSS),.VDD(VDD),.Y(g21343),.A(g16428));
  NOT NOT1_7282(.VSS(VSS),.VDD(VDD),.Y(I26925),.A(g27015));
  NOT NOT1_7283(.VSS(VSS),.VDD(VDD),.Y(g8390),.A(g3385));
  NOT NOT1_7284(.VSS(VSS),.VDD(VDD),.Y(g32927),.A(g30825));
  NOT NOT1_7285(.VSS(VSS),.VDD(VDD),.Y(g15345),.A(I17108));
  NOT NOT1_7286(.VSS(VSS),.VDD(VDD),.Y(g14432),.A(g12311));
  NOT NOT1_7287(.VSS(VSS),.VDD(VDD),.Y(g17680),.A(g14889));
  NOT NOT1_7288(.VSS(VSS),.VDD(VDD),.Y(g17144),.A(g14085));
  NOT NOT1_7289(.VSS(VSS),.VDD(VDD),.Y(g26634),.A(g25317));
  NOT NOT1_7290(.VSS(VSS),.VDD(VDD),.Y(g26851),.A(I25579));
  NOT NOT1_7291(.VSS(VSS),.VDD(VDD),.Y(g11447),.A(I14450));
  NOT NOT1_7292(.VSS(VSS),.VDD(VDD),.Y(g7926),.A(g3423));
  NOT NOT1_7293(.VSS(VSS),.VDD(VDD),.Y(I15162),.A(g10176));
  NOT NOT1_7294(.VSS(VSS),.VDD(VDD),.Y(g20546),.A(g18008));
  NOT NOT1_7295(.VSS(VSS),.VDD(VDD),.Y(g20089),.A(g17533));
  NOT NOT1_7296(.VSS(VSS),.VDD(VDD),.Y(g23971),.A(g20751));
  NOT NOT1_7297(.VSS(VSS),.VDD(VDD),.Y(I26378),.A(g26850));
  NOT NOT1_7298(.VSS(VSS),.VDD(VDD),.Y(g19720),.A(I20130));
  NOT NOT1_7299(.VSS(VSS),.VDD(VDD),.Y(g20211),.A(g16931));
  NOT NOT1_7300(.VSS(VSS),.VDD(VDD),.Y(I25369),.A(g24891));
  NOT NOT1_7301(.VSS(VSS),.VDD(VDD),.Y(g24089),.A(g19890));
  NOT NOT1_7302(.VSS(VSS),.VDD(VDD),.Y(I19851),.A(g16615));
  NOT NOT1_7303(.VSS(VSS),.VDD(VDD),.Y(g27597),.A(g26745));
  NOT NOT1_7304(.VSS(VSS),.VDD(VDD),.Y(g21369),.A(g16285));
  NOT NOT1_7305(.VSS(VSS),.VDD(VDD),.Y(I33291),.A(g34983));
  NOT NOT1_7306(.VSS(VSS),.VDD(VDD),.Y(g12077),.A(I14939));
  NOT NOT1_7307(.VSS(VSS),.VDD(VDD),.Y(g32649),.A(g30673));
  NOT NOT1_7308(.VSS(VSS),.VDD(VDD),.Y(g25553),.A(g22550));
  NOT NOT1_7309(.VSS(VSS),.VDD(VDD),.Y(g20088),.A(g17533));
  NOT NOT1_7310(.VSS(VSS),.VDD(VDD),.Y(I27391),.A(g27929));
  NOT NOT1_7311(.VSS(VSS),.VDD(VDD),.Y(g8356),.A(g54));
  NOT NOT1_7312(.VSS(VSS),.VDD(VDD),.Y(I20937),.A(g16967));
  NOT NOT1_7313(.VSS(VSS),.VDD(VDD),.Y(g9229),.A(g5052));
  NOT NOT1_7314(.VSS(VSS),.VDD(VDD),.Y(I13094),.A(g2724));
  NOT NOT1_7315(.VSS(VSS),.VDD(VDD),.Y(g14753),.A(g11317));
  NOT NOT1_7316(.VSS(VSS),.VDD(VDD),.Y(I33173),.A(g34887));
  NOT NOT1_7317(.VSS(VSS),.VDD(VDD),.Y(g24088),.A(g21209));
  NOT NOT1_7318(.VSS(VSS),.VDD(VDD),.Y(g19493),.A(g16349));
  NOT NOT1_7319(.VSS(VSS),.VDD(VDD),.Y(g24024),.A(g21193));
  NOT NOT1_7320(.VSS(VSS),.VDD(VDD),.Y(g14342),.A(g12163));
  NOT NOT1_7321(.VSS(VSS),.VDD(VDD),.Y(g34673),.A(I32803));
  NOT NOT1_7322(.VSS(VSS),.VDD(VDD),.Y(g34847),.A(I33067));
  NOT NOT1_7323(.VSS(VSS),.VDD(VDD),.Y(g31609),.A(I29211));
  NOT NOT1_7324(.VSS(VSS),.VDD(VDD),.Y(g29215),.A(I27561));
  NOT NOT1_7325(.VSS(VSS),.VDD(VDD),.Y(g10031),.A(I13552));
  NOT NOT1_7326(.VSS(VSS),.VDD(VDD),.Y(g32648),.A(g30614));
  NOT NOT1_7327(.VSS(VSS),.VDD(VDD),.Y(g32491),.A(g31566));
  NOT NOT1_7328(.VSS(VSS),.VDD(VDD),.Y(g32903),.A(g31376));
  NOT NOT1_7329(.VSS(VSS),.VDD(VDD),.Y(g25326),.A(g22228));
  NOT NOT1_7330(.VSS(VSS),.VDD(VDD),.Y(g14031),.A(I16289));
  NOT NOT1_7331(.VSS(VSS),.VDD(VDD),.Y(g9822),.A(g125));
  NOT NOT1_7332(.VSS(VSS),.VDD(VDD),.Y(g10199),.A(g1968));
  NOT NOT1_7333(.VSS(VSS),.VDD(VDD),.Y(I11801),.A(g6395));
  NOT NOT1_7334(.VSS(VSS),.VDD(VDD),.Y(I14455),.A(g10197));
  NOT NOT1_7335(.VSS(VSS),.VDD(VDD),.Y(g16605),.A(g13955));
  NOT NOT1_7336(.VSS(VSS),.VDD(VDD),.Y(g11472),.A(g7918));
  NOT NOT1_7337(.VSS(VSS),.VDD(VDD),.Y(I27579),.A(g28184));
  NOT NOT1_7338(.VSS(VSS),.VDD(VDD),.Y(I29371),.A(g30325));
  NOT NOT1_7339(.VSS(VSS),.VDD(VDD),.Y(g12923),.A(I15542));
  NOT NOT1_7340(.VSS(VSS),.VDD(VDD),.Y(g31608),.A(g29653));
  NOT NOT1_7341(.VSS(VSS),.VDD(VDD),.Y(g18527),.A(I19345));
  NOT NOT1_7342(.VSS(VSS),.VDD(VDD),.Y(g20497),.A(g18065));
  NOT NOT1_7343(.VSS(VSS),.VDD(VDD),.Y(g32604),.A(g31154));
  NOT NOT1_7344(.VSS(VSS),.VDD(VDD),.Y(g34062),.A(g33711));
  NOT NOT1_7345(.VSS(VSS),.VDD(VDD),.Y(I28588),.A(g29368));
  NOT NOT1_7346(.VSS(VSS),.VDD(VDD),.Y(g32755),.A(g31672));
  NOT NOT1_7347(.VSS(VSS),.VDD(VDD),.Y(I30959),.A(g32021));
  NOT NOT1_7348(.VSS(VSS),.VDD(VDD),.Y(g10198),.A(I13672));
  NOT NOT1_7349(.VSS(VSS),.VDD(VDD),.Y(g12300),.A(I15144));
  NOT NOT1_7350(.VSS(VSS),.VDD(VDD),.Y(g11911),.A(g10022));
  NOT NOT1_7351(.VSS(VSS),.VDD(VDD),.Y(g16812),.A(g13555));
  NOT NOT1_7352(.VSS(VSS),.VDD(VDD),.Y(g21412),.A(g15758));
  NOT NOT1_7353(.VSS(VSS),.VDD(VDD),.Y(g32770),.A(g31710));
  NOT NOT1_7354(.VSS(VSS),.VDD(VDD),.Y(g34933),.A(g34916));
  NOT NOT1_7355(.VSS(VSS),.VDD(VDD),.Y(g14198),.A(g12180));
  NOT NOT1_7356(.VSS(VSS),.VDD(VDD),.Y(g32563),.A(g31554));
  NOT NOT1_7357(.VSS(VSS),.VDD(VDD),.Y(I32089),.A(g33665));
  NOT NOT1_7358(.VSS(VSS),.VDD(VDD),.Y(I33134),.A(g34906));
  NOT NOT1_7359(.VSS(VSS),.VDD(VDD),.Y(g13246),.A(g10939));
  NOT NOT1_7360(.VSS(VSS),.VDD(VDD),.Y(g20700),.A(g17873));
  NOT NOT1_7361(.VSS(VSS),.VDD(VDD),.Y(g20659),.A(g17873));
  NOT NOT1_7362(.VSS(VSS),.VDD(VDD),.Y(g34851),.A(I33075));
  NOT NOT1_7363(.VSS(VSS),.VDD(VDD),.Y(g20625),.A(g15348));
  NOT NOT1_7364(.VSS(VSS),.VDD(VDD),.Y(g10393),.A(g6991));
  NOT NOT1_7365(.VSS(VSS),.VDD(VDD),.Y(g24126),.A(g19935));
  NOT NOT1_7366(.VSS(VSS),.VDD(VDD),.Y(g24625),.A(g23135));
  NOT NOT1_7367(.VSS(VSS),.VDD(VDD),.Y(g14330),.A(I16486));
  NOT NOT1_7368(.VSS(VSS),.VDD(VDD),.Y(g24987),.A(g23630));
  NOT NOT1_7369(.VSS(VSS),.VDD(VDD),.Y(g8954),.A(g1079));
  NOT NOT1_7370(.VSS(VSS),.VDD(VDD),.Y(g7543),.A(I12033));
  NOT NOT1_7371(.VSS(VSS),.VDD(VDD),.Y(g31799),.A(g29385));
  NOT NOT1_7372(.VSS(VSS),.VDD(VDD),.Y(g23896),.A(g19210));
  NOT NOT1_7373(.VSS(VSS),.VDD(VDD),.Y(g25564),.A(g22312));
  NOT NOT1_7374(.VSS(VSS),.VDD(VDD),.Y(g8363),.A(g239));
  NOT NOT1_7375(.VSS(VSS),.VDD(VDD),.Y(g18894),.A(g16000));
  NOT NOT1_7376(.VSS(VSS),.VDD(VDD),.Y(g31813),.A(g29385));
  NOT NOT1_7377(.VSS(VSS),.VDD(VDD),.Y(g21228),.A(g17531));
  NOT NOT1_7378(.VSS(VSS),.VDD(VDD),.Y(g33799),.A(g33299));
  NOT NOT1_7379(.VSS(VSS),.VDD(VDD),.Y(g10365),.A(g6867));
  NOT NOT1_7380(.VSS(VSS),.VDD(VDD),.Y(g22224),.A(g19277));
  NOT NOT1_7381(.VSS(VSS),.VDD(VDD),.Y(g33813),.A(I31659));
  NOT NOT1_7382(.VSS(VSS),.VDD(VDD),.Y(g8032),.A(I12355));
  NOT NOT1_7383(.VSS(VSS),.VDD(VDD),.Y(g19517),.A(g16777));
  NOT NOT1_7384(.VSS(VSS),.VDD(VDD),.Y(g23228),.A(g21070));
  NOT NOT1_7385(.VSS(VSS),.VDD(VDD),.Y(I18373),.A(g13011));
  NOT NOT1_7386(.VSS(VSS),.VDD(VDD),.Y(g29906),.A(g28793));
  NOT NOT1_7387(.VSS(VSS),.VDD(VDD),.Y(g29348),.A(g28194));
  NOT NOT1_7388(.VSS(VSS),.VDD(VDD),.Y(g16795),.A(I18009));
  NOT NOT1_7389(.VSS(VSS),.VDD(VDD),.Y(g10960),.A(g9007));
  NOT NOT1_7390(.VSS(VSS),.VDD(VDD),.Y(I17675),.A(g13394));
  NOT NOT1_7391(.VSS(VSS),.VDD(VDD),.Y(g23011),.A(g20330));
  NOT NOT1_7392(.VSS(VSS),.VDD(VDD),.Y(g31798),.A(g29385));
  NOT NOT1_7393(.VSS(VSS),.VDD(VDD),.Y(g32767),.A(g30735));
  NOT NOT1_7394(.VSS(VSS),.VDD(VDD),.Y(g32794),.A(g30937));
  NOT NOT1_7395(.VSS(VSS),.VDD(VDD),.Y(I14623),.A(g8925));
  NOT NOT1_7396(.VSS(VSS),.VDD(VDD),.Y(g11147),.A(g8417));
  NOT NOT1_7397(.VSS(VSS),.VDD(VDD),.Y(g11754),.A(g8229));
  NOT NOT1_7398(.VSS(VSS),.VDD(VDD),.Y(I17154),.A(g13605));
  NOT NOT1_7399(.VSS(VSS),.VDD(VDD),.Y(I23680),.A(g23219));
  NOT NOT1_7400(.VSS(VSS),.VDD(VDD),.Y(g25183),.A(g22763));
  NOT NOT1_7401(.VSS(VSS),.VDD(VDD),.Y(g32899),.A(g31021));
  NOT NOT1_7402(.VSS(VSS),.VDD(VDD),.Y(g7534),.A(g1367));
  NOT NOT1_7403(.VSS(VSS),.VDD(VDD),.Y(g31805),.A(g29385));
  NOT NOT1_7404(.VSS(VSS),.VDD(VDD),.Y(g17224),.A(I18248));
  NOT NOT1_7405(.VSS(VSS),.VDD(VDD),.Y(g16514),.A(g14139));
  NOT NOT1_7406(.VSS(VSS),.VDD(VDD),.Y(g12885),.A(g10382));
  NOT NOT1_7407(.VSS(VSS),.VDD(VDD),.Y(g22495),.A(g19801));
  NOT NOT1_7408(.VSS(VSS),.VDD(VDD),.Y(g17308),.A(g14876));
  NOT NOT1_7409(.VSS(VSS),.VDD(VDD),.Y(g23582),.A(I22729));
  NOT NOT1_7410(.VSS(VSS),.VDD(VDD),.Y(g32633),.A(g31154));
  NOT NOT1_7411(.VSS(VSS),.VDD(VDD),.Y(g32898),.A(g30825));
  NOT NOT1_7412(.VSS(VSS),.VDD(VDD),.Y(I32659),.A(g34391));
  NOT NOT1_7413(.VSS(VSS),.VDD(VDD),.Y(g15048),.A(I16969));
  NOT NOT1_7414(.VSS(VSS),.VDD(VDD),.Y(g9620),.A(g6187));
  NOT NOT1_7415(.VSS(VSS),.VDD(VDD),.Y(g9462),.A(g6215));
  NOT NOT1_7416(.VSS(VSS),.VDD(VDD),.Y(I23336),.A(g22721));
  NOT NOT1_7417(.VSS(VSS),.VDD(VDD),.Y(I19756),.A(g17812));
  NOT NOT1_7418(.VSS(VSS),.VDD(VDD),.Y(g19362),.A(g16072));
  NOT NOT1_7419(.VSS(VSS),.VDD(VDD),.Y(g7927),.A(g4064));
  NOT NOT1_7420(.VSS(VSS),.VDD(VDD),.Y(g34574),.A(I32648));
  NOT NOT1_7421(.VSS(VSS),.VDD(VDD),.Y(g32719),.A(g31672));
  NOT NOT1_7422(.VSS(VSS),.VDD(VDD),.Y(I12041),.A(g2741));
  NOT NOT1_7423(.VSS(VSS),.VDD(VDD),.Y(g20060),.A(g16540));
  NOT NOT1_7424(.VSS(VSS),.VDD(VDD),.Y(g34047),.A(g33637));
  NOT NOT1_7425(.VSS(VSS),.VDD(VDD),.Y(g18979),.A(g16136));
  NOT NOT1_7426(.VSS(VSS),.VDD(VDD),.Y(g19523),.A(g16100));
  NOT NOT1_7427(.VSS(VSS),.VDD(VDD),.Y(g24060),.A(g21256));
  NOT NOT1_7428(.VSS(VSS),.VDD(VDD),.Y(g8912),.A(g4180));
  NOT NOT1_7429(.VSS(VSS),.VDD(VDD),.Y(I16120),.A(g11868));
  NOT NOT1_7430(.VSS(VSS),.VDD(VDD),.Y(g33934),.A(I31814));
  NOT NOT1_7431(.VSS(VSS),.VDD(VDD),.Y(g10708),.A(g7836));
  NOT NOT1_7432(.VSS(VSS),.VDD(VDD),.Y(g20197),.A(g16987));
  NOT NOT1_7433(.VSS(VSS),.VDD(VDD),.Y(g6928),.A(I11716));
  NOT NOT1_7434(.VSS(VSS),.VDD(VDD),.Y(I12746),.A(g4087));
  NOT NOT1_7435(.VSS(VSS),.VDD(VDD),.Y(g21379),.A(g17873));
  NOT NOT1_7436(.VSS(VSS),.VDD(VDD),.Y(g34311),.A(g34097));
  NOT NOT1_7437(.VSS(VSS),.VDD(VDD),.Y(I12493),.A(g5002));
  NOT NOT1_7438(.VSS(VSS),.VDD(VDD),.Y(g22976),.A(I22149));
  NOT NOT1_7439(.VSS(VSS),.VDD(VDD),.Y(g22985),.A(g20330));
  NOT NOT1_7440(.VSS(VSS),.VDD(VDD),.Y(g32718),.A(g30825));
  NOT NOT1_7441(.VSS(VSS),.VDD(VDD),.Y(g32521),.A(g31376));
  NOT NOT1_7442(.VSS(VSS),.VDD(VDD),.Y(g10087),.A(I13597));
  NOT NOT1_7443(.VSS(VSS),.VDD(VDD),.Y(g23925),.A(g21514));
  NOT NOT1_7444(.VSS(VSS),.VDD(VDD),.Y(g8357),.A(I12538));
  NOT NOT1_7445(.VSS(VSS),.VDD(VDD),.Y(g18978),.A(g16000));
  NOT NOT1_7446(.VSS(VSS),.VDD(VDD),.Y(g7946),.A(I12314));
  NOT NOT1_7447(.VSS(VSS),.VDD(VDD),.Y(g7660),.A(I12144));
  NOT NOT1_7448(.VSS(VSS),.VDD(VDD),.Y(g29653),.A(I27927));
  NOT NOT1_7449(.VSS(VSS),.VDD(VDD),.Y(I22729),.A(g21308));
  NOT NOT1_7450(.VSS(VSS),.VDD(VDD),.Y(g26820),.A(I25534));
  NOT NOT1_7451(.VSS(VSS),.VDD(VDD),.Y(g21050),.A(g17873));
  NOT NOT1_7452(.VSS(VSS),.VDD(VDD),.Y(g20527),.A(g18008));
  NOT NOT1_7453(.VSS(VSS),.VDD(VDD),.Y(I13597),.A(g4417));
  NOT NOT1_7454(.VSS(VSS),.VDD(VDD),.Y(g11367),.A(I14381));
  NOT NOT1_7455(.VSS(VSS),.VDD(VDD),.Y(g28918),.A(g27832));
  NOT NOT1_7456(.VSS(VSS),.VDD(VDD),.Y(g32832),.A(g30735));
  NOT NOT1_7457(.VSS(VSS),.VDD(VDD),.Y(I20321),.A(g16920));
  NOT NOT1_7458(.VSS(VSS),.VDD(VDD),.Y(g23378),.A(g21070));
  NOT NOT1_7459(.VSS(VSS),.VDD(VDD),.Y(g13394),.A(I15915));
  NOT NOT1_7460(.VSS(VSS),.VDD(VDD),.Y(I31491),.A(g33283));
  NOT NOT1_7461(.VSS(VSS),.VDD(VDD),.Y(g33761),.A(I31616));
  NOT NOT1_7462(.VSS(VSS),.VDD(VDD),.Y(g24527),.A(g22670));
  NOT NOT1_7463(.VSS(VSS),.VDD(VDD),.Y(g7903),.A(g969));
  NOT NOT1_7464(.VSS(VSS),.VDD(VDD),.Y(g30072),.A(I28301));
  NOT NOT1_7465(.VSS(VSS),.VDD(VDD),.Y(g17687),.A(g15042));
  NOT NOT1_7466(.VSS(VSS),.VDD(VDD),.Y(I31604),.A(g33176));
  NOT NOT1_7467(.VSS(VSS),.VDD(VDD),.Y(g28079),.A(I26578));
  NOT NOT1_7468(.VSS(VSS),.VDD(VDD),.Y(g10043),.A(g1632));
  NOT NOT1_7469(.VSS(VSS),.VDD(VDD),.Y(I13280),.A(g6140));
  NOT NOT1_7470(.VSS(VSS),.VDD(VDD),.Y(g7513),.A(g6315));
  NOT NOT1_7471(.VSS(VSS),.VDD(VDD),.Y(g26731),.A(g25470));
  NOT NOT1_7472(.VSS(VSS),.VDD(VDD),.Y(g34592),.A(I32684));
  NOT NOT1_7473(.VSS(VSS),.VDD(VDD),.Y(I11688),.A(g70));
  NOT NOT1_7474(.VSS(VSS),.VDD(VDD),.Y(I16698),.A(g12077));
  NOT NOT1_7475(.VSS(VSS),.VDD(VDD),.Y(g29333),.A(g28167));
  NOT NOT1_7476(.VSS(VSS),.VDD(VDD),.Y(g16473),.A(g13977));
  NOT NOT1_7477(.VSS(VSS),.VDD(VDD),.Y(I31770),.A(g33197));
  NOT NOT1_7478(.VSS(VSS),.VDD(VDD),.Y(g32861),.A(g31376));
  NOT NOT1_7479(.VSS(VSS),.VDD(VDD),.Y(g9842),.A(g3274));
  NOT NOT1_7480(.VSS(VSS),.VDD(VDD),.Y(g23944),.A(g19147));
  NOT NOT1_7481(.VSS(VSS),.VDD(VDD),.Y(g32573),.A(g30825));
  NOT NOT1_7482(.VSS(VSS),.VDD(VDD),.Y(g18094),.A(I18888));
  NOT NOT1_7483(.VSS(VSS),.VDD(VDD),.Y(g31013),.A(g29679));
  NOT NOT1_7484(.VSS(VSS),.VDD(VDD),.Y(I14589),.A(g8818));
  NOT NOT1_7485(.VSS(VSS),.VDD(VDD),.Y(g25213),.A(g23293));
  NOT NOT1_7486(.VSS(VSS),.VDD(VDD),.Y(g19437),.A(g16349));
  NOT NOT1_7487(.VSS(VSS),.VDD(VDD),.Y(g20503),.A(g15373));
  NOT NOT1_7488(.VSS(VSS),.VDD(VDD),.Y(g9298),.A(g5080));
  NOT NOT1_7489(.VSS(VSS),.VDD(VDD),.Y(g28598),.A(g27717));
  NOT NOT1_7490(.VSS(VSS),.VDD(VDD),.Y(I18909),.A(g16873));
  NOT NOT1_7491(.VSS(VSS),.VDD(VDD),.Y(g9392),.A(g5869));
  NOT NOT1_7492(.VSS(VSS),.VDD(VDD),.Y(g32926),.A(g31376));
  NOT NOT1_7493(.VSS(VSS),.VDD(VDD),.Y(I32855),.A(g34540));
  NOT NOT1_7494(.VSS(VSS),.VDD(VDD),.Y(g7178),.A(g4392));
  NOT NOT1_7495(.VSS(VSS),.VDD(VDD),.Y(g7436),.A(g5276));
  NOT NOT1_7496(.VSS(VSS),.VDD(VDD),.Y(I14836),.A(g9688));
  NOT NOT1_7497(.VSS(VSS),.VDD(VDD),.Y(g8626),.A(g4040));
  NOT NOT1_7498(.VSS(VSS),.VDD(VDD),.Y(g21681),.A(I21242));
  NOT NOT1_7499(.VSS(VSS),.VDD(VDD),.Y(g29963),.A(g28931));
  NOT NOT1_7500(.VSS(VSS),.VDD(VDD),.Y(g16724),.A(g14079));
  NOT NOT1_7501(.VSS(VSS),.VDD(VDD),.Y(g22842),.A(g19875));
  NOT NOT1_7502(.VSS(VSS),.VDD(VDD),.Y(g23681),.A(g21012));
  NOT NOT1_7503(.VSS(VSS),.VDD(VDD),.Y(I18117),.A(g13302));
  NOT NOT1_7504(.VSS(VSS),.VDD(VDD),.Y(g32612),.A(g30614));
  NOT NOT1_7505(.VSS(VSS),.VDD(VDD),.Y(g16325),.A(g13223));
  NOT NOT1_7506(.VSS(VSS),.VDD(VDD),.Y(g18877),.A(g15224));
  NOT NOT1_7507(.VSS(VSS),.VDD(VDD),.Y(I23309),.A(g21677));
  NOT NOT1_7508(.VSS(VSS),.VDD(VDD),.Y(g25452),.A(g22228));
  NOT NOT1_7509(.VSS(VSS),.VDD(VDD),.Y(g15371),.A(I17114));
  NOT NOT1_7510(.VSS(VSS),.VDD(VDD),.Y(g25047),.A(g23733));
  NOT NOT1_7511(.VSS(VSS),.VDD(VDD),.Y(g32099),.A(g31009));
  NOT NOT1_7512(.VSS(VSS),.VDD(VDD),.Y(g10375),.A(g6941));
  NOT NOT1_7513(.VSS(VSS),.VDD(VDD),.Y(I21288),.A(g18216));
  NOT NOT1_7514(.VSS(VSS),.VDD(VDD),.Y(g34820),.A(I33034));
  NOT NOT1_7515(.VSS(VSS),.VDD(VDD),.Y(g16920),.A(I18086));
  NOT NOT1_7516(.VSS(VSS),.VDD(VDD),.Y(g20714),.A(g15277));
  NOT NOT1_7517(.VSS(VSS),.VDD(VDD),.Y(g20450),.A(g15277));
  NOT NOT1_7518(.VSS(VSS),.VDD(VDD),.Y(g23429),.A(g20453));
  NOT NOT1_7519(.VSS(VSS),.VDD(VDD),.Y(g32701),.A(g31376));
  NOT NOT1_7520(.VSS(VSS),.VDD(VDD),.Y(g12076),.A(g9280));
  NOT NOT1_7521(.VSS(VSS),.VDD(VDD),.Y(g7335),.A(g2287));
  NOT NOT1_7522(.VSS(VSS),.VDD(VDD),.Y(g7831),.A(I12227));
  NOT NOT1_7523(.VSS(VSS),.VDD(VDD),.Y(I14119),.A(g7824));
  NOT NOT1_7524(.VSS(VSS),.VDD(VDD),.Y(g32777),.A(g31710));
  NOT NOT1_7525(.VSS(VSS),.VDD(VDD),.Y(g32534),.A(g30673));
  NOT NOT1_7526(.VSS(VSS),.VDD(VDD),.Y(g12721),.A(g10061));
  NOT NOT1_7527(.VSS(VSS),.VDD(VDD),.Y(g34152),.A(I32109));
  NOT NOT1_7528(.VSS(VSS),.VDD(VDD),.Y(g20707),.A(g18008));
  NOT NOT1_7529(.VSS(VSS),.VDD(VDD),.Y(g21428),.A(g15758));
  NOT NOT1_7530(.VSS(VSS),.VDD(VDD),.Y(I22622),.A(g21209));
  NOT NOT1_7531(.VSS(VSS),.VDD(VDD),.Y(g20910),.A(g15171));
  NOT NOT1_7532(.VSS(VSS),.VDD(VDD),.Y(g34846),.A(I33064));
  NOT NOT1_7533(.VSS(VSS),.VDD(VDD),.Y(g23793),.A(g19074));
  NOT NOT1_7534(.VSS(VSS),.VDD(VDD),.Y(g12054),.A(g7690));
  NOT NOT1_7535(.VSS(VSS),.VDD(VDD),.Y(g17392),.A(g14924));
  NOT NOT1_7536(.VSS(VSS),.VDD(VDD),.Y(g19600),.A(g16164));
  NOT NOT1_7537(.VSS(VSS),.VDD(VDD),.Y(g10337),.A(g5016));
  NOT NOT1_7538(.VSS(VSS),.VDD(VDD),.Y(g24819),.A(I23998));
  NOT NOT1_7539(.VSS(VSS),.VDD(VDD),.Y(g19781),.A(g16489));
  NOT NOT1_7540(.VSS(VSS),.VDD(VDD),.Y(g17489),.A(g12955));
  NOT NOT1_7541(.VSS(VSS),.VDD(VDD),.Y(I24334),.A(g22976));
  NOT NOT1_7542(.VSS(VSS),.VDD(VDD),.Y(g20496),.A(g17929));
  NOT NOT1_7543(.VSS(VSS),.VDD(VDD),.Y(g7805),.A(g4366));
  NOT NOT1_7544(.VSS(VSS),.VDD(VDD),.Y(g7916),.A(I12300));
  NOT NOT1_7545(.VSS(VSS),.VDD(VDD),.Y(g25051),.A(I24215));
  NOT NOT1_7546(.VSS(VSS),.VDD(VDD),.Y(g25072),.A(g23630));
  NOT NOT1_7547(.VSS(VSS),.VDD(VDD),.Y(g24818),.A(g23191));
  NOT NOT1_7548(.VSS(VSS),.VDD(VDD),.Y(g32462),.A(g30673));
  NOT NOT1_7549(.VSS(VSS),.VDD(VDD),.Y(I14749),.A(g10031));
  NOT NOT1_7550(.VSS(VSS),.VDD(VDD),.Y(g24979),.A(g22369));
  NOT NOT1_7551(.VSS(VSS),.VDD(VDD),.Y(g21690),.A(g16540));
  NOT NOT1_7552(.VSS(VSS),.VDD(VDD),.Y(g22830),.A(g20283));
  NOT NOT1_7553(.VSS(VSS),.VDD(VDD),.Y(g19952),.A(g15915));
  NOT NOT1_7554(.VSS(VSS),.VDD(VDD),.Y(g24055),.A(g19968));
  NOT NOT1_7555(.VSS(VSS),.VDD(VDD),.Y(g7749),.A(g996));
  NOT NOT1_7556(.VSS(VSS),.VDD(VDD),.Y(g19351),.A(g17367));
  NOT NOT1_7557(.VSS(VSS),.VDD(VDD),.Y(I12523),.A(g3794));
  NOT NOT1_7558(.VSS(VSS),.VDD(VDD),.Y(g23549),.A(g18833));
  NOT NOT1_7559(.VSS(VSS),.VDD(VDD),.Y(g27773),.A(I26378));
  NOT NOT1_7560(.VSS(VSS),.VDD(VDD),.Y(g20070),.A(g16173));
  NOT NOT1_7561(.VSS(VSS),.VDD(VDD),.Y(g20978),.A(g15595));
  NOT NOT1_7562(.VSS(VSS),.VDD(VDD),.Y(g24111),.A(g19890));
  NOT NOT1_7563(.VSS(VSS),.VDD(VDD),.Y(g28656),.A(g27742));
  NOT NOT1_7564(.VSS(VSS),.VDD(VDD),.Y(g9708),.A(g2741));
  NOT NOT1_7565(.VSS(VSS),.VDD(VDD),.Y(g24070),.A(g20014));
  NOT NOT1_7566(.VSS(VSS),.VDD(VDD),.Y(g24978),.A(g22342));
  NOT NOT1_7567(.VSS(VSS),.VDD(VDD),.Y(g34691),.A(I32843));
  NOT NOT1_7568(.VSS(VSS),.VDD(VDD),.Y(g29312),.A(g28877));
  NOT NOT1_7569(.VSS(VSS),.VDD(VDD),.Y(g20590),.A(g15426));
  NOT NOT1_7570(.VSS(VSS),.VDD(VDD),.Y(g22544),.A(g19589));
  NOT NOT1_7571(.VSS(VSS),.VDD(VDD),.Y(g22865),.A(g20330));
  NOT NOT1_7572(.VSS(VSS),.VDD(VDD),.Y(g23548),.A(g18833));
  NOT NOT1_7573(.VSS(VSS),.VDD(VDD),.Y(g8778),.A(I12758));
  NOT NOT1_7574(.VSS(VSS),.VDD(VDD),.Y(g29115),.A(g27779));
  NOT NOT1_7575(.VSS(VSS),.VDD(VDD),.Y(g7947),.A(g1500));
  NOT NOT1_7576(.VSS(VSS),.VDD(VDD),.Y(I20216),.A(g15862));
  NOT NOT1_7577(.VSS(VSS),.VDD(VDD),.Y(g24986),.A(g23590));
  NOT NOT1_7578(.VSS(VSS),.VDD(VDD),.Y(I14305),.A(g8805));
  NOT NOT1_7579(.VSS(VSS),.VDD(VDD),.Y(g9252),.A(g4304));
  NOT NOT1_7580(.VSS(VSS),.VDD(VDD),.Y(I26880),.A(g27527));
  NOT NOT1_7581(.VSS(VSS),.VDD(VDD),.Y(g23504),.A(g21468));
  NOT NOT1_7582(.VSS(VSS),.VDD(VDD),.Y(g13902),.A(g11389));
  NOT NOT1_7583(.VSS(VSS),.VDD(VDD),.Y(g13301),.A(g10862));
  NOT NOT1_7584(.VSS(VSS),.VDD(VDD),.Y(g31771),.A(I29337));
  NOT NOT1_7585(.VSS(VSS),.VDD(VDD),.Y(g19264),.A(I19802));
  NOT NOT1_7586(.VSS(VSS),.VDD(VDD),.Y(g18917),.A(g16077));
  NOT NOT1_7587(.VSS(VSS),.VDD(VDD),.Y(g19790),.A(g16971));
  NOT NOT1_7588(.VSS(VSS),.VDD(VDD),.Y(g20384),.A(g18008));
  NOT NOT1_7589(.VSS(VSS),.VDD(VDD),.Y(g12180),.A(g9477));
  NOT NOT1_7590(.VSS(VSS),.VDD(VDD),.Y(g9958),.A(g6148));
  NOT NOT1_7591(.VSS(VSS),.VDD(VDD),.Y(g29921),.A(g28864));
  NOT NOT1_7592(.VSS(VSS),.VDD(VDD),.Y(g13120),.A(g10632));
  NOT NOT1_7593(.VSS(VSS),.VDD(VDD),.Y(I18293),.A(g1079));
  NOT NOT1_7594(.VSS(VSS),.VDD(VDD),.Y(g24384),.A(g22885));
  NOT NOT1_7595(.VSS(VSS),.VDD(VDD),.Y(g25820),.A(g25051));
  NOT NOT1_7596(.VSS(VSS),.VDD(VDD),.Y(I26512),.A(g26817));
  NOT NOT1_7597(.VSS(VSS),.VDD(VDD),.Y(I17653),.A(g14276));
  NOT NOT1_7598(.VSS(VSS),.VDD(VDD),.Y(g20067),.A(g17328));
  NOT NOT1_7599(.VSS(VSS),.VDD(VDD),.Y(g32766),.A(g31376));
  NOT NOT1_7600(.VSS(VSS),.VDD(VDD),.Y(g6955),.A(I11726));
  NOT NOT1_7601(.VSS(VSS),.VDD(VDD),.Y(g29745),.A(g28500));
  NOT NOT1_7602(.VSS(VSS),.VDD(VDD),.Y(g24067),.A(g21256));
  NOT NOT1_7603(.VSS(VSS),.VDD(VDD),.Y(g24094),.A(g21143));
  NOT NOT1_7604(.VSS(VSS),.VDD(VDD),.Y(g11562),.A(g7648));
  NOT NOT1_7605(.VSS(VSS),.VDD(VDD),.Y(g17713),.A(g12947));
  NOT NOT1_7606(.VSS(VSS),.VDD(VDD),.Y(I18265),.A(g13350));
  NOT NOT1_7607(.VSS(VSS),.VDD(VDD),.Y(g34929),.A(I33179));
  NOT NOT1_7608(.VSS(VSS),.VDD(VDD),.Y(g27930),.A(I26451));
  NOT NOT1_7609(.VSS(VSS),.VDD(VDD),.Y(I12437),.A(g4999));
  NOT NOT1_7610(.VSS(VSS),.VDD(VDD),.Y(g27993),.A(I26503));
  NOT NOT1_7611(.VSS(VSS),.VDD(VDD),.Y(g8075),.A(g3742));
  NOT NOT1_7612(.VSS(VSS),.VDD(VDD),.Y(g32871),.A(g30937));
  NOT NOT1_7613(.VSS(VSS),.VDD(VDD),.Y(g30020),.A(g29097));
  NOT NOT1_7614(.VSS(VSS),.VDD(VDD),.Y(g30928),.A(I28908));
  NOT NOT1_7615(.VSS(VSS),.VDD(VDD),.Y(g22189),.A(I21769));
  NOT NOT1_7616(.VSS(VSS),.VDD(VDD),.Y(g8475),.A(I12608));
  NOT NOT1_7617(.VSS(VSS),.VDD(VDD),.Y(g26105),.A(I25146));
  NOT NOT1_7618(.VSS(VSS),.VDD(VDD),.Y(g9829),.A(g2250));
  NOT NOT1_7619(.VSS(VSS),.VDD(VDD),.Y(g12839),.A(g10350));
  NOT NOT1_7620(.VSS(VSS),.VDD(VDD),.Y(g6814),.A(g632));
  NOT NOT1_7621(.VSS(VSS),.VDD(VDD),.Y(g12930),.A(g12347));
  NOT NOT1_7622(.VSS(VSS),.VDD(VDD),.Y(g7873),.A(g1266));
  NOT NOT1_7623(.VSS(VSS),.VDD(VDD),.Y(g26743),.A(g25476));
  NOT NOT1_7624(.VSS(VSS),.VDD(VDD),.Y(g26827),.A(g24819));
  NOT NOT1_7625(.VSS(VSS),.VDD(VDD),.Y(g34583),.A(I32665));
  NOT NOT1_7626(.VSS(VSS),.VDD(VDD),.Y(g7632),.A(I12117));
  NOT NOT1_7627(.VSS(VSS),.VDD(VDD),.Y(g34928),.A(I33176));
  NOT NOT1_7628(.VSS(VSS),.VDD(VDD),.Y(g7095),.A(g6545));
  NOT NOT1_7629(.VSS(VSS),.VDD(VDD),.Y(I17636),.A(g14252));
  NOT NOT1_7630(.VSS(VSS),.VDD(VDD),.Y(g21057),.A(g15426));
  NOT NOT1_7631(.VSS(VSS),.VDD(VDD),.Y(g23002),.A(I22177));
  NOT NOT1_7632(.VSS(VSS),.VDD(VDD),.Y(g10079),.A(g1950));
  NOT NOT1_7633(.VSS(VSS),.VDD(VDD),.Y(g11290),.A(I14326));
  NOT NOT1_7634(.VSS(VSS),.VDD(VDD),.Y(g24150),.A(g19268));
  NOT NOT1_7635(.VSS(VSS),.VDD(VDD),.Y(g23057),.A(g20453));
  NOT NOT1_7636(.VSS(VSS),.VDD(VDD),.Y(I28594),.A(g29379));
  NOT NOT1_7637(.VSS(VSS),.VDD(VDD),.Y(g9911),.A(g2384));
  NOT NOT1_7638(.VSS(VSS),.VDD(VDD),.Y(g7495),.A(g4375));
  NOT NOT1_7639(.VSS(VSS),.VDD(VDD),.Y(g14545),.A(g12768));
  NOT NOT1_7640(.VSS(VSS),.VDD(VDD),.Y(g7437),.A(g5666));
  NOT NOT1_7641(.VSS(VSS),.VDD(VDD),.Y(g17610),.A(g15008));
  NOT NOT1_7642(.VSS(VSS),.VDD(VDD),.Y(I27253),.A(g27996));
  NOT NOT1_7643(.VSS(VSS),.VDD(VDD),.Y(I30995),.A(g32449));
  NOT NOT1_7644(.VSS(VSS),.VDD(VDD),.Y(g12838),.A(g10353));
  NOT NOT1_7645(.VSS(VSS),.VDD(VDD),.Y(g23128),.A(g20283));
  NOT NOT1_7646(.VSS(VSS),.VDD(VDD),.Y(I20569),.A(g16486));
  NOT NOT1_7647(.VSS(VSS),.VDD(VDD),.Y(I17852),.A(g3625));
  NOT NOT1_7648(.VSS(VSS),.VDD(VDD),.Y(g10078),.A(g1854));
  NOT NOT1_7649(.VSS(VSS),.VDD(VDD),.Y(g21245),.A(I20982));
  NOT NOT1_7650(.VSS(VSS),.VDD(VDD),.Y(g24019),.A(g19968));
  NOT NOT1_7651(.VSS(VSS),.VDD(VDD),.Y(g17189),.A(g14708));
  NOT NOT1_7652(.VSS(VSS),.VDD(VDD),.Y(g23245),.A(g20785));
  NOT NOT1_7653(.VSS(VSS),.VDD(VDD),.Y(I13287),.A(g110));
  NOT NOT1_7654(.VSS(VSS),.VDD(VDD),.Y(g26769),.A(g25400));
  NOT NOT1_7655(.VSS(VSS),.VDD(VDD),.Y(g8526),.A(g1526));
  NOT NOT1_7656(.VSS(VSS),.VDD(VDD),.Y(g19208),.A(g17367));
  NOT NOT1_7657(.VSS(VSS),.VDD(VDD),.Y(g20695),.A(I20781));
  NOT NOT1_7658(.VSS(VSS),.VDD(VDD),.Y(I20747),.A(g17141));
  NOT NOT1_7659(.VSS(VSS),.VDD(VDD),.Y(I31701),.A(g33164));
  NOT NOT1_7660(.VSS(VSS),.VDD(VDD),.Y(g21299),.A(g16600));
  NOT NOT1_7661(.VSS(VSS),.VDD(VDD),.Y(g30113),.A(g29154));
  NOT NOT1_7662(.VSS(VSS),.VDD(VDD),.Y(g9733),.A(g5736));
  NOT NOT1_7663(.VSS(VSS),.VDD(VDD),.Y(g10086),.A(g2193));
  NOT NOT1_7664(.VSS(VSS),.VDD(VDD),.Y(g23323),.A(g20283));
  NOT NOT1_7665(.VSS(VSS),.VDD(VDD),.Y(g23299),.A(I22400));
  NOT NOT1_7666(.VSS(VSS),.VDD(VDD),.Y(g9974),.A(g2518));
  NOT NOT1_7667(.VSS(VSS),.VDD(VDD),.Y(I32067),.A(g33661));
  NOT NOT1_7668(.VSS(VSS),.VDD(VDD),.Y(g17188),.A(I18224));
  NOT NOT1_7669(.VSS(VSS),.VDD(VDD),.Y(I11721),.A(g4145));
  NOT NOT1_7670(.VSS(VSS),.VDD(VDD),.Y(g17124),.A(g14051));
  NOT NOT1_7671(.VSS(VSS),.VDD(VDD),.Y(g17678),.A(I18653));
  NOT NOT1_7672(.VSS(VSS),.VDD(VDD),.Y(g34787),.A(I32991));
  NOT NOT1_7673(.VSS(VSS),.VDD(VDD),.Y(g26803),.A(g25389));
  NOT NOT1_7674(.VSS(VSS),.VDD(VDD),.Y(g12487),.A(g9340));
  NOT NOT1_7675(.VSS(VSS),.VDD(VDD),.Y(g20526),.A(g15171));
  NOT NOT1_7676(.VSS(VSS),.VDD(VDD),.Y(I22576),.A(g21282));
  NOT NOT1_7677(.VSS(VSS),.VDD(VDD),.Y(I28185),.A(g28803));
  NOT NOT1_7678(.VSS(VSS),.VDD(VDD),.Y(I18835),.A(g6365));
  NOT NOT1_7679(.VSS(VSS),.VDD(VDD),.Y(I13054),.A(g6744));
  NOT NOT1_7680(.VSS(VSS),.VDD(VDD),.Y(g24526),.A(g22942));
  NOT NOT1_7681(.VSS(VSS),.VDD(VDD),.Y(g19542),.A(g16349));
  NOT NOT1_7682(.VSS(VSS),.VDD(VDD),.Y(g30302),.A(g28924));
  NOT NOT1_7683(.VSS(VSS),.VDD(VDD),.Y(g7752),.A(g1542));
  NOT NOT1_7684(.VSS(VSS),.VDD(VDD),.Y(I16181),.A(g3672));
  NOT NOT1_7685(.VSS(VSS),.VDD(VDD),.Y(g18102),.A(I18912));
  NOT NOT1_7686(.VSS(VSS),.VDD(VDD),.Y(g8439),.A(g3129));
  NOT NOT1_7687(.VSS(VSS),.VDD(VDD),.Y(g9073),.A(g150));
  NOT NOT1_7688(.VSS(VSS),.VDD(VDD),.Y(g32629),.A(g31376));
  NOT NOT1_7689(.VSS(VSS),.VDD(VDD),.Y(g34302),.A(I32305));
  NOT NOT1_7690(.VSS(VSS),.VDD(VDD),.Y(I26989),.A(g27277));
  NOT NOT1_7691(.VSS(VSS),.VDD(VDD),.Y(I32150),.A(g33923));
  NOT NOT1_7692(.VSS(VSS),.VDD(VDD),.Y(g30105),.A(I28336));
  NOT NOT1_7693(.VSS(VSS),.VDD(VDD),.Y(g6836),.A(g1322));
  NOT NOT1_7694(.VSS(VSS),.VDD(VDD),.Y(g7917),.A(g1157));
  NOT NOT1_7695(.VSS(VSS),.VDD(VDD),.Y(I14630),.A(g7717));
  NOT NOT1_7696(.VSS(VSS),.VDD(VDD),.Y(g27279),.A(g26330));
  NOT NOT1_7697(.VSS(VSS),.VDD(VDD),.Y(g32472),.A(g30825));
  NOT NOT1_7698(.VSS(VSS),.VDD(VDD),.Y(g10159),.A(g4477));
  NOT NOT1_7699(.VSS(VSS),.VDD(VDD),.Y(g34827),.A(I33041));
  NOT NOT1_7700(.VSS(VSS),.VDD(VDD),.Y(g10532),.A(g10233));
  NOT NOT1_7701(.VSS(VSS),.VDD(VDD),.Y(g32628),.A(g31542));
  NOT NOT1_7702(.VSS(VSS),.VDD(VDD),.Y(g17093),.A(I18165));
  NOT NOT1_7703(.VSS(VSS),.VDD(VDD),.Y(g6918),.A(g3639));
  NOT NOT1_7704(.VSS(VSS),.VDD(VDD),.Y(g32911),.A(g31376));
  NOT NOT1_7705(.VSS(VSS),.VDD(VDD),.Y(g14125),.A(I16345));
  NOT NOT1_7706(.VSS(VSS),.VDD(VDD),.Y(g15344),.A(g14851));
  NOT NOT1_7707(.VSS(VSS),.VDD(VDD),.Y(g10158),.A(g2461));
  NOT NOT1_7708(.VSS(VSS),.VDD(VDD),.Y(g11403),.A(g7595));
  NOT NOT1_7709(.VSS(VSS),.VDD(VDD),.Y(g11547),.A(I14505));
  NOT NOT1_7710(.VSS(VSS),.VDD(VDD),.Y(g13895),.A(I16193));
  NOT NOT1_7711(.VSS(VSS),.VDD(VDD),.Y(g20917),.A(g15224));
  NOT NOT1_7712(.VSS(VSS),.VDD(VDD),.Y(I33140),.A(g34884));
  NOT NOT1_7713(.VSS(VSS),.VDD(VDD),.Y(I28883),.A(g30105));
  NOT NOT1_7714(.VSS(VSS),.VDD(VDD),.Y(g23232),.A(I22331));
  NOT NOT1_7715(.VSS(VSS),.VDD(VDD),.Y(g24866),.A(I24038));
  NOT NOT1_7716(.VSS(VSS),.VDD(VDD),.Y(g19905),.A(g15885));
  NOT NOT1_7717(.VSS(VSS),.VDD(VDD),.Y(I12790),.A(g4340));
  NOT NOT1_7718(.VSS(VSS),.VDD(VDD),.Y(I17609),.A(g13510));
  NOT NOT1_7719(.VSS(VSS),.VDD(VDD),.Y(g34769),.A(I32953));
  NOT NOT1_7720(.VSS(VSS),.VDD(VDD),.Y(I11655),.A(g1246));
  NOT NOT1_7721(.VSS(VSS),.VDD(VDD),.Y(g18876),.A(g15373));
  NOT NOT1_7722(.VSS(VSS),.VDD(VDD),.Y(g18885),.A(g15979));
  NOT NOT1_7723(.VSS(VSS),.VDD(VDD),.Y(g10353),.A(g6803));
  NOT NOT1_7724(.VSS(VSS),.VDD(VDD),.Y(g25046),.A(g23729));
  NOT NOT1_7725(.VSS(VSS),.VDD(VDD),.Y(g6993),.A(g4859));
  NOT NOT1_7726(.VSS(VSS),.VDD(VDD),.Y(g10295),.A(I13723));
  NOT NOT1_7727(.VSS(VSS),.VDD(VDD),.Y(g8919),.A(I12896));
  NOT NOT1_7728(.VSS(VSS),.VDD(VDD),.Y(g21697),.A(I21258));
  NOT NOT1_7729(.VSS(VSS),.VDD(VDD),.Y(g29013),.A(I27368));
  NOT NOT1_7730(.VSS(VSS),.VDD(VDD),.Y(I29981),.A(g31591));
  NOT NOT1_7731(.VSS(VSS),.VDD(VDD),.Y(g34768),.A(I32950));
  NOT NOT1_7732(.VSS(VSS),.VDD(VDD),.Y(g12039),.A(I14899));
  NOT NOT1_7733(.VSS(VSS),.VDD(VDD),.Y(g13715),.A(g10573));
  NOT NOT1_7734(.VSS(VSS),.VDD(VDD),.Y(I22745),.A(g19458));
  NOT NOT1_7735(.VSS(VSS),.VDD(VDD),.Y(g29214),.A(I27558));
  NOT NOT1_7736(.VSS(VSS),.VDD(VDD),.Y(g27038),.A(g25932));
  NOT NOT1_7737(.VSS(VSS),.VDD(VDD),.Y(g9206),.A(g5164));
  NOT NOT1_7738(.VSS(VSS),.VDD(VDD),.Y(g32591),.A(g30614));
  NOT NOT1_7739(.VSS(VSS),.VDD(VDD),.Y(I15572),.A(g10499));
  NOT NOT1_7740(.VSS(VSS),.VDD(VDD),.Y(g23995),.A(g19277));
  NOT NOT1_7741(.VSS(VSS),.VDD(VDD),.Y(g32776),.A(g31672));
  NOT NOT1_7742(.VSS(VSS),.VDD(VDD),.Y(g32785),.A(g31710));
  NOT NOT1_7743(.VSS(VSS),.VDD(VDD),.Y(I30989),.A(g32441));
  NOT NOT1_7744(.VSS(VSS),.VDD(VDD),.Y(g19565),.A(g16000));
  NOT NOT1_7745(.VSS(VSS),.VDD(VDD),.Y(g24077),.A(g20720));
  NOT NOT1_7746(.VSS(VSS),.VDD(VDD),.Y(g20706),.A(g18008));
  NOT NOT1_7747(.VSS(VSS),.VDD(VDD),.Y(I11734),.A(g4473));
  NOT NOT1_7748(.VSS(VSS),.VDD(VDD),.Y(g23880),.A(g19210));
  NOT NOT1_7749(.VSS(VSS),.VDD(VDD),.Y(g12038),.A(I14896));
  NOT NOT1_7750(.VSS(VSS),.VDD(VDD),.Y(g20597),.A(g17847));
  NOT NOT1_7751(.VSS(VSS),.VDD(VDD),.Y(I21042),.A(g15824));
  NOT NOT1_7752(.VSS(VSS),.VDD(VDD),.Y(g32754),.A(g30825));
  NOT NOT1_7753(.VSS(VSS),.VDD(VDD),.Y(I14570),.A(g7932));
  NOT NOT1_7754(.VSS(VSS),.VDD(VDD),.Y(g33435),.A(I30959));
  NOT NOT1_7755(.VSS(VSS),.VDD(VDD),.Y(g25282),.A(g22763));
  NOT NOT1_7756(.VSS(VSS),.VDD(VDD),.Y(I21189),.A(g17475));
  NOT NOT1_7757(.VSS(VSS),.VDD(VDD),.Y(g14336),.A(I16498));
  NOT NOT1_7758(.VSS(VSS),.VDD(VDD),.Y(g27187),.A(I25882));
  NOT NOT1_7759(.VSS(VSS),.VDD(VDD),.Y(g7296),.A(g5313));
  NOT NOT1_7760(.VSS(VSS),.VDD(VDD),.Y(g23512),.A(g20248));
  NOT NOT1_7761(.VSS(VSS),.VDD(VDD),.Y(g8616),.A(g2803));
  NOT NOT1_7762(.VSS(VSS),.VDD(VDD),.Y(g28752),.A(I27232));
  NOT NOT1_7763(.VSS(VSS),.VDD(VDD),.Y(g20923),.A(g15277));
  NOT NOT1_7764(.VSS(VSS),.VDD(VDD),.Y(g27975),.A(g26694));
  NOT NOT1_7765(.VSS(VSS),.VDD(VDD),.Y(g32859),.A(g30614));
  NOT NOT1_7766(.VSS(VSS),.VDD(VDD),.Y(g32825),.A(g30735));
  NOT NOT1_7767(.VSS(VSS),.VDD(VDD),.Y(g32950),.A(g31672));
  NOT NOT1_7768(.VSS(VSS),.VDD(VDD),.Y(g28954),.A(g27830));
  NOT NOT1_7769(.VSS(VSS),.VDD(VDD),.Y(g26710),.A(g25349));
  NOT NOT1_7770(.VSS(VSS),.VDD(VDD),.Y(g18660),.A(I19484));
  NOT NOT1_7771(.VSS(VSS),.VDD(VDD),.Y(g20624),.A(g18065));
  NOT NOT1_7772(.VSS(VSS),.VDD(VDD),.Y(g22455),.A(g19801));
  NOT NOT1_7773(.VSS(VSS),.VDD(VDD),.Y(g12975),.A(g12752));
  NOT NOT1_7774(.VSS(VSS),.VDD(VDD),.Y(g7532),.A(g1157));
  NOT NOT1_7775(.VSS(VSS),.VDD(VDD),.Y(I13694),.A(g117));
  NOT NOT1_7776(.VSS(VSS),.VDD(VDD),.Y(I16024),.A(g11171));
  NOT NOT1_7777(.VSS(VSS),.VDD(VDD),.Y(g32858),.A(g31327));
  NOT NOT1_7778(.VSS(VSS),.VDD(VDD),.Y(g33744),.A(I31604));
  NOT NOT1_7779(.VSS(VSS),.VDD(VDD),.Y(g7553),.A(g1274));
  NOT NOT1_7780(.VSS(VSS),.VDD(VDD),.Y(g8404),.A(g5005));
  NOT NOT1_7781(.VSS(VSS),.VDD(VDD),.Y(g15506),.A(I17131));
  NOT NOT1_7782(.VSS(VSS),.VDD(VDD),.Y(g31849),.A(g29385));
  NOT NOT1_7783(.VSS(VSS),.VDD(VDD),.Y(g8647),.A(g3416));
  NOT NOT1_7784(.VSS(VSS),.VDD(VDD),.Y(g14631),.A(g12239));
  NOT NOT1_7785(.VSS(VSS),.VDD(VDD),.Y(g10364),.A(g6869));
  NOT NOT1_7786(.VSS(VSS),.VDD(VDD),.Y(g19409),.A(g16431));
  NOT NOT1_7787(.VSS(VSS),.VDD(VDD),.Y(I14567),.A(g9708));
  NOT NOT1_7788(.VSS(VSS),.VDD(VDD),.Y(g12143),.A(I14999));
  NOT NOT1_7789(.VSS(VSS),.VDD(VDD),.Y(g20102),.A(g17533));
  NOT NOT1_7790(.VSS(VSS),.VDD(VDD),.Y(g16767),.A(I17989));
  NOT NOT1_7791(.VSS(VSS),.VDD(VDD),.Y(g20157),.A(g16886));
  NOT NOT1_7792(.VSS(VSS),.VDD(VDD),.Y(g25640),.A(I24781));
  NOT NOT1_7793(.VSS(VSS),.VDD(VDD),.Y(g12937),.A(g12419));
  NOT NOT1_7794(.VSS(VSS),.VDD(VDD),.Y(g28669),.A(g27705));
  NOT NOT1_7795(.VSS(VSS),.VDD(VDD),.Y(g26081),.A(g24619));
  NOT NOT1_7796(.VSS(VSS),.VDD(VDD),.Y(g8764),.A(g4826));
  NOT NOT1_7797(.VSS(VSS),.VDD(VDD),.Y(g22201),.A(g19277));
  NOT NOT1_7798(.VSS(VSS),.VDD(VDD),.Y(g24102),.A(g21143));
  NOT NOT1_7799(.VSS(VSS),.VDD(VDD),.Y(g23445),.A(I22564));
  NOT NOT1_7800(.VSS(VSS),.VDD(VDD),.Y(g31848),.A(g29385));
  NOT NOT1_7801(.VSS(VSS),.VDD(VDD),.Y(g18916),.A(g16053));
  NOT NOT1_7802(.VSS(VSS),.VDD(VDD),.Y(g24157),.A(I23315));
  NOT NOT1_7803(.VSS(VSS),.VDD(VDD),.Y(g32844),.A(g30937));
  NOT NOT1_7804(.VSS(VSS),.VDD(VDD),.Y(g9898),.A(g6444));
//
  AND2 AND2_0(.VSS(VSS),.VDD(VDD),.Y(g33848),.A(g33261),.B(g20384));
  AND2 AND2_1(.VSS(VSS),.VDD(VDD),.Y(g28260),.A(g27703),.B(g26518));
  AND2 AND2_2(.VSS(VSS),.VDD(VDD),.Y(g17617),.A(g7885),.B(g13326));
  AND2 AND2_3(.VSS(VSS),.VDD(VDD),.Y(g18550),.A(g2819),.B(g15277));
  AND2 AND2_4(.VSS(VSS),.VDD(VDD),.Y(g25768),.A(g2912),.B(g24560));
  AND2 AND2_5(.VSS(VSS),.VDD(VDD),.Y(g25803),.A(g24798),.B(g21024));
  AND2 AND2_6(.VSS(VSS),.VDD(VDD),.Y(g31141),.A(g12224),.B(g30038));
  AND3 AND3_0(.VSS(VSS),.VDD(VDD),.Y(I26960),.A(g24995),.B(g26424),.C(g22698));
  AND2 AND2_7(.VSS(VSS),.VDD(VDD),.Y(g22075),.A(g6247),.B(g19210));
  AND2 AND2_8(.VSS(VSS),.VDD(VDD),.Y(g18314),.A(g1585),.B(g16931));
  AND2 AND2_9(.VSS(VSS),.VDD(VDD),.Y(g33652),.A(g33393),.B(g18889));
  AND2 AND2_10(.VSS(VSS),.VDD(VDD),.Y(g18287),.A(g1442),.B(g16449));
  AND2 AND2_11(.VSS(VSS),.VDD(VDD),.Y(g27410),.A(g26549),.B(g17527));
  AND2 AND2_12(.VSS(VSS),.VDD(VDD),.Y(g16633),.A(g5196),.B(g14921));
  AND2 AND2_13(.VSS(VSS),.VDD(VDD),.Y(g30248),.A(g28743),.B(g23938));
  AND2 AND2_14(.VSS(VSS),.VDD(VDD),.Y(g34482),.A(g34405),.B(g18917));
  AND2 AND2_15(.VSS(VSS),.VDD(VDD),.Y(g23498),.A(g20234),.B(g12998));
  AND2 AND2_16(.VSS(VSS),.VDD(VDD),.Y(g28489),.A(g27010),.B(g12417));
  AND2 AND2_17(.VSS(VSS),.VDD(VDD),.Y(g26356),.A(g15581),.B(g25523));
  AND2 AND2_18(.VSS(VSS),.VDD(VDD),.Y(g18307),.A(g1559),.B(g16931));
  AND2 AND2_19(.VSS(VSS),.VDD(VDD),.Y(g29771),.A(g28322),.B(g23242));
  AND2 AND2_20(.VSS(VSS),.VDD(VDD),.Y(g30003),.A(g28149),.B(g9021));
  AND2 AND2_21(.VSS(VSS),.VDD(VDD),.Y(g34710),.A(g34553),.B(g20903));
  AND2 AND2_22(.VSS(VSS),.VDD(VDD),.Y(g16191),.A(g5475),.B(g14262));
  AND2 AND2_23(.VSS(VSS),.VDD(VDD),.Y(g22623),.A(g19337),.B(g19470));
  AND2 AND2_24(.VSS(VSS),.VDD(VDD),.Y(g21989),.A(g5587),.B(g19074));
  AND2 AND2_25(.VSS(VSS),.VDD(VDD),.Y(g30204),.A(g28670),.B(g23868));
  AND2 AND2_26(.VSS(VSS),.VDD(VDD),.Y(g13671),.A(g4498),.B(g10532));
  AND2 AND2_27(.VSS(VSS),.VDD(VDD),.Y(g26826),.A(g24907),.B(g15747));
  AND2 AND2_28(.VSS(VSS),.VDD(VDD),.Y(g27666),.A(g26865),.B(g23521));
  AND4 AND4_0(.VSS(VSS),.VDD(VDD),.Y(I31246),.A(g31672),.B(g31839),.C(g32810),.D(g32811));
  AND2 AND2_29(.VSS(VSS),.VDD(VDD),.Y(g18721),.A(g15138),.B(g16077));
  AND2 AND2_30(.VSS(VSS),.VDD(VDD),.Y(g22037),.A(g5941),.B(g19147));
  AND2 AND2_31(.VSS(VSS),.VDD(VDD),.Y(g25881),.A(g3821),.B(g24685));
  AND2 AND2_32(.VSS(VSS),.VDD(VDD),.Y(g26380),.A(g19572),.B(g25547));
  AND2 AND2_33(.VSS(VSS),.VDD(VDD),.Y(g33263),.A(g32393),.B(g25481));
  AND2 AND2_34(.VSS(VSS),.VDD(VDD),.Y(g18596),.A(g2941),.B(g16349));
  AND2 AND2_35(.VSS(VSS),.VDD(VDD),.Y(g32420),.A(g31127),.B(g19533));
  AND2 AND2_36(.VSS(VSS),.VDD(VDD),.Y(g28488),.A(g27969),.B(g17713));
  AND2 AND2_37(.VSS(VSS),.VDD(VDD),.Y(g27363),.A(g10231),.B(g26812));
  AND2 AND2_38(.VSS(VSS),.VDD(VDD),.Y(g23056),.A(g16052),.B(g19860));
  AND3 AND3_1(.VSS(VSS),.VDD(VDD),.Y(g27217),.A(g26236),.B(g8418),.C(g2610));
  AND2 AND2_39(.VSS(VSS),.VDD(VDD),.Y(g29683),.A(g1821),.B(g29046));
  AND2 AND2_40(.VSS(VSS),.VDD(VDD),.Y(g18243),.A(g1189),.B(g16431));
  AND2 AND2_41(.VSS(VSS),.VDD(VDD),.Y(g33332),.A(g32217),.B(g20608));
  AND3 AND3_2(.VSS(VSS),.VDD(VDD),.Y(I17692),.A(g14988),.B(g11450),.C(g6756));
  AND2 AND2_42(.VSS(VSS),.VDD(VDD),.Y(g21988),.A(g5583),.B(g19074));
  AND2 AND2_43(.VSS(VSS),.VDD(VDD),.Y(g26090),.A(g1624),.B(g25081));
  AND2 AND2_44(.VSS(VSS),.VDD(VDD),.Y(g21924),.A(g5057),.B(g21468));
  AND2 AND2_45(.VSS(VSS),.VDD(VDD),.Y(g28558),.A(g7301),.B(g27046));
  AND2 AND2_46(.VSS(VSS),.VDD(VDD),.Y(g18431),.A(g2185),.B(g18008));
  AND2 AND2_47(.VSS(VSS),.VDD(VDD),.Y(g26233),.A(g2279),.B(g25309));
  AND4 AND4_1(.VSS(VSS),.VDD(VDD),.Y(I31071),.A(g31170),.B(g31808),.C(g32557),.D(g32558));
  AND2 AND2_48(.VSS(VSS),.VDD(VDD),.Y(g26182),.A(g9978),.B(g25317));
  AND2 AND2_49(.VSS(VSS),.VDD(VDD),.Y(g26651),.A(g22707),.B(g24425));
  AND2 AND2_50(.VSS(VSS),.VDD(VDD),.Y(g12015),.A(g1002),.B(g7567));
  AND2 AND2_51(.VSS(VSS),.VDD(VDD),.Y(g34081),.A(g33706),.B(g19552));
  AND2 AND2_52(.VSS(VSS),.VDD(VDD),.Y(g27486),.A(g26519),.B(g17645));
  AND2 AND2_53(.VSS(VSS),.VDD(VDD),.Y(g31962),.A(g8033),.B(g31013));
  AND2 AND2_54(.VSS(VSS),.VDD(VDD),.Y(g24763),.A(g17569),.B(g22457));
  AND2 AND2_55(.VSS(VSS),.VDD(VDD),.Y(g33406),.A(g32355),.B(g21399));
  AND2 AND2_56(.VSS(VSS),.VDD(VDD),.Y(g18269),.A(g15069),.B(g16031));
  AND2 AND2_57(.VSS(VSS),.VDD(VDD),.Y(g33361),.A(g32257),.B(g20911));
  AND2 AND2_58(.VSS(VSS),.VDD(VDD),.Y(g15903),.A(g13796),.B(g13223));
  AND2 AND2_59(.VSS(VSS),.VDD(VDD),.Y(g18773),.A(g5694),.B(g15615));
  AND4 AND4_2(.VSS(VSS),.VDD(VDD),.Y(I31147),.A(g32668),.B(g32669),.C(g32670),.D(g32671));
  AND2 AND2_60(.VSS(VSS),.VDD(VDD),.Y(g18341),.A(g1648),.B(g17873));
  AND2 AND2_61(.VSS(VSS),.VDD(VDD),.Y(g29515),.A(g28888),.B(g22342));
  AND2 AND2_62(.VSS(VSS),.VDD(VDD),.Y(g29882),.A(g2361),.B(g29151));
  AND2 AND2_63(.VSS(VSS),.VDD(VDD),.Y(g18268),.A(g1280),.B(g16000));
  AND2 AND2_64(.VSS(VSS),.VDD(VDD),.Y(g29991),.A(g29179),.B(g12922));
  AND2 AND2_65(.VSS(VSS),.VDD(VDD),.Y(g21753),.A(g3179),.B(g20785));
  AND2 AND2_66(.VSS(VSS),.VDD(VDD),.Y(g31500),.A(g29802),.B(g23449));
  AND2 AND2_67(.VSS(VSS),.VDD(VDD),.Y(g18156),.A(g572),.B(g17533));
  AND2 AND2_68(.VSS(VSS),.VDD(VDD),.Y(g18655),.A(g15106),.B(g14454));
  AND3 AND3_3(.VSS(VSS),.VDD(VDD),.Y(g33500),.A(g32744),.B(I31196),.C(I31197));
  AND2 AND2_69(.VSS(VSS),.VDD(VDD),.Y(g24660),.A(g22648),.B(g19737));
  AND2 AND2_70(.VSS(VSS),.VDD(VDD),.Y(g33833),.A(g33093),.B(g25852));
  AND2 AND2_71(.VSS(VSS),.VDD(VDD),.Y(g32203),.A(g4249),.B(g31327));
  AND2 AND2_72(.VSS(VSS),.VDD(VDD),.Y(g18180),.A(g767),.B(g17328));
  AND2 AND2_73(.VSS(VSS),.VDD(VDD),.Y(g26513),.A(g19501),.B(g24365));
  AND2 AND2_74(.VSS(VSS),.VDD(VDD),.Y(g17418),.A(g9618),.B(g14407));
  AND3 AND3_4(.VSS(VSS),.VDD(VDD),.Y(I27409),.A(g25556),.B(g26424),.C(g22698));
  AND2 AND2_75(.VSS(VSS),.VDD(VDD),.Y(g34999),.A(g34998),.B(g23085));
  AND2 AND2_76(.VSS(VSS),.VDD(VDD),.Y(g18670),.A(g4621),.B(g15758));
  AND2 AND2_77(.VSS(VSS),.VDD(VDD),.Y(g34380),.A(g34158),.B(g20571));
  AND3 AND3_5(.VSS(VSS),.VDD(VDD),.Y(g25482),.A(g5752),.B(g23816),.C(I24597));
  AND2 AND2_78(.VSS(VSS),.VDD(VDD),.Y(g32044),.A(g31483),.B(g20085));
  AND4 AND4_3(.VSS(VSS),.VDD(VDD),.Y(I24684),.A(g20014),.B(g24033),.C(g24034),.D(g24035));
  AND2 AND2_79(.VSS(VSS),.VDD(VDD),.Y(g16612),.A(g5603),.B(g14927));
  AND2 AND2_80(.VSS(VSS),.VDD(VDD),.Y(g21736),.A(g3065),.B(g20330));
  AND2 AND2_81(.VSS(VSS),.VDD(VDD),.Y(g11546),.A(g7289),.B(g4375));
  AND2 AND2_82(.VSS(VSS),.VDD(VDD),.Y(g21887),.A(g15101),.B(g19801));
  AND2 AND2_83(.VSS(VSS),.VDD(VDD),.Y(g30233),.A(g28720),.B(g23913));
  AND2 AND2_84(.VSS(VSS),.VDD(VDD),.Y(g18734),.A(g4966),.B(g16826));
  AND4 AND4_4(.VSS(VSS),.VDD(VDD),.Y(I31151),.A(g30825),.B(g31822),.C(g32673),.D(g32674));
  AND2 AND2_85(.VSS(VSS),.VDD(VDD),.Y(g16324),.A(g13657),.B(g182));
  AND4 AND4_5(.VSS(VSS),.VDD(VDD),.Y(I31172),.A(g32703),.B(g32704),.C(g32705),.D(g32706));
  AND2 AND2_86(.VSS(VSS),.VDD(VDD),.Y(g18335),.A(g1687),.B(g17873));
  AND2 AND2_87(.VSS(VSS),.VDD(VDD),.Y(g16701),.A(g5547),.B(g14845));
  AND2 AND2_88(.VSS(VSS),.VDD(VDD),.Y(g22589),.A(g19267),.B(g19451));
  AND2 AND2_89(.VSS(VSS),.VDD(VDD),.Y(g32281),.A(g31257),.B(g20500));
  AND2 AND2_90(.VSS(VSS),.VDD(VDD),.Y(g34182),.A(g33691),.B(g24384));
  AND2 AND2_91(.VSS(VSS),.VDD(VDD),.Y(g28255),.A(g8515),.B(g27983));
  AND2 AND2_92(.VSS(VSS),.VDD(VDD),.Y(g16534),.A(g5575),.B(g14665));
  AND2 AND2_93(.VSS(VSS),.VDD(VDD),.Y(g28679),.A(g27572),.B(g20638));
  AND2 AND2_94(.VSS(VSS),.VDD(VDD),.Y(g11024),.A(g5436),.B(g9070));
  AND2 AND2_95(.VSS(VSS),.VDD(VDD),.Y(g16098),.A(g5148),.B(g14238));
  AND3 AND3_6(.VSS(VSS),.VDD(VDD),.Y(I13937),.A(g7340),.B(g7293),.C(g7261));
  AND2 AND2_96(.VSS(VSS),.VDD(VDD),.Y(g18993),.A(g11224),.B(g16172));
  AND2 AND2_97(.VSS(VSS),.VDD(VDD),.Y(g24550),.A(g3684),.B(g23308));
  AND2 AND2_98(.VSS(VSS),.VDD(VDD),.Y(g32301),.A(g31276),.B(g20547));
  AND2 AND2_99(.VSS(VSS),.VDD(VDD),.Y(g14643),.A(g11998),.B(g12023));
  AND2 AND2_100(.VSS(VSS),.VDD(VDD),.Y(g24314),.A(g4515),.B(g22228));
  AND2 AND2_101(.VSS(VSS),.VDD(VDD),.Y(g22588),.A(g79),.B(g20078));
  AND2 AND2_102(.VSS(VSS),.VDD(VDD),.Y(g21843),.A(g3869),.B(g21070));
  AND2 AND2_103(.VSS(VSS),.VDD(VDD),.Y(g32120),.A(g31639),.B(g29941));
  AND2 AND2_104(.VSS(VSS),.VDD(VDD),.Y(g24287),.A(g4401),.B(g22550));
  AND2 AND2_105(.VSS(VSS),.VDD(VDD),.Y(g28124),.A(g27368),.B(g22842));
  AND2 AND2_106(.VSS(VSS),.VDD(VDD),.Y(g15794),.A(g3239),.B(g14008));
  AND2 AND2_107(.VSS(VSS),.VDD(VDD),.Y(g18667),.A(g4601),.B(g17367));
  AND2 AND2_108(.VSS(VSS),.VDD(VDD),.Y(g18694),.A(g4722),.B(g16053));
  AND2 AND2_109(.VSS(VSS),.VDD(VDD),.Y(g12179),.A(g9745),.B(g10027));
  AND2 AND2_110(.VSS(VSS),.VDD(VDD),.Y(g24307),.A(g4486),.B(g22228));
  AND2 AND2_111(.VSS(VSS),.VDD(VDD),.Y(g29584),.A(g1706),.B(g29018));
  AND2 AND2_112(.VSS(VSS),.VDD(VDD),.Y(g27178),.A(g25997),.B(g16652));
  AND2 AND2_113(.VSS(VSS),.VDD(VDD),.Y(g21764),.A(g3227),.B(g20785));
  AND2 AND2_114(.VSS(VSS),.VDD(VDD),.Y(g11497),.A(g6398),.B(g7192));
  AND2 AND2_115(.VSS(VSS),.VDD(VDD),.Y(g18131),.A(g482),.B(g16971));
  AND3 AND3_7(.VSS(VSS),.VDD(VDD),.Y(g29206),.A(g24124),.B(I27528),.C(I27529));
  AND2 AND2_116(.VSS(VSS),.VDD(VDD),.Y(g13497),.A(g2724),.B(g12155));
  AND2 AND2_117(.VSS(VSS),.VDD(VDD),.Y(g28686),.A(g27574),.B(g20650));
  AND2 AND2_118(.VSS(VSS),.VDD(VDD),.Y(g32146),.A(g31624),.B(g29978));
  AND4 AND4_6(.VSS(VSS),.VDD(VDD),.Y(g28939),.A(g17321),.B(g25184),.C(g26424),.D(g27421));
  AND2 AND2_119(.VSS(VSS),.VDD(VDD),.Y(g24721),.A(g17488),.B(g22369));
  AND2 AND2_120(.VSS(VSS),.VDD(VDD),.Y(g22119),.A(g6581),.B(g19277));
  AND2 AND2_121(.VSS(VSS),.VDD(VDD),.Y(g21869),.A(g4087),.B(g19801));
  AND3 AND3_8(.VSS(VSS),.VDD(VDD),.Y(g27186),.A(g26195),.B(g8316),.C(g2342));
  AND2 AND2_122(.VSS(VSS),.VDD(VDD),.Y(g31273),.A(g30143),.B(g27779));
  AND2 AND2_123(.VSS(VSS),.VDD(VDD),.Y(g34513),.A(g9003),.B(g34346));
  AND2 AND2_124(.VSS(VSS),.VDD(VDD),.Y(g21960),.A(g5421),.B(g21514));
  AND2 AND2_125(.VSS(VSS),.VDD(VDD),.Y(g27676),.A(g26377),.B(g20627));
  AND2 AND2_126(.VSS(VSS),.VDD(VDD),.Y(g27685),.A(g13032),.B(g25895));
  AND2 AND2_127(.VSS(VSS),.VDD(VDD),.Y(g15633),.A(g3841),.B(g13584));
  AND2 AND2_128(.VSS(VSS),.VDD(VDD),.Y(g33106),.A(g32408),.B(g18990));
  AND2 AND2_129(.VSS(VSS),.VDD(VDD),.Y(g18487),.A(g2441),.B(g15426));
  AND2 AND2_130(.VSS(VSS),.VDD(VDD),.Y(g27373),.A(g26488),.B(g17477));
  AND2 AND2_131(.VSS(VSS),.VDD(VDD),.Y(g29759),.A(g28308),.B(g23226));
  AND2 AND2_132(.VSS(VSS),.VDD(VDD),.Y(g22118),.A(g6605),.B(g19277));
  AND2 AND2_133(.VSS(VSS),.VDD(VDD),.Y(g32290),.A(g31267),.B(g20525));
  AND2 AND2_134(.VSS(VSS),.VDD(VDD),.Y(g11126),.A(g6035),.B(g10185));
  AND2 AND2_135(.VSS(VSS),.VDD(VDD),.Y(g12186),.A(g1178),.B(g7519));
  AND3 AND3_9(.VSS(VSS),.VDD(VDD),.Y(g28267),.A(g7328),.B(g2227),.C(g27421));
  AND2 AND2_136(.VSS(VSS),.VDD(VDD),.Y(g17401),.A(g1083),.B(g13143));
  AND2 AND2_137(.VSS(VSS),.VDD(VDD),.Y(g21868),.A(g4076),.B(g19801));
  AND2 AND2_138(.VSS(VSS),.VDD(VDD),.Y(g18619),.A(g3466),.B(g17062));
  AND2 AND2_139(.VSS(VSS),.VDD(VDD),.Y(g18502),.A(g2567),.B(g15509));
  AND2 AND2_140(.VSS(VSS),.VDD(VDD),.Y(g22022),.A(g5873),.B(g19147));
  AND2 AND2_141(.VSS(VSS),.VDD(VDD),.Y(g34961),.A(g34944),.B(g23019));
  AND2 AND2_142(.VSS(VSS),.VDD(VDD),.Y(g12953),.A(g411),.B(g11048));
  AND2 AND2_143(.VSS(VSS),.VDD(VDD),.Y(g18557),.A(g2771),.B(g15277));
  AND3 AND3_10(.VSS(VSS),.VDD(VDD),.Y(g33812),.A(g23088),.B(g33187),.C(g9104));
  AND2 AND2_144(.VSS(VSS),.VDD(VDD),.Y(g18210),.A(g936),.B(g15938));
  AND2 AND2_145(.VSS(VSS),.VDD(VDD),.Y(g29758),.A(g28306),.B(g23222));
  AND2 AND2_146(.VSS(VSS),.VDD(VDD),.Y(g17119),.A(g5272),.B(g14800));
  AND3 AND3_11(.VSS(VSS),.VDD(VDD),.Y(g33463),.A(g32477),.B(I31011),.C(I31012));
  AND4 AND4_7(.VSS(VSS),.VDD(VDD),.Y(I31227),.A(g32784),.B(g32785),.C(g32786),.D(g32787));
  AND2 AND2_147(.VSS(VSS),.VDD(VDD),.Y(g18618),.A(g3457),.B(g17062));
  AND2 AND2_148(.VSS(VSS),.VDD(VDD),.Y(g18443),.A(g2265),.B(g18008));
  AND2 AND2_149(.VSS(VSS),.VDD(VDD),.Y(g24773),.A(g22832),.B(g19872));
  AND2 AND2_150(.VSS(VSS),.VDD(VDD),.Y(g21709),.A(g283),.B(g20283));
  AND2 AND2_151(.VSS(VSS),.VDD(VDD),.Y(g18279),.A(g1361),.B(g16136));
  AND2 AND2_152(.VSS(VSS),.VDD(VDD),.Y(g30026),.A(g28476),.B(g25064));
  AND2 AND2_153(.VSS(VSS),.VDD(VDD),.Y(g33371),.A(g32280),.B(g21155));
  AND2 AND2_154(.VSS(VSS),.VDD(VDD),.Y(g30212),.A(g28687),.B(g23879));
  AND2 AND2_155(.VSS(VSS),.VDD(VDD),.Y(g16766),.A(g6649),.B(g12915));
  AND2 AND2_156(.VSS(VSS),.VDD(VDD),.Y(g26387),.A(g24813),.B(g20231));
  AND2 AND2_157(.VSS(VSS),.VDD(VDD),.Y(g27334),.A(g12539),.B(g26769));
  AND2 AND2_158(.VSS(VSS),.VDD(VDD),.Y(g34212),.A(g33761),.B(g22689));
  AND2 AND2_159(.VSS(VSS),.VDD(VDD),.Y(g28219),.A(g9316),.B(g27573));
  AND2 AND2_160(.VSS(VSS),.VDD(VDD),.Y(g21708),.A(g15049),.B(g20283));
  AND2 AND2_161(.VSS(VSS),.VDD(VDD),.Y(g18278),.A(g1345),.B(g16136));
  AND3 AND3_12(.VSS(VSS),.VDD(VDD),.Y(I16111),.A(g8691),.B(g11409),.C(g11381));
  AND4 AND4_8(.VSS(VSS),.VDD(VDD),.Y(g26148),.A(g25357),.B(g11724),.C(g11709),.D(g11686));
  AND2 AND2_162(.VSS(VSS),.VDD(VDD),.Y(g23708),.A(g19050),.B(g9104));
  AND2 AND2_163(.VSS(VSS),.VDD(VDD),.Y(g16871),.A(g6597),.B(g14908));
  AND2 AND2_164(.VSS(VSS),.VDD(VDD),.Y(g29345),.A(g4749),.B(g28376));
  AND2 AND2_165(.VSS(VSS),.VDD(VDD),.Y(g22053),.A(g6116),.B(g21611));
  AND2 AND2_166(.VSS(VSS),.VDD(VDD),.Y(g23471),.A(g20148),.B(g20523));
  AND2 AND2_167(.VSS(VSS),.VDD(VDD),.Y(g26097),.A(g5821),.B(g25092));
  AND2 AND2_168(.VSS(VSS),.VDD(VDD),.Y(g18469),.A(g2399),.B(g15224));
  AND2 AND2_169(.VSS(VSS),.VDD(VDD),.Y(g24670),.A(g5138),.B(g23590));
  AND2 AND2_170(.VSS(VSS),.VDD(VDD),.Y(g33795),.A(g33138),.B(g20782));
  AND2 AND2_171(.VSS(VSS),.VDD(VDD),.Y(g28218),.A(g27768),.B(g26645));
  AND2 AND2_172(.VSS(VSS),.VDD(VDD),.Y(g29940),.A(g1740),.B(g28758));
  AND2 AND2_173(.VSS(VSS),.VDD(VDD),.Y(g26104),.A(g2250),.B(g25101));
  AND2 AND2_174(.VSS(VSS),.VDD(VDD),.Y(g18286),.A(g1404),.B(g16164));
  AND2 AND2_175(.VSS(VSS),.VDD(VDD),.Y(g22900),.A(g17137),.B(g19697));
  AND4 AND4_9(.VSS(VSS),.VDD(VDD),.Y(g27762),.A(g22472),.B(g25226),.C(g26424),.D(g26218));
  AND2 AND2_176(.VSS(VSS),.VDD(VDD),.Y(g15861),.A(g3957),.B(g14170));
  AND2 AND2_177(.VSS(VSS),.VDD(VDD),.Y(g8690),.A(g2941),.B(g2936));
  AND2 AND2_178(.VSS(VSS),.VDD(VDD),.Y(g27964),.A(g25956),.B(g22492));
  AND2 AND2_179(.VSS(VSS),.VDD(VDD),.Y(g18468),.A(g2393),.B(g15224));
  AND3 AND3_13(.VSS(VSS),.VDD(VDD),.Y(g25331),.A(g5366),.B(g22194),.C(I24508));
  AND2 AND2_180(.VSS(VSS),.VDD(VDD),.Y(g18306),.A(g15074),.B(g16931));
  AND2 AND2_181(.VSS(VSS),.VDD(VDD),.Y(g12762),.A(g4358),.B(g8977));
  AND2 AND2_182(.VSS(VSS),.VDD(VDD),.Y(g22036),.A(g5937),.B(g19147));
  AND2 AND2_183(.VSS(VSS),.VDD(VDD),.Y(g25449),.A(g6946),.B(g22496));
  AND2 AND2_184(.VSS(VSS),.VDD(VDD),.Y(g13060),.A(g8587),.B(g11110));
  AND2 AND2_185(.VSS(VSS),.VDD(VDD),.Y(g31514),.A(g20041),.B(g29956));
  AND2 AND2_186(.VSS(VSS),.VDD(VDD),.Y(g32403),.A(g31117),.B(g15842));
  AND2 AND2_187(.VSS(VSS),.VDD(VDD),.Y(g27216),.A(g26055),.B(g16725));
  AND3 AND3_14(.VSS(VSS),.VDD(VDD),.Y(g33514),.A(g32844),.B(I31266),.C(I31267));
  AND2 AND2_188(.VSS(VSS),.VDD(VDD),.Y(g22101),.A(g6474),.B(g18833));
  AND2 AND2_189(.VSS(VSS),.VDD(VDD),.Y(g24930),.A(g4826),.B(g23948));
  AND2 AND2_190(.VSS(VSS),.VDD(VDD),.Y(g29652),.A(g2667),.B(g29157));
  AND2 AND2_191(.VSS(VSS),.VDD(VDD),.Y(g29804),.A(g1592),.B(g29014));
  AND2 AND2_192(.VSS(VSS),.VDD(VDD),.Y(g17809),.A(g7873),.B(g13125));
  AND4 AND4_10(.VSS(VSS),.VDD(VDD),.Y(I31281),.A(g30735),.B(g31845),.C(g32861),.D(g32862));
  AND2 AND2_193(.VSS(VSS),.VDD(VDD),.Y(g28160),.A(g26309),.B(g27463));
  AND2 AND2_194(.VSS(VSS),.VDD(VDD),.Y(g15612),.A(g3143),.B(g13530));
  AND2 AND2_195(.VSS(VSS),.VDD(VDD),.Y(g25448),.A(g11202),.B(g22680));
  AND2 AND2_196(.VSS(VSS),.VDD(VDD),.Y(g18815),.A(g6523),.B(g15483));
  AND2 AND2_197(.VSS(VSS),.VDD(VDD),.Y(g30149),.A(g28605),.B(g21248));
  AND2 AND2_198(.VSS(VSS),.VDD(VDD),.Y(g25961),.A(g25199),.B(g20682));
  AND3 AND3_15(.VSS(VSS),.VDD(VDD),.Y(I27381),.A(g25549),.B(g26424),.C(g22698));
  AND3 AND3_16(.VSS(VSS),.VDD(VDD),.Y(g33507),.A(g32795),.B(I31231),.C(I31232));
  AND4 AND4_11(.VSS(VSS),.VDD(VDD),.Y(I31301),.A(g31327),.B(g31849),.C(g32889),.D(g32890));
  AND2 AND2_199(.VSS(VSS),.VDD(VDD),.Y(g20131),.A(g15170),.B(g14309));
  AND2 AND2_200(.VSS(VSS),.VDD(VDD),.Y(g15701),.A(g3821),.B(g13584));
  AND3 AND3_17(.VSS(VSS),.VDD(VDD),.Y(g10705),.A(g6850),.B(g10219),.C(g2689));
  AND2 AND2_201(.VSS(VSS),.VDD(VDD),.Y(g18601),.A(g3106),.B(g16987));
  AND2 AND2_202(.VSS(VSS),.VDD(VDD),.Y(g13411),.A(g4955),.B(g11834));
  AND2 AND2_203(.VSS(VSS),.VDD(VDD),.Y(g18187),.A(g794),.B(g17328));
  AND2 AND2_204(.VSS(VSS),.VDD(VDD),.Y(g18677),.A(g4639),.B(g15758));
  AND2 AND2_205(.VSS(VSS),.VDD(VDD),.Y(g14610),.A(g1484),.B(g10935));
  AND2 AND2_206(.VSS(VSS),.VDD(VDD),.Y(g28455),.A(g27289),.B(g20103));
  AND2 AND2_207(.VSS(VSS),.VDD(VDD),.Y(g33421),.A(g32374),.B(g21455));
  AND2 AND2_208(.VSS(VSS),.VDD(VDD),.Y(g21810),.A(g3578),.B(g20924));
  AND2 AND2_209(.VSS(VSS),.VDD(VDD),.Y(g17177),.A(g6657),.B(g14984));
  AND2 AND2_210(.VSS(VSS),.VDD(VDD),.Y(g21774),.A(g3361),.B(g20391));
  AND2 AND2_211(.VSS(VSS),.VDD(VDD),.Y(g29332),.A(g29107),.B(g22170));
  AND2 AND2_212(.VSS(VSS),.VDD(VDD),.Y(g23657),.A(g19401),.B(g11941));
  AND2 AND2_213(.VSS(VSS),.VDD(VDD),.Y(g28617),.A(g27533),.B(g20552));
  AND3 AND3_18(.VSS(VSS),.VDD(VDD),.Y(g34097),.A(g33772),.B(g9104),.C(g18957));
  AND2 AND2_214(.VSS(VSS),.VDD(VDD),.Y(g21955),.A(g5385),.B(g21514));
  AND2 AND2_215(.VSS(VSS),.VDD(VDD),.Y(g23774),.A(g14867),.B(g21252));
  AND2 AND2_216(.VSS(VSS),.VDD(VDD),.Y(g22064),.A(g15162),.B(g19210));
  AND3 AND3_19(.VSS(VSS),.VDD(VDD),.Y(I24600),.A(g6077),.B(g6082),.C(g9946));
  AND4 AND4_12(.VSS(VSS),.VDD(VDD),.Y(I31146),.A(g30735),.B(g31821),.C(g32666),.D(g32667));
  AND2 AND2_217(.VSS(VSS),.VDD(VDD),.Y(g25026),.A(g22929),.B(g10503));
  AND2 AND2_218(.VSS(VSS),.VDD(VDD),.Y(g34104),.A(g33916),.B(g23639));
  AND2 AND2_219(.VSS(VSS),.VDD(VDD),.Y(g27117),.A(g26055),.B(g16528));
  AND2 AND2_220(.VSS(VSS),.VDD(VDD),.Y(g21879),.A(g4132),.B(g19801));
  AND2 AND2_221(.VSS(VSS),.VDD(VDD),.Y(g34811),.A(g14165),.B(g34766));
  AND2 AND2_222(.VSS(VSS),.VDD(VDD),.Y(g21970),.A(g5401),.B(g21514));
  AND2 AND2_223(.VSS(VSS),.VDD(VDD),.Y(g18143),.A(g586),.B(g17533));
  AND2 AND2_224(.VSS(VSS),.VDD(VDD),.Y(g24502),.A(g23428),.B(g13223));
  AND2 AND2_225(.VSS(VSS),.VDD(VDD),.Y(g28201),.A(g27499),.B(g16720));
  AND2 AND2_226(.VSS(VSS),.VDD(VDD),.Y(g19536),.A(g518),.B(g16768));
  AND2 AND2_227(.VSS(VSS),.VDD(VDD),.Y(g19948),.A(g17515),.B(g16320));
  AND2 AND2_228(.VSS(VSS),.VDD(VDD),.Y(g29962),.A(g23616),.B(g28959));
  AND2 AND2_229(.VSS(VSS),.VDD(VDD),.Y(g21878),.A(g4129),.B(g19801));
  AND3 AND3_20(.VSS(VSS),.VDD(VDD),.Y(I16695),.A(g10207),.B(g12523),.C(g12463));
  AND2 AND2_230(.VSS(VSS),.VDD(VDD),.Y(g32127),.A(g31624),.B(g29950));
  AND2 AND2_231(.VSS(VSS),.VDD(VDD),.Y(g31541),.A(g22536),.B(g29348));
  AND2 AND2_232(.VSS(VSS),.VDD(VDD),.Y(g24618),.A(g22625),.B(g19672));
  AND2 AND2_233(.VSS(VSS),.VDD(VDD),.Y(g26229),.A(g1724),.B(g25275));
  AND3 AND3_21(.VSS(VSS),.VDD(VDD),.Y(g33473),.A(g32549),.B(I31061),.C(I31062));
  AND2 AND2_234(.VSS(VSS),.VDD(VDD),.Y(g18169),.A(g676),.B(g17433));
  AND2 AND2_235(.VSS(VSS),.VDD(VDD),.Y(g21886),.A(g4153),.B(g19801));
  AND2 AND2_236(.VSS(VSS),.VDD(VDD),.Y(g27568),.A(g26576),.B(g17791));
  AND2 AND2_237(.VSS(VSS),.VDD(VDD),.Y(g18791),.A(g6044),.B(g15634));
  AND2 AND2_238(.VSS(VSS),.VDD(VDD),.Y(g31789),.A(g30201),.B(g24013));
  AND2 AND2_239(.VSS(VSS),.VDD(VDD),.Y(g28467),.A(g26993),.B(g12295));
  AND2 AND2_240(.VSS(VSS),.VDD(VDD),.Y(g28494),.A(g27973),.B(g17741));
  AND2 AND2_241(.VSS(VSS),.VDD(VDD),.Y(g33789),.A(g33159),.B(g23022));
  AND2 AND2_242(.VSS(VSS),.VDD(VDD),.Y(g21792),.A(g3396),.B(g20391));
  AND2 AND2_243(.VSS(VSS),.VDD(VDD),.Y(g16591),.A(g5256),.B(g14879));
  AND2 AND2_244(.VSS(VSS),.VDD(VDD),.Y(g22009),.A(g5782),.B(g21562));
  AND2 AND2_245(.VSS(VSS),.VDD(VDD),.Y(g22665),.A(g17174),.B(g20905));
  AND2 AND2_246(.VSS(VSS),.VDD(VDD),.Y(g18168),.A(g681),.B(g17433));
  AND2 AND2_247(.VSS(VSS),.VDD(VDD),.Y(g18410),.A(g2079),.B(g15373));
  AND2 AND2_248(.VSS(VSS),.VDD(VDD),.Y(g21967),.A(g5456),.B(g21514));
  AND2 AND2_249(.VSS(VSS),.VDD(VDD),.Y(g21994),.A(g5607),.B(g19074));
  AND2 AND2_250(.VSS(VSS),.VDD(VDD),.Y(g31788),.A(g21352),.B(g29385));
  AND2 AND2_251(.VSS(VSS),.VDD(VDD),.Y(g33724),.A(g14145),.B(g33258));
  AND2 AND2_252(.VSS(VSS),.VDD(VDD),.Y(g32376),.A(g2689),.B(g31710));
  AND2 AND2_253(.VSS(VSS),.VDD(VDD),.Y(g19564),.A(g17175),.B(g13976));
  AND2 AND2_254(.VSS(VSS),.VDD(VDD),.Y(g33359),.A(g32252),.B(g20853));
  AND2 AND2_255(.VSS(VSS),.VDD(VDD),.Y(g25149),.A(g14030),.B(g23546));
  AND2 AND2_256(.VSS(VSS),.VDD(VDD),.Y(g17693),.A(g1306),.B(g13291));
  AND2 AND2_257(.VSS(VSS),.VDD(VDD),.Y(g22008),.A(g5774),.B(g21562));
  AND2 AND2_258(.VSS(VSS),.VDD(VDD),.Y(g32103),.A(g31609),.B(g29905));
  AND2 AND2_259(.VSS(VSS),.VDD(VDD),.Y(g24286),.A(g4405),.B(g22550));
  AND2 AND2_260(.VSS(VSS),.VDD(VDD),.Y(g18479),.A(g2449),.B(g15426));
  AND2 AND2_261(.VSS(VSS),.VDD(VDD),.Y(g18666),.A(g4593),.B(g17367));
  AND2 AND2_262(.VSS(VSS),.VDD(VDD),.Y(g33829),.A(g33240),.B(g20164));
  AND2 AND2_263(.VSS(VSS),.VDD(VDD),.Y(g18363),.A(g1840),.B(g17955));
  AND2 AND2_264(.VSS(VSS),.VDD(VDD),.Y(g32095),.A(g7619),.B(g30825));
  AND2 AND2_265(.VSS(VSS),.VDD(VDD),.Y(g18217),.A(g15063),.B(g16100));
  AND2 AND2_266(.VSS(VSS),.VDD(VDD),.Y(g33434),.A(g32239),.B(g29702));
  AND2 AND2_267(.VSS(VSS),.VDD(VDD),.Y(g24306),.A(g4483),.B(g22228));
  AND2 AND2_268(.VSS(VSS),.VDD(VDD),.Y(g33358),.A(g32249),.B(g20778));
  AND2 AND2_269(.VSS(VSS),.VDD(VDD),.Y(g25148),.A(g16867),.B(g23545));
  AND2 AND2_270(.VSS(VSS),.VDD(VDD),.Y(g11496),.A(g4382),.B(g7495));
  AND2 AND2_271(.VSS(VSS),.VDD(VDD),.Y(g15871),.A(g3203),.B(g13951));
  AND2 AND2_272(.VSS(VSS),.VDD(VDD),.Y(g18478),.A(g2445),.B(g15426));
  AND2 AND2_273(.VSS(VSS),.VDD(VDD),.Y(g30133),.A(g28591),.B(g21179));
  AND2 AND2_274(.VSS(VSS),.VDD(VDD),.Y(g33828),.A(g33090),.B(g24411));
  AND2 AND2_275(.VSS(VSS),.VDD(VDD),.Y(g28352),.A(g10014),.B(g27705));
  AND4 AND4_13(.VSS(VSS),.VDD(VDD),.Y(g11111),.A(g5297),.B(g7004),.C(g5283),.D(g9780));
  AND2 AND2_276(.VSS(VSS),.VDD(VDD),.Y(g14875),.A(g1495),.B(g10939));
  AND2 AND2_277(.VSS(VSS),.VDD(VDD),.Y(g34133),.A(g33845),.B(g23958));
  AND2 AND2_278(.VSS(VSS),.VDD(VDD),.Y(g21919),.A(g15144),.B(g21468));
  AND2 AND2_279(.VSS(VSS),.VDD(VDD),.Y(g30229),.A(g28716),.B(g23904));
  AND2 AND2_280(.VSS(VSS),.VDD(VDD),.Y(g25104),.A(g16800),.B(g23504));
  AND2 AND2_281(.VSS(VSS),.VDD(VDD),.Y(g11978),.A(g2629),.B(g7462));
  AND2 AND2_282(.VSS(VSS),.VDD(VDD),.Y(g26310),.A(g2102),.B(g25389));
  AND2 AND2_283(.VSS(VSS),.VDD(VDD),.Y(g23919),.A(g4122),.B(g19546));
  AND2 AND2_284(.VSS(VSS),.VDD(VDD),.Y(g32181),.A(g31020),.B(g19912));
  AND2 AND2_285(.VSS(VSS),.VDD(VDD),.Y(g33121),.A(g8748),.B(g32212));
  AND2 AND2_286(.VSS(VSS),.VDD(VDD),.Y(g18486),.A(g2485),.B(g15426));
  AND2 AND2_287(.VSS(VSS),.VDD(VDD),.Y(g27230),.A(g25906),.B(g19558));
  AND2 AND2_288(.VSS(VSS),.VDD(VDD),.Y(g27293),.A(g9972),.B(g26655));
  AND2 AND2_289(.VSS(VSS),.VDD(VDD),.Y(g29613),.A(g28208),.B(g19763));
  AND2 AND2_290(.VSS(VSS),.VDD(VDD),.Y(g28266),.A(g23748),.B(g27714));
  AND2 AND2_291(.VSS(VSS),.VDD(VDD),.Y(g19062),.A(g446),.B(g16180));
  AND2 AND2_292(.VSS(VSS),.VDD(VDD),.Y(g33344),.A(g32228),.B(g20670));
  AND2 AND2_293(.VSS(VSS),.VDD(VDD),.Y(g14218),.A(g875),.B(g10632));
  AND2 AND2_294(.VSS(VSS),.VDD(VDD),.Y(g21918),.A(g5097),.B(g21468));
  AND2 AND2_295(.VSS(VSS),.VDD(VDD),.Y(g30228),.A(g28715),.B(g23903));
  AND2 AND2_296(.VSS(VSS),.VDD(VDD),.Y(g26379),.A(g19904),.B(g25546));
  AND2 AND2_297(.VSS(VSS),.VDD(VDD),.Y(g18556),.A(g2823),.B(g15277));
  AND2 AND2_298(.VSS(VSS),.VDD(VDD),.Y(g25971),.A(g1917),.B(g24992));
  AND2 AND2_299(.VSS(VSS),.VDD(VDD),.Y(g24187),.A(g305),.B(g22722));
  AND2 AND2_300(.VSS(VSS),.VDD(VDD),.Y(g34228),.A(g33750),.B(g22942));
  AND2 AND2_301(.VSS(VSS),.VDD(VDD),.Y(g30011),.A(g29183),.B(g12930));
  AND2 AND2_302(.VSS(VSS),.VDD(VDD),.Y(g27265),.A(g26785),.B(g26759));
  AND4 AND4_14(.VSS(VSS),.VDD(VDD),.Y(I31226),.A(g29385),.B(g32781),.C(g32782),.D(g32783));
  AND2 AND2_303(.VSS(VSS),.VDD(VDD),.Y(g16844),.A(g7212),.B(g13000));
  AND2 AND2_304(.VSS(VSS),.VDD(VDD),.Y(g18580),.A(g2907),.B(g16349));
  AND2 AND2_305(.VSS(VSS),.VDD(VDD),.Y(g26050),.A(g9630),.B(g25047));
  AND4 AND4_15(.VSS(VSS),.VDD(VDD),.Y(g27416),.A(g8046),.B(g26314),.C(g9187),.D(g504));
  AND2 AND2_306(.VSS(VSS),.VDD(VDD),.Y(g26378),.A(g19576),.B(g25544));
  AND2 AND2_307(.VSS(VSS),.VDD(VDD),.Y(g13384),.A(g4944),.B(g11804));
  AND2 AND2_308(.VSS(VSS),.VDD(VDD),.Y(g29605),.A(g2445),.B(g28973));
  AND2 AND2_309(.VSS(VSS),.VDD(VDD),.Y(g18223),.A(g1030),.B(g16100));
  AND2 AND2_310(.VSS(VSS),.VDD(VDD),.Y(g23599),.A(g19050),.B(g9104));
  AND2 AND2_311(.VSS(VSS),.VDD(VDD),.Y(g27992),.A(g26800),.B(g23964));
  AND2 AND2_312(.VSS(VSS),.VDD(VDD),.Y(g22074),.A(g6239),.B(g19210));
  AND2 AND2_313(.VSS(VSS),.VDD(VDD),.Y(g27391),.A(g26549),.B(g17505));
  AND2 AND2_314(.VSS(VSS),.VDD(VDD),.Y(g24143),.A(g17694),.B(g21659));
  AND2 AND2_315(.VSS(VSS),.VDD(VDD),.Y(g25368),.A(g6946),.B(g22408));
  AND2 AND2_316(.VSS(VSS),.VDD(VDD),.Y(g27510),.A(g26576),.B(g17687));
  AND2 AND2_317(.VSS(VSS),.VDD(VDD),.Y(g34582),.A(g7764),.B(g34313));
  AND2 AND2_318(.VSS(VSS),.VDD(VDD),.Y(g32190),.A(g142),.B(g31233));
  AND2 AND2_319(.VSS(VSS),.VDD(VDD),.Y(g26096),.A(g9733),.B(g25268));
  AND2 AND2_320(.VSS(VSS),.VDD(VDD),.Y(g29951),.A(g1874),.B(g28786));
  AND2 AND2_321(.VSS(VSS),.VDD(VDD),.Y(g18110),.A(g441),.B(g17015));
  AND2 AND2_322(.VSS(VSS),.VDD(VDD),.Y(g34310),.A(g14003),.B(g34162));
  AND2 AND2_323(.VSS(VSS),.VDD(VDD),.Y(g25850),.A(g3502),.B(g24636));
  AND2 AND2_324(.VSS(VSS),.VDD(VDD),.Y(g15911),.A(g3111),.B(g13530));
  AND2 AND2_325(.VSS(VSS),.VDD(VDD),.Y(g28588),.A(g27489),.B(g20499));
  AND2 AND2_326(.VSS(VSS),.VDD(VDD),.Y(g28524),.A(g6821),.B(g27084));
  AND4 AND4_16(.VSS(VSS),.VDD(VDD),.Y(I31127),.A(g32638),.B(g32639),.C(g32640),.D(g32641));
  AND2 AND2_327(.VSS(VSS),.VDD(VDD),.Y(g18321),.A(g1620),.B(g17873));
  AND3 AND3_22(.VSS(VSS),.VDD(VDD),.Y(g24884),.A(g3401),.B(g23555),.C(I24051));
  AND2 AND2_328(.VSS(VSS),.VDD(VDD),.Y(g30925),.A(g29908),.B(g23309));
  AND2 AND2_329(.VSS(VSS),.VDD(VDD),.Y(g21817),.A(g3606),.B(g20924));
  AND2 AND2_330(.VSS(VSS),.VDD(VDD),.Y(g11019),.A(g5092),.B(g9036));
  AND2 AND2_331(.VSS(VSS),.VDD(VDD),.Y(g18179),.A(g763),.B(g17328));
  AND2 AND2_332(.VSS(VSS),.VDD(VDD),.Y(g13019),.A(g194),.B(g11737));
  AND2 AND2_333(.VSS(VSS),.VDD(VDD),.Y(g18531),.A(g2719),.B(g15277));
  AND2 AND2_334(.VSS(VSS),.VDD(VDD),.Y(g30112),.A(g28566),.B(g20919));
  AND2 AND2_335(.VSS(VSS),.VDD(VDD),.Y(g28477),.A(g27966),.B(g17676));
  AND2 AND2_336(.VSS(VSS),.VDD(VDD),.Y(g33760),.A(g33143),.B(g20328));
  AND2 AND2_337(.VSS(VSS),.VDD(VDD),.Y(g24410),.A(g3817),.B(g23139));
  AND2 AND2_338(.VSS(VSS),.VDD(VDD),.Y(g32089),.A(g27261),.B(g31021));
  AND2 AND2_339(.VSS(VSS),.VDD(VDD),.Y(g25229),.A(g7636),.B(g22654));
  AND2 AND2_340(.VSS(VSS),.VDD(VDD),.Y(g30050),.A(g22545),.B(g28126));
  AND2 AND2_341(.VSS(VSS),.VDD(VDD),.Y(g29795),.A(g28344),.B(g23257));
  AND3 AND3_23(.VSS(VSS),.VDD(VDD),.Y(g34112),.A(g22957),.B(g9104),.C(g33778));
  AND3 AND3_24(.VSS(VSS),.VDD(VDD),.Y(g11018),.A(g7655),.B(g7643),.C(g7627));
  AND2 AND2_342(.VSS(VSS),.VDD(VDD),.Y(g18178),.A(g758),.B(g17328));
  AND2 AND2_343(.VSS(VSS),.VDD(VDD),.Y(g18740),.A(g4572),.B(g17384));
  AND2 AND2_344(.VSS(VSS),.VDD(VDD),.Y(g26857),.A(g25062),.B(g25049));
  AND2 AND2_345(.VSS(VSS),.VDD(VDD),.Y(g34050),.A(g33772),.B(g22942));
  AND2 AND2_346(.VSS(VSS),.VDD(VDD),.Y(g21977),.A(g5535),.B(g19074));
  AND2 AND2_347(.VSS(VSS),.VDD(VDD),.Y(g22092),.A(g6419),.B(g18833));
  AND2 AND2_348(.VSS(VSS),.VDD(VDD),.Y(g23532),.A(g19400),.B(g11852));
  AND2 AND2_349(.VSS(VSS),.VDD(VDD),.Y(g23901),.A(g19606),.B(g7963));
  AND2 AND2_350(.VSS(VSS),.VDD(VDD),.Y(g34378),.A(g13095),.B(g34053));
  AND2 AND2_351(.VSS(VSS),.VDD(VDD),.Y(g16025),.A(g446),.B(g14063));
  AND3 AND3_25(.VSS(VSS),.VDD(VDD),.Y(g33506),.A(g32788),.B(I31226),.C(I31227));
  AND3 AND3_26(.VSS(VSS),.VDD(VDD),.Y(I24530),.A(g9501),.B(g9733),.C(g5747));
  AND2 AND2_352(.VSS(VSS),.VDD(VDD),.Y(g32088),.A(g27241),.B(g31070));
  AND2 AND2_353(.VSS(VSS),.VDD(VDD),.Y(g24666),.A(g11753),.B(g22975));
  AND2 AND2_354(.VSS(VSS),.VDD(VDD),.Y(g22518),.A(g12982),.B(g19398));
  AND2 AND2_355(.VSS(VSS),.VDD(VDD),.Y(g21783),.A(g3419),.B(g20391));
  AND4 AND4_17(.VSS(VSS),.VDD(VDD),.Y(I31297),.A(g32884),.B(g32885),.C(g32886),.D(g32887));
  AND2 AND2_356(.VSS(VSS),.VDD(VDD),.Y(g24217),.A(g18200),.B(g22594));
  AND2 AND2_357(.VSS(VSS),.VDD(VDD),.Y(g18186),.A(g753),.B(g17328));
  AND2 AND2_358(.VSS(VSS),.VDD(VDD),.Y(g15785),.A(g3558),.B(g14107));
  AND2 AND2_359(.VSS(VSS),.VDD(VDD),.Y(g18676),.A(g4358),.B(g15758));
  AND2 AND2_360(.VSS(VSS),.VDD(VDD),.Y(g18685),.A(g4688),.B(g15885));
  AND2 AND2_361(.VSS(VSS),.VDD(VDD),.Y(g34386),.A(g10800),.B(g34060));
  AND2 AND2_362(.VSS(VSS),.VDD(VDD),.Y(g18373),.A(g1890),.B(g15171));
  AND2 AND2_363(.VSS(VSS),.VDD(VDD),.Y(g29514),.A(g1608),.B(g28780));
  AND2 AND2_364(.VSS(VSS),.VDD(VDD),.Y(g24015),.A(g19540),.B(g10951));
  AND2 AND2_365(.VSS(VSS),.VDD(VDD),.Y(g30096),.A(g28546),.B(g20770));
  AND2 AND2_366(.VSS(VSS),.VDD(VDD),.Y(g22637),.A(g19363),.B(g19489));
  AND2 AND2_367(.VSS(VSS),.VDD(VDD),.Y(g17176),.A(g8616),.B(g13008));
  AND2 AND2_368(.VSS(VSS),.VDD(VDD),.Y(g34742),.A(g9000),.B(g34698));
  AND2 AND2_369(.VSS(VSS),.VDD(VDD),.Y(g28616),.A(g27532),.B(g20551));
  AND3 AND3_27(.VSS(VSS),.VDD(VDD),.Y(g34096),.A(g22957),.B(g9104),.C(g33772));
  AND2 AND2_370(.VSS(VSS),.VDD(VDD),.Y(g18654),.A(g4146),.B(g16249));
  AND2 AND2_371(.VSS(VSS),.VDD(VDD),.Y(g16203),.A(g5821),.B(g14297));
  AND2 AND2_372(.VSS(VSS),.VDD(VDD),.Y(g28313),.A(g27231),.B(g19766));
  AND2 AND2_373(.VSS(VSS),.VDD(VDD),.Y(g27116),.A(g26026),.B(g16527));
  AND4 AND4_18(.VSS(VSS),.VDD(VDD),.Y(I27509),.A(g24084),.B(g24085),.C(g24086),.D(g24087));
  AND2 AND2_374(.VSS(VSS),.VDD(VDD),.Y(g21823),.A(g3731),.B(g20453));
  AND2 AND2_375(.VSS(VSS),.VDD(VDD),.Y(g27615),.A(g26789),.B(g26770));
  AND2 AND2_376(.VSS(VSS),.VDD(VDD),.Y(g18800),.A(g6187),.B(g15348));
  AND2 AND2_377(.VSS(VSS),.VDD(VDD),.Y(g15859),.A(g3610),.B(g13923));
  AND4 AND4_19(.VSS(VSS),.VDD(VDD),.Y(I31181),.A(g29385),.B(g32716),.C(g32717),.D(g32718));
  AND2 AND2_378(.VSS(VSS),.VDD(VDD),.Y(g18417),.A(g2116),.B(g15373));
  AND2 AND2_379(.VSS(VSS),.VDD(VDD),.Y(g24556),.A(g4035),.B(g23341));
  AND2 AND2_380(.VSS(VSS),.VDD(VDD),.Y(g28285),.A(g9657),.B(g27717));
  AND2 AND2_381(.VSS(VSS),.VDD(VDD),.Y(g34681),.A(g34491),.B(g19438));
  AND4 AND4_20(.VSS(VSS),.VDD(VDD),.Y(I27508),.A(g19935),.B(g24082),.C(g24083),.D(g28033));
  AND2 AND2_382(.VSS(VSS),.VDD(VDD),.Y(g15858),.A(g3542),.B(g14045));
  AND2 AND2_383(.VSS(VSS),.VDD(VDD),.Y(g27041),.A(g8519),.B(g26330));
  AND2 AND2_384(.VSS(VSS),.VDD(VDD),.Y(g32126),.A(g31601),.B(g29948));
  AND2 AND2_385(.VSS(VSS),.VDD(VDD),.Y(g18334),.A(g1696),.B(g17873));
  AND2 AND2_386(.VSS(VSS),.VDD(VDD),.Y(g27275),.A(g25945),.B(g19745));
  AND2 AND2_387(.VSS(VSS),.VDD(VDD),.Y(g19756),.A(g9899),.B(g17154));
  AND2 AND2_388(.VSS(VSS),.VDD(VDD),.Y(g33927),.A(g33094),.B(g21412));
  AND3 AND3_28(.VSS(VSS),.VDD(VDD),.Y(g28254),.A(g7268),.B(g1668),.C(g27395));
  AND2 AND2_389(.VSS(VSS),.VDD(VDD),.Y(g27430),.A(g26488),.B(g17579));
  AND2 AND2_390(.VSS(VSS),.VDD(VDD),.Y(g34857),.A(g16540),.B(g34813));
  AND2 AND2_391(.VSS(VSS),.VDD(VDD),.Y(g10822),.A(g4264),.B(g8514));
  AND2 AND2_392(.VSS(VSS),.VDD(VDD),.Y(g24223),.A(g239),.B(g22594));
  AND2 AND2_393(.VSS(VSS),.VDD(VDD),.Y(g27493),.A(g246),.B(g26837));
  AND2 AND2_394(.VSS(VSS),.VDD(VDD),.Y(g16957),.A(g13064),.B(g10418));
  AND2 AND2_395(.VSS(VSS),.VDD(VDD),.Y(g25959),.A(g1648),.B(g24963));
  AND2 AND2_396(.VSS(VSS),.VDD(VDD),.Y(g30730),.A(g26346),.B(g29778));
  AND2 AND2_397(.VSS(VSS),.VDD(VDD),.Y(g25925),.A(g24990),.B(g23234));
  AND2 AND2_398(.VSS(VSS),.VDD(VDD),.Y(g28466),.A(g27960),.B(g17637));
  AND2 AND2_399(.VSS(VSS),.VDD(VDD),.Y(g25112),.A(g10428),.B(g23510));
  AND2 AND2_400(.VSS(VSS),.VDD(VDD),.Y(g21966),.A(g5406),.B(g21514));
  AND2 AND2_401(.VSS(VSS),.VDD(VDD),.Y(g18762),.A(g5475),.B(g17929));
  AND2 AND2_402(.VSS(VSS),.VDD(VDD),.Y(g25050),.A(g13056),.B(g22312));
  AND2 AND2_403(.VSS(VSS),.VDD(VDD),.Y(g20084),.A(g11591),.B(g16609));
  AND2 AND2_404(.VSS(VSS),.VDD(VDD),.Y(g32339),.A(g31474),.B(g20672));
  AND2 AND2_405(.VSS(VSS),.VDD(VDD),.Y(g31240),.A(g14793),.B(g30206));
  AND2 AND2_406(.VSS(VSS),.VDD(VDD),.Y(g19350),.A(g15968),.B(g13505));
  AND2 AND2_407(.VSS(VSS),.VDD(VDD),.Y(g34765),.A(g34692),.B(g20057));
  AND2 AND2_408(.VSS(VSS),.VDD(VDD),.Y(g27340),.A(g10199),.B(g26784));
  AND2 AND2_409(.VSS(VSS),.VDD(VDD),.Y(g27035),.A(g26348),.B(g1500));
  AND2 AND2_410(.VSS(VSS),.VDD(VDD),.Y(g18423),.A(g12851),.B(g18008));
  AND2 AND2_411(.VSS(VSS),.VDD(VDD),.Y(g29789),.A(g28270),.B(g10233));
  AND2 AND2_412(.VSS(VSS),.VDD(VDD),.Y(g32338),.A(g31466),.B(g20668));
  AND3 AND3_29(.VSS(VSS),.VDD(VDD),.Y(g33491),.A(g32679),.B(I31151),.C(I31152));
  AND2 AND2_413(.VSS(VSS),.VDD(VDD),.Y(g33903),.A(g33447),.B(g19146));
  AND2 AND2_414(.VSS(VSS),.VDD(VDD),.Y(g24922),.A(g4831),.B(g23931));
  AND2 AND2_415(.VSS(VSS),.VDD(VDD),.Y(g26129),.A(g2384),.B(g25121));
  AND2 AND2_416(.VSS(VSS),.VDD(VDD),.Y(g18216),.A(g967),.B(g15979));
  AND2 AND2_417(.VSS(VSS),.VDD(VDD),.Y(g24321),.A(g4558),.B(g22228));
  AND2 AND2_418(.VSS(VSS),.VDD(VDD),.Y(g16699),.A(g7134),.B(g12933));
  AND2 AND2_419(.VSS(VSS),.VDD(VDD),.Y(g27684),.A(g26386),.B(g20657));
  AND2 AND2_420(.VSS(VSS),.VDD(VDD),.Y(g28642),.A(g27555),.B(g20598));
  AND2 AND2_421(.VSS(VSS),.VDD(VDD),.Y(g18587),.A(g2980),.B(g16349));
  AND2 AND2_422(.VSS(VSS),.VDD(VDD),.Y(g25096),.A(g23778),.B(g20560));
  AND2 AND2_423(.VSS(VSS),.VDD(VDD),.Y(g29788),.A(g28335),.B(g23250));
  AND2 AND2_424(.VSS(VSS),.VDD(VDD),.Y(g26128),.A(g2319),.B(g25120));
  AND2 AND2_425(.VSS(VSS),.VDD(VDD),.Y(g14589),.A(g10586),.B(g10569));
  AND2 AND2_426(.VSS(VSS),.VDD(VDD),.Y(g29535),.A(g2303),.B(g28871));
  AND4 AND4_21(.VSS(VSS),.VDD(VDD),.Y(I31211),.A(g31021),.B(g31833),.C(g32759),.D(g32760));
  AND2 AND2_427(.VSS(VSS),.VDD(VDD),.Y(g27517),.A(g26400),.B(g17707));
  AND2 AND2_428(.VSS(VSS),.VDD(VDD),.Y(g10588),.A(g7004),.B(g5297));
  AND2 AND2_429(.VSS(VSS),.VDD(VDD),.Y(g18909),.A(g16226),.B(g13570));
  AND2 AND2_430(.VSS(VSS),.VDD(VDD),.Y(g32197),.A(g31144),.B(g20088));
  AND2 AND2_431(.VSS(VSS),.VDD(VDD),.Y(g18543),.A(g2779),.B(g15277));
  AND2 AND2_432(.VSS(VSS),.VDD(VDD),.Y(g26323),.A(g10262),.B(g25273));
  AND2 AND2_433(.VSS(VSS),.VDD(VDD),.Y(g24186),.A(g18102),.B(g22722));
  AND2 AND2_434(.VSS(VSS),.VDD(VDD),.Y(g14588),.A(g11957),.B(g11974));
  AND2 AND2_435(.VSS(VSS),.VDD(VDD),.Y(g24676),.A(g2748),.B(g23782));
  AND3 AND3_30(.VSS(VSS),.VDD(VDD),.Y(I16721),.A(g10224),.B(g12589),.C(g12525));
  AND2 AND2_436(.VSS(VSS),.VDD(VDD),.Y(g18117),.A(g464),.B(g17015));
  AND2 AND2_437(.VSS(VSS),.VDD(VDD),.Y(g16427),.A(g5216),.B(g14876));
  AND2 AND2_438(.VSS(VSS),.VDD(VDD),.Y(g25802),.A(g8106),.B(g24586));
  AND2 AND2_439(.VSS(VSS),.VDD(VDD),.Y(g22083),.A(g6287),.B(g19210));
  AND2 AND2_440(.VSS(VSS),.VDD(VDD),.Y(g32411),.A(g31119),.B(g13469));
  AND2 AND2_441(.VSS(VSS),.VDD(VDD),.Y(g23023),.A(g650),.B(g20248));
  AND2 AND2_442(.VSS(VSS),.VDD(VDD),.Y(g19691),.A(g9614),.B(g17085));
  AND2 AND2_443(.VSS(VSS),.VDD(VDD),.Y(g24654),.A(g11735),.B(g22922));
  AND2 AND2_444(.VSS(VSS),.VDD(VDD),.Y(g28630),.A(g27544),.B(g20575));
  AND2 AND2_445(.VSS(VSS),.VDD(VDD),.Y(g29344),.A(g29168),.B(g18932));
  AND2 AND2_446(.VSS(VSS),.VDD(VDD),.Y(g18569),.A(g94),.B(g16349));
  AND2 AND2_447(.VSS(VSS),.VDD(VDD),.Y(g30002),.A(g28481),.B(g23487));
  AND2 AND2_448(.VSS(VSS),.VDD(VDD),.Y(g27130),.A(g26026),.B(g16585));
  AND2 AND2_449(.VSS(VSS),.VDD(VDD),.Y(g30057),.A(g29144),.B(g9462));
  AND2 AND2_450(.VSS(VSS),.VDD(VDD),.Y(g22622),.A(g19336),.B(g19469));
  AND2 AND2_451(.VSS(VSS),.VDD(VDD),.Y(g18568),.A(g37),.B(g16349));
  AND2 AND2_452(.VSS(VSS),.VDD(VDD),.Y(g18747),.A(g5138),.B(g17847));
  AND2 AND2_453(.VSS(VSS),.VDD(VDD),.Y(g25765),.A(g24989),.B(g24973));
  AND2 AND2_454(.VSS(VSS),.VDD(VDD),.Y(g27362),.A(g26080),.B(g20036));
  AND2 AND2_455(.VSS(VSS),.VDD(VDD),.Y(g31990),.A(g31772),.B(g18945));
  AND2 AND2_456(.VSS(VSS),.VDD(VDD),.Y(g33899),.A(g32132),.B(g33335));
  AND2 AND2_457(.VSS(VSS),.VDD(VDD),.Y(g18242),.A(g962),.B(g16431));
  AND2 AND2_458(.VSS(VSS),.VDD(VDD),.Y(g10616),.A(g7998),.B(g174));
  AND2 AND2_459(.VSS(VSS),.VDD(VDD),.Y(g27523),.A(g26549),.B(g17718));
  AND2 AND2_460(.VSS(VSS),.VDD(VDD),.Y(g30245),.A(g28733),.B(g23935));
  AND4 AND4_22(.VSS(VSS),.VDD(VDD),.Y(I31126),.A(g30673),.B(g31818),.C(g32636),.D(g32637));
  AND2 AND2_461(.VSS(VSS),.VDD(VDD),.Y(g26232),.A(g2193),.B(g25396));
  AND2 AND2_462(.VSS(VSS),.VDD(VDD),.Y(g33898),.A(g33419),.B(g15655));
  AND2 AND2_463(.VSS(VSS),.VDD(VDD),.Y(g21816),.A(g3602),.B(g20924));
  AND2 AND2_464(.VSS(VSS),.VDD(VDD),.Y(g18123),.A(g479),.B(g16886));
  AND2 AND2_465(.VSS(VSS),.VDD(VDD),.Y(g18814),.A(g6519),.B(g15483));
  AND2 AND2_466(.VSS(VSS),.VDD(VDD),.Y(g33719),.A(g33141),.B(g19433));
  AND2 AND2_467(.VSS(VSS),.VDD(VDD),.Y(g24762),.A(g655),.B(g23573));
  AND3 AND3_31(.VSS(VSS),.VDD(VDD),.Y(g10704),.A(g2145),.B(g10200),.C(g2130));
  AND2 AND2_468(.VSS(VSS),.VDD(VDD),.Y(g34533),.A(g34318),.B(g19731));
  AND2 AND2_469(.VSS(VSS),.VDD(VDD),.Y(g18751),.A(g5156),.B(g17847));
  AND2 AND2_470(.VSS(VSS),.VDD(VDD),.Y(g18807),.A(g6386),.B(g15656));
  AND2 AND2_471(.VSS(VSS),.VDD(VDD),.Y(g21976),.A(g5527),.B(g19074));
  AND2 AND2_472(.VSS(VSS),.VDD(VDD),.Y(g21985),.A(g5571),.B(g19074));
  AND2 AND2_473(.VSS(VSS),.VDD(VDD),.Y(g15902),.A(g441),.B(g13975));
  AND2 AND2_474(.VSS(VSS),.VDD(VDD),.Y(g18772),.A(g5689),.B(g15615));
  AND2 AND2_475(.VSS(VSS),.VDD(VDD),.Y(g28555),.A(g27429),.B(g20373));
  AND2 AND2_476(.VSS(VSS),.VDD(VDD),.Y(g33718),.A(g33147),.B(g19432));
  AND2 AND2_477(.VSS(VSS),.VDD(VDD),.Y(g34298),.A(g8679),.B(g34132));
  AND2 AND2_478(.VSS(VSS),.VDD(VDD),.Y(g28454),.A(g26976),.B(g12233));
  AND3 AND3_32(.VSS(VSS),.VDD(VDD),.Y(g33521),.A(g32895),.B(I31301),.C(I31302));
  AND2 AND2_479(.VSS(VSS),.VDD(VDD),.Y(g18974),.A(g174),.B(g16127));
  AND4 AND4_23(.VSS(VSS),.VDD(VDD),.Y(g26261),.A(g24688),.B(g10678),.C(g8778),.D(g8757));
  AND2 AND2_480(.VSS(VSS),.VDD(VDD),.Y(g32315),.A(g31306),.B(g23517));
  AND2 AND2_481(.VSS(VSS),.VDD(VDD),.Y(g24423),.A(g4950),.B(g22897));
  AND2 AND2_482(.VSS(VSS),.VDD(VDD),.Y(g21752),.A(g3171),.B(g20785));
  AND4 AND4_24(.VSS(VSS),.VDD(VDD),.Y(g27727),.A(g22432),.B(g25211),.C(g26424),.D(g26195));
  AND4 AND4_25(.VSS(VSS),.VDD(VDD),.Y(I31296),.A(g30937),.B(g31848),.C(g32882),.D(g32883));
  AND2 AND2_483(.VSS(VSS),.VDD(VDD),.Y(g18639),.A(g3831),.B(g17096));
  AND2 AND2_484(.VSS(VSS),.VDD(VDD),.Y(g28570),.A(g27456),.B(g20434));
  AND2 AND2_485(.VSS(VSS),.VDD(VDD),.Y(g28712),.A(g27590),.B(g20708));
  AND2 AND2_486(.VSS(VSS),.VDD(VDD),.Y(g21954),.A(g5381),.B(g21514));
  AND2 AND2_487(.VSS(VSS),.VDD(VDD),.Y(g27222),.A(g26055),.B(g13932));
  AND2 AND2_488(.VSS(VSS),.VDD(VDD),.Y(g29760),.A(g28309),.B(g23227));
  AND2 AND2_489(.VSS(VSS),.VDD(VDD),.Y(g33832),.A(g33088),.B(g27991));
  AND2 AND2_490(.VSS(VSS),.VDD(VDD),.Y(g18230),.A(g1111),.B(g16326));
  AND4 AND4_26(.VSS(VSS),.VDD(VDD),.Y(g29029),.A(g14506),.B(g25227),.C(g26424),.D(g27494));
  AND2 AND2_491(.VSS(VSS),.VDD(VDD),.Y(g17139),.A(g8635),.B(g12967));
  AND2 AND2_492(.VSS(VSS),.VDD(VDD),.Y(g18293),.A(g1484),.B(g16449));
  AND4 AND4_27(.VSS(VSS),.VDD(VDD),.Y(g17653),.A(g11547),.B(g11592),.C(g6789),.D(I18620));
  AND2 AND2_493(.VSS(VSS),.VDD(VDD),.Y(g15738),.A(g1111),.B(g13260));
  AND2 AND2_494(.VSS(VSS),.VDD(VDD),.Y(g18638),.A(g3827),.B(g17096));
  AND2 AND2_495(.VSS(VSS),.VDD(VDD),.Y(g27437),.A(g26576),.B(g17589));
  AND2 AND2_496(.VSS(VSS),.VDD(VDD),.Y(g33440),.A(g32250),.B(g29719));
  AND2 AND2_497(.VSS(VSS),.VDD(VDD),.Y(g32055),.A(g10999),.B(g30825));
  AND2 AND2_498(.VSS(VSS),.VDD(VDD),.Y(g17138),.A(g255),.B(g13239));
  AND2 AND2_499(.VSS(VSS),.VDD(VDD),.Y(g18265),.A(g1270),.B(g16000));
  AND2 AND2_500(.VSS(VSS),.VDD(VDD),.Y(g25129),.A(g17682),.B(g23527));
  AND2 AND2_501(.VSS(VSS),.VDD(VDD),.Y(g15699),.A(g1437),.B(g13861));
  AND2 AND2_502(.VSS(VSS),.VDD(VDD),.Y(g30232),.A(g28719),.B(g23912));
  AND2 AND2_503(.VSS(VSS),.VDD(VDD),.Y(g32111),.A(g31616),.B(g29922));
  AND2 AND2_504(.VSS(VSS),.VDD(VDD),.Y(g18416),.A(g2112),.B(g15373));
  AND2 AND2_505(.VSS(VSS),.VDD(VDD),.Y(g25057),.A(g23275),.B(g20511));
  AND2 AND2_506(.VSS(VSS),.VDD(VDD),.Y(g32070),.A(g10967),.B(g30825));
  AND2 AND2_507(.VSS(VSS),.VDD(VDD),.Y(g33861),.A(g33271),.B(g20502));
  AND2 AND2_508(.VSS(VSS),.VDD(VDD),.Y(g28239),.A(g27135),.B(g19659));
  AND2 AND2_509(.VSS(VSS),.VDD(VDD),.Y(g25128),.A(g17418),.B(g23525));
  AND2 AND2_510(.VSS(VSS),.VDD(VDD),.Y(g17636),.A(g10829),.B(g13463));
  AND2 AND2_511(.VSS(VSS),.VDD(VDD),.Y(g11916),.A(g2227),.B(g7328));
  AND2 AND2_512(.VSS(VSS),.VDD(VDD),.Y(g33247),.A(g32130),.B(g19980));
  AND2 AND2_513(.VSS(VSS),.VDD(VDD),.Y(g28567),.A(g6832),.B(g27101));
  AND4 AND4_28(.VSS(VSS),.VDD(VDD),.Y(I31197),.A(g32740),.B(g32741),.C(g32742),.D(g32743));
  AND2 AND2_514(.VSS(VSS),.VDD(VDD),.Y(g27347),.A(g26400),.B(g17390));
  AND2 AND2_515(.VSS(VSS),.VDD(VDD),.Y(g18992),.A(g8341),.B(g16171));
  AND2 AND2_516(.VSS(VSS),.VDD(VDD),.Y(g18391),.A(g1982),.B(g15171));
  AND3 AND3_33(.VSS(VSS),.VDD(VDD),.Y(g24908),.A(g3752),.B(g23239),.C(I24075));
  AND2 AND2_517(.VSS(VSS),.VDD(VDD),.Y(g28238),.A(g27133),.B(g19658));
  AND2 AND2_518(.VSS(VSS),.VDD(VDD),.Y(g21842),.A(g3863),.B(g21070));
  AND2 AND2_519(.VSS(VSS),.VDD(VDD),.Y(g18510),.A(g2625),.B(g15509));
  AND2 AND2_520(.VSS(VSS),.VDD(VDD),.Y(g30261),.A(g28772),.B(g23961));
  AND2 AND2_521(.VSS(VSS),.VDD(VDD),.Y(g23392),.A(g7247),.B(g21430));
  AND2 AND2_522(.VSS(VSS),.VDD(VDD),.Y(g24569),.A(g5115),.B(g23382));
  AND2 AND2_523(.VSS(VSS),.VDD(VDD),.Y(g25323),.A(g6888),.B(g22359));
  AND2 AND2_524(.VSS(VSS),.VDD(VDD),.Y(g31324),.A(g30171),.B(g27937));
  AND2 AND2_525(.VSS(VSS),.VDD(VDD),.Y(g33099),.A(g32395),.B(g18944));
  AND2 AND2_526(.VSS(VSS),.VDD(VDD),.Y(g13287),.A(g1221),.B(g11472));
  AND2 AND2_527(.VSS(VSS),.VDD(VDD),.Y(g27600),.A(g26755),.B(g26725));
  AND4 AND4_29(.VSS(VSS),.VDD(VDD),.Y(g10733),.A(g3639),.B(g6905),.C(g3625),.D(g8542));
  AND2 AND2_528(.VSS(VSS),.VDD(VDD),.Y(g18579),.A(g2984),.B(g16349));
  AND2 AND2_529(.VSS(VSS),.VDD(VDD),.Y(g31777),.A(g21343),.B(g29385));
  AND2 AND2_530(.VSS(VSS),.VDD(VDD),.Y(g33701),.A(g33162),.B(g16305));
  AND2 AND2_531(.VSS(VSS),.VDD(VDD),.Y(g24747),.A(g17510),.B(g22417));
  AND2 AND2_532(.VSS(VSS),.VDD(VDD),.Y(g32067),.A(g4727),.B(g30614));
  AND2 AND2_533(.VSS(VSS),.VDD(VDD),.Y(g21559),.A(g16236),.B(g10897));
  AND2 AND2_534(.VSS(VSS),.VDD(VDD),.Y(g31272),.A(g30117),.B(g27742));
  AND3 AND3_34(.VSS(VSS),.VDD(VDD),.Y(I16618),.A(g10124),.B(g12341),.C(g12293));
  AND2 AND2_535(.VSS(VSS),.VDD(VDD),.Y(g15632),.A(g3494),.B(g13555));
  AND2 AND2_536(.VSS(VSS),.VDD(VDD),.Y(g28185),.A(g27026),.B(g19435));
  AND3 AND3_35(.VSS(VSS),.VDD(VDD),.Y(g10874),.A(g7791),.B(g6219),.C(g6227));
  AND2 AND2_537(.VSS(VSS),.VDD(VDD),.Y(g18578),.A(g2873),.B(g16349));
  AND2 AND2_538(.VSS(VSS),.VDD(VDD),.Y(g25775),.A(g2922),.B(g24568));
  AND2 AND2_539(.VSS(VSS),.VDD(VDD),.Y(g23424),.A(g7345),.B(g21556));
  AND2 AND2_540(.VSS(VSS),.VDD(VDD),.Y(g27351),.A(g10218),.B(g26804));
  AND2 AND2_541(.VSS(VSS),.VDD(VDD),.Y(g27372),.A(g26488),.B(g17476));
  AND2 AND2_542(.VSS(VSS),.VDD(VDD),.Y(g19768),.A(g2803),.B(g15833));
  AND2 AND2_543(.VSS(VSS),.VDD(VDD),.Y(g14874),.A(g1099),.B(g10909));
  AND2 AND2_544(.VSS(VSS),.VDD(VDD),.Y(g16671),.A(g6275),.B(g14817));
  AND2 AND2_545(.VSS(VSS),.VDD(VDD),.Y(g21558),.A(g15904),.B(g13729));
  AND2 AND2_546(.VSS(VSS),.VDD(VDD),.Y(g27821),.A(g7680),.B(g25892));
  AND2 AND2_547(.VSS(VSS),.VDD(VDD),.Y(g32150),.A(g31624),.B(g29995));
  AND2 AND2_548(.VSS(VSS),.VDD(VDD),.Y(g28154),.A(g8492),.B(g27306));
  AND2 AND2_549(.VSS(VSS),.VDD(VDD),.Y(g18586),.A(g2886),.B(g16349));
  AND2 AND2_550(.VSS(VSS),.VDD(VDD),.Y(g29649),.A(g2241),.B(g28678));
  AND3 AND3_36(.VSS(VSS),.VDD(VDD),.Y(g33462),.A(g32470),.B(I31006),.C(I31007));
  AND2 AND2_551(.VSS(VSS),.VDD(VDD),.Y(g21830),.A(g3774),.B(g20453));
  AND2 AND2_552(.VSS(VSS),.VDD(VDD),.Y(g26611),.A(g24935),.B(g20580));
  AND2 AND2_553(.VSS(VSS),.VDD(VDD),.Y(g20751),.A(g16260),.B(g4836));
  AND2 AND2_554(.VSS(VSS),.VDD(VDD),.Y(g10665),.A(g209),.B(g8292));
  AND2 AND2_555(.VSS(VSS),.VDD(VDD),.Y(g28637),.A(g22399),.B(g27011));
  AND2 AND2_556(.VSS(VSS),.VDD(VDD),.Y(g18442),.A(g2259),.B(g18008));
  AND2 AND2_557(.VSS(VSS),.VDD(VDD),.Y(g32019),.A(g30579),.B(g22358));
  AND2 AND2_558(.VSS(VSS),.VDD(VDD),.Y(g24772),.A(g16287),.B(g23061));
  AND2 AND2_559(.VSS(VSS),.VDD(VDD),.Y(g29648),.A(g2112),.B(g29121));
  AND2 AND2_560(.VSS(VSS),.VDD(VDD),.Y(g27264),.A(g25941),.B(g19714));
  AND2 AND2_561(.VSS(VSS),.VDD(VDD),.Y(g22115),.A(g6573),.B(g19277));
  AND2 AND2_562(.VSS(VSS),.VDD(VDD),.Y(g27137),.A(g26026),.B(g16606));
  AND2 AND2_563(.VSS(VSS),.VDD(VDD),.Y(g21865),.A(g3965),.B(g21070));
  AND2 AND2_564(.VSS(VSS),.VDD(VDD),.Y(g31140),.A(g2102),.B(g30037));
  AND2 AND2_565(.VSS(VSS),.VDD(VDD),.Y(g32196),.A(g27587),.B(g31376));
  AND2 AND2_566(.VSS(VSS),.VDD(VDD),.Y(g13942),.A(g5897),.B(g12512));
  AND2 AND2_567(.VSS(VSS),.VDD(VDD),.Y(g24639),.A(g6181),.B(g23699));
  AND2 AND2_568(.VSS(VSS),.VDD(VDD),.Y(g32018),.A(g4146),.B(g30937));
  AND2 AND2_569(.VSS(VSS),.VDD(VDD),.Y(g26271),.A(g1992),.B(g25341));
  AND2 AND2_570(.VSS(VSS),.VDD(VDD),.Y(g29604),.A(g2315),.B(g28966));
  AND3 AND3_37(.VSS(VSS),.VDD(VDD),.Y(g30316),.A(g29199),.B(g7097),.C(g6682));
  AND2 AND2_571(.VSS(VSS),.VDD(VDD),.Y(g21713),.A(g298),.B(g20283));
  AND2 AND2_572(.VSS(VSS),.VDD(VDD),.Y(g34499),.A(g31288),.B(g34339));
  AND2 AND2_573(.VSS(VSS),.VDD(VDD),.Y(g24230),.A(g901),.B(g22594));
  AND3 AND3_38(.VSS(VSS),.VDD(VDD),.Y(g13156),.A(g10816),.B(g10812),.C(g10805));
  AND2 AND2_574(.VSS(VSS),.VDD(VDD),.Y(g18116),.A(g168),.B(g17015));
  AND2 AND2_575(.VSS(VSS),.VDD(VDD),.Y(g24293),.A(g4438),.B(g22550));
  AND2 AND2_576(.VSS(VSS),.VDD(VDD),.Y(g18615),.A(g3347),.B(g17200));
  AND2 AND2_577(.VSS(VSS),.VDD(VDD),.Y(g22052),.A(g6113),.B(g21611));
  AND3 AND3_39(.VSS(VSS),.VDD(VDD),.Y(g10476),.A(g7244),.B(g7259),.C(I13862));
  AND2 AND2_578(.VSS(VSS),.VDD(VDD),.Y(g24638),.A(g22763),.B(g19690));
  AND2 AND2_579(.VSS(VSS),.VDD(VDD),.Y(g29770),.A(g28320),.B(g23238));
  AND2 AND2_580(.VSS(VSS),.VDD(VDD),.Y(g16190),.A(g14626),.B(g11810));
  AND2 AND2_581(.VSS(VSS),.VDD(VDD),.Y(g29563),.A(g1616),.B(g28853));
  AND4 AND4_30(.VSS(VSS),.VDD(VDD),.Y(I31202),.A(g32747),.B(g32748),.C(g32749),.D(g32750));
  AND2 AND2_582(.VSS(VSS),.VDD(VDD),.Y(g34498),.A(g13888),.B(g34336));
  AND2 AND2_583(.VSS(VSS),.VDD(VDD),.Y(g18720),.A(g15137),.B(g16795));
  AND2 AND2_584(.VSS(VSS),.VDD(VDD),.Y(g26753),.A(g16024),.B(g24452));
  AND4 AND4_31(.VSS(VSS),.VDD(VDD),.Y(I31257),.A(g32826),.B(g32827),.C(g32828),.D(g32829));
  AND2 AND2_585(.VSS(VSS),.VDD(VDD),.Y(g25880),.A(g8443),.B(g24814));
  AND4 AND4_32(.VSS(VSS),.VDD(VDD),.Y(g14555),.A(g12521),.B(g12356),.C(g12307),.D(I16671));
  AND2 AND2_586(.VSS(VSS),.VDD(VDD),.Y(g24416),.A(g4939),.B(g22870));
  AND2 AND2_587(.VSS(VSS),.VDD(VDD),.Y(g16520),.A(g5909),.B(g14965));
  AND2 AND2_588(.VSS(VSS),.VDD(VDD),.Y(g21705),.A(g209),.B(g20283));
  AND2 AND2_589(.VSS(VSS),.VDD(VDD),.Y(g30056),.A(g29165),.B(g12659));
  AND2 AND2_590(.VSS(VSS),.VDD(VDD),.Y(g18275),.A(g15070),.B(g16136));
  AND2 AND2_591(.VSS(VSS),.VDD(VDD),.Y(g26145),.A(g11962),.B(g25131));
  AND4 AND4_33(.VSS(VSS),.VDD(VDD),.Y(I31111),.A(g31070),.B(g31815),.C(g32615),.D(g32616));
  AND2 AND2_592(.VSS(VSS),.VDD(VDD),.Y(g18430),.A(g2204),.B(g18008));
  AND2 AND2_593(.VSS(VSS),.VDD(VDD),.Y(g18746),.A(g5134),.B(g17847));
  AND3 AND3_40(.VSS(VSS),.VDD(VDD),.Y(g27209),.A(g26213),.B(g8365),.C(g2051));
  AND2 AND2_594(.VSS(VSS),.VDD(VDD),.Y(g32402),.A(g4888),.B(g30990));
  AND2 AND2_595(.VSS(VSS),.VDD(VDD),.Y(g18493),.A(g2514),.B(g15426));
  AND2 AND2_596(.VSS(VSS),.VDD(VDD),.Y(g33871),.A(g33281),.B(g20546));
  AND2 AND2_597(.VSS(VSS),.VDD(VDD),.Y(g30080),.A(g28121),.B(g20674));
  AND2 AND2_598(.VSS(VSS),.VDD(VDD),.Y(g28215),.A(g9264),.B(g27565));
  AND2 AND2_599(.VSS(VSS),.VDD(VDD),.Y(g26650),.A(g10796),.B(g24424));
  AND3 AND3_41(.VSS(VSS),.VDD(VDD),.Y(g34080),.A(g22957),.B(g9104),.C(g33750));
  AND2 AND2_600(.VSS(VSS),.VDD(VDD),.Y(g16211),.A(g5445),.B(g14215));
  AND2 AND2_601(.VSS(VSS),.VDD(VDD),.Y(g27208),.A(g9037),.B(g26598));
  AND2 AND2_602(.VSS(VSS),.VDD(VDD),.Y(g18465),.A(g2384),.B(g15224));
  AND2 AND2_603(.VSS(VSS),.VDD(VDD),.Y(g29767),.A(g28317),.B(g23236));
  AND2 AND2_604(.VSS(VSS),.VDD(VDD),.Y(g29794),.A(g28342),.B(g23256));
  AND2 AND2_605(.VSS(VSS),.VDD(VDD),.Y(g21188),.A(g7666),.B(g15705));
  AND2 AND2_606(.VSS(VSS),.VDD(VDD),.Y(g33360),.A(g32253),.B(g20869));
  AND2 AND2_607(.VSS(VSS),.VDD(VDD),.Y(g18237),.A(g1146),.B(g16326));
  AND2 AND2_608(.VSS(VSS),.VDD(VDD),.Y(g29845),.A(g28375),.B(g23291));
  AND2 AND2_609(.VSS(VSS),.VDD(VDD),.Y(g23188),.A(g13994),.B(g20025));
  AND3 AND3_42(.VSS(VSS),.VDD(VDD),.Y(I16143),.A(g8751),.B(g11491),.C(g11445));
  AND2 AND2_610(.VSS(VSS),.VDD(VDD),.Y(g28439),.A(g27273),.B(g10233));
  AND2 AND2_611(.VSS(VSS),.VDD(VDD),.Y(g18340),.A(g1720),.B(g17873));
  AND2 AND2_612(.VSS(VSS),.VDD(VDD),.Y(g29899),.A(g28428),.B(g23375));
  AND2 AND2_613(.VSS(VSS),.VDD(VDD),.Y(g29990),.A(g29007),.B(g9239));
  AND2 AND2_614(.VSS(VSS),.VDD(VDD),.Y(g21939),.A(g5224),.B(g18997));
  AND2 AND2_615(.VSS(VSS),.VDD(VDD),.Y(g25831),.A(g3151),.B(g24623));
  AND2 AND2_616(.VSS(VSS),.VDD(VDD),.Y(g15784),.A(g3235),.B(g13977));
  AND2 AND2_617(.VSS(VSS),.VDD(VDD),.Y(g18806),.A(g6381),.B(g15656));
  AND2 AND2_618(.VSS(VSS),.VDD(VDD),.Y(g18684),.A(g4681),.B(g15885));
  AND2 AND2_619(.VSS(VSS),.VDD(VDD),.Y(g26393),.A(g19467),.B(g25558));
  AND2 AND2_620(.VSS(VSS),.VDD(VDD),.Y(g14567),.A(g10568),.B(g10552));
  AND2 AND2_621(.VSS(VSS),.VDD(VDD),.Y(g24835),.A(g8720),.B(g23233));
  AND2 AND2_622(.VSS(VSS),.VDD(VDD),.Y(g29633),.A(g1978),.B(g29085));
  AND4 AND4_34(.VSS(VSS),.VDD(VDD),.Y(I31067),.A(g32552),.B(g32553),.C(g32554),.D(g32555));
  AND2 AND2_623(.VSS(VSS),.VDD(VDD),.Y(g24014),.A(g7933),.B(g19063));
  AND2 AND2_624(.VSS(VSS),.VDD(VDD),.Y(g15103),.A(g4180),.B(g14454));
  AND2 AND2_625(.VSS(VSS),.VDD(VDD),.Y(g34753),.A(g34676),.B(g19586));
  AND2 AND2_626(.VSS(VSS),.VDD(VDD),.Y(g21938),.A(g5216),.B(g18997));
  AND2 AND2_627(.VSS(VSS),.VDD(VDD),.Y(g18142),.A(g577),.B(g17533));
  AND2 AND2_628(.VSS(VSS),.VDD(VDD),.Y(g34342),.A(g34103),.B(g19998));
  AND2 AND2_629(.VSS(VSS),.VDD(VDD),.Y(g30145),.A(g28603),.B(g21247));
  AND2 AND2_630(.VSS(VSS),.VDD(VDD),.Y(g30031),.A(g29071),.B(g10540));
  AND2 AND2_631(.VSS(VSS),.VDD(VDD),.Y(g27614),.A(g26785),.B(g26759));
  AND2 AND2_632(.VSS(VSS),.VDD(VDD),.Y(g32256),.A(g31249),.B(g20382));
  AND2 AND2_633(.VSS(VSS),.VDD(VDD),.Y(g18517),.A(g2652),.B(g15509));
  AND2 AND2_634(.VSS(VSS),.VDD(VDD),.Y(g27436),.A(g26576),.B(g17588));
  AND2 AND2_635(.VSS(VSS),.VDD(VDD),.Y(g30199),.A(g28664),.B(g23861));
  AND2 AND2_636(.VSS(VSS),.VDD(VDD),.Y(g29718),.A(g28512),.B(g11136));
  AND2 AND2_637(.VSS(VSS),.VDD(VDD),.Y(g29521),.A(g1744),.B(g28824));
  AND2 AND2_638(.VSS(VSS),.VDD(VDD),.Y(g16700),.A(g5208),.B(g14838));
  AND2 AND2_639(.VSS(VSS),.VDD(VDD),.Y(g31220),.A(g30273),.B(g25202));
  AND3 AND3_43(.VSS(VSS),.VDD(VDD),.Y(g33472),.A(g32542),.B(I31056),.C(I31057));
  AND2 AND2_640(.VSS(VSS),.VDD(VDD),.Y(g16126),.A(g5495),.B(g14262));
  AND2 AND2_641(.VSS(VSS),.VDD(VDD),.Y(g28284),.A(g11398),.B(g27994));
  AND2 AND2_642(.VSS(VSS),.VDD(VDD),.Y(g10675),.A(g3436),.B(g8500));
  AND2 AND2_643(.VSS(VSS),.VDD(VDD),.Y(g25989),.A(g25258),.B(g21012));
  AND4 AND4_35(.VSS(VSS),.VDD(VDD),.Y(g27073),.A(g7121),.B(g3873),.C(g3881),.D(g26281));
  AND2 AND2_644(.VSS(VSS),.VDD(VDD),.Y(g30198),.A(g28662),.B(g23860));
  AND2 AND2_645(.VSS(VSS),.VDD(VDD),.Y(g32300),.A(g31274),.B(g20544));
  AND2 AND2_646(.VSS(VSS),.VDD(VDD),.Y(g14185),.A(g8686),.B(g11744));
  AND2 AND2_647(.VSS(VSS),.VDD(VDD),.Y(g25056),.A(g12779),.B(g23456));
  AND2 AND2_648(.VSS(VSS),.VDD(VDD),.Y(g28304),.A(g27226),.B(g19753));
  AND2 AND2_649(.VSS(VSS),.VDD(VDD),.Y(g33911),.A(g33137),.B(g10725));
  AND2 AND2_650(.VSS(VSS),.VDD(VDD),.Y(g34198),.A(g33688),.B(g24491));
  AND2 AND2_651(.VSS(VSS),.VDD(VDD),.Y(g26161),.A(g2518),.B(g25139));
  AND2 AND2_652(.VSS(VSS),.VDD(VDD),.Y(g34529),.A(g34306),.B(g19634));
  AND2 AND2_653(.VSS(VSS),.VDD(VDD),.Y(g21875),.A(g4116),.B(g19801));
  AND2 AND2_654(.VSS(VSS),.VDD(VDD),.Y(g25988),.A(g9510),.B(g25016));
  AND4 AND4_36(.VSS(VSS),.VDD(VDD),.Y(I31196),.A(g30825),.B(g31830),.C(g32738),.D(g32739));
  AND2 AND2_655(.VSS(VSS),.VDD(VDD),.Y(g25924),.A(g24976),.B(g16846));
  AND2 AND2_656(.VSS(VSS),.VDD(VDD),.Y(g27346),.A(g26400),.B(g17389));
  AND2 AND2_657(.VSS(VSS),.VDD(VDD),.Y(g34528),.A(g34305),.B(g19617));
  AND2 AND2_658(.VSS(VSS),.VDD(VDD),.Y(g17692),.A(g1124),.B(g13307));
  AND2 AND2_659(.VSS(VSS),.VDD(VDD),.Y(g18130),.A(g528),.B(g16971));
  AND2 AND2_660(.VSS(VSS),.VDD(VDD),.Y(g34696),.A(g34531),.B(g20004));
  AND2 AND2_661(.VSS(VSS),.VDD(VDD),.Y(g18193),.A(g837),.B(g17821));
  AND2 AND2_662(.VSS(VSS),.VDD(VDD),.Y(g22013),.A(g5802),.B(g21562));
  AND2 AND2_663(.VSS(VSS),.VDD(VDD),.Y(g32157),.A(g31646),.B(g30021));
  AND2 AND2_664(.VSS(VSS),.VDD(VDD),.Y(g34393),.A(g34189),.B(g21304));
  AND2 AND2_665(.VSS(VSS),.VDD(VDD),.Y(g26259),.A(g24430),.B(g25232));
  AND3 AND3_44(.VSS(VSS),.VDD(VDD),.Y(I24508),.A(g9434),.B(g9672),.C(g5401));
  AND2 AND2_666(.VSS(VSS),.VDD(VDD),.Y(g18362),.A(g1834),.B(g17955));
  AND2 AND2_667(.VSS(VSS),.VDD(VDD),.Y(g23218),.A(g20200),.B(g16530));
  AND2 AND2_668(.VSS(VSS),.VDD(VDD),.Y(g29861),.A(g28390),.B(g23313));
  AND2 AND2_669(.VSS(VSS),.VDD(VDD),.Y(g29573),.A(g1752),.B(g28892));
  AND2 AND2_670(.VSS(VSS),.VDD(VDD),.Y(g33071),.A(g31591),.B(g32404));
  AND2 AND2_671(.VSS(VSS),.VDD(VDD),.Y(g21837),.A(g3719),.B(g20453));
  AND2 AND2_672(.VSS(VSS),.VDD(VDD),.Y(g34764),.A(g34691),.B(g20009));
  AND2 AND2_673(.VSS(VSS),.VDD(VDD),.Y(g22329),.A(g11940),.B(g20329));
  AND2 AND2_674(.VSS(VSS),.VDD(VDD),.Y(g10883),.A(g3355),.B(g9061));
  AND2 AND2_675(.VSS(VSS),.VDD(VDD),.Y(g18165),.A(g650),.B(g17433));
  AND2 AND2_676(.VSS(VSS),.VDD(VDD),.Y(g23837),.A(g21160),.B(g10804));
  AND2 AND2_677(.VSS(VSS),.VDD(VDD),.Y(g18523),.A(g2675),.B(g15509));
  AND2 AND2_678(.VSS(VSS),.VDD(VDD),.Y(g26087),.A(g5475),.B(g25072));
  AND2 AND2_679(.VSS(VSS),.VDD(VDD),.Y(g27034),.A(g26328),.B(g8609));
  AND2 AND2_680(.VSS(VSS),.VDD(VDD),.Y(g13306),.A(g441),.B(g11048));
  AND2 AND2_681(.VSS(VSS),.VDD(VDD),.Y(g31776),.A(g21329),.B(g29385));
  AND2 AND2_682(.VSS(VSS),.VDD(VDD),.Y(g34365),.A(g34149),.B(g20451));
  AND2 AND2_683(.VSS(VSS),.VDD(VDD),.Y(g26258),.A(g12875),.B(g25231));
  AND2 AND2_684(.VSS(VSS),.VDD(VDD),.Y(g19651),.A(g1111),.B(g16119));
  AND2 AND2_685(.VSS(VSS),.VDD(VDD),.Y(g33785),.A(g33100),.B(g20550));
  AND2 AND2_686(.VSS(VSS),.VDD(VDD),.Y(g29926),.A(g1604),.B(g28736));
  AND2 AND2_687(.VSS(VSS),.VDD(VDD),.Y(g34869),.A(g34816),.B(g19869));
  AND2 AND2_688(.VSS(VSS),.VDD(VDD),.Y(g28139),.A(g27337),.B(g26054));
  AND2 AND2_689(.VSS(VSS),.VDD(VDD),.Y(g22005),.A(g5759),.B(g21562));
  AND2 AND2_690(.VSS(VSS),.VDD(VDD),.Y(g31147),.A(g12286),.B(g30054));
  AND2 AND2_691(.VSS(VSS),.VDD(VDD),.Y(g28653),.A(g7544),.B(g27014));
  AND2 AND2_692(.VSS(VSS),.VDD(VDD),.Y(g13038),.A(g8509),.B(g11034));
  AND2 AND2_693(.VSS(VSS),.VDD(VDD),.Y(g27292),.A(g1714),.B(g26654));
  AND2 AND2_694(.VSS(VSS),.VDD(VDD),.Y(g29612),.A(g27875),.B(g28633));
  AND2 AND2_695(.VSS(VSS),.VDD(VDD),.Y(g24465),.A(g3827),.B(g23139));
  AND3 AND3_45(.VSS(VSS),.VDD(VDD),.Y(g12641),.A(g10295),.B(g3171),.C(g3179));
  AND2 AND2_696(.VSS(VSS),.VDD(VDD),.Y(g22538),.A(g14035),.B(g20248));
  AND2 AND2_697(.VSS(VSS),.VDD(VDD),.Y(g27153),.A(g26055),.B(g16629));
  AND2 AND2_698(.VSS(VSS),.VDD(VDD),.Y(g33355),.A(g32243),.B(g20769));
  AND2 AND2_699(.VSS(VSS),.VDD(VDD),.Y(g29324),.A(g29078),.B(g18883));
  AND2 AND2_700(.VSS(VSS),.VDD(VDD),.Y(g34868),.A(g34813),.B(g19866));
  AND2 AND2_701(.VSS(VSS),.VDD(VDD),.Y(g7396),.A(g392),.B(g441));
  AND2 AND2_702(.VSS(VSS),.VDD(VDD),.Y(g25031),.A(g20675),.B(g23432));
  AND2 AND2_703(.VSS(VSS),.VDD(VDD),.Y(g30161),.A(g28614),.B(g21275));
  AND2 AND2_704(.VSS(VSS),.VDD(VDD),.Y(g18475),.A(g12853),.B(g15426));
  AND2 AND2_705(.VSS(VSS),.VDD(VDD),.Y(g33859),.A(g33426),.B(g10531));
  AND4 AND4_37(.VSS(VSS),.VDD(VDD),.Y(g26244),.A(g24688),.B(g8812),.C(g10658),.D(g8757));
  AND2 AND2_706(.VSS(VSS),.VDD(VDD),.Y(g29534),.A(g28965),.B(g22457));
  AND2 AND2_707(.VSS(VSS),.VDD(VDD),.Y(g33370),.A(g32279),.B(g21139));
  AND2 AND2_708(.VSS(VSS),.VDD(VDD),.Y(g24983),.A(g23217),.B(g20238));
  AND2 AND2_709(.VSS(VSS),.VDD(VDD),.Y(g27409),.A(g26519),.B(g17524));
  AND2 AND2_710(.VSS(VSS),.VDD(VDD),.Y(g16855),.A(g4392),.B(g13107));
  AND2 AND2_711(.VSS(VSS),.VDD(VDD),.Y(g18727),.A(g4931),.B(g16077));
  AND2 AND2_712(.VSS(VSS),.VDD(VDD),.Y(g28415),.A(g27250),.B(g19963));
  AND2 AND2_713(.VSS(VSS),.VDD(VDD),.Y(g24684),.A(g11769),.B(g22989));
  AND2 AND2_714(.VSS(VSS),.VDD(VDD),.Y(g28333),.A(g27239),.B(g19787));
  AND2 AND2_715(.VSS(VSS),.VDD(VDD),.Y(g33858),.A(g33268),.B(g20448));
  AND2 AND2_716(.VSS(VSS),.VDD(VDD),.Y(g34709),.A(g34549),.B(g17242));
  AND2 AND2_717(.VSS(VSS),.VDD(VDD),.Y(g18222),.A(g1024),.B(g16100));
  AND2 AND2_718(.VSS(VSS),.VDD(VDD),.Y(g10501),.A(g1233),.B(g9007));
  AND2 AND2_719(.VSS(VSS),.VDD(VDD),.Y(g16870),.A(g6625),.B(g14905));
  AND2 AND2_720(.VSS(VSS),.VDD(VDD),.Y(g27136),.A(g26026),.B(g16605));
  AND2 AND2_721(.VSS(VSS),.VDD(VDD),.Y(g27408),.A(g26519),.B(g17523));
  AND4 AND4_38(.VSS(VSS),.VDD(VDD),.Y(g27635),.A(g23032),.B(g26281),.C(g26424),.D(g24996));
  AND2 AND2_722(.VSS(VSS),.VDD(VDD),.Y(g21915),.A(g5080),.B(g21468));
  AND2 AND2_723(.VSS(VSS),.VDD(VDD),.Y(g30225),.A(g28705),.B(g23897));
  AND2 AND2_724(.VSS(VSS),.VDD(VDD),.Y(g31151),.A(g10037),.B(g30065));
  AND2 AND2_725(.VSS(VSS),.VDD(VDD),.Y(g18437),.A(g2241),.B(g18008));
  AND2 AND2_726(.VSS(VSS),.VDD(VDD),.Y(g24142),.A(g17700),.B(g21657));
  AND4 AND4_39(.VSS(VSS),.VDD(VDD),.Y(I31001),.A(g29385),.B(g32456),.C(g32457),.D(g32458));
  AND2 AND2_727(.VSS(VSS),.VDD(VDD),.Y(g31996),.A(g31779),.B(g18979));
  AND2 AND2_728(.VSS(VSS),.VDD(VDD),.Y(g34225),.A(g33744),.B(g22942));
  AND4 AND4_40(.VSS(VSS),.VDD(VDD),.Y(I31077),.A(g32566),.B(g32567),.C(g32568),.D(g32569));
  AND2 AND2_729(.VSS(VSS),.VDD(VDD),.Y(g26602),.A(g7487),.B(g24453));
  AND2 AND2_730(.VSS(VSS),.VDD(VDD),.Y(g30258),.A(g28751),.B(g23953));
  AND2 AND2_731(.VSS(VSS),.VDD(VDD),.Y(g11937),.A(g1936),.B(g7362));
  AND2 AND2_732(.VSS(VSS),.VDD(VDD),.Y(g15860),.A(g3889),.B(g14160));
  AND3 AND3_46(.VSS(VSS),.VDD(VDD),.Y(g34087),.A(g33766),.B(g9104),.C(g18957));
  AND2 AND2_733(.VSS(VSS),.VDD(VDD),.Y(g23201),.A(g14027),.B(g20040));
  AND2 AND2_734(.VSS(VSS),.VDD(VDD),.Y(g33844),.A(g33257),.B(g20327));
  AND2 AND2_735(.VSS(VSS),.VDD(VDD),.Y(g33367),.A(g32271),.B(g21053));
  AND4 AND4_41(.VSS(VSS),.VDD(VDD),.Y(I31256),.A(g31021),.B(g31841),.C(g32824),.D(g32825));
  AND2 AND2_736(.VSS(VSS),.VDD(VDD),.Y(g18703),.A(g4776),.B(g16782));
  AND2 AND2_737(.VSS(VSS),.VDD(VDD),.Y(g22100),.A(g6466),.B(g18833));
  AND2 AND2_738(.VSS(VSS),.VDD(VDD),.Y(g18347),.A(g1756),.B(g17955));
  AND2 AND2_739(.VSS(VSS),.VDD(VDD),.Y(g19717),.A(g6527),.B(g17122));
  AND2 AND2_740(.VSS(VSS),.VDD(VDD),.Y(g14438),.A(g1087),.B(g10726));
  AND2 AND2_741(.VSS(VSS),.VDD(VDD),.Y(g30043),.A(g29106),.B(g9392));
  AND2 AND2_742(.VSS(VSS),.VDD(VDD),.Y(g18253),.A(g1211),.B(g16897));
  AND2 AND2_743(.VSS(VSS),.VDD(VDD),.Y(g25132),.A(g10497),.B(g23528));
  AND2 AND2_744(.VSS(VSS),.VDD(VDD),.Y(g30244),.A(g28732),.B(g23930));
  AND4 AND4_42(.VSS(VSS),.VDD(VDD),.Y(g26171),.A(g25357),.B(g6856),.C(g11709),.D(g11686));
  AND2 AND2_745(.VSS(VSS),.VDD(VDD),.Y(g15700),.A(g3089),.B(g13483));
  AND3 AND3_47(.VSS(VSS),.VDD(VDD),.Y(I24051),.A(g3380),.B(g3385),.C(g8492));
  AND2 AND2_746(.VSS(VSS),.VDD(VDD),.Y(g18600),.A(g3111),.B(g16987));
  AND2 AND2_747(.VSS(VSS),.VDD(VDD),.Y(g20193),.A(g15578),.B(g17264));
  AND2 AND2_748(.VSS(VSS),.VDD(VDD),.Y(g18781),.A(g5831),.B(g18065));
  AND2 AND2_749(.VSS(VSS),.VDD(VDD),.Y(g28585),.A(g27063),.B(g10530));
  AND2 AND2_750(.VSS(VSS),.VDD(VDD),.Y(g24193),.A(g336),.B(g22722));
  AND4 AND4_43(.VSS(VSS),.VDD(VDD),.Y(g28484),.A(g27187),.B(g10290),.C(g21163),.D(I26972));
  AND2 AND2_751(.VSS(VSS),.VDD(VDD),.Y(g33420),.A(g32373),.B(g21454));
  AND2 AND2_752(.VSS(VSS),.VDD(VDD),.Y(g30069),.A(g29175),.B(g12708));
  AND2 AND2_753(.VSS(VSS),.VDD(VDD),.Y(g29766),.A(g28316),.B(g23235));
  AND2 AND2_754(.VSS(VSS),.VDD(VDD),.Y(g18236),.A(g15065),.B(g16326));
  AND2 AND2_755(.VSS(VSS),.VDD(VDD),.Y(g21782),.A(g3416),.B(g20391));
  AND2 AND2_756(.VSS(VSS),.VDD(VDD),.Y(g17771),.A(g13288),.B(g13190));
  AND2 AND2_757(.VSS(VSS),.VDD(VDD),.Y(g20165),.A(g5156),.B(g17733));
  AND2 AND2_758(.VSS(VSS),.VDD(VDD),.Y(g34069),.A(g8774),.B(g33797));
  AND2 AND2_759(.VSS(VSS),.VDD(VDD),.Y(g21984),.A(g5563),.B(g19074));
  AND4 AND4_44(.VSS(VSS),.VDD(VDD),.Y(I31102),.A(g32603),.B(g32604),.C(g32605),.D(g32606));
  AND4 AND4_45(.VSS(VSS),.VDD(VDD),.Y(g26994),.A(g23032),.B(g26226),.C(g26424),.D(g25557));
  AND4 AND4_46(.VSS(VSS),.VDD(VDD),.Y(g27474),.A(g8038),.B(g26314),.C(g518),.D(g504));
  AND2 AND2_760(.VSS(VSS),.VDD(VDD),.Y(g28554),.A(g27426),.B(g20372));
  AND4 AND4_47(.VSS(VSS),.VDD(VDD),.Y(I31157),.A(g32682),.B(g32683),.C(g32684),.D(g32685));
  AND2 AND2_761(.VSS(VSS),.VDD(VDD),.Y(g18351),.A(g1760),.B(g17955));
  AND2 AND2_762(.VSS(VSS),.VDD(VDD),.Y(g18372),.A(g1886),.B(g15171));
  AND2 AND2_763(.VSS(VSS),.VDD(VDD),.Y(g24523),.A(g22318),.B(g19468));
  AND2 AND2_764(.VSS(VSS),.VDD(VDD),.Y(g32314),.A(g31304),.B(g23516));
  AND2 AND2_765(.VSS(VSS),.VDD(VDD),.Y(g29871),.A(g28400),.B(g23332));
  AND2 AND2_766(.VSS(VSS),.VDD(VDD),.Y(g33446),.A(g32385),.B(g21607));
  AND4 AND4_48(.VSS(VSS),.VDD(VDD),.Y(g27711),.A(g22369),.B(g25193),.C(g26424),.D(g26166));
  AND2 AND2_767(.VSS(VSS),.VDD(VDD),.Y(g16707),.A(g6641),.B(g15033));
  AND2 AND2_768(.VSS(VSS),.VDD(VDD),.Y(g21419),.A(g16681),.B(g13595));
  AND2 AND2_769(.VSS(VSS),.VDD(VDD),.Y(g32287),.A(g2823),.B(g30578));
  AND2 AND2_770(.VSS(VSS),.VDD(VDD),.Y(g34774),.A(g34695),.B(g20180));
  AND2 AND2_771(.VSS(VSS),.VDD(VDD),.Y(g18175),.A(g744),.B(g17328));
  AND2 AND2_772(.VSS(VSS),.VDD(VDD),.Y(g18821),.A(g15168),.B(g15680));
  AND2 AND2_773(.VSS(VSS),.VDD(VDD),.Y(g34955),.A(g34931),.B(g34320));
  AND2 AND2_774(.VSS(VSS),.VDD(VDD),.Y(g27327),.A(g2116),.B(g26732));
  AND2 AND2_775(.VSS(VSS),.VDD(VDD),.Y(g34375),.A(g13077),.B(g34049));
  AND2 AND2_776(.VSS(VSS),.VDD(VDD),.Y(g16202),.A(g86),.B(g14197));
  AND2 AND2_777(.VSS(VSS),.VDD(VDD),.Y(g28312),.A(g27828),.B(g26608));
  AND2 AND2_778(.VSS(VSS),.VDD(VDD),.Y(g28200),.A(g27652),.B(g11383));
  AND2 AND2_779(.VSS(VSS),.VDD(VDD),.Y(g32307),.A(g31291),.B(g23500));
  AND2 AND2_780(.VSS(VSS),.VDD(VDD),.Y(g14566),.A(g10566),.B(g10551));
  AND2 AND2_781(.VSS(VSS),.VDD(VDD),.Y(g32085),.A(g27253),.B(g31021));
  AND4 AND4_49(.VSS(VSS),.VDD(VDD),.Y(I31066),.A(g31070),.B(g31807),.C(g32550),.D(g32551));
  AND2 AND2_782(.VSS(VSS),.VDD(VDD),.Y(g29360),.A(g27364),.B(g28294));
  AND2 AND2_783(.VSS(VSS),.VDD(VDD),.Y(g21822),.A(g3727),.B(g20453));
  AND2 AND2_784(.VSS(VSS),.VDD(VDD),.Y(g22515),.A(g12981),.B(g19395));
  AND4 AND4_50(.VSS(VSS),.VDD(VDD),.Y(I31231),.A(g31376),.B(g31836),.C(g32789),.D(g32790));
  AND2 AND2_785(.VSS(VSS),.VDD(VDD),.Y(g22991),.A(g645),.B(g20248));
  AND2 AND2_786(.VSS(VSS),.VDD(VDD),.Y(g27537),.A(g26549),.B(g17742));
  AND2 AND2_787(.VSS(VSS),.VDD(VDD),.Y(g28115),.A(g27354),.B(g22759));
  AND2 AND2_788(.VSS(VSS),.VDD(VDD),.Y(g31540),.A(g29904),.B(g23548));
  AND2 AND2_789(.VSS(VSS),.VDD(VDD),.Y(g25087),.A(g17307),.B(g23489));
  AND2 AND2_790(.VSS(VSS),.VDD(VDD),.Y(g32054),.A(g10890),.B(g30735));
  AND2 AND2_791(.VSS(VSS),.VDD(VDD),.Y(g24475),.A(g3831),.B(g23139));
  AND2 AND2_792(.VSS(VSS),.VDD(VDD),.Y(g7685),.A(g4382),.B(g4375));
  AND2 AND2_793(.VSS(VSS),.VDD(VDD),.Y(g18264),.A(g1263),.B(g16000));
  AND2 AND2_794(.VSS(VSS),.VDD(VDD),.Y(g18790),.A(g6040),.B(g15634));
  AND2 AND2_795(.VSS(VSS),.VDD(VDD),.Y(g18137),.A(g538),.B(g17249));
  AND4 AND4_51(.VSS(VSS),.VDD(VDD),.Y(I27513),.A(g19984),.B(g24089),.C(g24090),.D(g28034));
  AND2 AND2_796(.VSS(VSS),.VDD(VDD),.Y(g18516),.A(g2638),.B(g15509));
  AND2 AND2_797(.VSS(VSS),.VDD(VDD),.Y(g34337),.A(g34095),.B(g19881));
  AND2 AND2_798(.VSS(VSS),.VDD(VDD),.Y(g24727),.A(g13300),.B(g23016));
  AND2 AND2_799(.VSS(VSS),.VDD(VDD),.Y(g34171),.A(g33925),.B(g24360));
  AND2 AND2_800(.VSS(VSS),.VDD(VDD),.Y(g16590),.A(g5236),.B(g14683));
  AND2 AND2_801(.VSS(VSS),.VDD(VDD),.Y(g24222),.A(g262),.B(g22594));
  AND2 AND2_802(.VSS(VSS),.VDD(VDD),.Y(g16986),.A(g246),.B(g13142));
  AND2 AND2_803(.VSS(VSS),.VDD(VDD),.Y(g27303),.A(g11996),.B(g26681));
  AND2 AND2_804(.VSS(VSS),.VDD(VDD),.Y(g11223),.A(g8281),.B(g8505));
  AND2 AND2_805(.VSS(VSS),.VDD(VDD),.Y(g25043),.A(g20733),.B(g23447));
  AND2 AND2_806(.VSS(VSS),.VDD(VDD),.Y(g32269),.A(g31253),.B(g20443));
  AND2 AND2_807(.VSS(VSS),.VDD(VDD),.Y(g21853),.A(g3917),.B(g21070));
  AND4 AND4_52(.VSS(VSS),.VDD(VDD),.Y(g28799),.A(g21434),.B(g26424),.C(g25348),.D(g27445));
  AND2 AND2_808(.VSS(VSS),.VDD(VDD),.Y(g26079),.A(g6199),.B(g25060));
  AND2 AND2_809(.VSS(VSS),.VDD(VDD),.Y(g34967),.A(g34951),.B(g23189));
  AND2 AND2_810(.VSS(VSS),.VDD(VDD),.Y(g28813),.A(g4104),.B(g27038));
  AND2 AND2_811(.VSS(VSS),.VDD(VDD),.Y(g29629),.A(g28211),.B(g19779));
  AND2 AND2_812(.VSS(VSS),.VDD(VDD),.Y(g32341),.A(g31472),.B(g23610));
  AND2 AND2_813(.VSS(VSS),.VDD(VDD),.Y(g31281),.A(g30106),.B(g27742));
  AND2 AND2_814(.VSS(VSS),.VDD(VDD),.Y(g15870),.A(g3231),.B(g13948));
  AND2 AND2_815(.VSS(VSS),.VDD(VDD),.Y(g26078),.A(g5128),.B(g25055));
  AND2 AND2_816(.VSS(VSS),.VDD(VDD),.Y(g32156),.A(g31639),.B(g30018));
  AND2 AND2_817(.VSS(VSS),.VDD(VDD),.Y(g25069),.A(g23296),.B(g20535));
  AND2 AND2_818(.VSS(VSS),.VDD(VDD),.Y(g24703),.A(g17592),.B(g22369));
  AND2 AND2_819(.VSS(VSS),.VDD(VDD),.Y(g31301),.A(g30170),.B(g27907));
  AND2 AND2_820(.VSS(VSS),.VDD(VDD),.Y(g18209),.A(g921),.B(g15938));
  AND2 AND2_821(.VSS(VSS),.VDD(VDD),.Y(g29628),.A(g27924),.B(g28648));
  AND2 AND2_822(.VSS(VSS),.VDD(VDD),.Y(g33902),.A(g33085),.B(g13202));
  AND2 AND2_823(.VSS(VSS),.VDD(VDD),.Y(g21836),.A(g3805),.B(g20453));
  AND2 AND2_824(.VSS(VSS),.VDD(VDD),.Y(g31120),.A(g1700),.B(g29976));
  AND2 AND2_825(.VSS(VSS),.VDD(VDD),.Y(g32180),.A(g2791),.B(g31638));
  AND2 AND2_826(.VSS(VSS),.VDD(VDD),.Y(g23836),.A(g4129),.B(g19495));
  AND2 AND2_827(.VSS(VSS),.VDD(VDD),.Y(g26086),.A(g9672),.B(g25255));
  AND2 AND2_828(.VSS(VSS),.VDD(VDD),.Y(g28674),.A(g27569),.B(g20629));
  AND2 AND2_829(.VSS(VSS),.VDD(VDD),.Y(g13321),.A(g847),.B(g11048));
  AND2 AND2_830(.VSS(VSS),.VDD(VDD),.Y(g25068),.A(g17574),.B(g23477));
  AND2 AND2_831(.VSS(VSS),.VDD(VDD),.Y(g25955),.A(g24720),.B(g19580));
  AND2 AND2_832(.VSS(VSS),.VDD(VDD),.Y(g30919),.A(g29898),.B(g23286));
  AND2 AND2_833(.VSS(VSS),.VDD(VDD),.Y(g18208),.A(g930),.B(g15938));
  AND2 AND2_834(.VSS(VSS),.VDD(VDD),.Y(g16801),.A(g5120),.B(g14238));
  AND2 AND2_835(.VSS(VSS),.VDD(VDD),.Y(g16735),.A(g6235),.B(g15027));
  AND2 AND2_836(.VSS(VSS),.VDD(VDD),.Y(g23401),.A(g7262),.B(g21460));
  AND2 AND2_837(.VSS(VSS),.VDD(VDD),.Y(g25879),.A(g11135),.B(g24683));
  AND2 AND2_838(.VSS(VSS),.VDD(VDD),.Y(g24600),.A(g22591),.B(g19652));
  AND2 AND2_839(.VSS(VSS),.VDD(VDD),.Y(g25970),.A(g1792),.B(g24991));
  AND2 AND2_840(.VSS(VSS),.VDD(VDD),.Y(g31146),.A(g12285),.B(g30053));
  AND2 AND2_841(.VSS(VSS),.VDD(VDD),.Y(g30010),.A(g29035),.B(g9274));
  AND2 AND2_842(.VSS(VSS),.VDD(VDD),.Y(g30918),.A(g8681),.B(g29707));
  AND2 AND2_843(.VSS(VSS),.VDD(VDD),.Y(g32335),.A(g6199),.B(g31566));
  AND4 AND4_53(.VSS(VSS),.VDD(VDD),.Y(g11178),.A(g6682),.B(g7097),.C(g6668),.D(g10061));
  AND2 AND2_844(.VSS(VSS),.VDD(VDD),.Y(g11740),.A(g8769),.B(g703));
  AND2 AND2_845(.VSS(VSS),.VDD(VDD),.Y(g18542),.A(g2787),.B(g15277));
  AND3 AND3_48(.VSS(VSS),.VDD(VDD),.Y(I18803),.A(g13156),.B(g11450),.C(g6756));
  AND2 AND2_846(.VSS(VSS),.VDD(VDD),.Y(g18453),.A(g2315),.B(g15224));
  AND2 AND2_847(.VSS(VSS),.VDD(VDD),.Y(g29591),.A(g28552),.B(g11346));
  AND2 AND2_848(.VSS(VSS),.VDD(VDD),.Y(g29785),.A(g28332),.B(g23248));
  AND2 AND2_849(.VSS(VSS),.VDD(VDD),.Y(g31290),.A(g29734),.B(g23335));
  AND2 AND2_850(.VSS(VSS),.VDD(VDD),.Y(g22114),.A(g6565),.B(g19277));
  AND2 AND2_851(.VSS(VSS),.VDD(VDD),.Y(g26159),.A(g2370),.B(g25137));
  AND2 AND2_852(.VSS(VSS),.VDD(VDD),.Y(g26125),.A(g1894),.B(g25117));
  AND2 AND2_853(.VSS(VSS),.VDD(VDD),.Y(g21864),.A(g3961),.B(g21070));
  AND2 AND2_854(.VSS(VSS),.VDD(VDD),.Y(g34079),.A(g33703),.B(g19532));
  AND2 AND2_855(.VSS(VSS),.VDD(VDD),.Y(g22082),.A(g6283),.B(g19210));
  AND2 AND2_856(.VSS(VSS),.VDD(VDD),.Y(g27390),.A(g26549),.B(g17504));
  AND2 AND2_857(.VSS(VSS),.VDD(VDD),.Y(g18726),.A(g4927),.B(g16077));
  AND4 AND4_54(.VSS(VSS),.VDD(VDD),.Y(g26977),.A(g23032),.B(g26261),.C(g26424),.D(g25550));
  AND2 AND2_858(.VSS(VSS),.VDD(VDD),.Y(g30599),.A(g18911),.B(g29863));
  AND2 AND2_859(.VSS(VSS),.VDD(VDD),.Y(g22107),.A(g6411),.B(g18833));
  AND2 AND2_860(.VSS(VSS),.VDD(VDD),.Y(g30078),.A(g28526),.B(g20667));
  AND2 AND2_861(.VSS(VSS),.VDD(VDD),.Y(g21749),.A(g3155),.B(g20785));
  AND2 AND2_862(.VSS(VSS),.VDD(VDD),.Y(g26158),.A(g2255),.B(g25432));
  AND4 AND4_55(.VSS(VSS),.VDD(VDD),.Y(g17725),.A(g11547),.B(g11592),.C(g6789),.D(I18716));
  AND2 AND2_863(.VSS(VSS),.VDD(VDD),.Y(g26783),.A(g25037),.B(g21048));
  AND4 AND4_56(.VSS(VSS),.VDD(VDD),.Y(I31287),.A(g32870),.B(g32871),.C(g32872),.D(g32873));
  AND2 AND2_864(.VSS(VSS),.VDD(VDD),.Y(g18614),.A(g3343),.B(g17200));
  AND2 AND2_865(.VSS(VSS),.VDD(VDD),.Y(g28692),.A(g27578),.B(g20661));
  AND4 AND4_57(.VSS(VSS),.VDD(VDD),.Y(g28761),.A(g21434),.B(g26424),.C(g25299),.D(g27416));
  AND2 AND2_866(.VSS(VSS),.VDD(VDD),.Y(g34078),.A(g33699),.B(g19531));
  AND2 AND2_867(.VSS(VSS),.VDD(VDD),.Y(g18436),.A(g2227),.B(g18008));
  AND2 AND2_868(.VSS(VSS),.VDD(VDD),.Y(g25967),.A(g9373),.B(g24986));
  AND2 AND2_869(.VSS(VSS),.VDD(VDD),.Y(g30598),.A(g18898),.B(g29862));
  AND2 AND2_870(.VSS(VSS),.VDD(VDD),.Y(g14585),.A(g1141),.B(g10905));
  AND2 AND2_871(.VSS(VSS),.VDD(VDD),.Y(g29859),.A(g28388),.B(g23307));
  AND4 AND4_58(.VSS(VSS),.VDD(VDD),.Y(I31307),.A(g32898),.B(g32899),.C(g32900),.D(g32901));
  AND4 AND4_59(.VSS(VSS),.VDD(VDD),.Y(I31076),.A(g30614),.B(g31809),.C(g32564),.D(g32565));
  AND2 AND2_872(.VSS(VSS),.VDD(VDD),.Y(g30086),.A(g28536),.B(g20704));
  AND2 AND2_873(.VSS(VSS),.VDD(VDD),.Y(g21748),.A(g15089),.B(g20785));
  AND2 AND2_874(.VSS(VSS),.VDD(VDD),.Y(g15707),.A(g4082),.B(g13506));
  AND2 AND2_875(.VSS(VSS),.VDD(VDD),.Y(g15819),.A(g3251),.B(g14101));
  AND2 AND2_876(.VSS(VSS),.VDD(VDD),.Y(g18607),.A(g3139),.B(g16987));
  AND3 AND3_49(.VSS(VSS),.VDD(VDD),.Y(g34086),.A(g20114),.B(g33766),.C(g9104));
  AND2 AND2_877(.VSS(VSS),.VDD(VDD),.Y(g18320),.A(g1616),.B(g17873));
  AND2 AND2_878(.VSS(VSS),.VDD(VDD),.Y(g24790),.A(g7074),.B(g23681));
  AND2 AND2_879(.VSS(VSS),.VDD(VDD),.Y(g21276),.A(g10157),.B(g17625));
  AND2 AND2_880(.VSS(VSS),.VDD(VDD),.Y(g21285),.A(g7857),.B(g16027));
  AND2 AND2_881(.VSS(VSS),.VDD(VDD),.Y(g26295),.A(g13070),.B(g25266));
  AND2 AND2_882(.VSS(VSS),.VDD(VDD),.Y(g29858),.A(g28387),.B(g23306));
  AND2 AND2_883(.VSS(VSS),.VDD(VDD),.Y(g21704),.A(g164),.B(g20283));
  AND2 AND2_884(.VSS(VSS),.VDD(VDD),.Y(g18274),.A(g1311),.B(g16031));
  AND2 AND2_885(.VSS(VSS),.VDD(VDD),.Y(g22849),.A(g1227),.B(g19653));
  AND2 AND2_886(.VSS(VSS),.VDD(VDD),.Y(g33366),.A(g32268),.B(g21010));
  AND2 AND2_887(.VSS(VSS),.VDD(VDD),.Y(g27522),.A(g26549),.B(g17717));
  AND2 AND2_888(.VSS(VSS),.VDD(VDD),.Y(g26823),.A(g24401),.B(g13106));
  AND2 AND2_889(.VSS(VSS),.VDD(VDD),.Y(g15818),.A(g3941),.B(g14082));
  AND2 AND2_890(.VSS(VSS),.VDD(VDD),.Y(g18530),.A(g2715),.B(g15277));
  AND3 AND3_50(.VSS(VSS),.VDD(VDD),.Y(g25459),.A(g6058),.B(g23844),.C(I24582));
  AND2 AND2_891(.VSS(VSS),.VDD(VDD),.Y(g18593),.A(g2999),.B(g16349));
  AND2 AND2_892(.VSS(VSS),.VDD(VDD),.Y(g18346),.A(g1752),.B(g17955));
  AND2 AND2_893(.VSS(VSS),.VDD(VDD),.Y(g19716),.A(g12100),.B(g17121));
  AND2 AND2_894(.VSS(VSS),.VDD(VDD),.Y(g21809),.A(g3574),.B(g20924));
  AND2 AND2_895(.VSS(VSS),.VDD(VDD),.Y(g23254),.A(g20056),.B(g20110));
  AND2 AND2_896(.VSS(VSS),.VDD(VDD),.Y(g28214),.A(g27731),.B(g26625));
  AND2 AND2_897(.VSS(VSS),.VDD(VDD),.Y(g15111),.A(g4281),.B(g14454));
  AND2 AND2_898(.VSS(VSS),.VDD(VDD),.Y(g22848),.A(g19449),.B(g19649));
  AND2 AND2_899(.VSS(VSS),.VDD(VDD),.Y(g18122),.A(g15052),.B(g17015));
  AND2 AND2_900(.VSS(VSS),.VDD(VDD),.Y(g23900),.A(g1129),.B(g19408));
  AND2 AND2_901(.VSS(VSS),.VDD(VDD),.Y(g34322),.A(g14188),.B(g34174));
  AND4 AND4_60(.VSS(VSS),.VDD(VDD),.Y(g14608),.A(g12638),.B(g12476),.C(g12429),.D(I16721));
  AND2 AND2_902(.VSS(VSS),.VDD(VDD),.Y(g15978),.A(g246),.B(g14032));
  AND2 AND2_903(.VSS(VSS),.VDD(VDD),.Y(g18565),.A(g2852),.B(g16349));
  AND2 AND2_904(.VSS(VSS),.VDD(VDD),.Y(g26336),.A(g10307),.B(g25480));
  AND2 AND2_905(.VSS(VSS),.VDD(VDD),.Y(g30125),.A(g28581),.B(g21056));
  AND2 AND2_906(.VSS(VSS),.VDD(VDD),.Y(g18464),.A(g2370),.B(g15224));
  AND2 AND2_907(.VSS(VSS),.VDD(VDD),.Y(g21808),.A(g3570),.B(g20924));
  AND2 AND2_908(.VSS(VSS),.VDD(VDD),.Y(g29844),.A(g28374),.B(g23290));
  AND2 AND2_909(.VSS(VSS),.VDD(VDD),.Y(g34532),.A(g34314),.B(g19710));
  AND2 AND2_910(.VSS(VSS),.VDD(VDD),.Y(g15590),.A(g3139),.B(g13530));
  AND2 AND2_911(.VSS(VSS),.VDD(VDD),.Y(g29367),.A(g8575),.B(g28325));
  AND2 AND2_912(.VSS(VSS),.VDD(VDD),.Y(g28539),.A(g27187),.B(g12762));
  AND2 AND2_913(.VSS(VSS),.VDD(VDD),.Y(g10921),.A(g1548),.B(g8685));
  AND2 AND2_914(.VSS(VSS),.VDD(VDD),.Y(g27483),.A(g26488),.B(g17642));
  AND2 AND2_915(.VSS(VSS),.VDD(VDD),.Y(g30158),.A(g28613),.B(g21274));
  AND2 AND2_916(.VSS(VSS),.VDD(VDD),.Y(g33403),.A(g32352),.B(g21396));
  AND2 AND2_917(.VSS(VSS),.VDD(VDD),.Y(g24422),.A(g4771),.B(g22896));
  AND4 AND4_61(.VSS(VSS),.VDD(VDD),.Y(I31341),.A(g31710),.B(g31856),.C(g32947),.D(g32948));
  AND2 AND2_918(.VSS(VSS),.VDD(VDD),.Y(g32278),.A(g2811),.B(g30572));
  AND2 AND2_919(.VSS(VSS),.VDD(VDD),.Y(g27553),.A(g26293),.B(g23353));
  AND2 AND2_920(.VSS(VSS),.VDD(VDD),.Y(g18641),.A(g3841),.B(g17096));
  AND2 AND2_921(.VSS(VSS),.VDD(VDD),.Y(g18797),.A(g6173),.B(g15348));
  AND2 AND2_922(.VSS(VSS),.VDD(VDD),.Y(g25079),.A(g21011),.B(g23483));
  AND4 AND4_62(.VSS(VSS),.VDD(VDD),.Y(I31156),.A(g31070),.B(g31823),.C(g32680),.D(g32681));
  AND2 AND2_923(.VSS(VSS),.VDD(VDD),.Y(g18292),.A(g1472),.B(g16449));
  AND2 AND2_924(.VSS(VSS),.VDD(VDD),.Y(g16706),.A(g6621),.B(g14868));
  AND2 AND2_925(.VSS(VSS),.VDD(VDD),.Y(g31226),.A(g30282),.B(g25218));
  AND2 AND2_926(.VSS(VSS),.VDD(VDD),.Y(g32286),.A(g31658),.B(g29312));
  AND2 AND2_927(.VSS(VSS),.VDD(VDD),.Y(g34561),.A(g34368),.B(g17410));
  AND2 AND2_928(.VSS(VSS),.VDD(VDD),.Y(g16597),.A(g6263),.B(g15021));
  AND2 AND2_929(.VSS(VSS),.VDD(VDD),.Y(g18153),.A(g626),.B(g17533));
  AND2 AND2_930(.VSS(VSS),.VDD(VDD),.Y(g27326),.A(g12048),.B(g26731));
  AND2 AND2_931(.VSS(VSS),.VDD(VDD),.Y(g25078),.A(g23298),.B(g20538));
  AND2 AND2_932(.VSS(VSS),.VDD(VDD),.Y(g31481),.A(g29768),.B(g23417));
  AND2 AND2_933(.VSS(VSS),.VDD(VDD),.Y(g32039),.A(g31476),.B(g20070));
  AND2 AND2_934(.VSS(VSS),.VDD(VDD),.Y(g33715),.A(g33135),.B(g19416));
  AND2 AND2_935(.VSS(VSS),.VDD(VDD),.Y(g32306),.A(g31289),.B(g23499));
  AND2 AND2_936(.VSS(VSS),.VDD(VDD),.Y(g34295),.A(g34057),.B(g19370));
  AND3 AND3_51(.VSS(VSS),.VDD(VDD),.Y(g33481),.A(g32607),.B(I31101),.C(I31102));
  AND2 AND2_937(.VSS(VSS),.VDD(VDD),.Y(g22135),.A(g6657),.B(g19277));
  AND2 AND2_938(.VSS(VSS),.VDD(VDD),.Y(g27536),.A(g26519),.B(g17738));
  AND2 AND2_939(.VSS(VSS),.VDD(VDD),.Y(g18409),.A(g2084),.B(g15373));
  AND4 AND4_63(.VSS(VSS),.VDD(VDD),.Y(g27040),.A(g7812),.B(g6565),.C(g6573),.D(g26226));
  AND2 AND2_940(.VSS(VSS),.VDD(VDD),.Y(g25086),.A(g13941),.B(g23488));
  AND2 AND2_941(.VSS(VSS),.VDD(VDD),.Y(g21733),.A(g3034),.B(g20330));
  AND3 AND3_52(.VSS(VSS),.VDD(VDD),.Y(g10674),.A(g6841),.B(g10200),.C(g2130));
  AND2 AND2_942(.VSS(VSS),.VDD(VDD),.Y(g18136),.A(g550),.B(g17249));
  AND2 AND2_943(.VSS(VSS),.VDD(VDD),.Y(g18408),.A(g2070),.B(g15373));
  AND2 AND2_944(.VSS(VSS),.VDD(VDD),.Y(g18635),.A(g3808),.B(g17096));
  AND2 AND2_945(.VSS(VSS),.VDD(VDD),.Y(g24726),.A(g15965),.B(g23015));
  AND2 AND2_946(.VSS(VSS),.VDD(VDD),.Y(g27252),.A(g26733),.B(g26703));
  AND2 AND2_947(.VSS(VSS),.VDD(VDD),.Y(g24913),.A(g4821),.B(g23908));
  AND2 AND2_948(.VSS(VSS),.VDD(VDD),.Y(g21874),.A(g4112),.B(g19801));
  AND2 AND2_949(.VSS(VSS),.VDD(VDD),.Y(g25817),.A(g24807),.B(g21163));
  AND2 AND2_950(.VSS(VSS),.VDD(VDD),.Y(g32187),.A(g30672),.B(g25287));
  AND2 AND2_951(.VSS(VSS),.VDD(VDD),.Y(g26289),.A(g2551),.B(g25400));
  AND2 AND2_952(.VSS(VSS),.VDD(VDD),.Y(g24436),.A(g3125),.B(g23067));
  AND2 AND2_953(.VSS(VSS),.VDD(VDD),.Y(g25159),.A(g4907),.B(g22908));
  AND3 AND3_53(.VSS(VSS),.VDD(VDD),.Y(g10732),.A(g6850),.B(g2697),.C(g2689));
  AND2 AND2_954(.VSS(VSS),.VDD(VDD),.Y(g22049),.A(g6082),.B(g21611));
  AND2 AND2_955(.VSS(VSS),.VDD(VDD),.Y(g25125),.A(g20187),.B(g23520));
  AND2 AND2_956(.VSS(VSS),.VDD(VDD),.Y(g27564),.A(g26305),.B(g23378));
  AND2 AND2_957(.VSS(VSS),.VDD(VDD),.Y(g25901),.A(g24853),.B(g16290));
  AND2 AND2_958(.VSS(VSS),.VDD(VDD),.Y(g26023),.A(g9528),.B(g25036));
  AND4 AND4_64(.VSS(VSS),.VDD(VDD),.Y(I31131),.A(g31542),.B(g31819),.C(g32643),.D(g32644));
  AND2 AND2_959(.VSS(VSS),.VDD(VDD),.Y(g34966),.A(g34950),.B(g23170));
  AND2 AND2_960(.VSS(VSS),.VDD(VDD),.Y(g31490),.A(g29786),.B(g23429));
  AND2 AND2_961(.VSS(VSS),.VDD(VDD),.Y(g10934),.A(g9197),.B(g7918));
  AND2 AND2_962(.VSS(VSS),.VDD(VDD),.Y(g24607),.A(g5817),.B(g23666));
  AND2 AND2_963(.VSS(VSS),.VDD(VDD),.Y(g25977),.A(g25236),.B(g20875));
  AND2 AND2_964(.VSS(VSS),.VDD(VDD),.Y(g26288),.A(g2259),.B(g25309));
  AND3 AND3_54(.VSS(VSS),.VDD(VDD),.Y(g33490),.A(g32672),.B(I31146),.C(I31147));
  AND2 AND2_965(.VSS(VSS),.VDD(VDD),.Y(g19681),.A(g5835),.B(g17014));
  AND2 AND2_966(.VSS(VSS),.VDD(VDD),.Y(g24320),.A(g6973),.B(g22228));
  AND2 AND2_967(.VSS(VSS),.VDD(VDD),.Y(g28235),.A(g9467),.B(g27592));
  AND2 AND2_968(.VSS(VSS),.VDD(VDD),.Y(g26571),.A(g10472),.B(g24386));
  AND2 AND2_969(.VSS(VSS),.VDD(VDD),.Y(g23166),.A(g13959),.B(g19979));
  AND2 AND2_970(.VSS(VSS),.VDD(VDD),.Y(g23009),.A(g20196),.B(g14219));
  AND2 AND2_971(.VSS(VSS),.VDD(VDD),.Y(g22048),.A(g6052),.B(g21611));
  AND2 AND2_972(.VSS(VSS),.VDD(VDD),.Y(g26308),.A(g6961),.B(g25289));
  AND3 AND3_55(.VSS(VSS),.VDD(VDD),.Y(g29203),.A(g24095),.B(I27513),.C(I27514));
  AND2 AND2_973(.VSS(VSS),.VDD(VDD),.Y(g18164),.A(g699),.B(g17433));
  AND2 AND2_974(.VSS(VSS),.VDD(VDD),.Y(g28683),.A(g27876),.B(g20649));
  AND2 AND2_975(.VSS(VSS),.VDD(VDD),.Y(g32143),.A(g31646),.B(g29967));
  AND2 AND2_976(.VSS(VSS),.VDD(VDD),.Y(g31784),.A(g30176),.B(g24003));
  AND2 AND2_977(.VSS(VSS),.VDD(VDD),.Y(g34364),.A(g34048),.B(g24366));
  AND2 AND2_978(.VSS(VSS),.VDD(VDD),.Y(g33784),.A(g33107),.B(g20531));
  AND2 AND2_979(.VSS(VSS),.VDD(VDD),.Y(g31376),.A(g24952),.B(g29814));
  AND2 AND2_980(.VSS(VSS),.VDD(VDD),.Y(g31297),.A(g30144),.B(g27837));
  AND2 AND2_981(.VSS(VSS),.VDD(VDD),.Y(g27183),.A(g26055),.B(g16658));
  AND2 AND2_982(.VSS(VSS),.VDD(VDD),.Y(g33376),.A(g32294),.B(g21268));
  AND2 AND2_983(.VSS(VSS),.VDD(VDD),.Y(g27673),.A(g25769),.B(g23541));
  AND2 AND2_984(.VSS(VSS),.VDD(VDD),.Y(g22004),.A(g5742),.B(g21562));
  AND2 AND2_985(.VSS(VSS),.VDD(VDD),.Y(g23008),.A(g1570),.B(g19783));
  AND2 AND2_986(.VSS(VSS),.VDD(VDD),.Y(g33889),.A(g33303),.B(g20641));
  AND4 AND4_65(.VSS(VSS),.VDD(VDD),.Y(g11123),.A(g5644),.B(g7028),.C(g5630),.D(g9864));
  AND2 AND2_987(.VSS(VSS),.VDD(VDD),.Y(g24464),.A(g3480),.B(g23112));
  AND3 AND3_56(.VSS(VSS),.VDD(VDD),.Y(I24027),.A(g3029),.B(g3034),.C(g8426));
  AND2 AND2_988(.VSS(VSS),.VDD(VDD),.Y(g16885),.A(g6605),.B(g14950));
  AND2 AND2_989(.VSS(VSS),.VDD(VDD),.Y(g32169),.A(g31014),.B(g23046));
  AND2 AND2_990(.VSS(VSS),.VDD(VDD),.Y(g18575),.A(g2878),.B(g16349));
  AND2 AND2_991(.VSS(VSS),.VDD(VDD),.Y(g18474),.A(g2287),.B(g15224));
  AND2 AND2_992(.VSS(VSS),.VDD(VDD),.Y(g29902),.A(g28430),.B(g23377));
  AND2 AND2_993(.VSS(VSS),.VDD(VDD),.Y(g30289),.A(g28884),.B(g24000));
  AND2 AND2_994(.VSS(VSS),.VDD(VDD),.Y(g29377),.A(g28132),.B(g19387));
  AND2 AND2_995(.VSS(VSS),.VDD(VDD),.Y(g13807),.A(g4504),.B(g10606));
  AND2 AND2_996(.VSS(VSS),.VDD(VDD),.Y(g18711),.A(g15136),.B(g15915));
  AND2 AND2_997(.VSS(VSS),.VDD(VDD),.Y(g32168),.A(g30597),.B(g25185));
  AND2 AND2_998(.VSS(VSS),.VDD(VDD),.Y(g32410),.A(g4933),.B(g30997));
  AND4 AND4_66(.VSS(VSS),.VDD(VDD),.Y(g28991),.A(g14438),.B(g25209),.C(g26424),.D(g27469));
  AND2 AND2_999(.VSS(VSS),.VDD(VDD),.Y(g13974),.A(g6243),.B(g12578));
  AND2 AND2_1000(.VSS(VSS),.VDD(VDD),.Y(g18327),.A(g1636),.B(g17873));
  AND2 AND2_1001(.VSS(VSS),.VDD(VDD),.Y(g24797),.A(g22872),.B(g19960));
  AND2 AND2_1002(.VSS(VSS),.VDD(VDD),.Y(g30023),.A(g28508),.B(g20570));
  AND2 AND2_1003(.VSS(VSS),.VDD(VDD),.Y(g21712),.A(g294),.B(g20283));
  AND3 AND3_57(.VSS(VSS),.VDD(VDD),.Y(I24482),.A(g9364),.B(g9607),.C(g5057));
  AND2 AND2_1004(.VSS(VSS),.VDD(VDD),.Y(g18109),.A(g437),.B(g17015));
  AND2 AND2_1005(.VSS(VSS),.VDD(VDD),.Y(g27508),.A(g26549),.B(g17684));
  AND2 AND2_1006(.VSS(VSS),.VDD(VDD),.Y(g16763),.A(g6239),.B(g14937));
  AND2 AND2_1007(.VSS(VSS),.VDD(VDD),.Y(g27634),.A(g26805),.B(g26793));
  AND2 AND2_1008(.VSS(VSS),.VDD(VDD),.Y(g34309),.A(g13947),.B(g34147));
  AND2 AND2_1009(.VSS(VSS),.VDD(VDD),.Y(g21914),.A(g5077),.B(g21468));
  AND2 AND2_1010(.VSS(VSS),.VDD(VDD),.Y(g24292),.A(g4443),.B(g22550));
  AND2 AND2_1011(.VSS(VSS),.VDD(VDD),.Y(g30224),.A(g28704),.B(g23896));
  AND2 AND2_1012(.VSS(VSS),.VDD(VDD),.Y(g18537),.A(g6856),.B(g15277));
  AND4 AND4_67(.VSS(VSS),.VDD(VDD),.Y(I24710),.A(g24071),.B(g24072),.C(g24073),.D(g24074));
  AND2 AND2_1013(.VSS(VSS),.VDD(VDD),.Y(g34224),.A(g33736),.B(g22670));
  AND3 AND3_58(.VSS(VSS),.VDD(VDD),.Y(g30308),.A(g29178),.B(g7004),.C(g5297));
  AND2 AND2_1014(.VSS(VSS),.VDD(VDD),.Y(g22106),.A(g6497),.B(g18833));
  AND3 AND3_59(.VSS(VSS),.VDD(VDD),.Y(I24552),.A(g9733),.B(g9316),.C(g5747));
  AND2 AND2_1015(.VSS(VSS),.VDD(VDD),.Y(g29645),.A(g1714),.B(g29018));
  AND3 AND3_60(.VSS(VSS),.VDD(VDD),.Y(I24003),.A(g8097),.B(g8334),.C(g3045));
  AND4 AND4_68(.VSS(VSS),.VDD(VDD),.Y(g17613),.A(g11547),.B(g11592),.C(g11640),.D(I18568));
  AND2 AND2_1016(.VSS(VSS),.VDD(VDD),.Y(g34571),.A(g27225),.B(g34299));
  AND2 AND2_1017(.VSS(VSS),.VDD(VDD),.Y(g18108),.A(g433),.B(g17015));
  AND2 AND2_1018(.VSS(VSS),.VDD(VDD),.Y(g14207),.A(g8639),.B(g11793));
  AND2 AND2_1019(.VSS(VSS),.VDD(VDD),.Y(g21907),.A(g5033),.B(g21468));
  AND4 AND4_69(.VSS(VSS),.VDD(VDD),.Y(I31286),.A(g30825),.B(g31846),.C(g32868),.D(g32869));
  AND3 AND3_61(.VSS(VSS),.VDD(VDD),.Y(I13862),.A(g7232),.B(g7219),.C(g7258));
  AND2 AND2_1020(.VSS(VSS),.VDD(VDD),.Y(g15077),.A(g2138),.B(g12955));
  AND2 AND2_1021(.VSS(VSS),.VDD(VDD),.Y(g24409),.A(g3484),.B(g23112));
  AND2 AND2_1022(.VSS(VSS),.VDD(VDD),.Y(g25966),.A(g9364),.B(g24985));
  AND4 AND4_70(.VSS(VSS),.VDD(VDD),.Y(I31306),.A(g30614),.B(g31850),.C(g32896),.D(g32897));
  AND2 AND2_1023(.VSS(VSS),.VDD(VDD),.Y(g13265),.A(g9018),.B(g11493));
  AND2 AND2_1024(.VSS(VSS),.VDD(VDD),.Y(g18283),.A(g1384),.B(g16136));
  AND2 AND2_1025(.VSS(VSS),.VDD(VDD),.Y(g15706),.A(g13296),.B(g13484));
  AND2 AND2_1026(.VSS(VSS),.VDD(VDD),.Y(g18606),.A(g3133),.B(g16987));
  AND2 AND2_1027(.VSS(VSS),.VDD(VDD),.Y(g18492),.A(g2523),.B(g15426));
  AND2 AND2_1028(.VSS(VSS),.VDD(VDD),.Y(g18303),.A(g1536),.B(g16489));
  AND2 AND2_1029(.VSS(VSS),.VDD(VDD),.Y(g24408),.A(g23989),.B(g18946));
  AND2 AND2_1030(.VSS(VSS),.VDD(VDD),.Y(g24635),.A(g19874),.B(g22883));
  AND2 AND2_1031(.VSS(VSS),.VDD(VDD),.Y(g34495),.A(g34274),.B(g19365));
  AND2 AND2_1032(.VSS(VSS),.VDD(VDD),.Y(g22033),.A(g5925),.B(g19147));
  AND2 AND2_1033(.VSS(VSS),.VDD(VDD),.Y(g27213),.A(g26026),.B(g16721));
  AND2 AND2_1034(.VSS(VSS),.VDD(VDD),.Y(g18750),.A(g15145),.B(g17847));
  AND2 AND2_1035(.VSS(VSS),.VDD(VDD),.Y(g31520),.A(g29879),.B(g23507));
  AND4 AND4_71(.VSS(VSS),.VDD(VDD),.Y(I31187),.A(g32726),.B(g32727),.C(g32728),.D(g32729));
  AND3 AND3_62(.VSS(VSS),.VDD(VDD),.Y(g33520),.A(g32888),.B(I31296),.C(I31297));
  AND2 AND2_1036(.VSS(VSS),.VDD(VDD),.Y(g18982),.A(g3835),.B(g16159));
  AND2 AND2_1037(.VSS(VSS),.VDD(VDD),.Y(g18381),.A(g1882),.B(g15171));
  AND2 AND2_1038(.VSS(VSS),.VDD(VDD),.Y(g34687),.A(g14181),.B(g34543));
  AND2 AND2_1039(.VSS(VSS),.VDD(VDD),.Y(g21941),.A(g5232),.B(g18997));
  AND2 AND2_1040(.VSS(VSS),.VDD(VDD),.Y(g26842),.A(g2894),.B(g24522));
  AND3 AND3_63(.VSS(VSS),.VDD(VDD),.Y(I27429),.A(g25562),.B(g26424),.C(g22698));
  AND2 AND2_1041(.VSS(VSS),.VDD(VDD),.Y(g27452),.A(g26400),.B(g17600));
  AND2 AND2_1042(.VSS(VSS),.VDD(VDD),.Y(g21382),.A(g10086),.B(g17625));
  AND2 AND2_1043(.VSS(VSS),.VDD(VDD),.Y(g29632),.A(g28899),.B(g22417));
  AND2 AND2_1044(.VSS(VSS),.VDD(VDD),.Y(g31211),.A(g10156),.B(g30102));
  AND4 AND4_72(.VSS(VSS),.VDD(VDD),.Y(g26195),.A(g25357),.B(g6856),.C(g11709),.D(g7558));
  AND2 AND2_1045(.VSS(VSS),.VDD(VDD),.Y(g34752),.A(g34675),.B(g19544));
  AND2 AND2_1046(.VSS(VSS),.VDD(VDD),.Y(g23675),.A(g19050),.B(g9104));
  AND2 AND2_1047(.VSS(VSS),.VDD(VDD),.Y(g18174),.A(g739),.B(g17328));
  AND2 AND2_1048(.VSS(VSS),.VDD(VDD),.Y(g27311),.A(g12431),.B(g26693));
  AND2 AND2_1049(.VSS(VSS),.VDD(VDD),.Y(g18796),.A(g6167),.B(g15348));
  AND2 AND2_1050(.VSS(VSS),.VDD(VDD),.Y(g28725),.A(g27596),.B(g20779));
  AND2 AND2_1051(.VSS(VSS),.VDD(VDD),.Y(g32084),.A(g10948),.B(g30825));
  AND2 AND2_1052(.VSS(VSS),.VDD(VDD),.Y(g32110),.A(g31639),.B(g29921));
  AND2 AND2_1053(.VSS(VSS),.VDD(VDD),.Y(g16596),.A(g5941),.B(g14892));
  AND2 AND2_1054(.VSS(VSS),.VDD(VDD),.Y(g28114),.A(g25869),.B(g27051));
  AND2 AND2_1055(.VSS(VSS),.VDD(VDD),.Y(g25571),.A(I24694),.B(I24695));
  AND2 AND2_1056(.VSS(VSS),.VDD(VDD),.Y(g33860),.A(g33270),.B(g20501));
  AND2 AND2_1057(.VSS(VSS),.VDD(VDD),.Y(g32321),.A(g27613),.B(g31376));
  AND2 AND2_1058(.VSS(VSS),.VDD(VDD),.Y(g16243),.A(g6483),.B(g14275));
  AND2 AND2_1059(.VSS(VSS),.VDD(VDD),.Y(g29661),.A(g1687),.B(g29015));
  AND2 AND2_1060(.VSS(VSS),.VDD(VDD),.Y(g29547),.A(g1748),.B(g28857));
  AND2 AND2_1061(.VSS(VSS),.VDD(VDD),.Y(g29895),.A(g2495),.B(g29170));
  AND2 AND2_1062(.VSS(VSS),.VDD(VDD),.Y(g28107),.A(g27970),.B(g18874));
  AND2 AND2_1063(.VSS(VSS),.VDD(VDD),.Y(g10683),.A(g7289),.B(g4438));
  AND2 AND2_1064(.VSS(VSS),.VDD(VDD),.Y(g32179),.A(g31748),.B(g27907));
  AND2 AND2_1065(.VSS(VSS),.VDD(VDD),.Y(g21935),.A(g5196),.B(g18997));
  AND2 AND2_1066(.VSS(VSS),.VDD(VDD),.Y(g18390),.A(g1978),.B(g15171));
  AND2 AND2_1067(.VSS(VSS),.VDD(VDD),.Y(g31497),.A(g20041),.B(g29930));
  AND3 AND3_64(.VSS(VSS),.VDD(VDD),.Y(g33497),.A(g32723),.B(I31181),.C(I31182));
  AND2 AND2_1068(.VSS(VSS),.VDD(VDD),.Y(g20109),.A(g17954),.B(g17616));
  AND2 AND2_1069(.VSS(VSS),.VDD(VDD),.Y(g24327),.A(g4549),.B(g22228));
  AND2 AND2_1070(.VSS(VSS),.VDD(VDD),.Y(g21883),.A(g4141),.B(g19801));
  AND2 AND2_1071(.VSS(VSS),.VDD(VDD),.Y(g32178),.A(g31747),.B(g27886));
  AND2 AND2_1072(.VSS(VSS),.VDD(VDD),.Y(g15876),.A(g13512),.B(g13223));
  AND2 AND2_1073(.VSS(VSS),.VDD(VDD),.Y(g24537),.A(g22626),.B(g10851));
  AND2 AND2_1074(.VSS(VSS),.VDD(VDD),.Y(g11116),.A(g9960),.B(g6466));
  AND2 AND2_1075(.VSS(VSS),.VDD(VDD),.Y(g20108),.A(g15508),.B(g11048));
  AND2 AND2_1076(.VSS(VSS),.VDD(VDD),.Y(g34842),.A(g34762),.B(g20168));
  AND2 AND2_1077(.VSS(VSS),.VDD(VDD),.Y(g18192),.A(g817),.B(g17821));
  AND2 AND2_1078(.VSS(VSS),.VDD(VDD),.Y(g22012),.A(g5752),.B(g21562));
  AND2 AND2_1079(.VSS(VSS),.VDD(VDD),.Y(g26544),.A(g7446),.B(g24357));
  AND4 AND4_73(.VSS(VSS),.VDD(VDD),.Y(I27504),.A(g24077),.B(g24078),.C(g24079),.D(g24080));
  AND3 AND3_65(.VSS(VSS),.VDD(VDD),.Y(I18620),.A(g13156),.B(g11450),.C(g11498));
  AND2 AND2_1080(.VSS(VSS),.VDD(VDD),.Y(g25816),.A(g8164),.B(g24604));
  AND2 AND2_1081(.VSS(VSS),.VDD(VDD),.Y(g33700),.A(g33148),.B(g11012));
  AND2 AND2_1082(.VSS(VSS),.VDD(VDD),.Y(g33126),.A(g9044),.B(g32201));
  AND2 AND2_1083(.VSS(VSS),.VDD(VDD),.Y(g31987),.A(g31767),.B(g22198));
  AND2 AND2_1084(.VSS(VSS),.VDD(VDD),.Y(g29551),.A(g2173),.B(g28867));
  AND2 AND2_1085(.VSS(VSS),.VDD(VDD),.Y(g29572),.A(g1620),.B(g28885));
  AND2 AND2_1086(.VSS(VSS),.VDD(VDD),.Y(g26713),.A(g25447),.B(g20714));
  AND4 AND4_74(.VSS(VSS),.VDD(VDD),.Y(I31217),.A(g32768),.B(g32769),.C(g32770),.D(g32771));
  AND2 AND2_1087(.VSS(VSS),.VDD(VDD),.Y(g34489),.A(g34421),.B(g19068));
  AND2 AND2_1088(.VSS(VSS),.VDD(VDD),.Y(g24283),.A(g4411),.B(g22550));
  AND2 AND2_1089(.VSS(VSS),.VDD(VDD),.Y(g18522),.A(g2671),.B(g15509));
  AND2 AND2_1090(.VSS(VSS),.VDD(VDD),.Y(g27350),.A(g10217),.B(g26803));
  AND2 AND2_1091(.VSS(VSS),.VDD(VDD),.Y(g18663),.A(g4311),.B(g17367));
  AND2 AND2_1092(.VSS(VSS),.VDD(VDD),.Y(g24606),.A(g5489),.B(g23630));
  AND2 AND2_1093(.VSS(VSS),.VDD(VDD),.Y(g25976),.A(g9443),.B(g25000));
  AND2 AND2_1094(.VSS(VSS),.VDD(VDD),.Y(g24303),.A(g4369),.B(g22228));
  AND2 AND2_1095(.VSS(VSS),.VDD(VDD),.Y(g16670),.A(g5953),.B(g14999));
  AND2 AND2_1096(.VSS(VSS),.VDD(VDD),.Y(g27820),.A(g7670),.B(g25932));
  AND2 AND2_1097(.VSS(VSS),.VDD(VDD),.Y(g34525),.A(g34297),.B(g19528));
  AND4 AND4_75(.VSS(VSS),.VDD(VDD),.Y(g28141),.A(g10831),.B(g11797),.C(g11261),.D(g27163));
  AND2 AND2_1098(.VSS(VSS),.VDD(VDD),.Y(g34488),.A(g34417),.B(g18988));
  AND2 AND2_1099(.VSS(VSS),.VDD(VDD),.Y(g28652),.A(g27282),.B(g10288));
  AND2 AND2_1100(.VSS(VSS),.VDD(VDD),.Y(g13493),.A(g9880),.B(g11866));
  AND3 AND3_66(.VSS(VSS),.VDD(VDD),.Y(g25374),.A(g5366),.B(g23789),.C(I24527));
  AND2 AND2_1101(.VSS(VSS),.VDD(VDD),.Y(g31943),.A(g4717),.B(g30614));
  AND3 AND3_67(.VSS(VSS),.VDD(VDD),.Y(I24505),.A(g9607),.B(g9229),.C(g5057));
  AND2 AND2_1102(.VSS(VSS),.VDD(VDD),.Y(g21729),.A(g3021),.B(g20330));
  AND2 AND2_1103(.VSS(VSS),.VDD(VDD),.Y(g26610),.A(g14198),.B(g24405));
  AND2 AND2_1104(.VSS(VSS),.VDD(VDD),.Y(g33339),.A(g32221),.B(g20634));
  AND2 AND2_1105(.VSS(VSS),.VDD(VDD),.Y(g33943),.A(g33384),.B(g21609));
  AND2 AND2_1106(.VSS(VSS),.VDD(VDD),.Y(g31296),.A(g30119),.B(g27779));
  AND2 AND2_1107(.VSS(VSS),.VDD(VDD),.Y(g34558),.A(g34353),.B(g20578));
  AND2 AND2_1108(.VSS(VSS),.VDD(VDD),.Y(g16734),.A(g5961),.B(g14735));
  AND2 AND2_1109(.VSS(VSS),.VDD(VDD),.Y(g23577),.A(g19444),.B(g13033));
  AND2 AND2_1110(.VSS(VSS),.VDD(VDD),.Y(g18483),.A(g2453),.B(g15426));
  AND2 AND2_1111(.VSS(VSS),.VDD(VDD),.Y(g24750),.A(g17662),.B(g22472));
  AND2 AND2_1112(.VSS(VSS),.VDD(VDD),.Y(g32334),.A(g31375),.B(g23568));
  AND2 AND2_1113(.VSS(VSS),.VDD(VDD),.Y(g21728),.A(g3010),.B(g20330));
  AND2 AND2_1114(.VSS(VSS),.VDD(VDD),.Y(g33338),.A(g32220),.B(g20633));
  AND2 AND2_1115(.VSS(VSS),.VDD(VDD),.Y(g28263),.A(g23747),.B(g27711));
  AND2 AND2_1116(.VSS(VSS),.VDD(VDD),.Y(g16930),.A(g239),.B(g13132));
  AND2 AND2_1117(.VSS(VSS),.VDD(VDD),.Y(g23439),.A(g13771),.B(g20452));
  AND2 AND2_1118(.VSS(VSS),.VDD(VDD),.Y(g11035),.A(g5441),.B(g9800));
  AND2 AND2_1119(.VSS(VSS),.VDD(VDD),.Y(g18553),.A(g2827),.B(g15277));
  AND2 AND2_1120(.VSS(VSS),.VDD(VDD),.Y(g13035),.A(g8497),.B(g11033));
  AND2 AND2_1121(.VSS(VSS),.VDD(VDD),.Y(g26270),.A(g1700),.B(g25275));
  AND2 AND2_1122(.VSS(VSS),.VDD(VDD),.Y(g31969),.A(g31189),.B(g22139));
  AND2 AND2_1123(.VSS(VSS),.VDD(VDD),.Y(g29784),.A(g28331),.B(g23247));
  AND2 AND2_1124(.VSS(VSS),.VDD(VDD),.Y(g26124),.A(g1811),.B(g25116));
  AND2 AND2_1125(.VSS(VSS),.VDD(VDD),.Y(g22920),.A(g19764),.B(g19719));
  AND2 AND2_1126(.VSS(VSS),.VDD(VDD),.Y(g16667),.A(g5268),.B(g14659));
  AND2 AND2_1127(.VSS(VSS),.VDD(VDD),.Y(g20174),.A(g5503),.B(g17754));
  AND2 AND2_1128(.VSS(VSS),.VDD(VDD),.Y(g29376),.A(g14002),.B(g28504));
  AND2 AND2_1129(.VSS(VSS),.VDD(VDD),.Y(g27413),.A(g26576),.B(g17530));
  AND2 AND2_1130(.VSS(VSS),.VDD(VDD),.Y(g34865),.A(g16540),.B(g34836));
  AND2 AND2_1131(.VSS(VSS),.VDD(VDD),.Y(g16965),.A(g269),.B(g13140));
  AND2 AND2_1132(.VSS(VSS),.VDD(VDD),.Y(g18949),.A(g10183),.B(g17625));
  AND2 AND2_1133(.VSS(VSS),.VDD(VDD),.Y(g31968),.A(g31757),.B(g22168));
  AND2 AND2_1134(.VSS(VSS),.VDD(VDD),.Y(g18326),.A(g1664),.B(g17873));
  AND2 AND2_1135(.VSS(VSS),.VDD(VDD),.Y(g24796),.A(g7097),.B(g23714));
  AND2 AND2_1136(.VSS(VSS),.VDD(VDD),.Y(g11142),.A(g6381),.B(g10207));
  AND2 AND2_1137(.VSS(VSS),.VDD(VDD),.Y(g27691),.A(g25778),.B(g23609));
  AND4 AND4_76(.VSS(VSS),.VDD(VDD),.Y(g17724),.A(g11547),.B(g11592),.C(g11640),.D(I18713));
  AND2 AND2_1138(.VSS(VSS),.VDD(VDD),.Y(g29354),.A(g4961),.B(g28421));
  AND4 AND4_77(.VSS(VSS),.VDD(VDD),.Y(I27533),.A(g21143),.B(g24125),.C(g24126),.D(g24127));
  AND2 AND2_1139(.VSS(VSS),.VDD(VDD),.Y(g18536),.A(g2748),.B(g15277));
  AND2 AND2_1140(.VSS(VSS),.VDD(VDD),.Y(g23349),.A(g13662),.B(g20182));
  AND2 AND2_1141(.VSS(VSS),.VDD(VDD),.Y(g22121),.A(g6593),.B(g19277));
  AND2 AND2_1142(.VSS(VSS),.VDD(VDD),.Y(g29888),.A(g28418),.B(g23352));
  AND2 AND2_1143(.VSS(VSS),.VDD(VDD),.Y(g33855),.A(g33265),.B(g20441));
  AND2 AND2_1144(.VSS(VSS),.VDD(VDD),.Y(g14206),.A(g8655),.B(g11790));
  AND2 AND2_1145(.VSS(VSS),.VDD(VDD),.Y(g21906),.A(g5022),.B(g21468));
  AND2 AND2_1146(.VSS(VSS),.VDD(VDD),.Y(g18702),.A(g15133),.B(g16856));
  AND2 AND2_1147(.VSS(VSS),.VDD(VDD),.Y(g21348),.A(g10121),.B(g17625));
  AND2 AND2_1148(.VSS(VSS),.VDD(VDD),.Y(g18757),.A(g5352),.B(g15595));
  AND2 AND2_1149(.VSS(VSS),.VDD(VDD),.Y(g31527),.A(g7553),.B(g29343));
  AND2 AND2_1150(.VSS(VSS),.VDD(VDD),.Y(g23083),.A(g16076),.B(g19878));
  AND2 AND2_1151(.VSS(VSS),.VDD(VDD),.Y(g23348),.A(g15570),.B(g21393));
  AND2 AND2_1152(.VSS(VSS),.VDD(VDD),.Y(g15076),.A(g2130),.B(g12955));
  AND2 AND2_1153(.VSS(VSS),.VDD(VDD),.Y(g33870),.A(g33280),.B(g20545));
  AND2 AND2_1154(.VSS(VSS),.VDD(VDD),.Y(g33411),.A(g32361),.B(g21410));
  AND3 AND3_68(.VSS(VSS),.VDD(VDD),.Y(g33527),.A(g32939),.B(I31331),.C(I31332));
  AND2 AND2_1155(.VSS(VSS),.VDD(VDD),.Y(g26294),.A(g4245),.B(g25230));
  AND4 AND4_78(.VSS(VSS),.VDD(VDD),.Y(I31321),.A(g31376),.B(g31852),.C(g32919),.D(g32920));
  AND2 AND2_1156(.VSS(VSS),.VDD(VDD),.Y(g16619),.A(g6629),.B(g14947));
  AND2 AND2_1157(.VSS(VSS),.VDD(VDD),.Y(g30042),.A(g29142),.B(g12601));
  AND2 AND2_1158(.VSS(VSS),.VDD(VDD),.Y(g18252),.A(g990),.B(g16897));
  AND2 AND2_1159(.VSS(VSS),.VDD(VDD),.Y(g18621),.A(g3476),.B(g17062));
  AND2 AND2_1160(.VSS(VSS),.VDD(VDD),.Y(g25559),.A(g13004),.B(g22649));
  AND2 AND2_1161(.VSS(VSS),.VDD(VDD),.Y(g30255),.A(g28748),.B(g23946));
  AND3 AND3_69(.VSS(VSS),.VDD(VDD),.Y(g25488),.A(g6404),.B(g23865),.C(I24603));
  AND4 AND4_79(.VSS(VSS),.VDD(VDD),.Y(g28833),.A(g21434),.B(g26424),.C(g25388),.D(g27469));
  AND2 AND2_1162(.VSS(VSS),.VDD(VDD),.Y(g16618),.A(g6609),.B(g15039));
  AND2 AND2_1163(.VSS(VSS),.VDD(VDD),.Y(g34679),.A(g14093),.B(g34539));
  AND2 AND2_1164(.VSS(VSS),.VDD(VDD),.Y(g18564),.A(g2844),.B(g16349));
  AND2 AND2_1165(.VSS(VSS),.VDD(VDD),.Y(g30188),.A(g28644),.B(g23841));
  AND2 AND2_1166(.VSS(VSS),.VDD(VDD),.Y(g24192),.A(g311),.B(g22722));
  AND2 AND2_1167(.VSS(VSS),.VDD(VDD),.Y(g30124),.A(g28580),.B(g21055));
  AND2 AND2_1168(.VSS(VSS),.VDD(VDD),.Y(g16279),.A(g4512),.B(g14424));
  AND2 AND2_1169(.VSS(VSS),.VDD(VDD),.Y(g34678),.A(g34490),.B(g19431));
  AND2 AND2_1170(.VSS(VSS),.VDD(VDD),.Y(g27020),.A(g4601),.B(g25852));
  AND2 AND2_1171(.VSS(VSS),.VDD(VDD),.Y(g31503),.A(g20041),.B(g29945));
  AND3 AND3_70(.VSS(VSS),.VDD(VDD),.Y(I18716),.A(g13156),.B(g11450),.C(g6756));
  AND4 AND4_80(.VSS(VSS),.VDD(VDD),.Y(I31186),.A(g31376),.B(g31828),.C(g32724),.D(g32725));
  AND3 AND3_71(.VSS(VSS),.VDD(VDD),.Y(g33503),.A(g32765),.B(I31211),.C(I31212));
  AND2 AND2_1172(.VSS(VSS),.VDD(VDD),.Y(g24663),.A(g16621),.B(g22974));
  AND2 AND2_1173(.VSS(VSS),.VDD(VDD),.Y(g33867),.A(g33277),.B(g20529));
  AND2 AND2_1174(.VSS(VSS),.VDD(VDD),.Y(g17682),.A(g9742),.B(g14637));
  AND2 AND2_1175(.VSS(VSS),.VDD(VDD),.Y(g34686),.A(g34494),.B(g19494));
  AND2 AND2_1176(.VSS(VSS),.VDD(VDD),.Y(g13523),.A(g7046),.B(g12246));
  AND2 AND2_1177(.VSS(VSS),.VDD(VDD),.Y(g18183),.A(g781),.B(g17328));
  AND2 AND2_1178(.VSS(VSS),.VDD(VDD),.Y(g18673),.A(g4643),.B(g15758));
  AND2 AND2_1179(.VSS(VSS),.VDD(VDD),.Y(g25865),.A(g25545),.B(g18991));
  AND4 AND4_81(.VSS(VSS),.VDD(VDD),.Y(g26218),.A(g25357),.B(g6856),.C(g7586),.D(g11686));
  AND2 AND2_1180(.VSS(VSS),.VDD(VDD),.Y(g18397),.A(g2004),.B(g15373));
  AND2 AND2_1181(.VSS(VSS),.VDD(VDD),.Y(g30030),.A(g29198),.B(g12347));
  AND2 AND2_1182(.VSS(VSS),.VDD(VDD),.Y(g30267),.A(g28776),.B(g23967));
  AND3 AND3_72(.VSS(VSS),.VDD(VDD),.Y(g34093),.A(g20114),.B(g33755),.C(g9104));
  AND2 AND2_1183(.VSS(VSS),.VDD(VDD),.Y(g33450),.A(g32266),.B(g29737));
  AND2 AND2_1184(.VSS(VSS),.VDD(VDD),.Y(g22760),.A(g9360),.B(g20237));
  AND2 AND2_1185(.VSS(VSS),.VDD(VDD),.Y(g22134),.A(g6653),.B(g19277));
  AND2 AND2_1186(.VSS(VSS),.VDD(VDD),.Y(g27113),.A(g25997),.B(g16522));
  AND2 AND2_1187(.VSS(VSS),.VDD(VDD),.Y(g32242),.A(g31245),.B(g20324));
  AND2 AND2_1188(.VSS(VSS),.VDD(VDD),.Y(g18509),.A(g2587),.B(g15509));
  AND2 AND2_1189(.VSS(VSS),.VDD(VDD),.Y(g22029),.A(g5901),.B(g19147));
  AND2 AND2_1190(.VSS(VSS),.VDD(VDD),.Y(g31707),.A(g30081),.B(g23886));
  AND2 AND2_1191(.VSS(VSS),.VDD(VDD),.Y(g34065),.A(g33813),.B(g23148));
  AND3 AND3_73(.VSS(VSS),.VDD(VDD),.Y(g33819),.A(g23088),.B(g33176),.C(g9104));
  AND2 AND2_1192(.VSS(VSS),.VDD(VDD),.Y(g33707),.A(g33174),.B(g13346));
  AND2 AND2_1193(.VSS(VSS),.VDD(VDD),.Y(g18933),.A(g16237),.B(g13597));
  AND2 AND2_1194(.VSS(VSS),.VDD(VDD),.Y(g33910),.A(g33134),.B(g7836));
  AND2 AND2_1195(.VSS(VSS),.VDD(VDD),.Y(g24553),.A(g22983),.B(g19539));
  AND2 AND2_1196(.VSS(VSS),.VDD(VDD),.Y(g26160),.A(g2453),.B(g25138));
  AND2 AND2_1197(.VSS(VSS),.VDD(VDD),.Y(g28273),.A(g27927),.B(g23729));
  AND2 AND2_1198(.VSS(VSS),.VDD(VDD),.Y(g7696),.A(g2955),.B(g2950));
  AND2 AND2_1199(.VSS(VSS),.VDD(VDD),.Y(g18508),.A(g2606),.B(g15509));
  AND2 AND2_1200(.VSS(VSS),.VDD(VDD),.Y(g22028),.A(g5893),.B(g19147));
  AND2 AND2_1201(.VSS(VSS),.VDD(VDD),.Y(g27302),.A(g1848),.B(g26680));
  AND2 AND2_1202(.VSS(VSS),.VDD(VDD),.Y(g18634),.A(g3813),.B(g17096));
  AND2 AND2_1203(.VSS(VSS),.VDD(VDD),.Y(g21333),.A(g1300),.B(g15740));
  AND2 AND2_1204(.VSS(VSS),.VDD(VDD),.Y(g23415),.A(g20077),.B(g20320));
  AND2 AND2_1205(.VSS(VSS),.VDD(VDD),.Y(g27357),.A(g26400),.B(g17414));
  AND2 AND2_1206(.VSS(VSS),.VDD(VDD),.Y(g25042),.A(g23262),.B(g20496));
  AND2 AND2_1207(.VSS(VSS),.VDD(VDD),.Y(g31496),.A(g2338),.B(g30312));
  AND2 AND2_1208(.VSS(VSS),.VDD(VDD),.Y(g33818),.A(g33236),.B(g20113));
  AND2 AND2_1209(.VSS(VSS),.VDD(VDD),.Y(g24949),.A(g23796),.B(g20751));
  AND3 AND3_74(.VSS(VSS),.VDD(VDD),.Y(g33496),.A(g32714),.B(I31176),.C(I31177));
  AND2 AND2_1210(.VSS(VSS),.VDD(VDD),.Y(g19461),.A(g11708),.B(g16846));
  AND2 AND2_1211(.VSS(VSS),.VDD(VDD),.Y(g27105),.A(g26026),.B(g16511));
  AND2 AND2_1212(.VSS(VSS),.VDD(VDD),.Y(g24326),.A(g4552),.B(g22228));
  AND2 AND2_1213(.VSS(VSS),.VDD(VDD),.Y(g30219),.A(g28698),.B(g23887));
  AND2 AND2_1214(.VSS(VSS),.VDD(VDD),.Y(g17134),.A(g5619),.B(g14851));
  AND2 AND2_1215(.VSS(VSS),.VDD(VDD),.Y(g21852),.A(g3909),.B(g21070));
  AND2 AND2_1216(.VSS(VSS),.VDD(VDD),.Y(g15839),.A(g3929),.B(g13990));
  AND2 AND2_1217(.VSS(VSS),.VDD(VDD),.Y(g34875),.A(g34836),.B(g20073));
  AND2 AND2_1218(.VSS(VSS),.VDD(VDD),.Y(g28812),.A(g26972),.B(g13037));
  AND2 AND2_1219(.VSS(VSS),.VDD(VDD),.Y(g33111),.A(g24005),.B(g32421));
  AND2 AND2_1220(.VSS(VSS),.VDD(VDD),.Y(g34219),.A(g33736),.B(g22942));
  AND2 AND2_1221(.VSS(VSS),.VDD(VDD),.Y(g31070),.A(g29814),.B(g25985));
  AND2 AND2_1222(.VSS(VSS),.VDD(VDD),.Y(g19145),.A(g8450),.B(g16200));
  AND2 AND2_1223(.VSS(VSS),.VDD(VDD),.Y(g24536),.A(g19516),.B(g22635));
  AND2 AND2_1224(.VSS(VSS),.VDD(VDD),.Y(g29860),.A(g28389),.B(g23312));
  AND2 AND2_1225(.VSS(VSS),.VDD(VDD),.Y(g17506),.A(g9744),.B(g14505));
  AND2 AND2_1226(.VSS(VSS),.VDD(VDD),.Y(g25124),.A(g4917),.B(g22908));
  AND2 AND2_1227(.VSS(VSS),.VDD(VDD),.Y(g15694),.A(g457),.B(g13437));
  AND2 AND2_1228(.VSS(VSS),.VDD(VDD),.Y(g15838),.A(g3602),.B(g14133));
  AND2 AND2_1229(.VSS(VSS),.VDD(VDD),.Y(g21963),.A(g5436),.B(g21514));
  AND2 AND2_1230(.VSS(VSS),.VDD(VDD),.Y(g24702),.A(g17464),.B(g22342));
  AND2 AND2_1231(.VSS(VSS),.VDD(VDD),.Y(g34218),.A(g33744),.B(g22670));
  AND2 AND2_1232(.VSS(VSS),.VDD(VDD),.Y(g24757),.A(g7004),.B(g23563));
  AND2 AND2_1233(.VSS(VSS),.VDD(VDD),.Y(g31986),.A(g31766),.B(g22197));
  AND2 AND2_1234(.VSS(VSS),.VDD(VDD),.Y(g19736),.A(g12136),.B(g17136));
  AND2 AND2_1235(.VSS(VSS),.VDD(VDD),.Y(g24904),.A(g11761),.B(g23279));
  AND2 AND2_1236(.VSS(VSS),.VDD(VDD),.Y(g28234),.A(g27877),.B(g26686));
  AND2 AND2_1237(.VSS(VSS),.VDD(VDD),.Y(g32293),.A(g2827),.B(g30593));
  AND4 AND4_82(.VSS(VSS),.VDD(VDD),.Y(I31216),.A(g30937),.B(g31834),.C(g32766),.D(g32767));
  AND2 AND2_1238(.VSS(VSS),.VDD(VDD),.Y(g25939),.A(g24583),.B(g19490));
  AND2 AND2_1239(.VSS(VSS),.VDD(VDD),.Y(g26277),.A(g2547),.B(g25400));
  AND2 AND2_1240(.VSS(VSS),.VDD(VDD),.Y(g18213),.A(g952),.B(g15979));
  AND2 AND2_1241(.VSS(VSS),.VDD(VDD),.Y(g32265),.A(g2799),.B(g30567));
  AND2 AND2_1242(.VSS(VSS),.VDD(VDD),.Y(g25030),.A(g23251),.B(g20432));
  AND2 AND2_1243(.VSS(VSS),.VDD(VDD),.Y(g25938),.A(g8997),.B(g24953));
  AND2 AND2_1244(.VSS(VSS),.VDD(VDD),.Y(g25093),.A(g12831),.B(g23493));
  AND2 AND2_1245(.VSS(VSS),.VDD(VDD),.Y(g31067),.A(g29484),.B(g22868));
  AND2 AND2_1246(.VSS(VSS),.VDD(VDD),.Y(g24564),.A(g23198),.B(g21163));
  AND2 AND2_1247(.VSS(VSS),.VDD(VDD),.Y(g29625),.A(g28514),.B(g14226));
  AND3 AND3_75(.VSS(VSS),.VDD(VDD),.Y(g29987),.A(g29197),.B(g26424),.C(g22763));
  AND2 AND2_1248(.VSS(VSS),.VDD(VDD),.Y(g19393),.A(g691),.B(g16325));
  AND2 AND2_1249(.VSS(VSS),.VDD(VDD),.Y(g16884),.A(g6159),.B(g14321));
  AND2 AND2_1250(.VSS(VSS),.VDD(VDD),.Y(g18574),.A(g2882),.B(g16349));
  AND2 AND2_1251(.VSS(VSS),.VDD(VDD),.Y(g23484),.A(g20160),.B(g20541));
  AND2 AND2_1252(.VSS(VSS),.VDD(VDD),.Y(g18452),.A(g2311),.B(g15224));
  AND2 AND2_1253(.VSS(VSS),.VDD(VDD),.Y(g18205),.A(g904),.B(g15938));
  AND2 AND2_1254(.VSS(VSS),.VDD(VDD),.Y(g31150),.A(g1682),.B(g30063));
  AND2 AND2_1255(.VSS(VSS),.VDD(VDD),.Y(g23554),.A(g20390),.B(g13024));
  AND4 AND4_83(.VSS(VSS),.VDD(VDD),.Y(I31117),.A(g32624),.B(g32625),.C(g32626),.D(g32627));
  AND2 AND2_1256(.VSS(VSS),.VDD(VDD),.Y(g18311),.A(g1554),.B(g16931));
  AND2 AND2_1257(.VSS(VSS),.VDD(VDD),.Y(g33801),.A(g33437),.B(g25327));
  AND2 AND2_1258(.VSS(VSS),.VDD(VDD),.Y(g24673),.A(g22659),.B(g19748));
  AND2 AND2_1259(.VSS(VSS),.VDD(VDD),.Y(g33735),.A(g33118),.B(g19553));
  AND2 AND2_1260(.VSS(VSS),.VDD(VDD),.Y(g33877),.A(g33287),.B(g20563));
  AND3 AND3_76(.VSS(VSS),.VDD(VDD),.Y(I24582),.A(g9809),.B(g9397),.C(g6093));
  AND2 AND2_1261(.VSS(VSS),.VDD(VDD),.Y(g30915),.A(g29886),.B(g24778));
  AND2 AND2_1262(.VSS(VSS),.VDD(VDD),.Y(g29943),.A(g2165),.B(g28765));
  AND2 AND2_1263(.VSS(VSS),.VDD(VDD),.Y(g34470),.A(g7834),.B(g34325));
  AND2 AND2_1264(.VSS(VSS),.VDD(VDD),.Y(g16666),.A(g5200),.B(g14794));
  AND2 AND2_1265(.VSS(VSS),.VDD(VDD),.Y(g25875),.A(g8390),.B(g24809));
  AND2 AND2_1266(.VSS(VSS),.VDD(VDD),.Y(g31019),.A(g29481),.B(g22856));
  AND3 AND3_77(.VSS(VSS),.VDD(VDD),.Y(I18765),.A(g13156),.B(g11450),.C(g11498));
  AND2 AND2_1267(.VSS(VSS),.VDD(VDD),.Y(g29644),.A(g28216),.B(g19794));
  AND2 AND2_1268(.VSS(VSS),.VDD(VDD),.Y(g29338),.A(g29145),.B(g22181));
  AND2 AND2_1269(.VSS(VSS),.VDD(VDD),.Y(g30277),.A(g28817),.B(g23987));
  AND2 AND2_1270(.VSS(VSS),.VDD(VDD),.Y(g13063),.A(g8567),.B(g10808));
  AND2 AND2_1271(.VSS(VSS),.VDD(VDD),.Y(g31018),.A(g29480),.B(g22855));
  AND2 AND2_1272(.VSS(VSS),.VDD(VDD),.Y(g32014),.A(g8715),.B(g30673));
  AND2 AND2_1273(.VSS(VSS),.VDD(VDD),.Y(g29969),.A(g28121),.B(g20509));
  AND2 AND2_1274(.VSS(VSS),.VDD(VDD),.Y(g30075),.A(g28525),.B(g20662));
  AND2 AND2_1275(.VSS(VSS),.VDD(VDD),.Y(g26155),.A(g1945),.B(g25134));
  AND2 AND2_1276(.VSS(VSS),.VDD(VDD),.Y(g14221),.A(g8686),.B(g11823));
  AND2 AND2_1277(.VSS(VSS),.VDD(VDD),.Y(g21921),.A(g5109),.B(g21468));
  AND2 AND2_1278(.VSS(VSS),.VDD(VDD),.Y(g26822),.A(g24841),.B(g13116));
  AND4 AND4_84(.VSS(VSS),.VDD(VDD),.Y(I31242),.A(g32805),.B(g32806),.C(g32807),.D(g32808));
  AND4 AND4_85(.VSS(VSS),.VDD(VDD),.Y(g16486),.A(g6772),.B(g11592),.C(g6789),.D(I17692));
  AND2 AND2_1279(.VSS(VSS),.VDD(VDD),.Y(g18592),.A(g2994),.B(g16349));
  AND2 AND2_1280(.VSS(VSS),.VDD(VDD),.Y(g23921),.A(g19379),.B(g4146));
  AND2 AND2_1281(.VSS(VSS),.VDD(VDD),.Y(g18756),.A(g5348),.B(g15595));
  AND2 AND2_1282(.VSS(VSS),.VDD(VDD),.Y(g34075),.A(g33692),.B(g19517));
  AND2 AND2_1283(.VSS(VSS),.VDD(VDD),.Y(g31526),.A(g22521),.B(g29342));
  AND2 AND2_1284(.VSS(VSS),.VDD(VDD),.Y(g24634),.A(g22634),.B(g19685));
  AND2 AND2_1285(.VSS(VSS),.VDD(VDD),.Y(g30595),.A(g18911),.B(g29847));
  AND3 AND3_78(.VSS(VSS),.VDD(VDD),.Y(g33526),.A(g32932),.B(I31326),.C(I31327));
  AND2 AND2_1286(.VSS(VSS),.VDD(VDD),.Y(g24872),.A(g23088),.B(g9104));
  AND2 AND2_1287(.VSS(VSS),.VDD(VDD),.Y(g29968),.A(g2433),.B(g28843));
  AND2 AND2_1288(.VSS(VSS),.VDD(VDD),.Y(g21745),.A(g3017),.B(g20330));
  AND2 AND2_1289(.VSS(VSS),.VDD(VDD),.Y(g18780),.A(g5827),.B(g18065));
  AND2 AND2_1290(.VSS(VSS),.VDD(VDD),.Y(g12027),.A(g9499),.B(g9729));
  AND2 AND2_1291(.VSS(VSS),.VDD(VDD),.Y(g14613),.A(g10602),.B(g10585));
  AND2 AND2_1292(.VSS(VSS),.VDD(VDD),.Y(g27249),.A(g25929),.B(g19678));
  AND2 AND2_1293(.VSS(VSS),.VDD(VDD),.Y(g21799),.A(g3530),.B(g20924));
  AND2 AND2_1294(.VSS(VSS),.VDD(VDD),.Y(g29855),.A(g2287),.B(g29093));
  AND2 AND2_1295(.VSS(VSS),.VDD(VDD),.Y(g17770),.A(g7863),.B(g13189));
  AND2 AND2_1296(.VSS(VSS),.VDD(VDD),.Y(g21813),.A(g3590),.B(g20924));
  AND2 AND2_1297(.VSS(VSS),.VDD(VDD),.Y(g23799),.A(g14911),.B(g21279));
  AND2 AND2_1298(.VSS(VSS),.VDD(VDD),.Y(g27482),.A(g26488),.B(g17641));
  AND2 AND2_1299(.VSS(VSS),.VDD(VDD),.Y(g15815),.A(g3594),.B(g14075));
  AND2 AND2_1300(.VSS(VSS),.VDD(VDD),.Y(g28541),.A(g27403),.B(g20274));
  AND2 AND2_1301(.VSS(VSS),.VDD(VDD),.Y(g10947),.A(g9200),.B(g1430));
  AND2 AND2_1302(.VSS(VSS),.VDD(VDD),.Y(g18350),.A(g1779),.B(g17955));
  AND3 AND3_79(.VSS(VSS),.VDD(VDD),.Y(I24603),.A(g9892),.B(g9467),.C(g6439));
  AND2 AND2_1303(.VSS(VSS),.VDD(VDD),.Y(g33402),.A(g32351),.B(g21395));
  AND2 AND2_1304(.VSS(VSS),.VDD(VDD),.Y(g29870),.A(g2421),.B(g29130));
  AND2 AND2_1305(.VSS(VSS),.VDD(VDD),.Y(g29527),.A(g28945),.B(g22432));
  AND2 AND2_1306(.VSS(VSS),.VDD(VDD),.Y(g27710),.A(g26422),.B(g20904));
  AND2 AND2_1307(.VSS(VSS),.VDD(VDD),.Y(g21798),.A(g3522),.B(g20924));
  AND2 AND2_1308(.VSS(VSS),.VDD(VDD),.Y(g34782),.A(g34711),.B(g33888));
  AND4 AND4_86(.VSS(VSS),.VDD(VDD),.Y(I27529),.A(g28038),.B(g24121),.C(g24122),.D(g24123));
  AND2 AND2_1309(.VSS(VSS),.VDD(VDD),.Y(g18820),.A(g15166),.B(g15563));
  AND2 AND2_1310(.VSS(VSS),.VDD(VDD),.Y(g26853),.A(g94),.B(g24533));
  AND4 AND4_87(.VSS(VSS),.VDD(VDD),.Y(g28789),.A(g21434),.B(g26424),.C(g25340),.D(g27440));
  AND2 AND2_1311(.VSS(VSS),.VDD(VDD),.Y(g21973),.A(g5511),.B(g19074));
  AND2 AND2_1312(.VSS(VSS),.VDD(VDD),.Y(g32116),.A(g31658),.B(g29929));
  AND2 AND2_1313(.VSS(VSS),.VDD(VDD),.Y(g27204),.A(g26026),.B(g16689));
  AND2 AND2_1314(.VSS(VSS),.VDD(VDD),.Y(g33866),.A(g33276),.B(g20528));
  AND2 AND2_1315(.VSS(VSS),.VDD(VDD),.Y(g22899),.A(g19486),.B(g19695));
  AND2 AND2_1316(.VSS(VSS),.VDD(VDD),.Y(g21805),.A(g3550),.B(g20924));
  AND2 AND2_1317(.VSS(VSS),.VDD(VDD),.Y(g22990),.A(g19555),.B(g19760));
  AND4 AND4_88(.VSS(VSS),.VDD(VDD),.Y(I27528),.A(g20998),.B(g24118),.C(g24119),.D(g24120));
  AND2 AND2_1318(.VSS(VSS),.VDD(VDD),.Y(g18152),.A(g613),.B(g17533));
  AND2 AND2_1319(.VSS(VSS),.VDD(VDD),.Y(g25915),.A(g24926),.B(g9602));
  AND2 AND2_1320(.VSS(VSS),.VDD(VDD),.Y(g32041),.A(g13913),.B(g31262));
  AND2 AND2_1321(.VSS(VSS),.VDD(VDD),.Y(g18396),.A(g2008),.B(g15373));
  AND2 AND2_1322(.VSS(VSS),.VDD(VDD),.Y(g22633),.A(g19359),.B(g19479));
  AND4 AND4_89(.VSS(VSS),.VDD(VDD),.Y(g17767),.A(g6772),.B(g11592),.C(g6789),.D(I18765));
  AND2 AND2_1323(.VSS(VSS),.VDD(VDD),.Y(g18731),.A(g15140),.B(g16861));
  AND2 AND2_1324(.VSS(VSS),.VDD(VDD),.Y(g30266),.A(g28775),.B(g23966));
  AND2 AND2_1325(.VSS(VSS),.VDD(VDD),.Y(g28535),.A(g11981),.B(g27088));
  AND2 AND2_1326(.VSS(VSS),.VDD(VDD),.Y(g15937),.A(g11950),.B(g14387));
  AND2 AND2_1327(.VSS(VSS),.VDD(VDD),.Y(g25201),.A(g12346),.B(g23665));
  AND2 AND2_1328(.VSS(VSS),.VDD(VDD),.Y(g22191),.A(g8119),.B(g19875));
  AND2 AND2_1329(.VSS(VSS),.VDD(VDD),.Y(g16179),.A(g6187),.B(g14321));
  AND2 AND2_1330(.VSS(VSS),.VDD(VDD),.Y(g29867),.A(g1996),.B(g29117));
  AND2 AND2_1331(.VSS(VSS),.VDD(VDD),.Y(g29894),.A(g2070),.B(g29169));
  AND2 AND2_1332(.VSS(VSS),.VDD(VDD),.Y(g19069),.A(g8397),.B(g16186));
  AND2 AND2_1333(.VSS(VSS),.VDD(VDD),.Y(g21732),.A(g3004),.B(g20330));
  AND2 AND2_1334(.VSS(VSS),.VDD(VDD),.Y(g16531),.A(g5232),.B(g14656));
  AND2 AND2_1335(.VSS(VSS),.VDD(VDD),.Y(g13542),.A(g10053),.B(g11927));
  AND2 AND2_1336(.VSS(VSS),.VDD(VDD),.Y(g21934),.A(g5220),.B(g18997));
  AND2 AND2_1337(.VSS(VSS),.VDD(VDD),.Y(g18413),.A(g2089),.B(g15373));
  AND2 AND2_1338(.VSS(VSS),.VDD(VDD),.Y(g24912),.A(g23687),.B(g20682));
  AND2 AND2_1339(.VSS(VSS),.VDD(VDD),.Y(g26119),.A(g11944),.B(g25109));
  AND2 AND2_1340(.VSS(VSS),.VDD(VDD),.Y(g24311),.A(g4498),.B(g22228));
  AND2 AND2_1341(.VSS(VSS),.VDD(VDD),.Y(g16178),.A(g5845),.B(g14297));
  AND2 AND2_1342(.VSS(VSS),.VDD(VDD),.Y(g18691),.A(g4727),.B(g16053));
  AND2 AND2_1343(.VSS(VSS),.VDD(VDD),.Y(g15884),.A(g3901),.B(g14113));
  AND2 AND2_1344(.VSS(VSS),.VDD(VDD),.Y(g33689),.A(g33144),.B(g11006));
  AND2 AND2_1345(.VSS(VSS),.VDD(VDD),.Y(g32340),.A(g31468),.B(g23585));
  AND2 AND2_1346(.VSS(VSS),.VDD(VDD),.Y(g29581),.A(g28462),.B(g11796));
  AND2 AND2_1347(.VSS(VSS),.VDD(VDD),.Y(g32035),.A(g4176),.B(g30937));
  AND2 AND2_1348(.VSS(VSS),.VDD(VDD),.Y(g31280),.A(g29717),.B(g23305));
  AND2 AND2_1349(.VSS(VSS),.VDD(VDD),.Y(g17191),.A(g1384),.B(g13242));
  AND2 AND2_1350(.VSS(VSS),.VDD(VDD),.Y(g17719),.A(g9818),.B(g14675));
  AND2 AND2_1351(.VSS(VSS),.VDD(VDD),.Y(g21761),.A(g3215),.B(g20785));
  AND3 AND3_80(.VSS(VSS),.VDD(VDD),.Y(g29315),.A(g29188),.B(g7051),.C(g5990));
  AND4 AND4_90(.VSS(VSS),.VDD(VDD),.Y(g27999),.A(g23032),.B(g26200),.C(g26424),.D(g25529));
  AND2 AND2_1352(.VSS(VSS),.VDD(VDD),.Y(g26864),.A(g2907),.B(g24548));
  AND2 AND2_1353(.VSS(VSS),.VDD(VDD),.Y(g26022),.A(g25271),.B(g20751));
  AND2 AND2_1354(.VSS(VSS),.VDD(VDD),.Y(g13436),.A(g9721),.B(g11811));
  AND2 AND2_1355(.VSS(VSS),.VDD(VDD),.Y(g18405),.A(g2040),.B(g15373));
  AND2 AND2_1356(.VSS(VSS),.VDD(VDD),.Y(g31300),.A(g30148),.B(g27858));
  AND2 AND2_1357(.VSS(VSS),.VDD(VDD),.Y(g30167),.A(g28622),.B(g23793));
  AND2 AND2_1358(.VSS(VSS),.VDD(VDD),.Y(g30194),.A(g28651),.B(g23849));
  AND2 AND2_1359(.VSS(VSS),.VDD(VDD),.Y(g30589),.A(g18898),.B(g29811));
  AND4 AND4_91(.VSS(VSS),.VDD(VDD),.Y(I24690),.A(g24043),.B(g24044),.C(g24045),.D(g24046));
  AND3 AND3_81(.VSS(VSS),.VDD(VDD),.Y(I24549),.A(g5385),.B(g5390),.C(g9792));
  AND2 AND2_1360(.VSS(VSS),.VDD(VDD),.Y(g26749),.A(g24494),.B(g23578));
  AND2 AND2_1361(.VSS(VSS),.VDD(VDD),.Y(g27090),.A(g25997),.B(g16423));
  AND3 AND3_82(.VSS(VSS),.VDD(VDD),.Y(g29202),.A(g24088),.B(I27508),.C(I27509));
  AND2 AND2_1362(.VSS(VSS),.VDD(VDD),.Y(g25782),.A(g2936),.B(g24571));
  AND2 AND2_1363(.VSS(VSS),.VDD(VDD),.Y(g32142),.A(g31616),.B(g29965));
  AND2 AND2_1364(.VSS(VSS),.VDD(VDD),.Y(g13320),.A(g417),.B(g11048));
  AND2 AND2_1365(.VSS(VSS),.VDD(VDD),.Y(g26313),.A(g12645),.B(g25326));
  AND3 AND3_83(.VSS(VSS),.VDD(VDD),.Y(g28291),.A(g7411),.B(g2070),.C(g27469));
  AND2 AND2_1366(.VSS(VSS),.VDD(VDD),.Y(g29979),.A(g23655),.B(g28991));
  AND2 AND2_1367(.VSS(VSS),.VDD(VDD),.Y(g34588),.A(g26082),.B(g34323));
  AND2 AND2_1368(.VSS(VSS),.VDD(VDD),.Y(g22861),.A(g19792),.B(g19670));
  AND2 AND2_1369(.VSS(VSS),.VDD(VDD),.Y(g27651),.A(g22448),.B(g25781));
  AND2 AND2_1370(.VSS(VSS),.VDD(VDD),.Y(g34524),.A(g9083),.B(g34359));
  AND2 AND2_1371(.VSS(VSS),.VDD(VDD),.Y(g33102),.A(g32399),.B(g18978));
  AND4 AND4_92(.VSS(VSS),.VDD(VDD),.Y(I31007),.A(g32466),.B(g32467),.C(g32468),.D(g32469));
  AND2 AND2_1372(.VSS(VSS),.VDD(VDD),.Y(g26276),.A(g2461),.B(g25476));
  AND2 AND2_1373(.VSS(VSS),.VDD(VDD),.Y(g26285),.A(g1834),.B(g25300));
  AND2 AND2_1374(.VSS(VSS),.VDD(VDD),.Y(g34401),.A(g34199),.B(g21383));
  AND2 AND2_1375(.VSS(VSS),.VDD(VDD),.Y(g34477),.A(g26344),.B(g34328));
  AND2 AND2_1376(.VSS(VSS),.VDD(VDD),.Y(g22045),.A(g6069),.B(g21611));
  AND2 AND2_1377(.VSS(VSS),.VDD(VDD),.Y(g18583),.A(g2936),.B(g16349));
  AND2 AND2_1378(.VSS(VSS),.VDD(VDD),.Y(g29590),.A(g2625),.B(g28615));
  AND3 AND3_84(.VSS(VSS),.VDD(VDD),.Y(g34119),.A(g20516),.B(g9104),.C(g33755));
  AND2 AND2_1379(.VSS(VSS),.VDD(VDD),.Y(g26254),.A(g2413),.B(g25349));
  AND2 AND2_1380(.VSS(VSS),.VDD(VDD),.Y(g31066),.A(g29483),.B(g22865));
  AND2 AND2_1381(.VSS(VSS),.VDD(VDD),.Y(g31231),.A(g30290),.B(g25239));
  AND2 AND2_1382(.VSS(VSS),.VDD(VDD),.Y(g29986),.A(g28468),.B(g23473));
  AND2 AND2_1383(.VSS(VSS),.VDD(VDD),.Y(g22099),.A(g6462),.B(g18833));
  AND2 AND2_1384(.VSS(VSS),.VDD(VDD),.Y(g27932),.A(g25944),.B(g19369));
  AND2 AND2_1385(.VSS(VSS),.VDD(VDD),.Y(g27331),.A(g10177),.B(g26754));
  AND2 AND2_1386(.VSS(VSS),.VDD(VDD),.Y(g30118),.A(g28574),.B(g21050));
  AND2 AND2_1387(.VSS(VSS),.VDD(VDD),.Y(g24820),.A(g13944),.B(g23978));
  AND2 AND2_1388(.VSS(VSS),.VDD(VDD),.Y(g26808),.A(g25521),.B(g21185));
  AND2 AND2_1389(.VSS(VSS),.VDD(VDD),.Y(g16762),.A(g5901),.B(g14930));
  AND2 AND2_1390(.VSS(VSS),.VDD(VDD),.Y(g20152),.A(g11545),.B(g16727));
  AND2 AND2_1391(.VSS(VSS),.VDD(VDD),.Y(g22534),.A(g8766),.B(g21389));
  AND3 AND3_85(.VSS(VSS),.VDD(VDD),.Y(g29384),.A(g26424),.B(g22763),.C(g28179));
  AND2 AND2_1392(.VSS(VSS),.VDD(VDD),.Y(g22098),.A(g6459),.B(g18833));
  AND2 AND2_1393(.VSS(VSS),.VDD(VDD),.Y(g32193),.A(g30732),.B(g25410));
  AND4 AND4_93(.VSS(VSS),.VDD(VDD),.Y(I31116),.A(g31154),.B(g31816),.C(g32622),.D(g32623));
  AND3 AND3_86(.VSS(VSS),.VDD(VDD),.Y(g24846),.A(g3361),.B(g23555),.C(I24018));
  AND2 AND2_1394(.VSS(VSS),.VDD(VDD),.Y(g26101),.A(g1760),.B(g25098));
  AND2 AND2_1395(.VSS(VSS),.VDD(VDD),.Y(g33876),.A(g33286),.B(g20562));
  AND2 AND2_1396(.VSS(VSS),.VDD(VDD),.Y(g33885),.A(g33296),.B(g20609));
  AND2 AND2_1397(.VSS(VSS),.VDD(VDD),.Y(g26177),.A(g2079),.B(g25154));
  AND2 AND2_1398(.VSS(VSS),.VDD(VDD),.Y(g18113),.A(g405),.B(g17015));
  AND2 AND2_1399(.VSS(VSS),.VDD(VDD),.Y(g18787),.A(g15158),.B(g15634));
  AND2 AND2_1400(.VSS(VSS),.VDD(VDD),.Y(g32165),.A(g31669),.B(g27742));
  AND2 AND2_1401(.VSS(VSS),.VDD(VDD),.Y(g24731),.A(g6519),.B(g23733));
  AND4 AND4_94(.VSS(VSS),.VDD(VDD),.Y(I31041),.A(g31566),.B(g31803),.C(g32513),.D(g32514));
  AND2 AND2_1402(.VSS(VSS),.VDD(VDD),.Y(g18282),.A(g1379),.B(g16136));
  AND2 AND2_1403(.VSS(VSS),.VDD(VDD),.Y(g34748),.A(g34672),.B(g19529));
  AND2 AND2_1404(.VSS(VSS),.VDD(VDD),.Y(g27505),.A(g26519),.B(g17681));
  AND2 AND2_1405(.VSS(VSS),.VDD(VDD),.Y(g27404),.A(g26400),.B(g17518));
  AND2 AND2_1406(.VSS(VSS),.VDD(VDD),.Y(g31763),.A(g30127),.B(g23965));
  AND2 AND2_1407(.VSS(VSS),.VDD(VDD),.Y(g18302),.A(g1514),.B(g16489));
  AND3 AND3_87(.VSS(VSS),.VDD(VDD),.Y(g33511),.A(g32823),.B(I31251),.C(I31252));
  AND2 AND2_1408(.VSS(VSS),.VDD(VDD),.Y(g15084),.A(g2710),.B(g12983));
  AND2 AND2_1409(.VSS(VSS),.VDD(VDD),.Y(g18357),.A(g1816),.B(g17955));
  AND2 AND2_1410(.VSS(VSS),.VDD(VDD),.Y(g19545),.A(g3147),.B(g16769));
  AND2 AND2_1411(.VSS(VSS),.VDD(VDD),.Y(g29877),.A(g28405),.B(g23340));
  AND2 AND2_1412(.VSS(VSS),.VDD(VDD),.Y(g15110),.A(g4245),.B(g14454));
  AND2 AND2_1413(.VSS(VSS),.VDD(VDD),.Y(g18105),.A(g417),.B(g17015));
  AND2 AND2_1414(.VSS(VSS),.VDD(VDD),.Y(g10724),.A(g3689),.B(g8728));
  AND2 AND2_1415(.VSS(VSS),.VDD(VDD),.Y(g22032),.A(g5921),.B(g19147));
  AND2 AND2_1416(.VSS(VSS),.VDD(VDD),.Y(g30254),.A(g28747),.B(g23944));
  AND2 AND2_1417(.VSS(VSS),.VDD(VDD),.Y(g18743),.A(g5115),.B(g17847));
  AND2 AND2_1418(.VSS(VSS),.VDD(VDD),.Y(g27212),.A(g25997),.B(g16717));
  AND2 AND2_1419(.VSS(VSS),.VDD(VDD),.Y(g10829),.A(g7289),.B(g4375));
  AND4 AND4_95(.VSS(VSS),.VDD(VDD),.Y(I31237),.A(g32798),.B(g32799),.C(g32800),.D(g32801));
  AND2 AND2_1420(.VSS(VSS),.VDD(VDD),.Y(g21771),.A(g3255),.B(g20785));
  AND2 AND2_1421(.VSS(VSS),.VDD(VDD),.Y(g10828),.A(g6888),.B(g7640));
  AND2 AND2_1422(.VSS(VSS),.VDD(VDD),.Y(g18640),.A(g3835),.B(g17096));
  AND2 AND2_1423(.VSS(VSS),.VDD(VDD),.Y(g18769),.A(g15151),.B(g18062));
  AND2 AND2_1424(.VSS(VSS),.VDD(VDD),.Y(g22061),.A(g6065),.B(g21611));
  AND2 AND2_1425(.VSS(VSS),.VDD(VDD),.Y(g30101),.A(g28551),.B(g20780));
  AND2 AND2_1426(.VSS(VSS),.VDD(VDD),.Y(g30177),.A(g28631),.B(g23814));
  AND2 AND2_1427(.VSS(VSS),.VDD(VDD),.Y(g29526),.A(g28938),.B(g22384));
  AND2 AND2_1428(.VSS(VSS),.VDD(VDD),.Y(g17140),.A(g8616),.B(g12968));
  AND2 AND2_1429(.VSS(VSS),.VDD(VDD),.Y(g26630),.A(g7592),.B(g24419));
  AND2 AND2_1430(.VSS(VSS),.VDD(VDD),.Y(g34560),.A(g34366),.B(g17366));
  AND2 AND2_1431(.VSS(VSS),.VDD(VDD),.Y(g18768),.A(g5503),.B(g17929));
  AND2 AND2_1432(.VSS(VSS),.VDD(VDD),.Y(g18803),.A(g15161),.B(g15480));
  AND2 AND2_1433(.VSS(VSS),.VDD(VDD),.Y(g31480),.A(g1644),.B(g30296));
  AND4 AND4_96(.VSS(VSS),.VDD(VDD),.Y(I31142),.A(g32661),.B(g32662),.C(g32663),.D(g32664));
  AND3 AND3_88(.VSS(VSS),.VDD(VDD),.Y(g33480),.A(g32600),.B(I31096),.C(I31097));
  AND2 AND2_1434(.VSS(VSS),.VDD(VDD),.Y(g24929),.A(g23751),.B(g20875));
  AND2 AND2_1435(.VSS(VSS),.VDD(VDD),.Y(g22871),.A(g9523),.B(g20871));
  AND4 AND4_97(.VSS(VSS),.VDD(VDD),.Y(g26166),.A(g25357),.B(g11724),.C(g11709),.D(g7558));
  AND2 AND2_1436(.VSS(VSS),.VDD(VDD),.Y(g27723),.A(g26512),.B(g21049));
  AND2 AND2_1437(.VSS(VSS),.VDD(VDD),.Y(g15654),.A(g3845),.B(g13584));
  AND2 AND2_1438(.VSS(VSS),.VDD(VDD),.Y(g31314),.A(g30183),.B(g27937));
  AND2 AND2_1439(.VSS(VSS),.VDD(VDD),.Y(g28240),.A(g27356),.B(g17239));
  AND2 AND2_1440(.VSS(VSS),.VDD(VDD),.Y(g27149),.A(g25997),.B(g16623));
  AND2 AND2_1441(.VSS(VSS),.VDD(VDD),.Y(g30064),.A(g28517),.B(g20630));
  AND4 AND4_98(.VSS(VSS),.VDD(VDD),.Y(g17766),.A(g6772),.B(g11592),.C(g11640),.D(I18762));
  AND2 AND2_1442(.VSS(VSS),.VDD(VDD),.Y(g27433),.A(g26519),.B(g17583));
  AND2 AND2_1443(.VSS(VSS),.VDD(VDD),.Y(g27387),.A(g26488),.B(g17499));
  AND2 AND2_1444(.VSS(VSS),.VDD(VDD),.Y(g15936),.A(g475),.B(g13999));
  AND2 AND2_1445(.VSS(VSS),.VDD(VDD),.Y(g25285),.A(g22152),.B(g13061));
  AND2 AND2_1446(.VSS(VSS),.VDD(VDD),.Y(g29866),.A(g1906),.B(g29116));
  AND2 AND2_1447(.VSS(VSS),.VDD(VDD),.Y(g27148),.A(g25997),.B(g16622));
  AND2 AND2_1448(.VSS(VSS),.VDD(VDD),.Y(g21882),.A(g4057),.B(g19801));
  AND2 AND2_1449(.VSS(VSS),.VDD(VDD),.Y(g21991),.A(g5595),.B(g19074));
  AND2 AND2_1450(.VSS(VSS),.VDD(VDD),.Y(g26485),.A(g24968),.B(g10502));
  AND2 AND2_1451(.VSS(VSS),.VDD(VDD),.Y(g23991),.A(g19209),.B(g21428));
  AND2 AND2_1452(.VSS(VSS),.VDD(VDD),.Y(g27097),.A(g25867),.B(g22526));
  AND2 AND2_1453(.VSS(VSS),.VDD(VDD),.Y(g33721),.A(g33163),.B(g19440));
  AND2 AND2_1454(.VSS(VSS),.VDD(VDD),.Y(g19656),.A(g2807),.B(g15844));
  AND2 AND2_1455(.VSS(VSS),.VDD(VDD),.Y(g27104),.A(g25997),.B(g16510));
  AND2 AND2_1456(.VSS(VSS),.VDD(VDD),.Y(g16751),.A(g13155),.B(g13065));
  AND2 AND2_1457(.VSS(VSS),.VDD(VDD),.Y(g16807),.A(g6585),.B(g14978));
  AND2 AND2_1458(.VSS(VSS),.VDD(VDD),.Y(g27646),.A(g13094),.B(g25773));
  AND2 AND2_1459(.VSS(VSS),.VDD(VDD),.Y(g25900),.A(g24390),.B(g19368));
  AND2 AND2_1460(.VSS(VSS),.VDD(VDD),.Y(g34874),.A(g34833),.B(g20060));
  AND2 AND2_1461(.VSS(VSS),.VDD(VDD),.Y(g23407),.A(g9295),.B(g20273));
  AND2 AND2_1462(.VSS(VSS),.VDD(VDD),.Y(g33243),.A(g32124),.B(g19947));
  AND2 AND2_1463(.VSS(VSS),.VDD(VDD),.Y(g28563),.A(g11981),.B(g27100));
  AND2 AND2_1464(.VSS(VSS),.VDD(VDD),.Y(g25466),.A(g23574),.B(g21346));
  AND2 AND2_1465(.VSS(VSS),.VDD(VDD),.Y(g19680),.A(g12028),.B(g17013));
  AND2 AND2_1466(.VSS(VSS),.VDD(VDD),.Y(g33431),.A(g32364),.B(g32377));
  AND2 AND2_1467(.VSS(VSS),.VDD(VDD),.Y(g16639),.A(g6291),.B(g14974));
  AND2 AND2_1468(.VSS(VSS),.VDD(VDD),.Y(g26712),.A(g24508),.B(g24463));
  AND3 AND3_89(.VSS(VSS),.VDD(VDD),.Y(I17741),.A(g14988),.B(g11450),.C(g11498));
  AND2 AND2_1469(.VSS(VSS),.VDD(VDD),.Y(g18662),.A(g15126),.B(g17367));
  AND2 AND2_1470(.VSS(VSS),.VDD(VDD),.Y(g32175),.A(g31709),.B(g27858));
  AND2 AND2_1471(.VSS(VSS),.VDD(VDD),.Y(g30166),.A(g28621),.B(g23792));
  AND2 AND2_1472(.VSS(VSS),.VDD(VDD),.Y(g30009),.A(g29034),.B(g10518));
  AND2 AND2_1473(.VSS(VSS),.VDD(VDD),.Y(g24302),.A(g15124),.B(g22228));
  AND2 AND2_1474(.VSS(VSS),.VDD(VDD),.Y(g16638),.A(g6271),.B(g14773));
  AND2 AND2_1475(.VSS(VSS),.VDD(VDD),.Y(g33269),.A(g31970),.B(g15582));
  AND2 AND2_1476(.VSS(VSS),.VDD(VDD),.Y(g34665),.A(g34583),.B(g19067));
  AND3 AND3_90(.VSS(VSS),.VDD(VDD),.Y(g22472),.A(g7753),.B(g9285),.C(g21289));
  AND2 AND2_1477(.VSS(VSS),.VDD(VDD),.Y(g18890),.A(g10158),.B(g17625));
  AND2 AND2_1478(.VSS(VSS),.VDD(VDD),.Y(g13492),.A(g9856),.B(g11865));
  AND2 AND2_1479(.VSS(VSS),.VDD(VDD),.Y(g27369),.A(g25894),.B(g25324));
  AND2 AND2_1480(.VSS(VSS),.VDD(VDD),.Y(g24743),.A(g22708),.B(g19789));
  AND2 AND2_1481(.VSS(VSS),.VDD(VDD),.Y(g30008),.A(g29191),.B(g12297));
  AND2 AND2_1482(.VSS(VSS),.VDD(VDD),.Y(g18249),.A(g1216),.B(g16897));
  AND2 AND2_1483(.VSS(VSS),.VDD(VDD),.Y(g33942),.A(g33383),.B(g21608));
  AND2 AND2_1484(.VSS(VSS),.VDD(VDD),.Y(g33341),.A(g32223),.B(g20640));
  AND2 AND2_1485(.VSS(VSS),.VDD(VDD),.Y(g18482),.A(g2472),.B(g15426));
  AND2 AND2_1486(.VSS(VSS),.VDD(VDD),.Y(g14506),.A(g1430),.B(g10755));
  AND2 AND2_1487(.VSS(VSS),.VDD(VDD),.Y(g29688),.A(g2509),.B(g28713));
  AND4 AND4_99(.VSS(VSS),.VDD(VDD),.Y(I31006),.A(g31376),.B(g31796),.C(g32464),.D(g32465));
  AND2 AND2_1488(.VSS(VSS),.VDD(VDD),.Y(g29624),.A(g28491),.B(g8070));
  AND2 AND2_1489(.VSS(VSS),.VDD(VDD),.Y(g14028),.A(g8673),.B(g11797));
  AND2 AND2_1490(.VSS(VSS),.VDD(VDD),.Y(g18248),.A(g15067),.B(g16897));
  AND2 AND2_1491(.VSS(VSS),.VDD(VDD),.Y(g16841),.A(g5913),.B(g14858));
  AND2 AND2_1492(.VSS(VSS),.VDD(VDD),.Y(g18710),.A(g15135),.B(g17302));
  AND2 AND2_1493(.VSS(VSS),.VDD(VDD),.Y(g34476),.A(g34399),.B(g18891));
  AND2 AND2_1494(.VSS(VSS),.VDD(VDD),.Y(g34485),.A(g34411),.B(g18952));
  AND2 AND2_1495(.VSS(VSS),.VDD(VDD),.Y(g18552),.A(g2815),.B(g15277));
  AND2 AND2_1496(.VSS(VSS),.VDD(VDD),.Y(g24640),.A(g6509),.B(g23733));
  AND2 AND2_1497(.VSS(VSS),.VDD(VDD),.Y(g24769),.A(g19619),.B(g23058));
  AND2 AND2_1498(.VSS(VSS),.VDD(VDD),.Y(g19631),.A(g1484),.B(g16093));
  AND2 AND2_1499(.VSS(VSS),.VDD(VDD),.Y(g18204),.A(g914),.B(g15938));
  AND4 AND4_100(.VSS(VSS),.VDD(VDD),.Y(I31222),.A(g32775),.B(g32776),.C(g32777),.D(g32778));
  AND2 AND2_1500(.VSS(VSS),.VDD(VDD),.Y(g27412),.A(g26576),.B(g17529));
  AND2 AND2_1501(.VSS(VSS),.VDD(VDD),.Y(g34555),.A(g34349),.B(g20512));
  AND2 AND2_1502(.VSS(VSS),.VDD(VDD),.Y(g18779),.A(g5821),.B(g18065));
  AND2 AND2_1503(.VSS(VSS),.VDD(VDD),.Y(g22071),.A(g6251),.B(g19210));
  AND2 AND2_1504(.VSS(VSS),.VDD(VDD),.Y(g24803),.A(g22901),.B(g20005));
  AND3 AND3_91(.VSS(VSS),.VDD(VDD),.Y(g33734),.A(g7806),.B(g33136),.C(I31593));
  AND2 AND2_1505(.VSS(VSS),.VDD(VDD),.Y(g30914),.A(g29873),.B(g20887));
  AND2 AND2_1506(.VSS(VSS),.VDD(VDD),.Y(g21759),.A(g3199),.B(g20785));
  AND2 AND2_1507(.VSS(VSS),.VDD(VDD),.Y(g15117),.A(g4300),.B(g14454));
  AND2 AND2_1508(.VSS(VSS),.VDD(VDD),.Y(g23725),.A(g14772),.B(g21138));
  AND2 AND2_1509(.VSS(VSS),.VDD(VDD),.Y(g18778),.A(g5817),.B(g18065));
  AND2 AND2_1510(.VSS(VSS),.VDD(VDD),.Y(g25874),.A(g11118),.B(g24665));
  AND2 AND2_1511(.VSS(VSS),.VDD(VDD),.Y(g27229),.A(g26055),.B(g16774));
  AND2 AND2_1512(.VSS(VSS),.VDD(VDD),.Y(g31993),.A(g31774),.B(g22214));
  AND2 AND2_1513(.VSS(VSS),.VDD(VDD),.Y(g21758),.A(g3191),.B(g20785));
  AND2 AND2_1514(.VSS(VSS),.VDD(VDD),.Y(g26176),.A(g1964),.B(g25467));
  AND2 AND2_1515(.VSS(VSS),.VDD(VDD),.Y(g26092),.A(g9766),.B(g25083));
  AND2 AND2_1516(.VSS(VSS),.VDD(VDD),.Y(g18786),.A(g15156),.B(g15345));
  AND2 AND2_1517(.VSS(VSS),.VDD(VDD),.Y(g27228),.A(g26055),.B(g16773));
  AND3 AND3_92(.VSS(VSS),.VDD(VDD),.Y(g24881),.A(g3050),.B(g23211),.C(I24048));
  AND4 AND4_101(.VSS(VSS),.VDD(VDD),.Y(I31347),.A(g32956),.B(g32957),.C(g32958),.D(g32959));
  AND2 AND2_1518(.VSS(VSS),.VDD(VDD),.Y(g22859),.A(g9456),.B(g20734));
  AND2 AND2_1519(.VSS(VSS),.VDD(VDD),.Y(g26154),.A(g1830),.B(g25426));
  AND2 AND2_1520(.VSS(VSS),.VDD(VDD),.Y(g30239),.A(g28728),.B(g23923));
  AND2 AND2_1521(.VSS(VSS),.VDD(VDD),.Y(g17785),.A(g13341),.B(g10762));
  AND2 AND2_1522(.VSS(VSS),.VDD(VDD),.Y(g25166),.A(g17506),.B(g23571));
  AND2 AND2_1523(.VSS(VSS),.VDD(VDD),.Y(g31131),.A(g2393),.B(g30020));
  AND2 AND2_1524(.VSS(VSS),.VDD(VDD),.Y(g18647),.A(g4040),.B(g17271));
  AND2 AND2_1525(.VSS(VSS),.VDD(VDD),.Y(g34074),.A(g33685),.B(g19498));
  AND2 AND2_1526(.VSS(VSS),.VDD(VDD),.Y(g30594),.A(g18898),.B(g29846));
  AND2 AND2_1527(.VSS(VSS),.VDD(VDD),.Y(g18356),.A(g1802),.B(g17955));
  AND2 AND2_1528(.VSS(VSS),.VDD(VDD),.Y(g29876),.A(g28404),.B(g23339));
  AND2 AND2_1529(.VSS(VSS),.VDD(VDD),.Y(g29885),.A(g28416),.B(g23350));
  AND2 AND2_1530(.VSS(VSS),.VDD(VDD),.Y(g21744),.A(g3103),.B(g20330));
  AND2 AND2_1531(.VSS(VSS),.VDD(VDD),.Y(g30238),.A(g28727),.B(g23922));
  AND2 AND2_1532(.VSS(VSS),.VDD(VDD),.Y(g34567),.A(g34377),.B(g17491));
  AND3 AND3_93(.VSS(VSS),.VDD(VDD),.Y(I31600),.A(g31009),.B(g8400),.C(g7809));
  AND2 AND2_1533(.VSS(VSS),.VDD(VDD),.Y(g28440),.A(g27274),.B(g20059));
  AND2 AND2_1534(.VSS(VSS),.VDD(VDD),.Y(g18826),.A(g7097),.B(g15680));
  AND2 AND2_1535(.VSS(VSS),.VDD(VDD),.Y(g18380),.A(g1926),.B(g15171));
  AND2 AND2_1536(.VSS(VSS),.VDD(VDD),.Y(g19571),.A(g3498),.B(g16812));
  AND3 AND3_94(.VSS(VSS),.VDD(VDD),.Y(g33487),.A(g32649),.B(I31131),.C(I31132));
  AND2 AND2_1537(.VSS(VSS),.VDD(VDD),.Y(g22172),.A(g8064),.B(g19857));
  AND2 AND2_1538(.VSS(VSS),.VDD(VDD),.Y(g29854),.A(g2197),.B(g29092));
  AND2 AND2_1539(.VSS(VSS),.VDD(VDD),.Y(g21849),.A(g3889),.B(g21070));
  AND2 AND2_1540(.VSS(VSS),.VDD(VDD),.Y(g21940),.A(g5228),.B(g18997));
  AND4 AND4_102(.VSS(VSS),.VDD(VDD),.Y(I31236),.A(g30735),.B(g31837),.C(g32796),.D(g32797));
  AND2 AND2_1541(.VSS(VSS),.VDD(VDD),.Y(g15814),.A(g3574),.B(g13920));
  AND2 AND2_1542(.VSS(VSS),.VDD(VDD),.Y(g31502),.A(g2472),.B(g29311));
  AND2 AND2_1543(.VSS(VSS),.VDD(VDD),.Y(g28573),.A(g7349),.B(g27059));
  AND3 AND3_95(.VSS(VSS),.VDD(VDD),.Y(g25485),.A(g6098),.B(g22220),.C(I24600));
  AND3 AND3_96(.VSS(VSS),.VDD(VDD),.Y(g33502),.A(g32758),.B(I31206),.C(I31207));
  AND2 AND2_1544(.VSS(VSS),.VDD(VDD),.Y(g29511),.A(g1736),.B(g28783));
  AND2 AND2_1545(.VSS(VSS),.VDD(VDD),.Y(g31210),.A(g2509),.B(g30100));
  AND4 AND4_103(.VSS(VSS),.VDD(VDD),.Y(I31351),.A(g30937),.B(g31858),.C(g32961),.D(g32962));
  AND2 AND2_1546(.VSS(VSS),.VDD(VDD),.Y(g18233),.A(g1094),.B(g16326));
  AND2 AND2_1547(.VSS(VSS),.VDD(VDD),.Y(g28247),.A(g27147),.B(g19675));
  AND2 AND2_1548(.VSS(VSS),.VDD(VDD),.Y(g21848),.A(g3913),.B(g21070));
  AND2 AND2_1549(.VSS(VSS),.VDD(VDD),.Y(g15807),.A(g3570),.B(g13898));
  AND2 AND2_1550(.VSS(VSS),.VDD(VDD),.Y(g18182),.A(g776),.B(g17328));
  AND2 AND2_1551(.VSS(VSS),.VDD(VDD),.Y(g27310),.A(g26574),.B(g23059));
  AND2 AND2_1552(.VSS(VSS),.VDD(VDD),.Y(g18651),.A(g15102),.B(g16249));
  AND2 AND2_1553(.VSS(VSS),.VDD(VDD),.Y(g18672),.A(g15127),.B(g15758));
  AND2 AND2_1554(.VSS(VSS),.VDD(VDD),.Y(g34382),.A(g34167),.B(g20618));
  AND2 AND2_1555(.VSS(VSS),.VDD(VDD),.Y(g30185),.A(g28640),.B(g23838));
  AND2 AND2_1556(.VSS(VSS),.VDD(VDD),.Y(g34519),.A(g34293),.B(g19504));
  AND2 AND2_1557(.VSS(VSS),.VDD(VDD),.Y(g17151),.A(g8659),.B(g12996));
  AND2 AND2_1558(.VSS(VSS),.VDD(VDD),.Y(g21804),.A(g3542),.B(g20924));
  AND2 AND2_1559(.VSS(VSS),.VDD(VDD),.Y(g34185),.A(g33702),.B(g24389));
  AND2 AND2_1560(.VSS(VSS),.VDD(VDD),.Y(g27627),.A(g13266),.B(g25790));
  AND2 AND2_1561(.VSS(VSS),.VDD(VDD),.Y(g25570),.A(I24689),.B(I24690));
  AND2 AND2_1562(.VSS(VSS),.VDD(VDD),.Y(g27959),.A(g25948),.B(g19374));
  AND2 AND2_1563(.VSS(VSS),.VDD(VDD),.Y(g28612),.A(g27524),.B(g20539));
  AND3 AND3_97(.VSS(VSS),.VDD(VDD),.Y(g34092),.A(g33750),.B(g9104),.C(g18957));
  AND2 AND2_1564(.VSS(VSS),.VDD(VDD),.Y(g30154),.A(g28611),.B(g23769));
  AND2 AND2_1565(.VSS(VSS),.VDD(VDD),.Y(g28324),.A(g9875),.B(g27687));
  AND2 AND2_1566(.VSS(VSS),.VDD(VDD),.Y(g24482),.A(g6875),.B(g23055));
  AND2 AND2_1567(.VSS(VSS),.VDD(VDD),.Y(g31278),.A(g29716),.B(g23302));
  AND2 AND2_1568(.VSS(VSS),.VDD(VDD),.Y(g34518),.A(g34292),.B(g19503));
  AND2 AND2_1569(.VSS(VSS),.VDD(VDD),.Y(g32274),.A(g31256),.B(g20447));
  AND2 AND2_1570(.VSS(VSS),.VDD(VDD),.Y(g27050),.A(g25789),.B(g22338));
  AND2 AND2_1571(.VSS(VSS),.VDD(VDD),.Y(g27958),.A(g25950),.B(g22449));
  AND2 AND2_1572(.VSS(VSS),.VDD(VDD),.Y(g25907),.A(g24799),.B(g22519));
  AND2 AND2_1573(.VSS(VSS),.VDD(VDD),.Y(g24710),.A(g22679),.B(g19771));
  AND2 AND2_1574(.VSS(VSS),.VDD(VDD),.Y(g27378),.A(g26089),.B(g20052));
  AND4 AND4_104(.VSS(VSS),.VDD(VDD),.Y(I31137),.A(g32654),.B(g32655),.C(g32656),.D(g32657));
  AND2 AND2_1575(.VSS(VSS),.VDD(VDD),.Y(g18331),.A(g1682),.B(g17873));
  AND3 AND3_98(.VSS(VSS),.VDD(VDD),.Y(I27364),.A(g25541),.B(g26424),.C(g22698));
  AND2 AND2_1576(.VSS(VSS),.VDD(VDD),.Y(g24552),.A(g22487),.B(g19538));
  AND3 AND3_99(.VSS(VSS),.VDD(VDD),.Y(g33469),.A(g32519),.B(I31041),.C(I31042));
  AND2 AND2_1577(.VSS(VSS),.VDD(VDD),.Y(g28251),.A(g27826),.B(g23662));
  AND2 AND2_1578(.VSS(VSS),.VDD(VDD),.Y(g30935),.A(g8808),.B(g29745));
  AND2 AND2_1579(.VSS(VSS),.VDD(VDD),.Y(g28272),.A(g27721),.B(g26548));
  AND2 AND2_1580(.VSS(VSS),.VDD(VDD),.Y(g31286),.A(g30159),.B(g27858));
  AND2 AND2_1581(.VSS(VSS),.VDD(VDD),.Y(g32122),.A(g31646),.B(g29944));
  AND2 AND2_1582(.VSS(VSS),.VDD(VDD),.Y(g18513),.A(g2575),.B(g15509));
  AND2 AND2_1583(.VSS(VSS),.VDD(VDD),.Y(g21332),.A(g996),.B(g15739));
  AND2 AND2_1584(.VSS(VSS),.VDD(VDD),.Y(g18449),.A(g12852),.B(g15224));
  AND3 AND3_100(.VSS(VSS),.VDD(VDD),.Y(I26972),.A(g25011),.B(g26424),.C(g22698));
  AND2 AND2_1585(.VSS(VSS),.VDD(VDD),.Y(g27386),.A(g26488),.B(g17498));
  AND2 AND2_1586(.VSS(VSS),.VDD(VDD),.Y(g19752),.A(g2771),.B(g15864));
  AND3 AND3_101(.VSS(VSS),.VDD(VDD),.Y(g33468),.A(g32512),.B(I31036),.C(I31037));
  AND2 AND2_1587(.VSS(VSS),.VDD(VDD),.Y(g15841),.A(g4273),.B(g13868));
  AND2 AND2_1588(.VSS(VSS),.VDD(VDD),.Y(g25567),.A(I24674),.B(I24675));
  AND2 AND2_1589(.VSS(VSS),.VDD(VDD),.Y(g27096),.A(g26026),.B(g16475));
  AND2 AND2_1590(.VSS(VSS),.VDD(VDD),.Y(g18448),.A(g2153),.B(g18008));
  AND2 AND2_1591(.VSS(VSS),.VDD(VDD),.Y(g29550),.A(g28990),.B(g22457));
  AND2 AND2_1592(.VSS(VSS),.VDD(VDD),.Y(g32034),.A(g14124),.B(g31239));
  AND2 AND2_1593(.VSS(VSS),.VDD(VDD),.Y(g25238),.A(g12466),.B(g23732));
  AND2 AND2_1594(.VSS(VSS),.VDD(VDD),.Y(g16806),.A(g6247),.B(g14971));
  AND2 AND2_1595(.VSS(VSS),.VDD(VDD),.Y(g29314),.A(g29005),.B(g22144));
  AND2 AND2_1596(.VSS(VSS),.VDD(VDD),.Y(g22059),.A(g6148),.B(g21611));
  AND2 AND2_1597(.VSS(VSS),.VDD(VDD),.Y(g21962),.A(g5428),.B(g21514));
  AND2 AND2_1598(.VSS(VSS),.VDD(VDD),.Y(g18505),.A(g2583),.B(g15509));
  AND2 AND2_1599(.VSS(VSS),.VDD(VDD),.Y(g21361),.A(g7869),.B(g16066));
  AND2 AND2_1600(.VSS(VSS),.VDD(VDD),.Y(g22025),.A(g5905),.B(g19147));
  AND2 AND2_1601(.VSS(VSS),.VDD(VDD),.Y(g18404),.A(g2066),.B(g15373));
  AND2 AND2_1602(.VSS(VSS),.VDD(VDD),.Y(g24786),.A(g661),.B(g23654));
  AND2 AND2_1603(.VSS(VSS),.VDD(VDD),.Y(g33815),.A(g33449),.B(g12911));
  AND2 AND2_1604(.VSS(VSS),.VDD(VDD),.Y(g32292),.A(g31269),.B(g20530));
  AND2 AND2_1605(.VSS(VSS),.VDD(VDD),.Y(g10898),.A(g3706),.B(g9100));
  AND2 AND2_1606(.VSS(VSS),.VDD(VDD),.Y(g18717),.A(g4849),.B(g15915));
  AND2 AND2_1607(.VSS(VSS),.VDD(VDD),.Y(g22058),.A(g6098),.B(g21611));
  AND2 AND2_1608(.VSS(VSS),.VDD(VDD),.Y(g31187),.A(g10118),.B(g30090));
  AND2 AND2_1609(.VSS(VSS),.VDD(VDD),.Y(g32153),.A(g31646),.B(g29999));
  AND2 AND2_1610(.VSS(VSS),.VDD(VDD),.Y(g24647),.A(g19903),.B(g22907));
  AND2 AND2_1611(.VSS(VSS),.VDD(VDD),.Y(g33677),.A(g33443),.B(g31937));
  AND2 AND2_1612(.VSS(VSS),.VDD(VDD),.Y(g31975),.A(g31761),.B(g22177));
  AND4 AND4_105(.VSS(VSS),.VDD(VDD),.Y(g13252),.A(g11561),.B(g11511),.C(g11469),.D(g699));
  AND2 AND2_1613(.VSS(VSS),.VDD(VDD),.Y(g18212),.A(g947),.B(g15979));
  AND2 AND2_1614(.VSS(VSS),.VDD(VDD),.Y(g29596),.A(g27823),.B(g28620));
  AND2 AND2_1615(.VSS(VSS),.VDD(VDD),.Y(g24945),.A(g23183),.B(g20197));
  AND3 AND3_102(.VSS(VSS),.VDD(VDD),.Y(g10719),.A(g6841),.B(g2138),.C(g2130));
  AND2 AND2_1616(.VSS(VSS),.VDD(VDD),.Y(g16517),.A(g5248),.B(g14797));
  AND2 AND2_1617(.VSS(VSS),.VDD(VDD),.Y(g21833),.A(g15096),.B(g20453));
  AND2 AND2_1618(.VSS(VSS),.VDD(VDD),.Y(g30215),.A(g28690),.B(g23881));
  AND2 AND2_1619(.VSS(VSS),.VDD(VDD),.Y(g32409),.A(g4754),.B(g30996));
  AND2 AND2_1620(.VSS(VSS),.VDD(VDD),.Y(g14719),.A(g4392),.B(g10830));
  AND2 AND2_1621(.VSS(VSS),.VDD(VDD),.Y(g34215),.A(g33778),.B(g22670));
  AND2 AND2_1622(.VSS(VSS),.VDD(VDD),.Y(g30577),.A(g26267),.B(g29679));
  AND2 AND2_1623(.VSS(VSS),.VDD(VDD),.Y(g34577),.A(g24577),.B(g34307));
  AND3 AND3_103(.VSS(VSS),.VDD(VDD),.Y(g25518),.A(g6444),.B(g23865),.C(I24625));
  AND2 AND2_1624(.VSS(VSS),.VDD(VDD),.Y(g27428),.A(g26400),.B(g17576));
  AND2 AND2_1625(.VSS(VSS),.VDD(VDD),.Y(g13564),.A(g4480),.B(g12820));
  AND2 AND2_1626(.VSS(VSS),.VDD(VDD),.Y(g22044),.A(g6058),.B(g21611));
  AND2 AND2_1627(.VSS(VSS),.VDD(VDD),.Y(g26304),.A(g2697),.B(g25246));
  AND2 AND2_1628(.VSS(VSS),.VDD(VDD),.Y(g31143),.A(g29506),.B(g22999));
  AND4 AND4_106(.VSS(VSS),.VDD(VDD),.Y(I24709),.A(g21256),.B(g24068),.C(g24069),.D(g24070));
  AND4 AND4_107(.VSS(VSS),.VDD(VDD),.Y(I31021),.A(g31070),.B(g31799),.C(g32485),.D(g32486));
  AND2 AND2_1629(.VSS(VSS),.VDD(VDD),.Y(g24998),.A(g17412),.B(g23408));
  AND2 AND2_1630(.VSS(VSS),.VDD(VDD),.Y(g12730),.A(g9024),.B(g4349));
  AND2 AND2_1631(.VSS(VSS),.VDD(VDD),.Y(g27765),.A(g4146),.B(g25886));
  AND2 AND2_1632(.VSS(VSS),.VDD(VDD),.Y(g24651),.A(g2741),.B(g23472));
  AND2 AND2_1633(.VSS(VSS),.VDD(VDD),.Y(g24672),.A(g19534),.B(g22981));
  AND2 AND2_1634(.VSS(VSS),.VDD(VDD),.Y(g14832),.A(g1489),.B(g10939));
  AND2 AND2_1635(.VSS(VSS),.VDD(VDD),.Y(g29773),.A(g28203),.B(g10233));
  AND2 AND2_1636(.VSS(VSS),.VDD(VDD),.Y(g27690),.A(g25784),.B(g23607));
  AND2 AND2_1637(.VSS(VSS),.VDD(VDD),.Y(g16193),.A(g6533),.B(g14348));
  AND2 AND2_1638(.VSS(VSS),.VDD(VDD),.Y(g27549),.A(g26576),.B(g14785));
  AND2 AND2_1639(.VSS(VSS),.VDD(VDD),.Y(g31169),.A(g10083),.B(g30079));
  AND2 AND2_1640(.VSS(VSS),.VDD(VDD),.Y(g11397),.A(g5360),.B(g7139));
  AND2 AND2_1641(.VSS(VSS),.VDD(VDD),.Y(g18723),.A(g4922),.B(g16077));
  AND2 AND2_1642(.VSS(VSS),.VDD(VDD),.Y(g25883),.A(g13728),.B(g24699));
  AND2 AND2_1643(.VSS(VSS),.VDD(VDD),.Y(g28360),.A(g27401),.B(g19861));
  AND2 AND2_1644(.VSS(VSS),.VDD(VDD),.Y(g22120),.A(g6585),.B(g19277));
  AND2 AND2_1645(.VSS(VSS),.VDD(VDD),.Y(g33884),.A(g33295),.B(g20590));
  AND2 AND2_1646(.VSS(VSS),.VDD(VDD),.Y(g15116),.A(g4297),.B(g14454));
  AND2 AND2_1647(.VSS(VSS),.VDD(VDD),.Y(g18149),.A(g608),.B(g17533));
  AND2 AND2_1648(.VSS(VSS),.VDD(VDD),.Y(g27548),.A(g26576),.B(g17763));
  AND2 AND2_1649(.VSS(VSS),.VDD(VDD),.Y(g31168),.A(g2241),.B(g30077));
  AND2 AND2_1650(.VSS(VSS),.VDD(VDD),.Y(g32164),.A(g30733),.B(g25171));
  AND2 AND2_1651(.VSS(VSS),.VDD(VDD),.Y(g18433),.A(g2197),.B(g18008));
  AND2 AND2_1652(.VSS(VSS),.VDD(VDD),.Y(g33410),.A(g32360),.B(g21409));
  AND2 AND2_1653(.VSS(VSS),.VDD(VDD),.Y(g18387),.A(g1955),.B(g15171));
  AND2 AND2_1654(.VSS(VSS),.VDD(VDD),.Y(g24331),.A(g6977),.B(g22228));
  AND2 AND2_1655(.VSS(VSS),.VDD(VDD),.Y(g30083),.A(g28533),.B(g20698));
  AND2 AND2_1656(.VSS(VSS),.VDD(VDD),.Y(g13509),.A(g9951),.B(g11889));
  AND2 AND2_1657(.VSS(VSS),.VDD(VDD),.Y(g27504),.A(g26519),.B(g17680));
  AND2 AND2_1658(.VSS(VSS),.VDD(VDD),.Y(g18620),.A(g3470),.B(g17062));
  AND2 AND2_1659(.VSS(VSS),.VDD(VDD),.Y(g18148),.A(g562),.B(g17533));
  AND2 AND2_1660(.VSS(VSS),.VDD(VDD),.Y(g21947),.A(g5256),.B(g18997));
  AND2 AND2_1661(.VSS(VSS),.VDD(VDD),.Y(g30284),.A(g28852),.B(g23994));
  AND2 AND2_1662(.VSS(VSS),.VDD(VDD),.Y(g34083),.A(g33714),.B(g19573));
  AND2 AND2_1663(.VSS(VSS),.VDD(VDD),.Y(g34348),.A(g34125),.B(g20128));
  AND3 AND3_104(.VSS(VSS),.VDD(VDD),.Y(I31593),.A(g31003),.B(g8350),.C(g7788));
  AND3 AND3_105(.VSS(VSS),.VDD(VDD),.Y(g33479),.A(g32593),.B(I31091),.C(I31092));
  AND2 AND2_1664(.VSS(VSS),.VDD(VDD),.Y(g34284),.A(g34046),.B(g19351));
  AND2 AND2_1665(.VSS(VSS),.VDD(VDD),.Y(g21605),.A(g13005),.B(g15695));
  AND4 AND4_108(.VSS(VSS),.VDD(VDD),.Y(I31346),.A(g31021),.B(g31857),.C(g32954),.D(g32955));
  AND2 AND2_1666(.VSS(VSS),.VDD(VDD),.Y(g33363),.A(g32262),.B(g20918));
  AND2 AND2_1667(.VSS(VSS),.VDD(VDD),.Y(g13508),.A(g9927),.B(g11888));
  AND2 AND2_1668(.VSS(VSS),.VDD(VDD),.Y(g18104),.A(g392),.B(g17015));
  AND2 AND2_1669(.VSS(VSS),.VDD(VDD),.Y(g18811),.A(g6500),.B(g15483));
  AND2 AND2_1670(.VSS(VSS),.VDD(VDD),.Y(g18646),.A(g4031),.B(g17271));
  AND4 AND4_109(.VSS(VSS),.VDD(VDD),.Y(I31122),.A(g32631),.B(g32632),.C(g32633),.D(g32634));
  AND2 AND2_1671(.VSS(VSS),.VDD(VDD),.Y(g14612),.A(g11971),.B(g11993));
  AND2 AND2_1672(.VSS(VSS),.VDD(VDD),.Y(g31478),.A(g29764),.B(g23410));
  AND2 AND2_1673(.VSS(VSS),.VDD(VDD),.Y(g8234),.A(g4515),.B(g4521));
  AND2 AND2_1674(.VSS(VSS),.VDD(VDD),.Y(g31015),.A(g29476),.B(g22758));
  AND2 AND2_1675(.VSS(VSS),.VDD(VDD),.Y(g18343),.A(g12847),.B(g17955));
  AND3 AND3_106(.VSS(VSS),.VDD(VDD),.Y(g24897),.A(g3401),.B(g23223),.C(I24064));
  AND2 AND2_1676(.VSS(VSS),.VDD(VDD),.Y(g29839),.A(g1728),.B(g29045));
  AND2 AND2_1677(.VSS(VSS),.VDD(VDD),.Y(g30566),.A(g26247),.B(g29507));
  AND3 AND3_107(.VSS(VSS),.VDD(VDD),.Y(g33478),.A(g32584),.B(I31086),.C(I31087));
  AND2 AND2_1678(.VSS(VSS),.VDD(VDD),.Y(g24961),.A(g23193),.B(g20209));
  AND2 AND2_1679(.VSS(VSS),.VDD(VDD),.Y(g21812),.A(g3586),.B(g20924));
  AND2 AND2_1680(.VSS(VSS),.VDD(VDD),.Y(g17146),.A(g5965),.B(g14895));
  AND2 AND2_1681(.VSS(VSS),.VDD(VDD),.Y(g34566),.A(g34376),.B(g17489));
  AND2 AND2_1682(.VSS(VSS),.VDD(VDD),.Y(g28451),.A(g27283),.B(g20090));
  AND2 AND2_1683(.VSS(VSS),.VDD(VDD),.Y(g16222),.A(g6513),.B(g14348));
  AND2 AND2_1684(.VSS(VSS),.VDD(VDD),.Y(g31486),.A(g29777),.B(g23422));
  AND2 AND2_1685(.VSS(VSS),.VDD(VDD),.Y(g32327),.A(g31319),.B(g23544));
  AND2 AND2_1686(.VSS(VSS),.VDD(VDD),.Y(g29667),.A(g2671),.B(g29157));
  AND2 AND2_1687(.VSS(VSS),.VDD(VDD),.Y(g29838),.A(g1636),.B(g29044));
  AND2 AND2_1688(.VSS(VSS),.VDD(VDD),.Y(g27129),.A(g26026),.B(g16584));
  AND3 AND3_108(.VSS(VSS),.VDD(VDD),.Y(g33486),.A(g32642),.B(I31126),.C(I31127));
  AND2 AND2_1689(.VSS(VSS),.VDD(VDD),.Y(g32109),.A(g31609),.B(g29920));
  AND2 AND2_1690(.VSS(VSS),.VDD(VDD),.Y(g21951),.A(g5272),.B(g18997));
  AND2 AND2_1691(.VSS(VSS),.VDD(VDD),.Y(g26852),.A(g24975),.B(g24958));
  AND2 AND2_1692(.VSS(VSS),.VDD(VDD),.Y(g21972),.A(g15152),.B(g19074));
  AND4 AND4_110(.VSS(VSS),.VDD(VDD),.Y(g27057),.A(g7791),.B(g6219),.C(g6227),.D(g26261));
  AND2 AND2_1693(.VSS(VSS),.VDD(VDD),.Y(g19610),.A(g1141),.B(g16069));
  AND2 AND2_1694(.VSS(VSS),.VDD(VDD),.Y(g18369),.A(g12848),.B(g15171));
  AND2 AND2_1695(.VSS(VSS),.VDD(VDD),.Y(g24717),.A(g22684),.B(g19777));
  AND2 AND2_1696(.VSS(VSS),.VDD(VDD),.Y(g27128),.A(g25997),.B(g16583));
  AND2 AND2_1697(.VSS(VSS),.VDD(VDD),.Y(g28246),.A(g8572),.B(g27976));
  AND4 AND4_111(.VSS(VSS),.VDD(VDD),.Y(I31292),.A(g32877),.B(g32878),.C(g32879),.D(g32880));
  AND2 AND2_1698(.VSS(VSS),.VDD(VDD),.Y(g32108),.A(g31631),.B(g29913));
  AND2 AND2_1699(.VSS(VSS),.VDD(VDD),.Y(g30139),.A(g28596),.B(g21184));
  AND2 AND2_1700(.VSS(VSS),.VDD(VDD),.Y(g18368),.A(g1728),.B(g17955));
  AND2 AND2_1701(.VSS(VSS),.VDD(VDD),.Y(g34139),.A(g33827),.B(g23314));
  AND2 AND2_1702(.VSS(VSS),.VDD(VDD),.Y(g16703),.A(g5889),.B(g15002));
  AND2 AND2_1703(.VSS(VSS),.VDD(VDD),.Y(g22632),.A(g19356),.B(g19476));
  AND2 AND2_1704(.VSS(VSS),.VDD(VDD),.Y(g31223),.A(g20028),.B(g29689));
  AND2 AND2_1705(.VSS(VSS),.VDD(VDD),.Y(g21795),.A(g3506),.B(g20924));
  AND2 AND2_1706(.VSS(VSS),.VDD(VDD),.Y(g32283),.A(g31259),.B(g20506));
  AND2 AND2_1707(.VSS(VSS),.VDD(VDD),.Y(g27323),.A(g26268),.B(g23086));
  AND2 AND2_1708(.VSS(VSS),.VDD(VDD),.Y(g30138),.A(g28595),.B(g21182));
  AND2 AND2_1709(.VSS(VSS),.VDD(VDD),.Y(g27299),.A(g26546),.B(g23028));
  AND2 AND2_1710(.VSS(VSS),.VDD(VDD),.Y(g29619),.A(g2269),.B(g29060));
  AND2 AND2_1711(.VSS(VSS),.VDD(VDD),.Y(g32303),.A(g27550),.B(g31376));
  AND2 AND2_1712(.VSS(VSS),.VDD(VDD),.Y(g34138),.A(g33929),.B(g23828));
  AND2 AND2_1713(.VSS(VSS),.VDD(VDD),.Y(g11047),.A(g6474),.B(g9212));
  AND2 AND2_1714(.VSS(VSS),.VDD(VDD),.Y(g18412),.A(g2098),.B(g15373));
  AND4 AND4_112(.VSS(VSS),.VDD(VDD),.Y(I31136),.A(g29385),.B(g32651),.C(g32652),.D(g32653));
  AND2 AND2_1715(.VSS(VSS),.VDD(VDD),.Y(g11205),.A(g8217),.B(g8439));
  AND2 AND2_1716(.VSS(VSS),.VDD(VDD),.Y(g13047),.A(g8534),.B(g11042));
  AND2 AND2_1717(.VSS(VSS),.VDD(VDD),.Y(g27298),.A(g26573),.B(g23026));
  AND2 AND2_1718(.VSS(VSS),.VDD(VDD),.Y(g29618),.A(g28870),.B(g22384));
  AND2 AND2_1719(.VSS(VSS),.VDD(VDD),.Y(g19383),.A(g16893),.B(g13223));
  AND2 AND2_1720(.VSS(VSS),.VDD(VDD),.Y(g34415),.A(g34207),.B(g21458));
  AND2 AND2_1721(.VSS(VSS),.VDD(VDD),.Y(g18133),.A(g15055),.B(g17249));
  AND2 AND2_1722(.VSS(VSS),.VDD(VDD),.Y(g23514),.A(g20149),.B(g11829));
  AND2 AND2_1723(.VSS(VSS),.VDD(VDD),.Y(g26484),.A(g24946),.B(g8841));
  AND2 AND2_1724(.VSS(VSS),.VDD(VDD),.Y(g33110),.A(g32404),.B(g32415));
  AND2 AND2_1725(.VSS(VSS),.VDD(VDD),.Y(g13912),.A(g5551),.B(g12450));
  AND2 AND2_1726(.VSS(VSS),.VDD(VDD),.Y(g34333),.A(g9984),.B(g34192));
  AND2 AND2_1727(.VSS(VSS),.VDD(VDD),.Y(g24723),.A(g17490),.B(g22384));
  AND2 AND2_1728(.VSS(VSS),.VDD(VDD),.Y(g31321),.A(g30146),.B(g27886));
  AND2 AND2_1729(.VSS(VSS),.VDD(VDD),.Y(g18229),.A(g1099),.B(g16326));
  AND2 AND2_1730(.VSS(VSS),.VDD(VDD),.Y(g33922),.A(g33448),.B(g7202));
  AND2 AND2_1731(.VSS(VSS),.VDD(VDD),.Y(g14061),.A(g8715),.B(g11834));
  AND3 AND3_109(.VSS(VSS),.VDD(VDD),.Y(g33531),.A(g32967),.B(I31351),.C(I31352));
  AND2 AND2_1732(.VSS(VSS),.VDD(VDD),.Y(g18228),.A(g1061),.B(g16129));
  AND2 AND2_1733(.VSS(VSS),.VDD(VDD),.Y(g24387),.A(g3457),.B(g22761));
  AND2 AND2_1734(.VSS(VSS),.VDD(VDD),.Y(g26312),.A(g2704),.B(g25264));
  AND2 AND2_1735(.VSS(VSS),.VDD(VDD),.Y(g34963),.A(g34946),.B(g23041));
  AND4 AND4_113(.VSS(VSS),.VDD(VDD),.Y(g26200),.A(g24688),.B(g10678),.C(g10658),.D(g10627));
  AND2 AND2_1736(.VSS(VSS),.VDD(VDD),.Y(g32174),.A(g31708),.B(g27837));
  AND2 AND2_1737(.VSS(VSS),.VDD(VDD),.Y(g21163),.A(g16321),.B(g4878));
  AND2 AND2_1738(.VSS(VSS),.VDD(VDD),.Y(g21012),.A(g16304),.B(g4688));
  AND2 AND2_1739(.VSS(VSS),.VDD(VDD),.Y(g28151),.A(g8426),.B(g27295));
  AND2 AND2_1740(.VSS(VSS),.VDD(VDD),.Y(g18716),.A(g4878),.B(g15915));
  AND2 AND2_1741(.VSS(VSS),.VDD(VDD),.Y(g31186),.A(g2375),.B(g30088));
  AND2 AND2_1742(.VSS(VSS),.VDD(VDD),.Y(g33186),.A(g32037),.B(g22830));
  AND2 AND2_1743(.VSS(VSS),.VDD(VDD),.Y(g24646),.A(g22640),.B(g19711));
  AND2 AND2_1744(.VSS(VSS),.VDD(VDD),.Y(g33676),.A(g33125),.B(g7970));
  AND2 AND2_1745(.VSS(VSS),.VDD(VDD),.Y(g33373),.A(g32288),.B(g21205));
  AND2 AND2_1746(.VSS(VSS),.VDD(VDD),.Y(g16516),.A(g5228),.B(g14627));
  AND2 AND2_1747(.VSS(VSS),.VDD(VDD),.Y(g27697),.A(g25785),.B(g23649));
  AND2 AND2_1748(.VSS(VSS),.VDD(VDD),.Y(g18582),.A(g2922),.B(g16349));
  AND2 AND2_1749(.VSS(VSS),.VDD(VDD),.Y(g27995),.A(g26809),.B(g23985));
  AND2 AND2_1750(.VSS(VSS),.VDD(VDD),.Y(g31654),.A(g29325),.B(g13062));
  AND2 AND2_1751(.VSS(VSS),.VDD(VDD),.Y(g30576),.A(g18898),.B(g29800));
  AND2 AND2_1752(.VSS(VSS),.VDD(VDD),.Y(g22127),.A(g6625),.B(g19277));
  AND2 AND2_1753(.VSS(VSS),.VDD(VDD),.Y(g34585),.A(g24705),.B(g34316));
  AND2 AND2_1754(.VSS(VSS),.VDD(VDD),.Y(g34484),.A(g34407),.B(g18939));
  AND2 AND2_1755(.VSS(VSS),.VDD(VDD),.Y(g18310),.A(g1333),.B(g16931));
  AND2 AND2_1756(.VSS(VSS),.VDD(VDD),.Y(g29601),.A(g1890),.B(g28955));
  AND2 AND2_1757(.VSS(VSS),.VDD(VDD),.Y(g31936),.A(g31213),.B(g24005));
  AND2 AND2_1758(.VSS(VSS),.VDD(VDD),.Y(g33417),.A(g32371),.B(g21424));
  AND4 AND4_114(.VSS(VSS),.VDD(VDD),.Y(I31327),.A(g32928),.B(g32929),.C(g32930),.D(g32931));
  AND2 AND2_1759(.VSS(VSS),.VDD(VDD),.Y(g21789),.A(g3451),.B(g20391));
  AND2 AND2_1760(.VSS(VSS),.VDD(VDD),.Y(g26799),.A(g25247),.B(g21068));
  AND2 AND2_1761(.VSS(VSS),.VDD(VDD),.Y(g29975),.A(g28986),.B(g10420));
  AND2 AND2_1762(.VSS(VSS),.VDD(VDD),.Y(g34554),.A(g34347),.B(g20495));
  AND2 AND2_1763(.VSS(VSS),.VDD(VDD),.Y(g18627),.A(g15093),.B(g17093));
  AND2 AND2_1764(.VSS(VSS),.VDD(VDD),.Y(g15863),.A(g13762),.B(g13223));
  AND2 AND2_1765(.VSS(VSS),.VDD(VDD),.Y(g18379),.A(g1906),.B(g15171));
  AND2 AND2_1766(.VSS(VSS),.VDD(VDD),.Y(g30200),.A(g28665),.B(g23862));
  AND2 AND2_1767(.VSS(VSS),.VDD(VDD),.Y(g21788),.A(g3401),.B(g20391));
  AND2 AND2_1768(.VSS(VSS),.VDD(VDD),.Y(g33334),.A(g32219),.B(g20613));
  AND2 AND2_1769(.VSS(VSS),.VDD(VDD),.Y(g18112),.A(g182),.B(g17015));
  AND2 AND2_1770(.VSS(VSS),.VDD(VDD),.Y(g16422),.A(g8216),.B(g13627));
  AND2 AND2_1771(.VSS(VSS),.VDD(VDD),.Y(g23724),.A(g14767),.B(g21123));
  AND2 AND2_1772(.VSS(VSS),.VDD(VDD),.Y(g25852),.A(g4593),.B(g24411));
  AND2 AND2_1773(.VSS(VSS),.VDD(VDD),.Y(g18378),.A(g1932),.B(g15171));
  AND2 AND2_1774(.VSS(VSS),.VDD(VDD),.Y(g22103),.A(g15164),.B(g18833));
  AND3 AND3_110(.VSS(VSS),.VDD(VDD),.Y(g34115),.A(g20516),.B(g9104),.C(g33750));
  AND2 AND2_1775(.VSS(VSS),.VDD(VDD),.Y(g21829),.A(g3770),.B(g20453));
  AND2 AND2_1776(.VSS(VSS),.VDD(VDD),.Y(g29937),.A(g13044),.B(g29196));
  AND2 AND2_1777(.VSS(VSS),.VDD(VDD),.Y(g14220),.A(g8612),.B(g11820));
  AND2 AND2_1778(.VSS(VSS),.VDD(VDD),.Y(g21920),.A(g5062),.B(g21468));
  AND2 AND2_1779(.VSS(VSS),.VDD(VDD),.Y(g23920),.A(g4135),.B(g19549));
  AND2 AND2_1780(.VSS(VSS),.VDD(VDD),.Y(g22095),.A(g6428),.B(g18833));
  AND2 AND2_1781(.VSS(VSS),.VDD(VDD),.Y(g16208),.A(g3965),.B(g14085));
  AND2 AND2_1782(.VSS(VSS),.VDD(VDD),.Y(g25963),.A(g1657),.B(g24978));
  AND2 AND2_1783(.VSS(VSS),.VDD(VDD),.Y(g28318),.A(g27233),.B(g19770));
  AND2 AND2_1784(.VSS(VSS),.VDD(VDD),.Y(g18386),.A(g1964),.B(g15171));
  AND2 AND2_1785(.VSS(VSS),.VDD(VDD),.Y(g30921),.A(g29900),.B(g24789));
  AND2 AND2_1786(.VSS(VSS),.VDD(VDD),.Y(g28227),.A(g9397),.B(g27583));
  AND2 AND2_1787(.VSS(VSS),.VDD(VDD),.Y(g21828),.A(g3767),.B(g20453));
  AND2 AND2_1788(.VSS(VSS),.VDD(VDD),.Y(g15703),.A(g452),.B(g13437));
  AND2 AND2_1789(.VSS(VSS),.VDD(VDD),.Y(g17784),.A(g1152),.B(g13215));
  AND2 AND2_1790(.VSS(VSS),.VDD(VDD),.Y(g23828),.A(g9104),.B(g19128));
  AND2 AND2_1791(.VSS(VSS),.VDD(VDD),.Y(g18603),.A(g3119),.B(g16987));
  AND2 AND2_1792(.VSS(VSS),.VDD(VDD),.Y(g21946),.A(g5252),.B(g18997));
  AND2 AND2_1793(.VSS(VSS),.VDD(VDD),.Y(g18742),.A(g5120),.B(g17847));
  AND4 AND4_115(.VSS(VSS),.VDD(VDD),.Y(g27445),.A(g8038),.B(g26314),.C(g9187),.D(g504));
  AND2 AND2_1794(.VSS(VSS),.VDD(VDD),.Y(g33423),.A(g32225),.B(g29657));
  AND2 AND2_1795(.VSS(VSS),.VDD(VDD),.Y(g29884),.A(g2555),.B(g29153));
  AND2 AND2_1796(.VSS(VSS),.VDD(VDD),.Y(g23121),.A(g19128),.B(g9104));
  AND2 AND2_1797(.VSS(VSS),.VDD(VDD),.Y(g24229),.A(g896),.B(g22594));
  AND2 AND2_1798(.VSS(VSS),.VDD(VDD),.Y(g34745),.A(g34669),.B(g19482));
  AND2 AND2_1799(.VSS(VSS),.VDD(VDD),.Y(g27316),.A(g2407),.B(g26710));
  AND2 AND2_1800(.VSS(VSS),.VDD(VDD),.Y(g24228),.A(g862),.B(g22594));
  AND2 AND2_1801(.VSS(VSS),.VDD(VDD),.Y(g18681),.A(g4653),.B(g15885));
  AND4 AND4_116(.VSS(VSS),.VDD(VDD),.Y(I31091),.A(g29385),.B(g32586),.C(g32587),.D(g32588));
  AND2 AND2_1802(.VSS(VSS),.VDD(VDD),.Y(g24011),.A(g7939),.B(g19524));
  AND2 AND2_1803(.VSS(VSS),.VDD(VDD),.Y(g32326),.A(g31317),.B(g23539));
  AND2 AND2_1804(.VSS(VSS),.VDD(VDD),.Y(g29666),.A(g28980),.B(g22498));
  AND2 AND2_1805(.VSS(VSS),.VDD(VDD),.Y(g17181),.A(g1945),.B(g13014));
  AND2 AND2_1806(.VSS(VSS),.VDD(VDD),.Y(g16614),.A(g5945),.B(g14933));
  AND2 AND2_1807(.VSS(VSS),.VDD(VDD),.Y(g17671),.A(g7685),.B(g13485));
  AND2 AND2_1808(.VSS(VSS),.VDD(VDD),.Y(g29363),.A(g8458),.B(g28444));
  AND2 AND2_1809(.VSS(VSS),.VDD(VDD),.Y(g23682),.A(g16970),.B(g20874));
  AND2 AND2_1810(.VSS(VSS),.VDD(VDD),.Y(g18802),.A(g6195),.B(g15348));
  AND2 AND2_1811(.VSS(VSS),.VDD(VDD),.Y(g18429),.A(g2193),.B(g18008));
  AND2 AND2_1812(.VSS(VSS),.VDD(VDD),.Y(g32040),.A(g14122),.B(g31243));
  AND2 AND2_1813(.VSS(VSS),.VDD(VDD),.Y(g24716),.A(g15935),.B(g23004));
  AND4 AND4_117(.VSS(VSS),.VDD(VDD),.Y(I24680),.A(g24029),.B(g24030),.C(g24031),.D(g24032));
  AND2 AND2_1814(.VSS(VSS),.VDD(VDD),.Y(g33909),.A(g33131),.B(g10708));
  AND2 AND2_1815(.VSS(VSS),.VDD(VDD),.Y(g34184),.A(g33698),.B(g24388));
  AND2 AND2_1816(.VSS(VSS),.VDD(VDD),.Y(g18730),.A(g4950),.B(g16861));
  AND2 AND2_1817(.VSS(VSS),.VDD(VDD),.Y(g15821),.A(g3598),.B(g14110));
  AND2 AND2_1818(.VSS(VSS),.VDD(VDD),.Y(g27988),.A(g26781),.B(g23941));
  AND2 AND2_1819(.VSS(VSS),.VDD(VDD),.Y(g18793),.A(g6159),.B(g15348));
  AND2 AND2_1820(.VSS(VSS),.VDD(VDD),.Y(g18428),.A(g2169),.B(g18008));
  AND2 AND2_1821(.VSS(VSS),.VDD(VDD),.Y(g24582),.A(g5808),.B(g23402));
  AND2 AND2_1822(.VSS(VSS),.VDD(VDD),.Y(g33908),.A(g33092),.B(g18935));
  AND3 AND3_111(.VSS(VSS),.VDD(VDD),.Y(g28281),.A(g7362),.B(g1936),.C(g27440));
  AND2 AND2_1823(.VSS(VSS),.VDD(VDD),.Y(g16593),.A(g5599),.B(g14885));
  AND2 AND2_1824(.VSS(VSS),.VDD(VDD),.Y(g12924),.A(g1570),.B(g10980));
  AND2 AND2_1825(.VSS(VSS),.VDD(VDD),.Y(g27432),.A(g26519),.B(g17582));
  AND2 AND2_1826(.VSS(VSS),.VDD(VDD),.Y(g13020),.A(g401),.B(g11048));
  AND2 AND2_1827(.VSS(VSS),.VDD(VDD),.Y(g18765),.A(g5489),.B(g17929));
  AND2 AND2_1828(.VSS(VSS),.VDD(VDD),.Y(g28301),.A(g27224),.B(g19750));
  AND2 AND2_1829(.VSS(VSS),.VDD(VDD),.Y(g24310),.A(g4495),.B(g22228));
  AND2 AND2_1830(.VSS(VSS),.VDD(VDD),.Y(g16122),.A(g9491),.B(g14291));
  AND2 AND2_1831(.VSS(VSS),.VDD(VDD),.Y(g18690),.A(g15130),.B(g16053));
  AND4 AND4_118(.VSS(VSS),.VDD(VDD),.Y(g28739),.A(g21434),.B(g26424),.C(g25274),.D(g27395));
  AND2 AND2_1832(.VSS(VSS),.VDD(VDD),.Y(g18549),.A(g2799),.B(g15277));
  AND2 AND2_1833(.VSS(VSS),.VDD(VDD),.Y(g11046),.A(g9889),.B(g6120));
  AND2 AND2_1834(.VSS(VSS),.VDD(VDD),.Y(g25921),.A(g24936),.B(g9664));
  AND2 AND2_1835(.VSS(VSS),.VDD(VDD),.Y(g13046),.A(g6870),.B(g11270));
  AND2 AND2_1836(.VSS(VSS),.VDD(VDD),.Y(g26207),.A(g2638),.B(g25170));
  AND2 AND2_1837(.VSS(VSS),.VDD(VDD),.Y(g24627),.A(g22763),.B(g19679));
  AND2 AND2_1838(.VSS(VSS),.VDD(VDD),.Y(g29580),.A(g28519),.B(g14186));
  AND2 AND2_1839(.VSS(VSS),.VDD(VDD),.Y(g21760),.A(g3207),.B(g20785));
  AND2 AND2_1840(.VSS(VSS),.VDD(VDD),.Y(g20112),.A(g13540),.B(g16661));
  AND2 AND2_1841(.VSS(VSS),.VDD(VDD),.Y(g31242),.A(g29373),.B(g25409));
  AND2 AND2_1842(.VSS(VSS),.VDD(VDD),.Y(g22089),.A(g6311),.B(g19210));
  AND2 AND2_1843(.VSS(VSS),.VDD(VDD),.Y(g27461),.A(g26576),.B(g17611));
  AND2 AND2_1844(.VSS(VSS),.VDD(VDD),.Y(g33242),.A(g32123),.B(g19931));
  AND2 AND2_1845(.VSS(VSS),.VDD(VDD),.Y(g18548),.A(g2807),.B(g15277));
  AND2 AND2_1846(.VSS(VSS),.VDD(VDD),.Y(g15873),.A(g3550),.B(g14072));
  AND2 AND2_1847(.VSS(VSS),.VDD(VDD),.Y(g28645),.A(g27556),.B(g20599));
  AND4 AND4_119(.VSS(VSS),.VDD(VDD),.Y(I31192),.A(g32733),.B(g32734),.C(g32735),.D(g32736));
  AND2 AND2_1848(.VSS(VSS),.VDD(VDD),.Y(g27342),.A(g12592),.B(g26792));
  AND2 AND2_1849(.VSS(VSS),.VDD(VDD),.Y(g24378),.A(g3106),.B(g22718));
  AND2 AND2_1850(.VSS(VSS),.VDD(VDD),.Y(g16641),.A(g6613),.B(g14782));
  AND2 AND2_1851(.VSS(VSS),.VDD(VDD),.Y(g27145),.A(g14121),.B(g26382));
  AND2 AND2_1852(.VSS(VSS),.VDD(VDD),.Y(g22088),.A(g6307),.B(g19210));
  AND2 AND2_1853(.VSS(VSS),.VDD(VDD),.Y(g18504),.A(g2579),.B(g15509));
  AND2 AND2_1854(.VSS(VSS),.VDD(VDD),.Y(g22024),.A(g5897),.B(g19147));
  AND2 AND2_1855(.VSS(VSS),.VDD(VDD),.Y(g31123),.A(g1834),.B(g29994));
  AND2 AND2_1856(.VSS(VSS),.VDD(VDD),.Y(g32183),.A(g2795),.B(g31653));
  AND2 AND2_1857(.VSS(VSS),.VDD(VDD),.Y(g19266),.A(g246),.B(g16214));
  AND2 AND2_1858(.VSS(VSS),.VDD(VDD),.Y(g33814),.A(g33098),.B(g28144));
  AND2 AND2_1859(.VSS(VSS),.VDD(VDD),.Y(g28290),.A(g23780),.B(g27759));
  AND2 AND2_1860(.VSS(VSS),.VDD(VDD),.Y(g32397),.A(g31068),.B(g15830));
  AND2 AND2_1861(.VSS(VSS),.VDD(VDD),.Y(g13282),.A(g3546),.B(g11480));
  AND2 AND2_1862(.VSS(VSS),.VDD(VDD),.Y(g27650),.A(g26519),.B(g15479));
  AND4 AND4_120(.VSS(VSS),.VDD(VDD),.Y(g29110),.A(g27187),.B(g12687),.C(g20751),.D(I27429));
  AND2 AND2_1863(.VSS(VSS),.VDD(VDD),.Y(g25973),.A(g2342),.B(g24994));
  AND2 AND2_1864(.VSS(VSS),.VDD(VDD),.Y(g18317),.A(g12846),.B(g17873));
  AND2 AND2_1865(.VSS(VSS),.VDD(VDD),.Y(g33807),.A(g33112),.B(g25452));
  AND2 AND2_1866(.VSS(VSS),.VDD(VDD),.Y(g31974),.A(g31760),.B(g22176));
  AND2 AND2_1867(.VSS(VSS),.VDD(VDD),.Y(g29321),.A(g29033),.B(g22148));
  AND2 AND2_1868(.VSS(VSS),.VDD(VDD),.Y(g33639),.A(g33386),.B(g18829));
  AND4 AND4_121(.VSS(VSS),.VDD(VDD),.Y(g26241),.A(g24688),.B(g10678),.C(g8778),.D(g10627));
  AND2 AND2_1869(.VSS(VSS),.VDD(VDD),.Y(g34214),.A(g33772),.B(g22689));
  AND2 AND2_1870(.VSS(VSS),.VDD(VDD),.Y(g29531),.A(g1664),.B(g28559));
  AND2 AND2_1871(.VSS(VSS),.VDD(VDD),.Y(g31230),.A(g30285),.B(g20751));
  AND2 AND2_1872(.VSS(VSS),.VDD(VDD),.Y(g18129),.A(g518),.B(g16971));
  AND2 AND2_1873(.VSS(VSS),.VDD(VDD),.Y(g30207),.A(g28680),.B(g23874));
  AND2 AND2_1874(.VSS(VSS),.VDD(VDD),.Y(g16635),.A(g5607),.B(g14959));
  AND2 AND2_1875(.VSS(VSS),.VDD(VDD),.Y(g27696),.A(g25800),.B(g23647));
  AND2 AND2_1876(.VSS(VSS),.VDD(VDD),.Y(g34329),.A(g14511),.B(g34181));
  AND2 AND2_1877(.VSS(VSS),.VDD(VDD),.Y(g27330),.A(g2541),.B(g26744));
  AND2 AND2_1878(.VSS(VSS),.VDD(VDD),.Y(g27393),.A(g26099),.B(g20066));
  AND2 AND2_1879(.VSS(VSS),.VDD(VDD),.Y(g28427),.A(g27258),.B(g20008));
  AND2 AND2_1880(.VSS(VSS),.VDD(VDD),.Y(g24681),.A(g16653),.B(g22988));
  AND2 AND2_1881(.VSS(VSS),.VDD(VDD),.Y(g29178),.A(g27163),.B(g12687));
  AND2 AND2_1882(.VSS(VSS),.VDD(VDD),.Y(g29740),.A(g2648),.B(g29154));
  AND2 AND2_1883(.VSS(VSS),.VDD(VDD),.Y(g30005),.A(g28230),.B(g24394));
  AND2 AND2_1884(.VSS(VSS),.VDD(VDD),.Y(g22126),.A(g6621),.B(g19277));
  AND2 AND2_1885(.VSS(VSS),.VDD(VDD),.Y(g18128),.A(g504),.B(g16971));
  AND2 AND2_1886(.VSS(VSS),.VDD(VDD),.Y(g21927),.A(g5164),.B(g18997));
  AND2 AND2_1887(.VSS(VSS),.VDD(VDD),.Y(g26100),.A(g1677),.B(g25097));
  AND2 AND2_1888(.VSS(VSS),.VDD(VDD),.Y(g19588),.A(g3849),.B(g16853));
  AND2 AND2_1889(.VSS(VSS),.VDD(VDD),.Y(g33416),.A(g32370),.B(g21423));
  AND2 AND2_1890(.VSS(VSS),.VDD(VDD),.Y(g29685),.A(g2084),.B(g28711));
  AND4 AND4_122(.VSS(VSS),.VDD(VDD),.Y(I31326),.A(g30735),.B(g31853),.C(g32926),.D(g32927));
  AND2 AND2_1891(.VSS(VSS),.VDD(VDD),.Y(g18245),.A(g1193),.B(g16431));
  AND2 AND2_1892(.VSS(VSS),.VDD(VDD),.Y(g27132),.A(g26055),.B(g16589));
  AND2 AND2_1893(.VSS(VSS),.VDD(VDD),.Y(g34538),.A(g34330),.B(g20054));
  AND2 AND2_1894(.VSS(VSS),.VDD(VDD),.Y(g18626),.A(g3498),.B(g17062));
  AND2 AND2_1895(.VSS(VSS),.VDD(VDD),.Y(g15913),.A(g3933),.B(g14021));
  AND2 AND2_1896(.VSS(VSS),.VDD(VDD),.Y(g24730),.A(g6177),.B(g23699));
  AND2 AND2_1897(.VSS(VSS),.VDD(VDD),.Y(g31992),.A(g31773),.B(g22213));
  AND2 AND2_1898(.VSS(VSS),.VDD(VDD),.Y(g18323),.A(g1632),.B(g17873));
  AND2 AND2_1899(.VSS(VSS),.VDD(VDD),.Y(g33841),.A(g33254),.B(g20268));
  AND2 AND2_1900(.VSS(VSS),.VDD(VDD),.Y(g18299),.A(g1526),.B(g16489));
  AND2 AND2_1901(.VSS(VSS),.VDD(VDD),.Y(g18533),.A(g2729),.B(g15277));
  AND2 AND2_1902(.VSS(VSS),.VDD(VDD),.Y(g28547),.A(g6821),.B(g27091));
  AND3 AND3_112(.VSS(VSS),.VDD(VDD),.Y(g33510),.A(g32816),.B(I31246),.C(I31247));
  AND2 AND2_1903(.VSS(VSS),.VDD(VDD),.Y(g24765),.A(g17699),.B(g22498));
  AND2 AND2_1904(.VSS(VSS),.VDD(VDD),.Y(g18298),.A(g15073),.B(g16489));
  AND3 AND3_113(.VSS(VSS),.VDD(VDD),.Y(g27161),.A(g26166),.B(g8241),.C(g1783));
  AND2 AND2_1905(.VSS(VSS),.VDD(VDD),.Y(g30241),.A(g28729),.B(g23926));
  AND4 AND4_123(.VSS(VSS),.VDD(VDD),.Y(I31252),.A(g32819),.B(g32820),.C(g32821),.D(g32822));
  AND2 AND2_1906(.VSS(VSS),.VDD(VDD),.Y(g31579),.A(g19128),.B(g29814));
  AND2 AND2_1907(.VSS(VSS),.VDD(VDD),.Y(g18775),.A(g7028),.B(g15615));
  AND2 AND2_1908(.VSS(VSS),.VDD(VDD),.Y(g24549),.A(g23162),.B(g20887));
  AND2 AND2_1909(.VSS(VSS),.VDD(VDD),.Y(g28226),.A(g27825),.B(g26667));
  AND2 AND2_1910(.VSS(VSS),.VDD(VDD),.Y(g21755),.A(g3203),.B(g20785));
  AND2 AND2_1911(.VSS(VSS),.VDD(VDD),.Y(g29334),.A(g29148),.B(g18908));
  AND2 AND2_1912(.VSS(VSS),.VDD(VDD),.Y(g16474),.A(g8280),.B(g13666));
  AND2 AND2_1913(.VSS(VSS),.VDD(VDD),.Y(g23755),.A(g14821),.B(g21204));
  AND2 AND2_1914(.VSS(VSS),.VDD(VDD),.Y(g27259),.A(g26755),.B(g26725));
  AND2 AND2_1915(.VSS(VSS),.VDD(VDD),.Y(g19749),.A(g732),.B(g16646));
  AND2 AND2_1916(.VSS(VSS),.VDD(VDD),.Y(g32047),.A(g27248),.B(g31070));
  AND2 AND2_1917(.VSS(VSS),.VDD(VDD),.Y(g33835),.A(g4340),.B(g33413));
  AND2 AND2_1918(.VSS(VSS),.VDD(VDD),.Y(g9968),.A(g1339),.B(g1500));
  AND2 AND2_1919(.VSS(VSS),.VDD(VDD),.Y(g21770),.A(g3251),.B(g20785));
  AND2 AND2_1920(.VSS(VSS),.VDD(VDD),.Y(g32205),.A(g30922),.B(g28463));
  AND2 AND2_1921(.VSS(VSS),.VDD(VDD),.Y(g21981),.A(g5543),.B(g19074));
  AND2 AND2_1922(.VSS(VSS),.VDD(VDD),.Y(g22060),.A(g6151),.B(g21611));
  AND2 AND2_1923(.VSS(VSS),.VDD(VDD),.Y(g10902),.A(g7858),.B(g1129));
  AND2 AND2_1924(.VSS(VSS),.VDD(VDD),.Y(g18737),.A(g4975),.B(g16826));
  AND2 AND2_1925(.VSS(VSS),.VDD(VDD),.Y(g27087),.A(g13872),.B(g26284));
  AND2 AND2_1926(.VSS(VSS),.VDD(VDD),.Y(g28572),.A(g27829),.B(g15669));
  AND2 AND2_1927(.VSS(VSS),.VDD(VDD),.Y(g12259),.A(g9480),.B(g640));
  AND2 AND2_1928(.VSS(VSS),.VDD(VDD),.Y(g24504),.A(g22226),.B(g19410));
  AND2 AND2_1929(.VSS(VSS),.VDD(VDD),.Y(g32311),.A(g31295),.B(g20582));
  AND2 AND2_1930(.VSS(VSS),.VDD(VDD),.Y(g25207),.A(g22513),.B(g10621));
  AND2 AND2_1931(.VSS(VSS),.VDD(VDD),.Y(g29762),.A(g28298),.B(g10233));
  AND2 AND2_1932(.VSS(VSS),.VDD(VDD),.Y(g18232),.A(g1124),.B(g16326));
  AND2 AND2_1933(.VSS(VSS),.VDD(VDD),.Y(g34771),.A(g34693),.B(g20147));
  AND2 AND2_1934(.VSS(VSS),.VDD(VDD),.Y(g29964),.A(g2008),.B(g28830));
  AND2 AND2_1935(.VSS(VSS),.VDD(VDD),.Y(g16537),.A(g5937),.B(g14855));
  AND2 AND2_1936(.VSS(VSS),.VDD(VDD),.Y(g11027),.A(g5097),.B(g9724));
  AND2 AND2_1937(.VSS(VSS),.VDD(VDD),.Y(g30235),.A(g28723),.B(g23915));
  AND3 AND3_114(.VSS(VSS),.VDD(VDD),.Y(I18713),.A(g13156),.B(g6767),.C(g6756));
  AND3 AND3_115(.VSS(VSS),.VDD(VDD),.Y(g25328),.A(g5022),.B(g23764),.C(I24505));
  AND2 AND2_1938(.VSS(VSS),.VDD(VDD),.Y(g11890),.A(g7499),.B(g9155));
  AND2 AND2_1939(.VSS(VSS),.VDD(VDD),.Y(g24317),.A(g4534),.B(g22228));
  AND2 AND2_1940(.VSS(VSS),.VDD(VDD),.Y(g15797),.A(g3909),.B(g14139));
  AND2 AND2_1941(.VSS(VSS),.VDD(VDD),.Y(g18697),.A(g4749),.B(g16777));
  AND2 AND2_1942(.VSS(VSS),.VDD(VDD),.Y(g27043),.A(g26335),.B(g8632));
  AND2 AND2_1943(.VSS(VSS),.VDD(VDD),.Y(g32051),.A(g31506),.B(g10831));
  AND4 AND4_124(.VSS(VSS),.VDD(VDD),.Y(g16283),.A(g11547),.B(g11592),.C(g6789),.D(I17606));
  AND2 AND2_1944(.VSS(VSS),.VDD(VDD),.Y(g29587),.A(g2181),.B(g28935));
  AND4 AND4_125(.VSS(VSS),.VDD(VDD),.Y(I31062),.A(g32545),.B(g32546),.C(g32547),.D(g32548));
  AND2 AND2_1945(.VSS(VSS),.VDD(VDD),.Y(g18261),.A(g1256),.B(g16000));
  AND2 AND2_1946(.VSS(VSS),.VDD(VDD),.Y(g21767),.A(g3239),.B(g20785));
  AND2 AND2_1947(.VSS(VSS),.VDD(VDD),.Y(g21794),.A(g15094),.B(g20924));
  AND2 AND2_1948(.VSS(VSS),.VDD(VDD),.Y(g21845),.A(g3881),.B(g21070));
  AND2 AND2_1949(.VSS(VSS),.VDD(VDD),.Y(g12043),.A(g1345),.B(g7601));
  AND2 AND2_1950(.VSS(VSS),.VDD(VDD),.Y(g16303),.A(g4527),.B(g12921));
  AND2 AND2_1951(.VSS(VSS),.VDD(VDD),.Y(g10290),.A(g4358),.B(g4349));
  AND2 AND2_1952(.VSS(VSS),.VDD(VDD),.Y(g24002),.A(g19613),.B(g10971));
  AND2 AND2_1953(.VSS(VSS),.VDD(VDD),.Y(g21990),.A(g5591),.B(g19074));
  AND2 AND2_1954(.VSS(VSS),.VDD(VDD),.Y(g11003),.A(g7880),.B(g1300));
  AND2 AND2_1955(.VSS(VSS),.VDD(VDD),.Y(g18512),.A(g2619),.B(g15509));
  AND2 AND2_1956(.VSS(VSS),.VDD(VDD),.Y(g23990),.A(g19610),.B(g10951));
  AND4 AND4_126(.VSS(VSS),.VDD(VDD),.Y(I27524),.A(g28037),.B(g24114),.C(g24115),.D(g24116));
  AND2 AND2_1957(.VSS(VSS),.VDD(VDD),.Y(g33720),.A(g33161),.B(g19439));
  AND3 AND3_116(.VSS(VSS),.VDD(VDD),.Y(g19560),.A(g15832),.B(g1157),.C(g10893));
  AND2 AND2_1958(.VSS(VSS),.VDD(VDD),.Y(g29909),.A(g28435),.B(g23388));
  AND4 AND4_127(.VSS(VSS),.VDD(VDD),.Y(g27602),.A(g23032),.B(g26244),.C(g26424),.D(g24966));
  AND2 AND2_1959(.VSS(VSS),.VDD(VDD),.Y(g31275),.A(g30147),.B(g27800));
  AND2 AND2_1960(.VSS(VSS),.VDD(VDD),.Y(g34515),.A(g34288),.B(g19491));
  AND2 AND2_1961(.VSS(VSS),.VDD(VDD),.Y(g34414),.A(g34206),.B(g21457));
  AND4 AND4_128(.VSS(VSS),.VDD(VDD),.Y(g28889),.A(g17292),.B(g25169),.C(g26424),.D(g27395));
  AND2 AND2_1962(.VSS(VSS),.VDD(VDD),.Y(g31746),.A(g30093),.B(g23905));
  AND2 AND2_1963(.VSS(VSS),.VDD(VDD),.Y(g27375),.A(g26519),.B(g17479));
  AND2 AND2_1964(.VSS(VSS),.VDD(VDD),.Y(g26206),.A(g2523),.B(g25495));
  AND2 AND2_1965(.VSS(VSS),.VDD(VDD),.Y(g31493),.A(g29791),.B(g23434));
  AND2 AND2_1966(.VSS(VSS),.VDD(VDD),.Y(g32350),.A(g2697),.B(g31710));
  AND2 AND2_1967(.VSS(VSS),.VDD(VDD),.Y(g21719),.A(g358),.B(g21037));
  AND3 AND3_117(.VSS(VSS),.VDD(VDD),.Y(g33493),.A(g32693),.B(I31161),.C(I31162));
  AND2 AND2_1968(.VSS(VSS),.VDD(VDD),.Y(g24323),.A(g4546),.B(g22228));
  AND2 AND2_1969(.VSS(VSS),.VDD(VDD),.Y(g24299),.A(g4456),.B(g22550));
  AND2 AND2_1970(.VSS(VSS),.VDD(VDD),.Y(g13778),.A(g4540),.B(g10597));
  AND2 AND2_1971(.VSS(VSS),.VDD(VDD),.Y(g13081),.A(g8626),.B(g11122));
  AND2 AND2_1972(.VSS(VSS),.VDD(VDD),.Y(g29569),.A(g29028),.B(g22498));
  AND2 AND2_1973(.VSS(VSS),.VDD(VDD),.Y(g21718),.A(g370),.B(g21037));
  AND3 AND3_118(.VSS(VSS),.VDD(VDD),.Y(g33465),.A(g32491),.B(I31021),.C(I31022));
  AND2 AND2_1974(.VSS(VSS),.VDD(VDD),.Y(g31237),.A(g29366),.B(g25325));
  AND3 AND3_119(.VSS(VSS),.VDD(VDD),.Y(g10632),.A(g7475),.B(g7441),.C(g890));
  AND2 AND2_1975(.VSS(VSS),.VDD(VDD),.Y(g24298),.A(g4392),.B(g22550));
  AND2 AND2_1976(.VSS(VSS),.VDD(VDD),.Y(g33237),.A(g32394),.B(g25198));
  AND2 AND2_1977(.VSS(VSS),.VDD(VDD),.Y(g32152),.A(g31631),.B(g29998));
  AND2 AND2_1978(.VSS(VSS),.VDD(VDD),.Y(g18445),.A(g2273),.B(g18008));
  AND2 AND2_1979(.VSS(VSS),.VDD(VDD),.Y(g24775),.A(g17594),.B(g22498));
  AND2 AND2_1980(.VSS(VSS),.VDD(VDD),.Y(g29568),.A(g2571),.B(g28950));
  AND2 AND2_1981(.VSS(VSS),.VDD(VDD),.Y(g29747),.A(g28286),.B(g23196));
  AND2 AND2_1982(.VSS(VSS),.VDD(VDD),.Y(g32396),.A(g4698),.B(g30983));
  AND2 AND2_1983(.VSS(VSS),.VDD(VDD),.Y(g33340),.A(g32222),.B(g20639));
  AND2 AND2_1984(.VSS(VSS),.VDD(VDD),.Y(g21832),.A(g3787),.B(g20453));
  AND2 AND2_1985(.VSS(VSS),.VDD(VDD),.Y(g18499),.A(g2476),.B(g15426));
  AND2 AND2_1986(.VSS(VSS),.VDD(VDD),.Y(g18316),.A(g1564),.B(g16931));
  AND2 AND2_1987(.VSS(VSS),.VDD(VDD),.Y(g33684),.A(g33139),.B(g13565));
  AND2 AND2_1988(.VSS(VSS),.VDD(VDD),.Y(g16840),.A(g5467),.B(g14262));
  AND2 AND2_1989(.VSS(VSS),.VDD(VDD),.Y(g31142),.A(g2527),.B(g30039));
  AND2 AND2_1990(.VSS(VSS),.VDD(VDD),.Y(g22055),.A(g6128),.B(g21611));
  AND2 AND2_1991(.VSS(VSS),.VDD(VDD),.Y(g18498),.A(g2547),.B(g15426));
  AND2 AND2_1992(.VSS(VSS),.VDD(VDD),.Y(g32413),.A(g31121),.B(g19518));
  AND2 AND2_1993(.VSS(VSS),.VDD(VDD),.Y(g19693),.A(g6181),.B(g17087));
  AND2 AND2_1994(.VSS(VSS),.VDD(VDD),.Y(g22111),.A(g6549),.B(g19277));
  AND4 AND4_129(.VSS(VSS),.VDD(VDD),.Y(I31047),.A(g32524),.B(g32525),.C(g32526),.D(g32527));
  AND2 AND2_1995(.VSS(VSS),.VDD(VDD),.Y(g21861),.A(g3949),.B(g21070));
  AND2 AND2_1996(.VSS(VSS),.VDD(VDD),.Y(g34584),.A(g24653),.B(g34315));
  AND2 AND2_1997(.VSS(VSS),.VDD(VDD),.Y(g22070),.A(g6243),.B(g19210));
  AND2 AND2_1998(.VSS(VSS),.VDD(VDD),.Y(g13998),.A(g6589),.B(g12629));
  AND2 AND2_1999(.VSS(VSS),.VDD(VDD),.Y(g31517),.A(g29849),.B(g23482));
  AND2 AND2_2000(.VSS(VSS),.VDD(VDD),.Y(g26345),.A(g13051),.B(g25505));
  AND2 AND2_2001(.VSS(VSS),.VDD(VDD),.Y(g28426),.A(g27257),.B(g20006));
  AND3 AND3_120(.VSS(VSS),.VDD(VDD),.Y(g33517),.A(g32867),.B(I31281),.C(I31282));
  AND2 AND2_2002(.VSS(VSS),.VDD(VDD),.Y(g29751),.A(g28297),.B(g23216));
  AND2 AND2_2003(.VSS(VSS),.VDD(VDD),.Y(g29807),.A(g28359),.B(g23272));
  AND4 AND4_130(.VSS(VSS),.VDD(VDD),.Y(I31311),.A(g30673),.B(g31851),.C(g32903),.D(g32904));
  AND2 AND2_2004(.VSS(VSS),.VDD(VDD),.Y(g29772),.A(g28323),.B(g23243));
  AND2 AND2_2005(.VSS(VSS),.VDD(VDD),.Y(g22590),.A(g19274),.B(g19452));
  AND2 AND2_2006(.VSS(VSS),.VDD(VDD),.Y(g16192),.A(g6191),.B(g14321));
  AND2 AND2_2007(.VSS(VSS),.VDD(VDD),.Y(g26849),.A(g2994),.B(g24527));
  AND2 AND2_2008(.VSS(VSS),.VDD(VDD),.Y(g29974),.A(g29173),.B(g12914));
  AND2 AND2_2009(.VSS(VSS),.VDD(VDD),.Y(g15711),.A(g460),.B(g13437));
  AND2 AND2_2010(.VSS(VSS),.VDD(VDD),.Y(g18611),.A(g15090),.B(g17200));
  AND2 AND2_2011(.VSS(VSS),.VDD(VDD),.Y(g27459),.A(g26549),.B(g17609));
  AND2 AND2_2012(.VSS(VSS),.VDD(VDD),.Y(g21926),.A(g15147),.B(g18997));
  AND2 AND2_2013(.VSS(VSS),.VDD(VDD),.Y(g18722),.A(g4917),.B(g16077));
  AND2 AND2_2014(.VSS(VSS),.VDD(VDD),.Y(g26399),.A(g15572),.B(g25566));
  AND3 AND3_121(.VSS(VSS),.VDD(VDD),.Y(g25414),.A(g5406),.B(g22194),.C(I24549));
  AND2 AND2_2015(.VSS(VSS),.VDD(VDD),.Y(g25991),.A(g2060),.B(g25023));
  AND2 AND2_2016(.VSS(VSS),.VDD(VDD),.Y(g23389),.A(g9072),.B(g19757));
  AND2 AND2_2017(.VSS(VSS),.VDD(VDD),.Y(g29639),.A(g28510),.B(g11618));
  AND2 AND2_2018(.VSS(VSS),.VDD(VDD),.Y(g15109),.A(g4269),.B(g14454));
  AND2 AND2_2019(.VSS(VSS),.VDD(VDD),.Y(g26848),.A(g2950),.B(g24526));
  AND3 AND3_122(.VSS(VSS),.VDD(VDD),.Y(I16646),.A(g10160),.B(g12413),.C(g12343));
  AND2 AND2_2020(.VSS(VSS),.VDD(VDD),.Y(g26398),.A(g24946),.B(g10474));
  AND3 AND3_123(.VSS(VSS),.VDD(VDD),.Y(g22384),.A(g9354),.B(g9285),.C(g20784));
  AND2 AND2_2021(.VSS(VSS),.VDD(VDD),.Y(g18432),.A(g2223),.B(g18008));
  AND4 AND4_131(.VSS(VSS),.VDD(VDD),.Y(I24705),.A(g24064),.B(g24065),.C(g24066),.D(g24067));
  AND2 AND2_2022(.VSS(VSS),.VDD(VDD),.Y(g29638),.A(g2583),.B(g29025));
  AND4 AND4_132(.VSS(VSS),.VDD(VDD),.Y(I31051),.A(g31376),.B(g31804),.C(g32529),.D(g32530));
  AND2 AND2_2023(.VSS(VSS),.VDD(VDD),.Y(g21701),.A(g153),.B(g20283));
  AND4 AND4_133(.VSS(VSS),.VDD(VDD),.Y(I31072),.A(g32559),.B(g32560),.C(g32561),.D(g32562));
  AND2 AND2_2024(.VSS(VSS),.VDD(VDD),.Y(g18271),.A(g1296),.B(g16031));
  AND2 AND2_2025(.VSS(VSS),.VDD(VDD),.Y(g30082),.A(g29181),.B(g12752));
  AND2 AND2_2026(.VSS(VSS),.VDD(VDD),.Y(g34114),.A(g33920),.B(g23742));
  AND2 AND2_2027(.VSS(VSS),.VDD(VDD),.Y(g15108),.A(g4264),.B(g14454));
  AND2 AND2_2028(.VSS(VSS),.VDD(VDD),.Y(g21777),.A(g3380),.B(g20391));
  AND2 AND2_2029(.VSS(VSS),.VDD(VDD),.Y(g34758),.A(g34683),.B(g19657));
  AND2 AND2_2030(.VSS(VSS),.VDD(VDD),.Y(g26652),.A(g10799),.B(g24426));
  AND2 AND2_2031(.VSS(VSS),.VDD(VDD),.Y(g31130),.A(g12191),.B(g30019));
  AND2 AND2_2032(.VSS(VSS),.VDD(VDD),.Y(g22067),.A(g6215),.B(g19210));
  AND2 AND2_2033(.VSS(VSS),.VDD(VDD),.Y(g22094),.A(g6398),.B(g18833));
  AND2 AND2_2034(.VSS(VSS),.VDD(VDD),.Y(g34082),.A(g33709),.B(g19554));
  AND2 AND2_2035(.VSS(VSS),.VDD(VDD),.Y(g30107),.A(g28560),.B(g20909));
  AND2 AND2_2036(.VSS(VSS),.VDD(VDD),.Y(g21251),.A(g13969),.B(g17470));
  AND4 AND4_134(.VSS(VSS),.VDD(VDD),.Y(I24679),.A(g19968),.B(g24026),.C(g24027),.D(g24028));
  AND2 AND2_2037(.VSS(VSS),.VDD(VDD),.Y(g33362),.A(g32259),.B(g20914));
  AND2 AND2_2038(.VSS(VSS),.VDD(VDD),.Y(g11449),.A(g6052),.B(g7175));
  AND2 AND2_2039(.VSS(VSS),.VDD(VDD),.Y(g27545),.A(g26519),.B(g17756));
  AND2 AND2_2040(.VSS(VSS),.VDD(VDD),.Y(g16483),.A(g5224),.B(g14915));
  AND2 AND2_2041(.VSS(VSS),.VDD(VDD),.Y(g18753),.A(g15148),.B(g15595));
  AND2 AND2_2042(.VSS(VSS),.VDD(VDD),.Y(g18461),.A(g2307),.B(g15224));
  AND2 AND2_2043(.VSS(VSS),.VDD(VDD),.Y(g31523),.A(g7528),.B(g29333));
  AND2 AND2_2044(.VSS(VSS),.VDD(VDD),.Y(g32020),.A(g4157),.B(g30937));
  AND2 AND2_2045(.VSS(VSS),.VDD(VDD),.Y(g18342),.A(g1592),.B(g17873));
  AND3 AND3_124(.VSS(VSS),.VDD(VDD),.Y(g33523),.A(g32909),.B(I31311),.C(I31312));
  AND2 AND2_2046(.VSS(VSS),.VDD(VDD),.Y(g29841),.A(g28371),.B(g23283));
  AND2 AND2_2047(.VSS(VSS),.VDD(VDD),.Y(g19914),.A(g2815),.B(g15853));
  AND2 AND2_2048(.VSS(VSS),.VDD(VDD),.Y(g29992),.A(g29012),.B(g10490));
  AND2 AND2_2049(.VSS(VSS),.VDD(VDD),.Y(g27599),.A(g26337),.B(g20033));
  AND2 AND2_2050(.VSS(VSS),.VDD(VDD),.Y(g34744),.A(g34668),.B(g19481));
  AND2 AND2_2051(.VSS(VSS),.VDD(VDD),.Y(g18145),.A(g582),.B(g17533));
  AND2 AND2_2052(.VSS(VSS),.VDD(VDD),.Y(g29510),.A(g28856),.B(g22342));
  AND2 AND2_2053(.VSS(VSS),.VDD(VDD),.Y(g32046),.A(g10925),.B(g30735));
  AND2 AND2_2054(.VSS(VSS),.VDD(VDD),.Y(g18199),.A(g832),.B(g17821));
  AND2 AND2_2055(.VSS(VSS),.VDD(VDD),.Y(g22019),.A(g5857),.B(g19147));
  AND2 AND2_2056(.VSS(VSS),.VDD(VDD),.Y(g27598),.A(g25899),.B(g10475));
  AND2 AND2_2057(.VSS(VSS),.VDD(VDD),.Y(g18650),.A(g6928),.B(g17271));
  AND2 AND2_2058(.VSS(VSS),.VDD(VDD),.Y(g18736),.A(g4991),.B(g16826));
  AND2 AND2_2059(.VSS(VSS),.VDD(VDD),.Y(g27086),.A(g25836),.B(g22495));
  AND2 AND2_2060(.VSS(VSS),.VDD(VDD),.Y(g31475),.A(g29756),.B(g23406));
  AND2 AND2_2061(.VSS(VSS),.VDD(VDD),.Y(g29579),.A(g28457),.B(g7964));
  AND2 AND2_2062(.VSS(VSS),.VDD(VDD),.Y(g17150),.A(g8579),.B(g12995));
  AND3 AND3_125(.VSS(VSS),.VDD(VDD),.Y(I24030),.A(g8390),.B(g8016),.C(g3396));
  AND3 AND3_126(.VSS(VSS),.VDD(VDD),.Y(g33475),.A(g32563),.B(I31071),.C(I31072));
  AND2 AND2_2063(.VSS(VSS),.VDD(VDD),.Y(g16536),.A(g5917),.B(g14996));
  AND2 AND2_2064(.VSS(VSS),.VDD(VDD),.Y(g18198),.A(g15059),.B(g17821));
  AND2 AND2_2065(.VSS(VSS),.VDD(VDD),.Y(g22018),.A(g15157),.B(g19147));
  AND2 AND2_2066(.VSS(VSS),.VDD(VDD),.Y(g18529),.A(g2712),.B(g15277));
  AND2 AND2_2067(.VSS(VSS),.VDD(VDD),.Y(g21997),.A(g5619),.B(g19074));
  AND2 AND2_2068(.VSS(VSS),.VDD(VDD),.Y(g32113),.A(g31601),.B(g29925));
  AND2 AND2_2069(.VSS(VSS),.VDD(VDD),.Y(g34398),.A(g7684),.B(g34070));
  AND4 AND4_135(.VSS(VSS),.VDD(VDD),.Y(I31152),.A(g32675),.B(g32676),.C(g32677),.D(g32678));
  AND2 AND2_2070(.VSS(VSS),.VDD(VDD),.Y(g33727),.A(g33115),.B(g19499));
  AND2 AND2_2071(.VSS(VSS),.VDD(VDD),.Y(g24499),.A(g22217),.B(g19394));
  AND2 AND2_2072(.VSS(VSS),.VDD(VDD),.Y(g29578),.A(g2491),.B(g28606));
  AND2 AND2_2073(.VSS(VSS),.VDD(VDD),.Y(g33863),.A(g33273),.B(g20505));
  AND2 AND2_2074(.VSS(VSS),.VDD(VDD),.Y(g19594),.A(g11913),.B(g17268));
  AND2 AND2_2075(.VSS(VSS),.VDD(VDD),.Y(g29835),.A(g28326),.B(g24866));
  AND2 AND2_2076(.VSS(VSS),.VDD(VDD),.Y(g34141),.A(g33932),.B(g23828));
  AND2 AND2_2077(.VSS(VSS),.VDD(VDD),.Y(g16702),.A(g5615),.B(g14691));
  AND2 AND2_2078(.VSS(VSS),.VDD(VDD),.Y(g24316),.A(g4527),.B(g22228));
  AND2 AND2_2079(.VSS(VSS),.VDD(VDD),.Y(g31222),.A(g2643),.B(g30113));
  AND2 AND2_2080(.VSS(VSS),.VDD(VDD),.Y(g32282),.A(g31258),.B(g20503));
  AND4 AND4_136(.VSS(VSS),.VDD(VDD),.Y(g27817),.A(g22498),.B(g25245),.C(g26424),.D(g26236));
  AND2 AND2_2081(.VSS(VSS),.VDD(VDD),.Y(g15796),.A(g3586),.B(g14015));
  AND2 AND2_2082(.VSS(VSS),.VDD(VDD),.Y(g18696),.A(g4741),.B(g16053));
  AND2 AND2_2083(.VSS(VSS),.VDD(VDD),.Y(g18330),.A(g1668),.B(g17873));
  AND2 AND2_2084(.VSS(VSS),.VDD(VDD),.Y(g32302),.A(g31279),.B(g23485));
  AND2 AND2_2085(.VSS(VSS),.VDD(VDD),.Y(g18393),.A(g1917),.B(g15171));
  AND2 AND2_2086(.VSS(VSS),.VDD(VDD),.Y(g24498),.A(g14036),.B(g23850));
  AND2 AND2_2087(.VSS(VSS),.VDD(VDD),.Y(g29586),.A(g1886),.B(g28927));
  AND2 AND2_2088(.VSS(VSS),.VDD(VDD),.Y(g16621),.A(g8278),.B(g13821));
  AND2 AND2_2089(.VSS(VSS),.VDD(VDD),.Y(g12817),.A(g1351),.B(g7601));
  AND2 AND2_2090(.VSS(VSS),.VDD(VDD),.Y(g21766),.A(g3235),.B(g20785));
  AND2 AND2_2091(.VSS(VSS),.VDD(VDD),.Y(g26833),.A(g2852),.B(g24509));
  AND2 AND2_2092(.VSS(VSS),.VDD(VDD),.Y(g26049),.A(g9621),.B(g25046));
  AND2 AND2_2093(.VSS(VSS),.VDD(VDD),.Y(g30263),.A(g28773),.B(g23962));
  AND2 AND2_2094(.VSS(VSS),.VDD(VDD),.Y(g32105),.A(g4922),.B(g30673));
  AND2 AND2_2095(.VSS(VSS),.VDD(VDD),.Y(g28658),.A(g27563),.B(g20611));
  AND2 AND2_2096(.VSS(VSS),.VDD(VDD),.Y(g18764),.A(g5485),.B(g17929));
  AND4 AND4_137(.VSS(VSS),.VDD(VDD),.Y(g20056),.A(g16291),.B(g9007),.C(g8954),.D(g8903));
  AND2 AND2_2097(.VSS(VSS),.VDD(VDD),.Y(g18365),.A(g1848),.B(g17955));
  AND2 AND2_2098(.VSS(VSS),.VDD(VDD),.Y(g27158),.A(g26609),.B(g16645));
  AND2 AND2_2099(.VSS(VSS),.VDD(VDD),.Y(g21871),.A(g4108),.B(g19801));
  AND2 AND2_2100(.VSS(VSS),.VDD(VDD),.Y(g25107),.A(g17643),.B(g23508));
  AND3 AND3_127(.VSS(VSS),.VDD(VDD),.Y(g22457),.A(g7753),.B(g7717),.C(g21288));
  AND2 AND2_2101(.VSS(VSS),.VDD(VDD),.Y(g15840),.A(g3949),.B(g14142));
  AND2 AND2_2102(.VSS(VSS),.VDD(VDD),.Y(g18132),.A(g513),.B(g16971));
  AND2 AND2_2103(.VSS(VSS),.VDD(VDD),.Y(g26048),.A(g5853),.B(g25044));
  AND2 AND2_2104(.VSS(VSS),.VDD(VDD),.Y(g28339),.A(g9946),.B(g27693));
  AND2 AND2_2105(.VSS(VSS),.VDD(VDD),.Y(g30135),.A(g28592),.B(g21180));
  AND2 AND2_2106(.VSS(VSS),.VDD(VDD),.Y(g24722),.A(g17618),.B(g22417));
  AND2 AND2_2107(.VSS(VSS),.VDD(VDD),.Y(g34135),.A(g33926),.B(g23802));
  AND3 AND3_128(.VSS(VSS),.VDD(VDD),.Y(I18782),.A(g13156),.B(g11450),.C(g6756));
  AND2 AND2_2108(.VSS(VSS),.VDD(VDD),.Y(g7948),.A(g1548),.B(g1430));
  AND2 AND2_2109(.VSS(VSS),.VDD(VDD),.Y(g29615),.A(g1844),.B(g29049));
  AND2 AND2_2110(.VSS(VSS),.VDD(VDD),.Y(g16673),.A(g6617),.B(g14822));
  AND2 AND2_2111(.VSS(VSS),.VDD(VDD),.Y(g18161),.A(g691),.B(g17433));
  AND2 AND2_2112(.VSS(VSS),.VDD(VDD),.Y(g34962),.A(g34945),.B(g23020));
  AND2 AND2_2113(.VSS(VSS),.VDD(VDD),.Y(g19637),.A(g5142),.B(g16958));
  AND2 AND2_2114(.VSS(VSS),.VDD(VDD),.Y(g26613),.A(g1361),.B(g24518));
  AND2 AND2_2115(.VSS(VSS),.VDD(VDD),.Y(g18709),.A(g59),.B(g17302));
  AND2 AND2_2116(.VSS(VSS),.VDD(VDD),.Y(g22001),.A(g5731),.B(g21562));
  AND2 AND2_2117(.VSS(VSS),.VDD(VDD),.Y(g22077),.A(g6263),.B(g19210));
  AND2 AND2_2118(.VSS(VSS),.VDD(VDD),.Y(g25848),.A(g25539),.B(g18977));
  AND2 AND2_2119(.VSS(VSS),.VDD(VDD),.Y(g14190),.A(g859),.B(g10632));
  AND2 AND2_2120(.VSS(VSS),.VDD(VDD),.Y(g27336),.A(g2675),.B(g26777));
  AND2 AND2_2121(.VSS(VSS),.VDD(VDD),.Y(g30049),.A(g13114),.B(g28167));
  AND2 AND2_2122(.VSS(VSS),.VDD(VDD),.Y(g18259),.A(g15068),.B(g16000));
  AND2 AND2_2123(.VSS(VSS),.VDD(VDD),.Y(g29746),.A(g28279),.B(g20037));
  AND2 AND2_2124(.VSS(VSS),.VDD(VDD),.Y(g34500),.A(g34276),.B(g30568));
  AND2 AND2_2125(.VSS(VSS),.VDD(VDD),.Y(g18225),.A(g1041),.B(g16100));
  AND2 AND2_2126(.VSS(VSS),.VDD(VDD),.Y(g33351),.A(g32236),.B(g20707));
  AND2 AND2_2127(.VSS(VSS),.VDD(VDD),.Y(g33372),.A(g32285),.B(g21183));
  AND2 AND2_2128(.VSS(VSS),.VDD(VDD),.Y(g18708),.A(g4818),.B(g16782));
  AND2 AND2_2129(.VSS(VSS),.VDD(VDD),.Y(g28197),.A(g27647),.B(g11344));
  AND2 AND2_2130(.VSS(VSS),.VDD(VDD),.Y(g25804),.A(g8069),.B(g24587));
  AND2 AND2_2131(.VSS(VSS),.VDD(VDD),.Y(g18471),.A(g2407),.B(g15224));
  AND2 AND2_2132(.VSS(VSS),.VDD(VDD),.Y(g33821),.A(g33238),.B(g20153));
  AND2 AND2_2133(.VSS(VSS),.VDD(VDD),.Y(g26273),.A(g2122),.B(g25389));
  AND2 AND2_2134(.VSS(VSS),.VDD(VDD),.Y(g30048),.A(g29193),.B(g12945));
  AND2 AND2_2135(.VSS(VSS),.VDD(VDD),.Y(g22689),.A(g18918),.B(g9104));
  AND2 AND2_2136(.VSS(VSS),.VDD(VDD),.Y(g18258),.A(g1221),.B(g16897));
  AND2 AND2_2137(.VSS(VSS),.VDD(VDD),.Y(g16634),.A(g5264),.B(g14953));
  AND2 AND2_2138(.VSS(VSS),.VDD(VDD),.Y(g20887),.A(g16282),.B(g4864));
  AND2 AND2_2139(.VSS(VSS),.VDD(VDD),.Y(g23451),.A(g13805),.B(g20510));
  AND2 AND2_2140(.VSS(VSS),.VDD(VDD),.Y(g24199),.A(g355),.B(g22722));
  AND2 AND2_2141(.VSS(VSS),.VDD(VDD),.Y(g24650),.A(g22641),.B(g19718));
  AND2 AND2_2142(.VSS(VSS),.VDD(VDD),.Y(g23220),.A(g19417),.B(g20067));
  AND3 AND3_129(.VSS(VSS),.VDD(VDD),.Y(g24887),.A(g3712),.B(g23239),.C(I24054));
  AND2 AND2_2143(.VSS(VSS),.VDD(VDD),.Y(g30004),.A(g28521),.B(g25837));
  AND4 AND4_138(.VSS(VSS),.VDD(VDD),.Y(I31046),.A(g29385),.B(g32521),.C(g32522),.D(g32523));
  AND2 AND2_2144(.VSS(VSS),.VDD(VDD),.Y(g22624),.A(g19344),.B(g19471));
  AND2 AND2_2145(.VSS(VSS),.VDD(VDD),.Y(g21911),.A(g5046),.B(g21468));
  AND2 AND2_2146(.VSS(VSS),.VDD(VDD),.Y(g30221),.A(g28700),.B(g23893));
  AND2 AND2_2147(.VSS(VSS),.VDD(VDD),.Y(g31790),.A(g21299),.B(g29385));
  AND2 AND2_2148(.VSS(VSS),.VDD(VDD),.Y(g33264),.A(g31965),.B(g21306));
  AND2 AND2_2149(.VSS(VSS),.VDD(VDD),.Y(g31516),.A(g29848),.B(g23476));
  AND2 AND2_2150(.VSS(VSS),.VDD(VDD),.Y(g24198),.A(g351),.B(g22722));
  AND2 AND2_2151(.VSS(VSS),.VDD(VDD),.Y(g33790),.A(g33108),.B(g20643));
  AND3 AND3_130(.VSS(VSS),.VDD(VDD),.Y(g33516),.A(g32860),.B(I31276),.C(I31277));
  AND2 AND2_2152(.VSS(VSS),.VDD(VDD),.Y(g29806),.A(g28358),.B(g23271));
  AND2 AND2_2153(.VSS(VSS),.VDD(VDD),.Y(g29684),.A(g1982),.B(g29085));
  AND2 AND2_2154(.VSS(VSS),.VDD(VDD),.Y(g18244),.A(g1171),.B(g16431));
  AND2 AND2_2155(.VSS(VSS),.VDD(VDD),.Y(g26234),.A(g2657),.B(g25514));
  AND2 AND2_2156(.VSS(VSS),.VDD(VDD),.Y(g22102),.A(g6479),.B(g18833));
  AND3 AND3_131(.VSS(VSS),.VDD(VDD),.Y(g24843),.A(g3010),.B(g23211),.C(I24015));
  AND2 AND2_2157(.VSS(VSS),.VDD(VDD),.Y(g33873),.A(g33291),.B(g20549));
  AND2 AND2_2158(.VSS(VSS),.VDD(VDD),.Y(g24330),.A(g18661),.B(g22228));
  AND2 AND2_2159(.VSS(VSS),.VDD(VDD),.Y(g22157),.A(g14608),.B(g18892));
  AND2 AND2_2160(.VSS(VSS),.VDD(VDD),.Y(g24393),.A(g3808),.B(g22844));
  AND3 AND3_132(.VSS(VSS),.VDD(VDD),.Y(I24075),.A(g3736),.B(g3742),.C(g8553));
  AND4 AND4_139(.VSS(VSS),.VDD(VDD),.Y(I31282),.A(g32863),.B(g32864),.C(g32865),.D(g32866));
  AND2 AND2_2161(.VSS(VSS),.VDD(VDD),.Y(g25962),.A(g9258),.B(g24971));
  AND4 AND4_140(.VSS(VSS),.VDD(VDD),.Y(g16213),.A(g6772),.B(g6782),.C(g11640),.D(I17552));
  AND2 AND2_2162(.VSS(VSS),.VDD(VDD),.Y(g24764),.A(g17570),.B(g22472));
  AND2 AND2_2163(.VSS(VSS),.VDD(VDD),.Y(g29517),.A(g1870),.B(g28827));
  AND4 AND4_141(.VSS(VSS),.VDD(VDD),.Y(I31302),.A(g32891),.B(g32892),.C(g32893),.D(g32894));
  AND4 AND4_142(.VSS(VSS),.VDD(VDD),.Y(I31357),.A(g32970),.B(g32971),.C(g32972),.D(g32973));
  AND2 AND2_2164(.VSS(VSS),.VDD(VDD),.Y(g21776),.A(g3376),.B(g20391));
  AND2 AND2_2165(.VSS(VSS),.VDD(VDD),.Y(g21785),.A(g3431),.B(g20391));
  AND4 AND4_143(.VSS(VSS),.VDD(VDD),.Y(I27519),.A(g28036),.B(g24107),.C(g24108),.D(g24109));
  AND2 AND2_2166(.VSS(VSS),.VDD(VDD),.Y(g18602),.A(g3115),.B(g16987));
  AND2 AND2_2167(.VSS(VSS),.VDD(VDD),.Y(g18810),.A(g6505),.B(g15483));
  AND2 AND2_2168(.VSS(VSS),.VDD(VDD),.Y(g15757),.A(g3207),.B(g14066));
  AND2 AND2_2169(.VSS(VSS),.VDD(VDD),.Y(g18657),.A(g4308),.B(g17128));
  AND2 AND2_2170(.VSS(VSS),.VDD(VDD),.Y(g22066),.A(g6209),.B(g19210));
  AND2 AND2_2171(.VSS(VSS),.VDD(VDD),.Y(g18774),.A(g5698),.B(g15615));
  AND2 AND2_2172(.VSS(VSS),.VDD(VDD),.Y(g7918),.A(g1205),.B(g1087));
  AND2 AND2_2173(.VSS(VSS),.VDD(VDD),.Y(g18375),.A(g1902),.B(g15171));
  AND2 AND2_2174(.VSS(VSS),.VDD(VDD),.Y(g31209),.A(g2084),.B(g30097));
  AND2 AND2_2175(.VSS(VSS),.VDD(VDD),.Y(g33422),.A(g32375),.B(g21456));
  AND2 AND2_2176(.VSS(VSS),.VDD(VDD),.Y(g34106),.A(g33917),.B(g23675));
  AND2 AND2_2177(.VSS(VSS),.VDD(VDD),.Y(g32248),.A(g31616),.B(g30299));
  AND2 AND2_2178(.VSS(VSS),.VDD(VDD),.Y(g21754),.A(g3195),.B(g20785));
  AND4 AND4_144(.VSS(VSS),.VDD(VDD),.Y(I27518),.A(g20720),.B(g24104),.C(g24105),.D(g24106));
  AND2 AND2_2179(.VSS(VSS),.VDD(VDD),.Y(g10625),.A(g3431),.B(g7926));
  AND2 AND2_2180(.VSS(VSS),.VDD(VDD),.Y(g27309),.A(g26603),.B(g23057));
  AND2 AND2_2181(.VSS(VSS),.VDD(VDD),.Y(g23754),.A(g14816),.B(g21189));
  AND2 AND2_2182(.VSS(VSS),.VDD(VDD),.Y(g28714),.A(g27591),.B(g20711));
  AND3 AND3_133(.VSS(VSS),.VDD(VDD),.Y(g16047),.A(g13322),.B(g1500),.C(g10699));
  AND2 AND2_2183(.VSS(VSS),.VDD(VDD),.Y(g25833),.A(g8228),.B(g24626));
  AND2 AND2_2184(.VSS(VSS),.VDD(VDD),.Y(g14126),.A(g881),.B(g10632));
  AND4 AND4_145(.VSS(VSS),.VDD(VDD),.Y(g16205),.A(g11547),.B(g6782),.C(g11640),.D(I17542));
  AND2 AND2_2185(.VSS(VSS),.VDD(VDD),.Y(g27288),.A(g26515),.B(g23013));
  AND2 AND2_2186(.VSS(VSS),.VDD(VDD),.Y(g28315),.A(g27232),.B(g19769));
  AND2 AND2_2187(.VSS(VSS),.VDD(VDD),.Y(g33834),.A(g33095),.B(g29172));
  AND2 AND2_2188(.VSS(VSS),.VDD(VDD),.Y(g31208),.A(g30262),.B(g25188));
  AND2 AND2_2189(.VSS(VSS),.VDD(VDD),.Y(g32204),.A(g4245),.B(g31327));
  AND2 AND2_2190(.VSS(VSS),.VDD(VDD),.Y(g21859),.A(g3941),.B(g21070));
  AND2 AND2_2191(.VSS(VSS),.VDD(VDD),.Y(g21825),.A(g3736),.B(g20453));
  AND2 AND2_2192(.VSS(VSS),.VDD(VDD),.Y(g21950),.A(g5268),.B(g18997));
  AND2 AND2_2193(.VSS(VSS),.VDD(VDD),.Y(g26514),.A(g7400),.B(g25564));
  AND2 AND2_2194(.VSS(VSS),.VDD(VDD),.Y(g22876),.A(g20136),.B(g9104));
  AND2 AND2_2195(.VSS(VSS),.VDD(VDD),.Y(g18337),.A(g1706),.B(g17873));
  AND2 AND2_2196(.VSS(VSS),.VDD(VDD),.Y(g28202),.A(g27659),.B(g11413));
  AND2 AND2_2197(.VSS(VSS),.VDD(VDD),.Y(g30033),.A(g29189),.B(g12937));
  AND2 AND2_2198(.VSS(VSS),.VDD(VDD),.Y(g28257),.A(g27179),.B(g19686));
  AND2 AND2_2199(.VSS(VSS),.VDD(VDD),.Y(g21858),.A(g3937),.B(g21070));
  AND2 AND2_2200(.VSS(VSS),.VDD(VDD),.Y(g29362),.A(g27379),.B(g28307));
  AND2 AND2_2201(.VSS(VSS),.VDD(VDD),.Y(g18171),.A(g728),.B(g17433));
  AND2 AND2_2202(.VSS(VSS),.VDD(VDD),.Y(g30234),.A(g28721),.B(g23914));
  AND2 AND2_2203(.VSS(VSS),.VDD(VDD),.Y(g34371),.A(g7450),.B(g34044));
  AND2 AND2_2204(.VSS(VSS),.VDD(VDD),.Y(g24709),.A(g16690),.B(g23000));
  AND2 AND2_2205(.VSS(VSS),.VDD(VDD),.Y(g31542),.A(g19050),.B(g29814));
  AND2 AND2_2206(.VSS(VSS),.VDD(VDD),.Y(g31021),.A(g26025),.B(g29814));
  AND2 AND2_2207(.VSS(VSS),.VDD(VDD),.Y(g29523),.A(g28930),.B(g22417));
  AND2 AND2_2208(.VSS(VSS),.VDD(VDD),.Y(g23151),.A(g18994),.B(g7162));
  AND2 AND2_2209(.VSS(VSS),.VDD(VDD),.Y(g28111),.A(g27343),.B(g22716));
  AND2 AND2_2210(.VSS(VSS),.VDD(VDD),.Y(g14296),.A(g2638),.B(g11897));
  AND2 AND2_2211(.VSS(VSS),.VDD(VDD),.Y(g21996),.A(g5615),.B(g19074));
  AND2 AND2_2212(.VSS(VSS),.VDD(VDD),.Y(g24225),.A(g246),.B(g22594));
  AND2 AND2_2213(.VSS(VSS),.VDD(VDD),.Y(g15673),.A(g182),.B(g13437));
  AND2 AND2_2214(.VSS(VSS),.VDD(VDD),.Y(g18792),.A(g7051),.B(g15634));
  AND2 AND2_2215(.VSS(VSS),.VDD(VDD),.Y(g15847),.A(g3191),.B(g14005));
  AND2 AND2_2216(.VSS(VSS),.VDD(VDD),.Y(g23996),.A(g19596),.B(g10951));
  AND2 AND2_2217(.VSS(VSS),.VDD(VDD),.Y(g24708),.A(g16474),.B(g22998));
  AND2 AND2_2218(.VSS(VSS),.VDD(VDD),.Y(g14644),.A(g10610),.B(g10605));
  AND3 AND3_134(.VSS(VSS),.VDD(VDD),.Y(g33913),.A(g23088),.B(g33204),.C(g9104));
  AND2 AND2_2219(.VSS(VSS),.VDD(VDD),.Y(g16592),.A(g5579),.B(g14688));
  AND2 AND2_2220(.VSS(VSS),.VDD(VDD),.Y(g21844),.A(g3873),.B(g21070));
  AND2 AND2_2221(.VSS(VSS),.VDD(VDD),.Y(g21394),.A(g13335),.B(g15799));
  AND2 AND2_2222(.VSS(VSS),.VDD(VDD),.Y(g32356),.A(g2704),.B(g31710));
  AND2 AND2_2223(.VSS(VSS),.VDD(VDD),.Y(g29475),.A(g14033),.B(g28500));
  AND2 AND2_2224(.VSS(VSS),.VDD(VDD),.Y(g18459),.A(g2331),.B(g15224));
  AND2 AND2_2225(.VSS(VSS),.VDD(VDD),.Y(g18425),.A(g2161),.B(g18008));
  AND2 AND2_2226(.VSS(VSS),.VDD(VDD),.Y(g33905),.A(g33089),.B(g15574));
  AND2 AND2_2227(.VSS(VSS),.VDD(VDD),.Y(g33073),.A(g32386),.B(g18828));
  AND2 AND2_2228(.VSS(VSS),.VDD(VDD),.Y(g12687),.A(g9024),.B(g8977));
  AND2 AND2_2229(.VSS(VSS),.VDD(VDD),.Y(g25106),.A(g17391),.B(g23506));
  AND2 AND2_2230(.VSS(VSS),.VDD(VDD),.Y(g26541),.A(g319),.B(g24375));
  AND2 AND2_2231(.VSS(VSS),.VDD(VDD),.Y(g34514),.A(g34286),.B(g19480));
  AND2 AND2_2232(.VSS(VSS),.VDD(VDD),.Y(g15851),.A(g3953),.B(g14157));
  AND2 AND2_2233(.VSS(VSS),.VDD(VDD),.Y(g15872),.A(g9095),.B(g14234));
  AND2 AND2_2234(.VSS(VSS),.VDD(VDD),.Y(g18458),.A(g2357),.B(g15224));
  AND2 AND2_2235(.VSS(VSS),.VDD(VDD),.Y(g19139),.A(g452),.B(g16195));
  AND2 AND2_2236(.VSS(VSS),.VDD(VDD),.Y(g27374),.A(g26519),.B(g17478));
  AND3 AND3_135(.VSS(VSS),.VDD(VDD),.Y(g33530),.A(g32960),.B(I31346),.C(I31347));
  AND2 AND2_2237(.VSS(VSS),.VDD(VDD),.Y(g21420),.A(g16093),.B(g13596));
  AND2 AND2_2238(.VSS(VSS),.VDD(VDD),.Y(g34507),.A(g34280),.B(g19454));
  AND2 AND2_2239(.VSS(VSS),.VDD(VDD),.Y(g31122),.A(g12144),.B(g29993));
  AND2 AND2_2240(.VSS(VSS),.VDD(VDD),.Y(g32182),.A(g31753),.B(g27937));
  AND4 AND4_146(.VSS(VSS),.VDD(VDD),.Y(g20069),.A(g16312),.B(g9051),.C(g9011),.D(g8955));
  AND2 AND2_2241(.VSS(VSS),.VDD(VDD),.Y(g33122),.A(g8859),.B(g32192));
  AND2 AND2_2242(.VSS(VSS),.VDD(VDD),.Y(g8530),.A(g2902),.B(g2907));
  AND4 AND4_147(.VSS(VSS),.VDD(VDD),.Y(I31027),.A(g32494),.B(g32495),.C(g32496),.D(g32497));
  AND3 AND3_136(.VSS(VSS),.VDD(VDD),.Y(I24524),.A(g5041),.B(g5046),.C(g9716));
  AND3 AND3_137(.VSS(VSS),.VDD(VDD),.Y(g33464),.A(g32484),.B(I31016),.C(I31017));
  AND3 AND3_138(.VSS(VSS),.VDD(VDD),.Y(I16129),.A(g8728),.B(g11443),.C(g11411));
  AND2 AND2_2243(.VSS(VSS),.VDD(VDD),.Y(g20602),.A(g10803),.B(g15580));
  AND4 AND4_148(.VSS(VSS),.VDD(VDD),.Y(g28150),.A(g10862),.B(g11834),.C(g11283),.D(g27187));
  AND3 AND3_139(.VSS(VSS),.VDD(VDD),.Y(g16846),.A(g14034),.B(g12591),.C(g11185));
  AND2 AND2_2244(.VSS(VSS),.VDD(VDD),.Y(g18545),.A(g2783),.B(g15277));
  AND2 AND2_2245(.VSS(VSS),.VDD(VDD),.Y(g25951),.A(g24500),.B(g19565));
  AND2 AND2_2246(.VSS(VSS),.VDD(VDD),.Y(g26325),.A(g12644),.B(g25370));
  AND2 AND2_2247(.VSS(VSS),.VDD(VDD),.Y(g24602),.A(g16507),.B(g22854));
  AND2 AND2_2248(.VSS(VSS),.VDD(VDD),.Y(g25972),.A(g2217),.B(g24993));
  AND2 AND2_2249(.VSS(VSS),.VDD(VDD),.Y(g18444),.A(g2269),.B(g18008));
  AND2 AND2_2250(.VSS(VSS),.VDD(VDD),.Y(g25033),.A(g17500),.B(g23433));
  AND3 AND3_140(.VSS(VSS),.VDD(VDD),.Y(g25371),.A(g5062),.B(g22173),.C(I24524));
  AND2 AND2_2251(.VSS(VSS),.VDD(VDD),.Y(g20375),.A(g671),.B(g16846));
  AND2 AND2_2252(.VSS(VSS),.VDD(VDD),.Y(g24657),.A(g22644),.B(g19730));
  AND2 AND2_2253(.VSS(VSS),.VDD(VDD),.Y(g24774),.A(g718),.B(g23614));
  AND2 AND2_2254(.VSS(VSS),.VDD(VDD),.Y(g16731),.A(g7153),.B(g12941));
  AND2 AND2_2255(.VSS(VSS),.VDD(VDD),.Y(g26829),.A(g2844),.B(g24505));
  AND2 AND2_2256(.VSS(VSS),.VDD(VDD),.Y(g27669),.A(g26840),.B(g13278));
  AND2 AND2_2257(.VSS(VSS),.VDD(VDD),.Y(g17480),.A(g9683),.B(g14433));
  AND2 AND2_2258(.VSS(VSS),.VDD(VDD),.Y(g19333),.A(g464),.B(g16223));
  AND2 AND2_2259(.VSS(VSS),.VDD(VDD),.Y(g29347),.A(g29176),.B(g22201));
  AND2 AND2_2260(.VSS(VSS),.VDD(VDD),.Y(g18599),.A(g2955),.B(g16349));
  AND2 AND2_2261(.VSS(VSS),.VDD(VDD),.Y(g22307),.A(g20027),.B(g21163));
  AND2 AND2_2262(.VSS(VSS),.VDD(VDD),.Y(g22076),.A(g6255),.B(g19210));
  AND2 AND2_2263(.VSS(VSS),.VDD(VDD),.Y(g22085),.A(g6295),.B(g19210));
  AND2 AND2_2264(.VSS(VSS),.VDD(VDD),.Y(g26358),.A(g19522),.B(g25528));
  AND3 AND3_141(.VSS(VSS),.VDD(VDD),.Y(I27349),.A(g25534),.B(g26424),.C(g22698));
  AND2 AND2_2265(.VSS(VSS),.VDD(VDD),.Y(g23025),.A(g16021),.B(g19798));
  AND2 AND2_2266(.VSS(VSS),.VDD(VDD),.Y(g27260),.A(g26766),.B(g26737));
  AND2 AND2_2267(.VSS(VSS),.VDD(VDD),.Y(g32331),.A(g31322),.B(g20637));
  AND2 AND2_2268(.VSS(VSS),.VDD(VDD),.Y(g31292),.A(g29735),.B(g23338));
  AND2 AND2_2269(.VSS(VSS),.VDD(VDD),.Y(g26828),.A(g24919),.B(g15756));
  AND2 AND2_2270(.VSS(VSS),.VDD(VDD),.Y(g27668),.A(g1367),.B(g25917));
  AND2 AND2_2271(.VSS(VSS),.VDD(VDD),.Y(g23540),.A(g16866),.B(g20622));
  AND2 AND2_2272(.VSS(VSS),.VDD(VDD),.Y(g18598),.A(g3003),.B(g16349));
  AND2 AND2_2273(.VSS(VSS),.VDD(VDD),.Y(g22054),.A(g6120),.B(g21611));
  AND2 AND2_2274(.VSS(VSS),.VDD(VDD),.Y(g28695),.A(g27580),.B(g20666));
  AND2 AND2_2275(.VSS(VSS),.VDD(VDD),.Y(g31153),.A(g12336),.B(g30068));
  AND2 AND2_2276(.VSS(VSS),.VDD(VDD),.Y(g27392),.A(g26576),.B(g17507));
  AND2 AND2_2277(.VSS(VSS),.VDD(VDD),.Y(g29600),.A(g1840),.B(g29049));
  AND2 AND2_2278(.VSS(VSS),.VDD(VDD),.Y(g26121),.A(g6167),.B(g25111));
  AND2 AND2_2279(.VSS(VSS),.VDD(VDD),.Y(g20171),.A(g16479),.B(g10476));
  AND2 AND2_2280(.VSS(VSS),.VDD(VDD),.Y(g34541),.A(g34331),.B(g20087));
  AND2 AND2_2281(.VSS(VSS),.VDD(VDD),.Y(g17307),.A(g9498),.B(g14343));
  AND2 AND2_2282(.VSS(VSS),.VDD(VDD),.Y(g15574),.A(g4311),.B(g13202));
  AND2 AND2_2283(.VSS(VSS),.VDD(VDD),.Y(g33409),.A(g32359),.B(g21408));
  AND3 AND3_142(.VSS(VSS),.VDD(VDD),.Y(I24616),.A(g6082),.B(g6088),.C(g9946));
  AND2 AND2_2284(.VSS(VSS),.VDD(VDD),.Y(g29952),.A(g23576),.B(g28939));
  AND2 AND2_2285(.VSS(VSS),.VDD(VDD),.Y(g27559),.A(g26576),.B(g17777));
  AND2 AND2_2286(.VSS(VSS),.VDD(VDD),.Y(g29351),.A(g4771),.B(g28406));
  AND2 AND2_2287(.VSS(VSS),.VDD(VDD),.Y(g27525),.A(g26576),.B(g17720));
  AND2 AND2_2288(.VSS(VSS),.VDD(VDD),.Y(g27488),.A(g26549),.B(g17648));
  AND2 AND2_2289(.VSS(VSS),.VDD(VDD),.Y(g18817),.A(g6533),.B(g15483));
  AND2 AND2_2290(.VSS(VSS),.VDD(VDD),.Y(g15912),.A(g3562),.B(g14018));
  AND4 AND4_149(.VSS(VSS),.VDD(VDD),.Y(g14581),.A(g12587),.B(g12428),.C(g12357),.D(I16695));
  AND2 AND2_2291(.VSS(VSS),.VDD(VDD),.Y(g18322),.A(g1608),.B(g17873));
  AND2 AND2_2292(.VSS(VSS),.VDD(VDD),.Y(g33408),.A(g32358),.B(g21407));
  AND4 AND4_150(.VSS(VSS),.VDD(VDD),.Y(I31081),.A(g30673),.B(g31810),.C(g32571),.D(g32572));
  AND2 AND2_2293(.VSS(VSS),.VDD(VDD),.Y(g24967),.A(g23197),.B(g20213));
  AND2 AND2_2294(.VSS(VSS),.VDD(VDD),.Y(g10707),.A(g3787),.B(g8561));
  AND2 AND2_2295(.VSS(VSS),.VDD(VDD),.Y(g18159),.A(g671),.B(g17433));
  AND2 AND2_2296(.VSS(VSS),.VDD(VDD),.Y(g27558),.A(g26576),.B(g17776));
  AND3 AND3_143(.VSS(VSS),.VDD(VDD),.Y(g25507),.A(g6098),.B(g23844),.C(I24616));
  AND2 AND2_2297(.VSS(VSS),.VDD(VDD),.Y(g22942),.A(g9104),.B(g20219));
  AND2 AND2_2298(.VSS(VSS),.VDD(VDD),.Y(g18125),.A(g15053),.B(g16886));
  AND2 AND2_2299(.VSS(VSS),.VDD(VDD),.Y(g18532),.A(g2724),.B(g15277));
  AND2 AND2_2300(.VSS(VSS),.VDD(VDD),.Y(g26291),.A(g2681),.B(g25439));
  AND2 AND2_2301(.VSS(VSS),.VDD(VDD),.Y(g30920),.A(g29889),.B(g21024));
  AND4 AND4_151(.VSS(VSS),.VDD(VDD),.Y(I24704),.A(g21193),.B(g24061),.C(g24062),.D(g24063));
  AND2 AND2_2302(.VSS(VSS),.VDD(VDD),.Y(g19585),.A(g17180),.B(g14004));
  AND2 AND2_2303(.VSS(VSS),.VDD(VDD),.Y(g14202),.A(g869),.B(g10632));
  AND2 AND2_2304(.VSS(VSS),.VDD(VDD),.Y(g16929),.A(g6505),.B(g14348));
  AND2 AND2_2305(.VSS(VSS),.VDD(VDD),.Y(g18158),.A(g667),.B(g17433));
  AND2 AND2_2306(.VSS(VSS),.VDD(VDD),.Y(g14257),.A(g8612),.B(g11878));
  AND2 AND2_2307(.VSS(VSS),.VDD(VDD),.Y(g21957),.A(g5390),.B(g21514));
  AND2 AND2_2308(.VSS(VSS),.VDD(VDD),.Y(g18783),.A(g5841),.B(g18065));
  AND2 AND2_2309(.VSS(VSS),.VDD(VDD),.Y(g23957),.A(g4138),.B(g19589));
  AND2 AND2_2310(.VSS(VSS),.VDD(VDD),.Y(g29516),.A(g28895),.B(g22369));
  AND4 AND4_152(.VSS(VSS),.VDD(VDD),.Y(g14496),.A(g12411),.B(g12244),.C(g12197),.D(I16618));
  AND2 AND2_2311(.VSS(VSS),.VDD(VDD),.Y(g22670),.A(g20114),.B(g9104));
  AND2 AND2_2312(.VSS(VSS),.VDD(VDD),.Y(g21739),.A(g3080),.B(g20330));
  AND4 AND4_153(.VSS(VSS),.VDD(VDD),.Y(I31356),.A(g31327),.B(g31859),.C(g32968),.D(g32969));
  AND2 AND2_2313(.VSS(VSS),.VDD(VDD),.Y(g25163),.A(g20217),.B(g23566));
  AND2 AND2_2314(.VSS(VSS),.VDD(VDD),.Y(g18561),.A(g2841),.B(g15277));
  AND2 AND2_2315(.VSS(VSS),.VDD(VDD),.Y(g18656),.A(g15120),.B(g17128));
  AND2 AND2_2316(.VSS(VSS),.VDD(VDD),.Y(g30121),.A(g28577),.B(g21052));
  AND2 AND2_2317(.VSS(VSS),.VDD(VDD),.Y(g25012),.A(g20644),.B(g23419));
  AND2 AND2_2318(.VSS(VSS),.VDD(VDD),.Y(g18353),.A(g1772),.B(g17955));
  AND2 AND2_2319(.VSS(VSS),.VDD(VDD),.Y(g18295),.A(g1489),.B(g16449));
  AND2 AND2_2320(.VSS(VSS),.VDD(VDD),.Y(g21738),.A(g3072),.B(g20330));
  AND3 AND3_144(.VSS(VSS),.VDD(VDD),.Y(g10590),.A(g7246),.B(g7392),.C(I13937));
  AND2 AND2_2321(.VSS(VSS),.VDD(VDD),.Y(g17156),.A(g305),.B(g13385));
  AND2 AND2_2322(.VSS(VSS),.VDD(VDD),.Y(g17655),.A(g7897),.B(g13342));
  AND2 AND2_2323(.VSS(VSS),.VDD(VDD),.Y(g18680),.A(g15128),.B(g15885));
  AND2 AND2_2324(.VSS(VSS),.VDD(VDD),.Y(g18144),.A(g590),.B(g17533));
  AND2 AND2_2325(.VSS(VSS),.VDD(VDD),.Y(g18823),.A(g6727),.B(g15680));
  AND2 AND2_2326(.VSS(VSS),.VDD(VDD),.Y(g34344),.A(g34107),.B(g20038));
  AND2 AND2_2327(.VSS(VSS),.VDD(VDD),.Y(g21699),.A(g142),.B(g20283));
  AND2 AND2_2328(.VSS(VSS),.VDD(VDD),.Y(g28706),.A(g27584),.B(g20681));
  AND2 AND2_2329(.VSS(VSS),.VDD(VDD),.Y(g28597),.A(g27515),.B(g20508));
  AND4 AND4_154(.VSS(VSS),.VDD(VDD),.Y(I31182),.A(g32719),.B(g32720),.C(g32721),.D(g32722));
  AND2 AND2_2330(.VSS(VSS),.VDD(VDD),.Y(g18336),.A(g1700),.B(g17873));
  AND2 AND2_2331(.VSS(VSS),.VDD(VDD),.Y(g24545),.A(g3333),.B(g23285));
  AND3 AND3_145(.VSS(VSS),.VDD(VDD),.Y(g33474),.A(g32556),.B(I31066),.C(I31067));
  AND2 AND2_2332(.VSS(VSS),.VDD(VDD),.Y(g28256),.A(g11398),.B(g27984));
  AND2 AND2_2333(.VSS(VSS),.VDD(VDD),.Y(g15820),.A(g3578),.B(g13955));
  AND2 AND2_2334(.VSS(VSS),.VDD(VDD),.Y(g28689),.A(g27575),.B(g20651));
  AND2 AND2_2335(.VSS(VSS),.VDD(VDD),.Y(g32149),.A(g31658),.B(g29983));
  AND2 AND2_2336(.VSS(VSS),.VDD(VDD),.Y(g27042),.A(g25774),.B(g19343));
  AND3 AND3_146(.VSS(VSS),.VDD(VDD),.Y(g33711),.A(g33176),.B(g10727),.C(g22332));
  AND2 AND2_2337(.VSS(VSS),.VDD(VDD),.Y(g30173),.A(g28118),.B(g13082));
  AND2 AND2_2338(.VSS(VSS),.VDD(VDD),.Y(g34291),.A(g34055),.B(g19366));
  AND2 AND2_2339(.VSS(VSS),.VDD(VDD),.Y(g31327),.A(g19200),.B(g29814));
  AND2 AND2_2340(.VSS(VSS),.VDD(VDD),.Y(g27255),.A(g25936),.B(g19689));
  AND2 AND2_2341(.VSS(VSS),.VDD(VDD),.Y(g28280),.A(g23761),.B(g27724));
  AND2 AND2_2342(.VSS(VSS),.VDD(VDD),.Y(g22131),.A(g6641),.B(g19277));
  AND2 AND2_2343(.VSS(VSS),.VDD(VDD),.Y(g29834),.A(g28368),.B(g23278));
  AND2 AND2_2344(.VSS(VSS),.VDD(VDD),.Y(g33327),.A(g32208),.B(g20561));
  AND2 AND2_2345(.VSS(VSS),.VDD(VDD),.Y(g34173),.A(g33679),.B(g24368));
  AND3 AND3_147(.VSS(VSS),.VDD(VDD),.Y(I24064),.A(g3385),.B(g3391),.C(g8492));
  AND3 AND3_148(.VSS(VSS),.VDD(VDD),.Y(g29208),.A(g24138),.B(I27538),.C(I27539));
  AND2 AND2_2346(.VSS(VSS),.VDD(VDD),.Y(g25788),.A(g8010),.B(g24579));
  AND2 AND2_2347(.VSS(VSS),.VDD(VDD),.Y(g32148),.A(g31631),.B(g29981));
  AND2 AND2_2348(.VSS(VSS),.VDD(VDD),.Y(g28624),.A(g22357),.B(g27009));
  AND2 AND2_2349(.VSS(VSS),.VDD(VDD),.Y(g28300),.A(g27771),.B(g26605));
  AND2 AND2_2350(.VSS(VSS),.VDD(VDD),.Y(g27270),.A(g26805),.B(g26793));
  AND2 AND2_2351(.VSS(VSS),.VDD(VDD),.Y(g32097),.A(g25960),.B(g31021));
  AND4 AND4_155(.VSS(VSS),.VDD(VDD),.Y(I31331),.A(g30825),.B(g31854),.C(g32933),.D(g32934));
  AND2 AND2_2352(.VSS(VSS),.VDD(VDD),.Y(g27678),.A(g947),.B(g25830));
  AND2 AND2_2353(.VSS(VSS),.VDD(VDD),.Y(g18631),.A(g3694),.B(g17226));
  AND2 AND2_2354(.VSS(VSS),.VDD(VDD),.Y(g32104),.A(g31616),.B(g29906));
  AND3 AND3_149(.VSS(VSS),.VDD(VDD),.Y(g7520),.A(g2704),.B(g2697),.C(g2689));
  AND2 AND2_2355(.VSS(VSS),.VDD(VDD),.Y(g18364),.A(g1844),.B(g17955));
  AND2 AND2_2356(.VSS(VSS),.VDD(VDD),.Y(g32343),.A(g31473),.B(g20710));
  AND2 AND2_2357(.VSS(VSS),.VDD(VDD),.Y(g31283),.A(g30156),.B(g27837));
  AND2 AND2_2358(.VSS(VSS),.VDD(VDD),.Y(g27460),.A(g26549),.B(g17610));
  AND2 AND2_2359(.VSS(VSS),.VDD(VDD),.Y(g27686),.A(g1291),.B(g25849));
  AND2 AND2_2360(.VSS(VSS),.VDD(VDD),.Y(g25946),.A(g24496),.B(g19537));
  AND2 AND2_2361(.VSS(VSS),.VDD(VDD),.Y(g31492),.A(g29790),.B(g23431));
  AND2 AND2_2362(.VSS(VSS),.VDD(VDD),.Y(g24817),.A(g22929),.B(g7235));
  AND2 AND2_2363(.VSS(VSS),.VDD(VDD),.Y(g30029),.A(g29164),.B(g12936));
  AND3 AND3_150(.VSS(VSS),.VDD(VDD),.Y(g33492),.A(g32686),.B(I31156),.C(I31157));
  AND2 AND2_2364(.VSS(VSS),.VDD(VDD),.Y(g19674),.A(g2819),.B(g15867));
  AND2 AND2_2365(.VSS(VSS),.VDD(VDD),.Y(g24322),.A(g4423),.B(g22228));
  AND2 AND2_2366(.VSS(VSS),.VDD(VDD),.Y(g12939),.A(g405),.B(g11048));
  AND2 AND2_2367(.VSS(VSS),.VDD(VDD),.Y(g27030),.A(g26343),.B(g7947));
  AND2 AND2_2368(.VSS(VSS),.VDD(VDD),.Y(g20977),.A(g10123),.B(g17301));
  AND2 AND2_2369(.VSS(VSS),.VDD(VDD),.Y(g13299),.A(g437),.B(g11048));
  AND2 AND2_2370(.VSS(VSS),.VDD(VDD),.Y(g24532),.A(g22331),.B(g19478));
  AND2 AND2_2371(.VSS(VSS),.VDD(VDD),.Y(g32369),.A(g2130),.B(g31672));
  AND2 AND2_2372(.VSS(VSS),.VDD(VDD),.Y(g27267),.A(g26026),.B(g17124));
  AND2 AND2_2373(.VSS(VSS),.VDD(VDD),.Y(g27294),.A(g9975),.B(g26656));
  AND2 AND2_2374(.VSS(VSS),.VDD(VDD),.Y(g29614),.A(g28860),.B(g22369));
  AND2 AND2_2375(.VSS(VSS),.VDD(VDD),.Y(g30028),.A(g29069),.B(g9311));
  AND3 AND3_151(.VSS(VSS),.VDD(VDD),.Y(g28231),.A(g27187),.B(g22763),.C(g27074));
  AND2 AND2_2376(.VSS(VSS),.VDD(VDD),.Y(g24977),.A(g23209),.B(g20232));
  AND2 AND2_2377(.VSS(VSS),.VDD(VDD),.Y(g34506),.A(g8833),.B(g34354));
  AND2 AND2_2378(.VSS(VSS),.VDD(VDD),.Y(g16803),.A(g5933),.B(g14810));
  AND2 AND2_2379(.VSS(VSS),.VDD(VDD),.Y(g31750),.A(g30103),.B(g23925));
  AND2 AND2_2380(.VSS(VSS),.VDD(VDD),.Y(g29607),.A(g28509),.B(g14208));
  AND2 AND2_2381(.VSS(VSS),.VDD(VDD),.Y(g18289),.A(g1448),.B(g16449));
  AND4 AND4_156(.VSS(VSS),.VDD(VDD),.Y(I31026),.A(g31194),.B(g31800),.C(g32492),.D(g32493));
  AND2 AND2_2382(.VSS(VSS),.VDD(VDD),.Y(g29320),.A(g29068),.B(g22147));
  AND2 AND2_2383(.VSS(VSS),.VDD(VDD),.Y(g33381),.A(g11842),.B(g32318));
  AND4 AND4_157(.VSS(VSS),.VDD(VDD),.Y(I31212),.A(g32761),.B(g32762),.C(g32763),.D(g32764));
  AND4 AND4_158(.VSS(VSS),.VDD(VDD),.Y(g29073),.A(g27163),.B(g10290),.C(g21012),.D(I27409));
  AND2 AND2_2384(.VSS(VSS),.VDD(VDD),.Y(g12065),.A(g9557),.B(g9805));
  AND2 AND2_2385(.VSS(VSS),.VDD(VDD),.Y(g18309),.A(g1339),.B(g16931));
  AND2 AND2_2386(.VSS(VSS),.VDD(VDD),.Y(g29530),.A(g1612),.B(g28820));
  AND2 AND2_2387(.VSS(VSS),.VDD(VDD),.Y(g24656),.A(g11736),.B(g22926));
  AND2 AND2_2388(.VSS(VSS),.VDD(VDD),.Y(g29593),.A(g28470),.B(g7985));
  AND2 AND2_2389(.VSS(VSS),.VDD(VDD),.Y(g33091),.A(g32392),.B(g18897));
  AND2 AND2_2390(.VSS(VSS),.VDD(VDD),.Y(g18288),.A(g1454),.B(g16449));
  AND2 AND2_2391(.VSS(VSS),.VDD(VDD),.Y(g18224),.A(g1036),.B(g16100));
  AND2 AND2_2392(.VSS(VSS),.VDD(VDD),.Y(g21715),.A(g160),.B(g20283));
  AND2 AND2_2393(.VSS(VSS),.VDD(VDD),.Y(g22039),.A(g5949),.B(g19147));
  AND2 AND2_2394(.VSS(VSS),.VDD(VDD),.Y(g29346),.A(g4894),.B(g28381));
  AND2 AND2_2395(.VSS(VSS),.VDD(VDD),.Y(g25173),.A(g12234),.B(g23589));
  AND2 AND2_2396(.VSS(VSS),.VDD(VDD),.Y(g24295),.A(g4434),.B(g22550));
  AND2 AND2_2397(.VSS(VSS),.VDD(VDD),.Y(g18571),.A(g2856),.B(g16349));
  AND2 AND2_2398(.VSS(VSS),.VDD(VDD),.Y(g18308),.A(g6832),.B(g16931));
  AND2 AND2_2399(.VSS(VSS),.VDD(VDD),.Y(g24680),.A(g16422),.B(g22986));
  AND2 AND2_2400(.VSS(VSS),.VDD(VDD),.Y(g27219),.A(g26026),.B(g16742));
  AND2 AND2_2401(.VSS(VSS),.VDD(VDD),.Y(g32412),.A(g4765),.B(g30998));
  AND2 AND2_2402(.VSS(VSS),.VDD(VDD),.Y(g24144),.A(g17727),.B(g21660));
  AND2 AND2_2403(.VSS(VSS),.VDD(VDD),.Y(g33796),.A(g33117),.B(g25267));
  AND2 AND2_2404(.VSS(VSS),.VDD(VDD),.Y(g19692),.A(g12066),.B(g17086));
  AND3 AND3_152(.VSS(VSS),.VDD(VDD),.Y(I24555),.A(g9559),.B(g9809),.C(g6093));
  AND2 AND2_2405(.VSS(VSS),.VDD(VDD),.Y(g29565),.A(g1932),.B(g28590));
  AND2 AND2_2406(.VSS(VSS),.VDD(VDD),.Y(g26604),.A(g13248),.B(g25051));
  AND2 AND2_2407(.VSS(VSS),.VDD(VDD),.Y(g17469),.A(g4076),.B(g13217));
  AND2 AND2_2408(.VSS(VSS),.VDD(VDD),.Y(g13737),.A(g4501),.B(g10571));
  AND2 AND2_2409(.VSS(VSS),.VDD(VDD),.Y(g22038),.A(g5945),.B(g19147));
  AND2 AND2_2410(.VSS(VSS),.VDD(VDD),.Y(g23551),.A(g10793),.B(g18948));
  AND2 AND2_2411(.VSS(VSS),.VDD(VDD),.Y(g23572),.A(g20230),.B(g20656));
  AND2 AND2_2412(.VSS(VSS),.VDD(VDD),.Y(g10917),.A(g9174),.B(g1087));
  AND2 AND2_2413(.VSS(VSS),.VDD(VDD),.Y(g12219),.A(g1189),.B(g7532));
  AND2 AND2_2414(.VSS(VSS),.VDD(VDD),.Y(g27218),.A(g25997),.B(g16740));
  AND2 AND2_2415(.VSS(VSS),.VDD(VDD),.Y(g30927),.A(g29910),.B(g24795));
  AND2 AND2_2416(.VSS(VSS),.VDD(VDD),.Y(g18495),.A(g2533),.B(g15426));
  AND2 AND2_2417(.VSS(VSS),.VDD(VDD),.Y(g33840),.A(g33253),.B(g20267));
  AND2 AND2_2418(.VSS(VSS),.VDD(VDD),.Y(g29641),.A(g28520),.B(g14237));
  AND2 AND2_2419(.VSS(VSS),.VDD(VDD),.Y(g29797),.A(g28347),.B(g23259));
  AND2 AND2_2420(.VSS(VSS),.VDD(VDD),.Y(g16662),.A(g4552),.B(g14753));
  AND2 AND2_2421(.VSS(VSS),.VDD(VDD),.Y(g13697),.A(g11166),.B(g8608));
  AND2 AND2_2422(.VSS(VSS),.VDD(VDD),.Y(g28660),.A(g27824),.B(g20623));
  AND2 AND2_2423(.VSS(VSS),.VDD(VDD),.Y(g18816),.A(g6527),.B(g15483));
  AND2 AND2_2424(.VSS(VSS),.VDD(VDD),.Y(g32011),.A(g8287),.B(g31134));
  AND2 AND2_2425(.VSS(VSS),.VDD(VDD),.Y(g27160),.A(g14163),.B(g26340));
  AND2 AND2_2426(.VSS(VSS),.VDD(VDD),.Y(g10706),.A(g3338),.B(g8691));
  AND2 AND2_2427(.VSS(VSS),.VDD(VDD),.Y(g15113),.A(g4291),.B(g14454));
  AND2 AND2_2428(.VSS(VSS),.VDD(VDD),.Y(g19207),.A(g7803),.B(g15992));
  AND2 AND2_2429(.VSS(VSS),.VDD(VDD),.Y(g18687),.A(g4664),.B(g15885));
  AND2 AND2_2430(.VSS(VSS),.VDD(VDD),.Y(g28456),.A(g27290),.B(g20104));
  AND4 AND4_159(.VSS(VSS),.VDD(VDD),.Y(I31097),.A(g32596),.B(g32597),.C(g32598),.D(g32599));
  AND2 AND2_2431(.VSS(VSS),.VDD(VDD),.Y(g17601),.A(g9616),.B(g14572));
  AND2 AND2_2432(.VSS(VSS),.VDD(VDD),.Y(g22143),.A(g19568),.B(g10971));
  AND2 AND2_2433(.VSS(VSS),.VDD(VDD),.Y(g21784),.A(g3423),.B(g20391));
  AND2 AND2_2434(.VSS(VSS),.VDD(VDD),.Y(g22937),.A(g753),.B(g20540));
  AND2 AND2_2435(.VSS(VSS),.VDD(VDD),.Y(g26845),.A(g24391),.B(g21426));
  AND2 AND2_2436(.VSS(VSS),.VDD(VDD),.Y(g14256),.A(g2079),.B(g11872));
  AND2 AND2_2437(.VSS(VSS),.VDD(VDD),.Y(g21956),.A(g5360),.B(g21514));
  AND2 AND2_2438(.VSS(VSS),.VDD(VDD),.Y(g18752),.A(g15146),.B(g17926));
  AND2 AND2_2439(.VSS(VSS),.VDD(VDD),.Y(g27455),.A(g26488),.B(g17603));
  AND2 AND2_2440(.VSS(VSS),.VDD(VDD),.Y(g26395),.A(g22547),.B(g25561));
  AND2 AND2_2441(.VSS(VSS),.VDD(VDD),.Y(g30604),.A(g18911),.B(g29878));
  AND3 AND3_153(.VSS(VSS),.VDD(VDD),.Y(g33522),.A(g32902),.B(I31306),.C(I31307));
  AND2 AND2_2442(.VSS(VSS),.VDD(VDD),.Y(g18374),.A(g1878),.B(g15171));
  AND2 AND2_2443(.VSS(VSS),.VDD(VDD),.Y(g29635),.A(g28910),.B(g22432));
  AND2 AND2_2444(.VSS(VSS),.VDD(VDD),.Y(g21889),.A(g4169),.B(g19801));
  AND2 AND2_2445(.VSS(VSS),.VDD(VDD),.Y(g23103),.A(g10143),.B(g20765));
  AND4 AND4_160(.VSS(VSS),.VDD(VDD),.Y(g27617),.A(g23032),.B(g26264),.C(g26424),.D(g24982));
  AND2 AND2_2446(.VSS(VSS),.VDD(VDD),.Y(g15105),.A(g4235),.B(g14454));
  AND2 AND2_2447(.VSS(VSS),.VDD(VDD),.Y(g21980),.A(g5567),.B(g19074));
  AND2 AND2_2448(.VSS(VSS),.VDD(VDD),.Y(g10624),.A(g8387),.B(g3072));
  AND2 AND2_2449(.VSS(VSS),.VDD(VDD),.Y(g28550),.A(g12009),.B(g27092));
  AND2 AND2_2450(.VSS(VSS),.VDD(VDD),.Y(g18643),.A(g3849),.B(g17096));
  AND2 AND2_2451(.VSS(VSS),.VDD(VDD),.Y(g7469),.A(g4382),.B(g4438));
  AND2 AND2_2452(.VSS(VSS),.VDD(VDD),.Y(g32310),.A(g27577),.B(g31376));
  AND2 AND2_2453(.VSS(VSS),.VDD(VDD),.Y(g16204),.A(g6537),.B(g14348));
  AND2 AND2_2454(.VSS(VSS),.VDD(VDD),.Y(g28314),.A(g27552),.B(g14205));
  AND2 AND2_2455(.VSS(VSS),.VDD(VDD),.Y(g21888),.A(g4165),.B(g19801));
  AND2 AND2_2456(.VSS(VSS),.VDD(VDD),.Y(g21824),.A(g3706),.B(g20453));
  AND2 AND2_2457(.VSS(VSS),.VDD(VDD),.Y(g26633),.A(g24964),.B(g20616));
  AND2 AND2_2458(.VSS(VSS),.VDD(VDD),.Y(g34563),.A(g34372),.B(g17465));
  AND3 AND3_154(.VSS(VSS),.VDD(VDD),.Y(I17542),.A(g13156),.B(g6767),.C(g6756));
  AND2 AND2_2459(.VSS(VSS),.VDD(VDD),.Y(g27201),.A(g25997),.B(g16685));
  AND2 AND2_2460(.VSS(VSS),.VDD(VDD),.Y(g27277),.A(g26359),.B(g14191));
  AND4 AND4_161(.VSS(VSS),.VDD(VDD),.Y(I24675),.A(g24022),.B(g24023),.C(g24024),.D(g24025));
  AND3 AND3_155(.VSS(VSS),.VDD(VDD),.Y(g33483),.A(g32621),.B(I31111),.C(I31112));
  AND2 AND2_2461(.VSS(VSS),.VDD(VDD),.Y(g26719),.A(g10709),.B(g24438));
  AND2 AND2_2462(.VSS(VSS),.VDD(VDD),.Y(g24289),.A(g4427),.B(g22550));
  AND2 AND2_2463(.VSS(VSS),.VDD(VDD),.Y(g18669),.A(g4608),.B(g17367));
  AND2 AND2_2464(.VSS(VSS),.VDD(VDD),.Y(g32112),.A(g31646),.B(g29923));
  AND2 AND2_2465(.VSS(VSS),.VDD(VDD),.Y(g25927),.A(g25004),.B(g20375));
  AND2 AND2_2466(.VSS(VSS),.VDD(VDD),.Y(g32050),.A(g11003),.B(g30825));
  AND2 AND2_2467(.VSS(VSS),.VDD(VDD),.Y(g24309),.A(g4480),.B(g22228));
  AND2 AND2_2468(.VSS(VSS),.VDD(VDD),.Y(g33862),.A(g33272),.B(g20504));
  AND2 AND2_2469(.VSS(VSS),.VDD(VDD),.Y(g18260),.A(g1252),.B(g16000));
  AND2 AND2_2470(.VSS(VSS),.VDD(VDD),.Y(g28243),.A(g27879),.B(g23423));
  AND2 AND2_2471(.VSS(VSS),.VDD(VDD),.Y(g24288),.A(g4417),.B(g22550));
  AND2 AND2_2472(.VSS(VSS),.VDD(VDD),.Y(g27595),.A(g26733),.B(g26703));
  AND2 AND2_2473(.VSS(VSS),.VDD(VDD),.Y(g24224),.A(g269),.B(g22594));
  AND2 AND2_2474(.VSS(VSS),.VDD(VDD),.Y(g18668),.A(g4322),.B(g17367));
  AND2 AND2_2475(.VSS(VSS),.VDD(VDD),.Y(g27467),.A(g269),.B(g26832));
  AND4 AND4_162(.VSS(VSS),.VDD(VDD),.Y(g27494),.A(g8038),.B(g26314),.C(g518),.D(g9077));
  AND2 AND2_2476(.VSS(VSS),.VDD(VDD),.Y(g31949),.A(g1287),.B(g30825));
  AND2 AND2_2477(.VSS(VSS),.VDD(VDD),.Y(g18392),.A(g1988),.B(g15171));
  AND2 AND2_2478(.VSS(VSS),.VDD(VDD),.Y(g29891),.A(g28420),.B(g23356));
  AND2 AND2_2479(.VSS(VSS),.VDD(VDD),.Y(g24308),.A(g4489),.B(g22228));
  AND2 AND2_2480(.VSS(VSS),.VDD(VDD),.Y(g21931),.A(g5188),.B(g18997));
  AND2 AND2_2481(.VSS(VSS),.VDD(VDD),.Y(g18195),.A(g847),.B(g17821));
  AND2 AND2_2482(.VSS(VSS),.VDD(VDD),.Y(g22015),.A(g5719),.B(g21562));
  AND2 AND2_2483(.VSS(VSS),.VDD(VDD),.Y(g18489),.A(g2509),.B(g15426));
  AND2 AND2_2484(.VSS(VSS),.VDD(VDD),.Y(g34395),.A(g34193),.B(g21336));
  AND2 AND2_2485(.VSS(VSS),.VDD(VDD),.Y(g31948),.A(g30670),.B(g18884));
  AND2 AND2_2486(.VSS(VSS),.VDD(VDD),.Y(g32096),.A(g31601),.B(g29893));
  AND2 AND2_2487(.VSS(VSS),.VDD(VDD),.Y(g28269),.A(g27205),.B(g19712));
  AND2 AND2_2488(.VSS(VSS),.VDD(VDD),.Y(g29575),.A(g2066),.B(g28604));
  AND2 AND2_2489(.VSS(VSS),.VDD(VDD),.Y(g15881),.A(g3582),.B(g13983));
  AND2 AND2_2490(.VSS(VSS),.VDD(VDD),.Y(g18559),.A(g12856),.B(g15277));
  AND2 AND2_2491(.VSS(VSS),.VDD(VDD),.Y(g25491),.A(g23615),.B(g21355));
  AND2 AND2_2492(.VSS(VSS),.VDD(VDD),.Y(g18525),.A(g2610),.B(g15509));
  AND2 AND2_2493(.VSS(VSS),.VDD(VDD),.Y(g18488),.A(g2495),.B(g15426));
  AND2 AND2_2494(.VSS(VSS),.VDD(VDD),.Y(g18424),.A(g2165),.B(g18008));
  AND2 AND2_2495(.VSS(VSS),.VDD(VDD),.Y(g28341),.A(g27240),.B(g19790));
  AND2 AND2_2496(.VSS(VSS),.VDD(VDD),.Y(g29711),.A(g2541),.B(g29134));
  AND2 AND2_2497(.VSS(VSS),.VDD(VDD),.Y(g33904),.A(g33321),.B(g21059));
  AND2 AND2_2498(.VSS(VSS),.VDD(VDD),.Y(g24495),.A(g6928),.B(g23127));
  AND2 AND2_2499(.VSS(VSS),.VDD(VDD),.Y(g28268),.A(g8572),.B(g27990));
  AND2 AND2_2500(.VSS(VSS),.VDD(VDD),.Y(g31252),.A(g29643),.B(g20101));
  AND2 AND2_2501(.VSS(VSS),.VDD(VDD),.Y(g29327),.A(g29070),.B(g22156));
  AND2 AND2_2502(.VSS(VSS),.VDD(VDD),.Y(g26861),.A(g25021),.B(g25003));
  AND2 AND2_2503(.VSS(VSS),.VDD(VDD),.Y(g33252),.A(g32155),.B(g20064));
  AND2 AND2_2504(.VSS(VSS),.VDD(VDD),.Y(g13080),.A(g6923),.B(g11357));
  AND2 AND2_2505(.VSS(VSS),.VDD(VDD),.Y(g18558),.A(g2803),.B(g15277));
  AND2 AND2_2506(.VSS(VSS),.VDD(VDD),.Y(g28655),.A(g27561),.B(g20603));
  AND2 AND2_2507(.VSS(VSS),.VDD(VDD),.Y(g30191),.A(g28647),.B(g23843));
  AND2 AND2_2508(.VSS(VSS),.VDD(VDD),.Y(g16233),.A(g6137),.B(g14251));
  AND2 AND2_2509(.VSS(VSS),.VDD(VDD),.Y(g29537),.A(g28976),.B(g22472));
  AND2 AND2_2510(.VSS(VSS),.VDD(VDD),.Y(g34191),.A(g33713),.B(g24404));
  AND2 AND2_2511(.VSS(VSS),.VDD(VDD),.Y(g16672),.A(g6295),.B(g15008));
  AND2 AND2_2512(.VSS(VSS),.VDD(VDD),.Y(g27822),.A(g4157),.B(g25893));
  AND4 AND4_163(.VSS(VSS),.VDD(VDD),.Y(I27539),.A(g28040),.B(g24135),.C(g24136),.D(g24137));
  AND2 AND2_2513(.VSS(VSS),.VDD(VDD),.Y(g26389),.A(g19949),.B(g25553));
  AND2 AND2_2514(.VSS(VSS),.VDD(VDD),.Y(g18893),.A(g16215),.B(g16030));
  AND2 AND2_2515(.VSS(VSS),.VDD(VDD),.Y(g25981),.A(g2051),.B(g25007));
  AND2 AND2_2516(.VSS(VSS),.VDD(VDD),.Y(g24687),.A(g5827),.B(g23666));
  AND4 AND4_164(.VSS(VSS),.VDD(VDD),.Y(I31011),.A(g30735),.B(g31797),.C(g32471),.D(g32472));
  AND2 AND2_2517(.VSS(VSS),.VDD(VDD),.Y(g27266),.A(g26789),.B(g26770));
  AND2 AND2_2518(.VSS(VSS),.VDD(VDD),.Y(g26612),.A(g901),.B(g24407));
  AND4 AND4_165(.VSS(VSS),.VDD(VDD),.Y(I27538),.A(g21209),.B(g24132),.C(g24133),.D(g24134));
  AND2 AND2_2519(.VSS(VSS),.VDD(VDD),.Y(g26388),.A(g19595),.B(g25552));
  AND2 AND2_2520(.VSS(VSS),.VDD(VDD),.Y(g18544),.A(g2791),.B(g15277));
  AND2 AND2_2521(.VSS(VSS),.VDD(VDD),.Y(g26324),.A(g2661),.B(g25439));
  AND2 AND2_2522(.VSS(VSS),.VDD(VDD),.Y(g32428),.A(g31133),.B(g16261));
  AND2 AND2_2523(.VSS(VSS),.VDD(VDD),.Y(g29606),.A(g28480),.B(g8011));
  AND2 AND2_2524(.VSS(VSS),.VDD(VDD),.Y(g21024),.A(g16306),.B(g4871));
  AND2 AND2_2525(.VSS(VSS),.VDD(VDD),.Y(g18713),.A(g4836),.B(g15915));
  AND2 AND2_2526(.VSS(VSS),.VDD(VDD),.Y(g13461),.A(g2719),.B(g11819));
  AND2 AND2_2527(.VSS(VSS),.VDD(VDD),.Y(g22084),.A(g6291),.B(g19210));
  AND2 AND2_2528(.VSS(VSS),.VDD(VDD),.Y(g31183),.A(g30249),.B(g25174));
  AND2 AND2_2529(.VSS(VSS),.VDD(VDD),.Y(g26251),.A(g1988),.B(g25341));
  AND2 AND2_2530(.VSS(VSS),.VDD(VDD),.Y(g22110),.A(g15167),.B(g19277));
  AND2 AND2_2531(.VSS(VSS),.VDD(VDD),.Y(g24643),.A(g22636),.B(g19696));
  AND2 AND2_2532(.VSS(VSS),.VDD(VDD),.Y(g26272),.A(g2036),.B(g25470));
  AND2 AND2_2533(.VSS(VSS),.VDD(VDD),.Y(g33847),.A(g33260),.B(g20383));
  AND2 AND2_2534(.VSS(VSS),.VDD(VDD),.Y(g21860),.A(g3945),.B(g21070));
  AND2 AND2_2535(.VSS(VSS),.VDD(VDD),.Y(g16513),.A(g8345),.B(g13708));
  AND2 AND2_2536(.VSS(VSS),.VDD(VDD),.Y(g28694),.A(g27579),.B(g20664));
  AND2 AND2_2537(.VSS(VSS),.VDD(VDD),.Y(g29750),.A(g28296),.B(g23215));
  AND2 AND2_2538(.VSS(VSS),.VDD(VDD),.Y(g29982),.A(g23656),.B(g28998));
  AND2 AND2_2539(.VSS(VSS),.VDD(VDD),.Y(g29381),.A(g28135),.B(g19399));
  AND2 AND2_2540(.VSS(VSS),.VDD(VDD),.Y(g18610),.A(g15088),.B(g17059));
  AND2 AND2_2541(.VSS(VSS),.VDD(VDD),.Y(g34861),.A(g16540),.B(g34827));
  AND2 AND2_2542(.VSS(VSS),.VDD(VDD),.Y(g30247),.A(g28735),.B(g23937));
  AND2 AND2_2543(.VSS(VSS),.VDD(VDD),.Y(g18705),.A(g4801),.B(g16782));
  AND2 AND2_2544(.VSS(VSS),.VDD(VDD),.Y(g13887),.A(g5204),.B(g12402));
  AND2 AND2_2545(.VSS(VSS),.VDD(VDD),.Y(g25990),.A(g9461),.B(g25017));
  AND2 AND2_2546(.VSS(VSS),.VDD(VDD),.Y(g23497),.A(g20169),.B(g20569));
  AND3 AND3_156(.VSS(VSS),.VDD(VDD),.Y(g33509),.A(g32809),.B(I31241),.C(I31242));
  AND2 AND2_2547(.VSS(VSS),.VDD(VDD),.Y(g24669),.A(g22653),.B(g19742));
  AND2 AND2_2548(.VSS(VSS),.VDD(VDD),.Y(g31933),.A(g939),.B(g30735));
  AND2 AND2_2549(.VSS(VSS),.VDD(VDD),.Y(g30926),.A(g29903),.B(g21163));
  AND2 AND2_2550(.VSS(VSS),.VDD(VDD),.Y(g30045),.A(g29200),.B(g12419));
  AND2 AND2_2551(.VSS(VSS),.VDD(VDD),.Y(g18255),.A(g1087),.B(g16897));
  AND2 AND2_2552(.VSS(VSS),.VDD(VDD),.Y(g18189),.A(g812),.B(g17821));
  AND2 AND2_2553(.VSS(VSS),.VDD(VDD),.Y(g27588),.A(g26690),.B(g26673));
  AND2 AND2_2554(.VSS(VSS),.VDD(VDD),.Y(g15779),.A(g13909),.B(g11214));
  AND2 AND2_2555(.VSS(VSS),.VDD(VDD),.Y(g18679),.A(g4633),.B(g15758));
  AND2 AND2_2556(.VSS(VSS),.VDD(VDD),.Y(g31508),.A(g29813),.B(g23459));
  AND2 AND2_2557(.VSS(VSS),.VDD(VDD),.Y(g34389),.A(g34170),.B(g20715));
  AND2 AND2_2558(.VSS(VSS),.VDD(VDD),.Y(g17321),.A(g1418),.B(g13105));
  AND4 AND4_166(.VSS(VSS),.VDD(VDD),.Y(I31112),.A(g32617),.B(g32618),.C(g32619),.D(g32620));
  AND2 AND2_2559(.VSS(VSS),.VDD(VDD),.Y(g34045),.A(g33766),.B(g22942));
  AND2 AND2_2560(.VSS(VSS),.VDD(VDD),.Y(g30612),.A(g26338),.B(g29597));
  AND3 AND3_157(.VSS(VSS),.VDD(VDD),.Y(g33508),.A(g32802),.B(I31236),.C(I31237));
  AND2 AND2_2561(.VSS(VSS),.VDD(VDD),.Y(g24668),.A(g11754),.B(g22979));
  AND2 AND2_2562(.VSS(VSS),.VDD(VDD),.Y(g21700),.A(g150),.B(g20283));
  AND2 AND2_2563(.VSS(VSS),.VDD(VDD),.Y(g30099),.A(g28549),.B(g20776));
  AND2 AND2_2564(.VSS(VSS),.VDD(VDD),.Y(g33872),.A(g33282),.B(g20548));
  AND2 AND2_2565(.VSS(VSS),.VDD(VDD),.Y(g18270),.A(g1291),.B(g16031));
  AND2 AND2_2566(.VSS(VSS),.VDD(VDD),.Y(g29796),.A(g28345),.B(g23258));
  AND2 AND2_2567(.VSS(VSS),.VDD(VDD),.Y(g17179),.A(g1041),.B(g13211));
  AND2 AND2_2568(.VSS(VSS),.VDD(VDD),.Y(g24392),.A(g3115),.B(g23067));
  AND2 AND2_2569(.VSS(VSS),.VDD(VDD),.Y(g22685),.A(g11891),.B(g20192));
  AND2 AND2_2570(.VSS(VSS),.VDD(VDD),.Y(g18188),.A(g807),.B(g17328));
  AND2 AND2_2571(.VSS(VSS),.VDD(VDD),.Y(g18124),.A(g102),.B(g16886));
  AND2 AND2_2572(.VSS(VSS),.VDD(VDD),.Y(g21987),.A(g5579),.B(g19074));
  AND2 AND2_2573(.VSS(VSS),.VDD(VDD),.Y(g18678),.A(g66),.B(g15758));
  AND2 AND2_2574(.VSS(VSS),.VDD(VDD),.Y(g34388),.A(g10802),.B(g34062));
  AND2 AND2_2575(.VSS(VSS),.VDD(VDD),.Y(g16026),.A(g854),.B(g14065));
  AND2 AND2_2576(.VSS(VSS),.VDD(VDD),.Y(g28557),.A(g27772),.B(g15647));
  AND2 AND2_2577(.VSS(VSS),.VDD(VDD),.Y(g34324),.A(g14064),.B(g34161));
  AND2 AND2_2578(.VSS(VSS),.VDD(VDD),.Y(g15081),.A(g2689),.B(g12983));
  AND2 AND2_2579(.VSS(VSS),.VDD(VDD),.Y(g13393),.A(g703),.B(g11048));
  AND2 AND2_2580(.VSS(VSS),.VDD(VDD),.Y(g16212),.A(g6167),.B(g14321));
  AND2 AND2_2581(.VSS(VSS),.VDD(VDD),.Y(g24195),.A(g74),.B(g22722));
  AND2 AND2_2582(.VSS(VSS),.VDD(VDD),.Y(g28210),.A(g9229),.B(g27554));
  AND2 AND2_2583(.VSS(VSS),.VDD(VDD),.Y(g32317),.A(g5507),.B(g31542));
  AND2 AND2_2584(.VSS(VSS),.VDD(VDD),.Y(g27119),.A(g25877),.B(g22542));
  AND2 AND2_2585(.VSS(VSS),.VDD(VDD),.Y(g30098),.A(g28548),.B(g20774));
  AND2 AND2_2586(.VSS(VSS),.VDD(VDD),.Y(g34701),.A(g34536),.B(g20179));
  AND4 AND4_167(.VSS(VSS),.VDD(VDD),.Y(g10721),.A(g3288),.B(g6875),.C(g3274),.D(g8481));
  AND2 AND2_2587(.VSS(VSS),.VDD(VDD),.Y(g20559),.A(g336),.B(g15831));
  AND2 AND2_2588(.VSS(VSS),.VDD(VDD),.Y(g30251),.A(g28745),.B(g23940));
  AND2 AND2_2589(.VSS(VSS),.VDD(VDD),.Y(g34534),.A(g34321),.B(g19743));
  AND2 AND2_2590(.VSS(VSS),.VDD(VDD),.Y(g23658),.A(g14687),.B(g20852));
  AND2 AND2_2591(.VSS(VSS),.VDD(VDD),.Y(g30272),.A(g28814),.B(g23982));
  AND3 AND3_158(.VSS(VSS),.VDD(VDD),.Y(g34098),.A(g33744),.B(g9104),.C(g18957));
  AND2 AND2_2592(.VSS(VSS),.VDD(VDD),.Y(g19206),.A(g460),.B(g16206));
  AND2 AND2_2593(.VSS(VSS),.VDD(VDD),.Y(g15786),.A(g13940),.B(g11233));
  AND2 AND2_2594(.VSS(VSS),.VDD(VDD),.Y(g18460),.A(g2351),.B(g15224));
  AND2 AND2_2595(.VSS(VSS),.VDD(VDD),.Y(g18686),.A(g4659),.B(g15885));
  AND2 AND2_2596(.VSS(VSS),.VDD(VDD),.Y(g24559),.A(g22993),.B(g19567));
  AND2 AND2_2597(.VSS(VSS),.VDD(VDD),.Y(g18383),.A(g1950),.B(g15171));
  AND2 AND2_2598(.VSS(VSS),.VDD(VDD),.Y(g29840),.A(g2153),.B(g29056));
  AND2 AND2_2599(.VSS(VSS),.VDD(VDD),.Y(g24488),.A(g6905),.B(g23082));
  AND4 AND4_168(.VSS(VSS),.VDD(VDD),.Y(I31096),.A(g31376),.B(g31812),.C(g32594),.D(g32595));
  AND2 AND2_2600(.VSS(VSS),.VDD(VDD),.Y(g24016),.A(g14528),.B(g21610));
  AND2 AND2_2601(.VSS(VSS),.VDD(VDD),.Y(g27118),.A(g26055),.B(g16529));
  AND3 AND3_159(.VSS(VSS),.VDD(VDD),.Y(g22417),.A(g7753),.B(g9285),.C(g21186));
  AND2 AND2_2602(.VSS(VSS),.VDD(VDD),.Y(g11960),.A(g2495),.B(g7424));
  AND2 AND2_2603(.VSS(VSS),.VDD(VDD),.Y(g32129),.A(g31658),.B(g29955));
  AND2 AND2_2604(.VSS(VSS),.VDD(VDD),.Y(g21943),.A(g5240),.B(g18997));
  AND2 AND2_2605(.VSS(VSS),.VDD(VDD),.Y(g25832),.A(g8219),.B(g24625));
  AND2 AND2_2606(.VSS(VSS),.VDD(VDD),.Y(g21296),.A(g7879),.B(g16072));
  AND2 AND2_2607(.VSS(VSS),.VDD(VDD),.Y(g24558),.A(g22516),.B(g19566));
  AND2 AND2_2608(.VSS(VSS),.VDD(VDD),.Y(g18267),.A(g1266),.B(g16000));
  AND2 AND2_2609(.VSS(VSS),.VDD(VDD),.Y(g18294),.A(g15072),.B(g16449));
  AND2 AND2_2610(.VSS(VSS),.VDD(VDD),.Y(g27616),.A(g26349),.B(g20449));
  AND2 AND2_2611(.VSS(VSS),.VDD(VDD),.Y(g26871),.A(g25038),.B(g25020));
  AND2 AND2_2612(.VSS(VSS),.VDD(VDD),.Y(g17654),.A(g962),.B(g13284));
  AND2 AND2_2613(.VSS(VSS),.VDD(VDD),.Y(g32128),.A(g31631),.B(g29953));
  AND3 AND3_160(.VSS(VSS),.VDD(VDD),.Y(I17575),.A(g13156),.B(g11450),.C(g6756));
  AND2 AND2_2614(.VSS(VSS),.VDD(VDD),.Y(g27313),.A(g1982),.B(g26701));
  AND2 AND2_2615(.VSS(VSS),.VDD(VDD),.Y(g29192),.A(g27163),.B(g10290));
  AND2 AND2_2616(.VSS(VSS),.VDD(VDD),.Y(g30032),.A(g29072),.B(g9326));
  AND2 AND2_2617(.VSS(VSS),.VDD(VDD),.Y(g21969),.A(g5373),.B(g21514));
  AND2 AND2_2618(.VSS(VSS),.VDD(VDD),.Y(g26360),.A(g10589),.B(g25533));
  AND2 AND2_2619(.VSS(VSS),.VDD(VDD),.Y(g25573),.A(I24704),.B(I24705));
  AND2 AND2_2620(.VSS(VSS),.VDD(VDD),.Y(g30140),.A(g28600),.B(g23749));
  AND2 AND2_2621(.VSS(VSS),.VDD(VDD),.Y(g27276),.A(g9750),.B(g26607));
  AND2 AND2_2622(.VSS(VSS),.VDD(VDD),.Y(g27285),.A(g9912),.B(g26632));
  AND2 AND2_2623(.VSS(VSS),.VDD(VDD),.Y(g29522),.A(g28923),.B(g22369));
  AND2 AND2_2624(.VSS(VSS),.VDD(VDD),.Y(g32323),.A(g31311),.B(g20610));
  AND2 AND2_2625(.VSS(VSS),.VDD(VDD),.Y(g24865),.A(g11323),.B(g23253));
  AND2 AND2_2626(.VSS(VSS),.VDD(VDD),.Y(g29663),.A(g1950),.B(g28693));
  AND2 AND2_2627(.VSS(VSS),.VDD(VDD),.Y(g34140),.A(g33931),.B(g23802));
  AND2 AND2_2628(.VSS(VSS),.VDD(VDD),.Y(g22762),.A(g9305),.B(g20645));
  AND2 AND2_2629(.VSS(VSS),.VDD(VDD),.Y(g15651),.A(g429),.B(g13414));
  AND2 AND2_2630(.VSS(VSS),.VDD(VDD),.Y(g21968),.A(g5459),.B(g21514));
  AND2 AND2_2631(.VSS(VSS),.VDD(VDD),.Y(g10655),.A(g8440),.B(g3423));
  AND2 AND2_2632(.VSS(VSS),.VDD(VDD),.Y(g15672),.A(g433),.B(g13458));
  AND2 AND2_2633(.VSS(VSS),.VDD(VDD),.Y(g27305),.A(g10041),.B(g26683));
  AND2 AND2_2634(.VSS(VSS),.VDD(VDD),.Y(g25926),.A(g25005),.B(g24839));
  AND2 AND2_2635(.VSS(VSS),.VDD(VDD),.Y(g24713),.A(g5831),.B(g23666));
  AND2 AND2_2636(.VSS(VSS),.VDD(VDD),.Y(g25045),.A(g17525),.B(g23448));
  AND2 AND2_2637(.VSS(VSS),.VDD(VDD),.Y(g18219),.A(g969),.B(g16100));
  AND2 AND2_2638(.VSS(VSS),.VDD(VDD),.Y(g27254),.A(g25935),.B(g19688));
  AND2 AND2_2639(.VSS(VSS),.VDD(VDD),.Y(g30061),.A(g1036),.B(g28188));
  AND2 AND2_2640(.VSS(VSS),.VDD(VDD),.Y(g33311),.A(g31942),.B(g12925));
  AND2 AND2_2641(.VSS(VSS),.VDD(VDD),.Y(g21855),.A(g3925),.B(g21070));
  AND2 AND2_2642(.VSS(VSS),.VDD(VDD),.Y(g34061),.A(g33800),.B(g23076));
  AND2 AND2_2643(.VSS(VSS),.VDD(VDD),.Y(g14180),.A(g872),.B(g10632));
  AND2 AND2_2644(.VSS(VSS),.VDD(VDD),.Y(g23855),.A(g4112),.B(g19455));
  AND2 AND2_2645(.VSS(VSS),.VDD(VDD),.Y(g22216),.A(g13660),.B(g20000));
  AND2 AND2_2646(.VSS(VSS),.VDD(VDD),.Y(g18218),.A(g1008),.B(g16100));
  AND2 AND2_2647(.VSS(VSS),.VDD(VDD),.Y(g21870),.A(g4093),.B(g19801));
  AND3 AND3_161(.VSS(VSS),.VDD(VDD),.Y(I17606),.A(g14988),.B(g11450),.C(g6756));
  AND2 AND2_2648(.VSS(VSS),.VDD(VDD),.Y(g28601),.A(g27506),.B(g20514));
  AND2 AND2_2649(.VSS(VSS),.VDD(VDD),.Y(g28677),.A(g27571),.B(g20635));
  AND2 AND2_2650(.VSS(VSS),.VDD(VDD),.Y(g27036),.A(g26329),.B(g11038));
  AND2 AND2_2651(.VSS(VSS),.VDD(VDD),.Y(g29553),.A(g2437),.B(g28911));
  AND2 AND2_2652(.VSS(VSS),.VDD(VDD),.Y(g26629),.A(g14173),.B(g24418));
  AND2 AND2_2653(.VSS(VSS),.VDD(VDD),.Y(g27177),.A(g25997),.B(g16651));
  AND2 AND2_2654(.VSS(VSS),.VDD(VDD),.Y(g27560),.A(g26299),.B(g20191));
  AND2 AND2_2655(.VSS(VSS),.VDD(VDD),.Y(g34871),.A(g34823),.B(g19908));
  AND2 AND2_2656(.VSS(VSS),.VDD(VDD),.Y(g24189),.A(g324),.B(g22722));
  AND2 AND2_2657(.VSS(VSS),.VDD(VDD),.Y(g31756),.A(g30114),.B(g23942));
  AND2 AND2_2658(.VSS(VSS),.VDD(VDD),.Y(g24679),.A(g13289),.B(g22985));
  AND2 AND2_2659(.VSS(VSS),.VDD(VDD),.Y(g11244),.A(g8346),.B(g8566));
  AND2 AND2_2660(.VSS(VSS),.VDD(VDD),.Y(g29949),.A(g23575),.B(g28924));
  AND2 AND2_2661(.VSS(VSS),.VDD(VDD),.Y(g32232),.A(g31241),.B(g20266));
  AND2 AND2_2662(.VSS(VSS),.VDD(VDD),.Y(g20188),.A(g5849),.B(g17772));
  AND2 AND2_2663(.VSS(VSS),.VDD(VDD),.Y(g18160),.A(g645),.B(g17433));
  AND2 AND2_2664(.VSS(VSS),.VDD(VDD),.Y(g29326),.A(g29105),.B(g22155));
  AND3 AND3_162(.VSS(VSS),.VDD(VDD),.Y(g10838),.A(g7738),.B(g5527),.C(g5535));
  AND2 AND2_2665(.VSS(VSS),.VDD(VDD),.Y(g28143),.A(g27344),.B(g26083));
  AND2 AND2_2666(.VSS(VSS),.VDD(VDD),.Y(g31780),.A(g30163),.B(g23999));
  AND3 AND3_163(.VSS(VSS),.VDD(VDD),.Y(g25462),.A(g6404),.B(g22300),.C(I24585));
  AND2 AND2_2667(.VSS(VSS),.VDD(VDD),.Y(g24188),.A(g316),.B(g22722));
  AND2 AND2_2668(.VSS(VSS),.VDD(VDD),.Y(g22117),.A(g6597),.B(g19277));
  AND2 AND2_2669(.VSS(VSS),.VDD(VDD),.Y(g29536),.A(g28969),.B(g22432));
  AND2 AND2_2670(.VSS(VSS),.VDD(VDD),.Y(g22000),.A(g5727),.B(g21562));
  AND2 AND2_2671(.VSS(VSS),.VDD(VDD),.Y(g21867),.A(g4082),.B(g19801));
  AND2 AND2_2672(.VSS(VSS),.VDD(VDD),.Y(g18455),.A(g2327),.B(g15224));
  AND2 AND2_2673(.VSS(VSS),.VDD(VDD),.Y(g24686),.A(g5485),.B(g23630));
  AND2 AND2_2674(.VSS(VSS),.VDD(VDD),.Y(g24939),.A(g23771),.B(g21012));
  AND2 AND2_2675(.VSS(VSS),.VDD(VDD),.Y(g29757),.A(g28305),.B(g23221));
  AND4 AND4_169(.VSS(VSS),.VDD(VDD),.Y(I31317),.A(g32914),.B(g32915),.C(g32916),.D(g32917));
  AND2 AND2_2676(.VSS(VSS),.VDD(VDD),.Y(g33350),.A(g32235),.B(g20702));
  AND2 AND2_2677(.VSS(VSS),.VDD(VDD),.Y(g32261),.A(g31251),.B(g20386));
  AND2 AND2_2678(.VSS(VSS),.VDD(VDD),.Y(g18617),.A(g3462),.B(g17062));
  AND2 AND2_2679(.VSS(VSS),.VDD(VDD),.Y(g18470),.A(g2403),.B(g15224));
  AND2 AND2_2680(.VSS(VSS),.VDD(VDD),.Y(g20093),.A(g15372),.B(g14584));
  AND2 AND2_2681(.VSS(VSS),.VDD(VDD),.Y(g33820),.A(g33075),.B(g26830));
  AND2 AND2_2682(.VSS(VSS),.VDD(VDD),.Y(g29621),.A(g2449),.B(g28994));
  AND3 AND3_164(.VSS(VSS),.VDD(VDD),.Y(I24576),.A(g5390),.B(g5396),.C(g9792));
  AND3 AND3_165(.VSS(VSS),.VDD(VDD),.Y(I24585),.A(g9621),.B(g9892),.C(g6439));
  AND2 AND2_2683(.VSS(VSS),.VDD(VDD),.Y(g10619),.A(g3080),.B(g7907));
  AND2 AND2_2684(.VSS(VSS),.VDD(VDD),.Y(g21714),.A(g278),.B(g20283));
  AND2 AND2_2685(.VSS(VSS),.VDD(VDD),.Y(g23581),.A(g20183),.B(g11900));
  AND2 AND2_2686(.VSS(VSS),.VDD(VDD),.Y(g24294),.A(g4452),.B(g22550));
  AND2 AND2_2687(.VSS(VSS),.VDD(VDD),.Y(g31152),.A(g10039),.B(g30067));
  AND2 AND2_2688(.VSS(VSS),.VDD(VDD),.Y(g25061),.A(g17586),.B(g23461));
  AND4 AND4_170(.VSS(VSS),.VDD(VDD),.Y(I31002),.A(g32459),.B(g32460),.C(g32461),.D(g32462));
  AND2 AND2_2689(.VSS(VSS),.VDD(VDD),.Y(g18201),.A(g15061),.B(g15938));
  AND2 AND2_2690(.VSS(VSS),.VDD(VDD),.Y(g33846),.A(g33259),.B(g20380));
  AND4 AND4_171(.VSS(VSS),.VDD(VDD),.Y(I31057),.A(g32538),.B(g32539),.C(g32540),.D(g32541));
  AND2 AND2_2691(.VSS(VSS),.VDD(VDD),.Y(g21707),.A(g191),.B(g20283));
  AND2 AND2_2692(.VSS(VSS),.VDD(VDD),.Y(g21819),.A(g3614),.B(g20924));
  AND2 AND2_2693(.VSS(VSS),.VDD(VDD),.Y(g29564),.A(g1882),.B(g28896));
  AND2 AND2_2694(.VSS(VSS),.VDD(VDD),.Y(g18277),.A(g1312),.B(g16136));
  AND2 AND2_2695(.VSS(VSS),.VDD(VDD),.Y(g14210),.A(g4392),.B(g10590));
  AND2 AND2_2696(.VSS(VSS),.VDD(VDD),.Y(g21910),.A(g5016),.B(g21468));
  AND2 AND2_2697(.VSS(VSS),.VDD(VDD),.Y(g26147),.A(g6513),.B(g25133));
  AND2 AND2_2698(.VSS(VSS),.VDD(VDD),.Y(g30220),.A(g28699),.B(g23888));
  AND2 AND2_2699(.VSS(VSS),.VDD(VDD),.Y(g28666),.A(g27567),.B(g20625));
  AND2 AND2_2700(.VSS(VSS),.VDD(VDD),.Y(g33731),.A(g33116),.B(g19520));
  AND2 AND2_2701(.VSS(VSS),.VDD(VDD),.Y(g28217),.A(g27733),.B(g23391));
  AND2 AND2_2702(.VSS(VSS),.VDD(VDD),.Y(g22123),.A(g6609),.B(g19277));
  AND2 AND2_2703(.VSS(VSS),.VDD(VDD),.Y(g21818),.A(g3610),.B(g20924));
  AND4 AND4_172(.VSS(VSS),.VDD(VDD),.Y(g17747),.A(g6772),.B(g11592),.C(g11640),.D(I18740));
  AND2 AND2_2704(.VSS(VSS),.VDD(VDD),.Y(g21979),.A(g5559),.B(g19074));
  AND2 AND2_2705(.VSS(VSS),.VDD(VDD),.Y(g16896),.A(g262),.B(g13120));
  AND2 AND2_2706(.VSS(VSS),.VDD(VDD),.Y(g27665),.A(g26872),.B(g23519));
  AND2 AND2_2707(.VSS(VSS),.VDD(VDD),.Y(g30246),.A(g28734),.B(g23936));
  AND2 AND2_2708(.VSS(VSS),.VDD(VDD),.Y(g25871),.A(g8334),.B(g24804));
  AND2 AND2_2709(.VSS(VSS),.VDD(VDD),.Y(g20875),.A(g16281),.B(g4681));
  AND2 AND2_2710(.VSS(VSS),.VDD(VDD),.Y(g18595),.A(g2927),.B(g16349));
  AND2 AND2_2711(.VSS(VSS),.VDD(VDD),.Y(g28478),.A(g27007),.B(g12345));
  AND2 AND2_2712(.VSS(VSS),.VDD(VDD),.Y(g18467),.A(g2380),.B(g15224));
  AND2 AND2_2713(.VSS(VSS),.VDD(VDD),.Y(g18494),.A(g2527),.B(g15426));
  AND2 AND2_2714(.VSS(VSS),.VDD(VDD),.Y(g19500),.A(g504),.B(g16712));
  AND2 AND2_2715(.VSS(VSS),.VDD(VDD),.Y(g24219),.A(g225),.B(g22594));
  AND2 AND2_2716(.VSS(VSS),.VDD(VDD),.Y(g26858),.A(g2970),.B(g24540));
  AND2 AND2_2717(.VSS(VSS),.VDD(VDD),.Y(g21978),.A(g5551),.B(g19074));
  AND2 AND2_2718(.VSS(VSS),.VDD(VDD),.Y(g11967),.A(g311),.B(g7802));
  AND2 AND2_2719(.VSS(VSS),.VDD(VDD),.Y(g18623),.A(g3484),.B(g17062));
  AND2 AND2_2720(.VSS(VSS),.VDD(VDD),.Y(g20218),.A(g6541),.B(g17815));
  AND2 AND2_2721(.VSS(VSS),.VDD(VDD),.Y(g30071),.A(g29184),.B(g12975));
  AND2 AND2_2722(.VSS(VSS),.VDD(VDD),.Y(g17123),.A(g225),.B(g13209));
  AND2 AND2_2723(.VSS(VSS),.VDD(VDD),.Y(g24218),.A(g872),.B(g22594));
  AND2 AND2_2724(.VSS(VSS),.VDD(VDD),.Y(g21986),.A(g5575),.B(g19074));
  AND2 AND2_2725(.VSS(VSS),.VDD(VDD),.Y(g34071),.A(g8854),.B(g33799));
  AND2 AND2_2726(.VSS(VSS),.VDD(VDD),.Y(g18782),.A(g5835),.B(g18065));
  AND2 AND2_2727(.VSS(VSS),.VDD(VDD),.Y(g27485),.A(g26519),.B(g17644));
  AND2 AND2_2728(.VSS(VSS),.VDD(VDD),.Y(g28556),.A(g27431),.B(g20374));
  AND2 AND2_2729(.VSS(VSS),.VDD(VDD),.Y(g29509),.A(g1600),.B(g28755));
  AND2 AND2_2730(.VSS(VSS),.VDD(VDD),.Y(g32316),.A(g31307),.B(g23522));
  AND2 AND2_2731(.VSS(VSS),.VDD(VDD),.Y(g33405),.A(g32354),.B(g21398));
  AND2 AND2_2732(.VSS(VSS),.VDD(VDD),.Y(g21741),.A(g15086),.B(g20330));
  AND2 AND2_2733(.VSS(VSS),.VDD(VDD),.Y(g26844),.A(g25261),.B(g21418));
  AND2 AND2_2734(.VSS(VSS),.VDD(VDD),.Y(g18419),.A(g2051),.B(g15373));
  AND2 AND2_2735(.VSS(VSS),.VDD(VDD),.Y(g27454),.A(g26488),.B(g17602));
  AND2 AND2_2736(.VSS(VSS),.VDD(VDD),.Y(g26394),.A(g22530),.B(g25560));
  AND2 AND2_2737(.VSS(VSS),.VDD(VDD),.Y(g18352),.A(g1798),.B(g17955));
  AND2 AND2_2738(.VSS(VSS),.VDD(VDD),.Y(g29634),.A(g2108),.B(g29121));
  AND2 AND2_2739(.VSS(VSS),.VDD(VDD),.Y(g29851),.A(g1668),.B(g29079));
  AND2 AND2_2740(.VSS(VSS),.VDD(VDD),.Y(g29872),.A(g28401),.B(g23333));
  AND2 AND2_2741(.VSS(VSS),.VDD(VDD),.Y(g28223),.A(g27338),.B(g17194));
  AND2 AND2_2742(.VSS(VSS),.VDD(VDD),.Y(g15104),.A(g6955),.B(g14454));
  AND2 AND2_2743(.VSS(VSS),.VDD(VDD),.Y(g34754),.A(g34677),.B(g19602));
  AND2 AND2_2744(.VSS(VSS),.VDD(VDD),.Y(g18155),.A(g15056),.B(g17533));
  AND2 AND2_2745(.VSS(VSS),.VDD(VDD),.Y(g21067),.A(g10085),.B(g17625));
  AND2 AND2_2746(.VSS(VSS),.VDD(VDD),.Y(g18418),.A(g2122),.B(g15373));
  AND2 AND2_2747(.VSS(VSS),.VDD(VDD),.Y(g18822),.A(g6723),.B(g15680));
  AND2 AND2_2748(.VSS(VSS),.VDD(VDD),.Y(g30825),.A(g29814),.B(g22332));
  AND2 AND2_2749(.VSS(VSS),.VDD(VDD),.Y(g19613),.A(g1437),.B(g16713));
  AND2 AND2_2750(.VSS(VSS),.VDD(VDD),.Y(g32056),.A(g27271),.B(g31021));
  AND2 AND2_2751(.VSS(VSS),.VDD(VDD),.Y(g18266),.A(g1274),.B(g16000));
  AND2 AND2_2752(.VSS(VSS),.VDD(VDD),.Y(g11010),.A(g4698),.B(g8933));
  AND2 AND2_2753(.VSS(VSS),.VDD(VDD),.Y(g34859),.A(g16540),.B(g34820));
  AND2 AND2_2754(.VSS(VSS),.VDD(VDD),.Y(g18170),.A(g661),.B(g17433));
  AND4 AND4_173(.VSS(VSS),.VDD(VDD),.Y(I31232),.A(g32791),.B(g32792),.C(g32793),.D(g32794));
  AND2 AND2_2755(.VSS(VSS),.VDD(VDD),.Y(g10677),.A(g4141),.B(g7611));
  AND2 AND2_2756(.VSS(VSS),.VDD(VDD),.Y(g22992),.A(g1227),.B(g19765));
  AND2 AND2_2757(.VSS(VSS),.VDD(VDD),.Y(g34370),.A(g34067),.B(g10554));
  AND4 AND4_174(.VSS(VSS),.VDD(VDD),.Y(I24674),.A(g19919),.B(g24019),.C(g24020),.D(g24021));
  AND2 AND2_2758(.VSS(VSS),.VDD(VDD),.Y(g21801),.A(g3554),.B(g20924));
  AND2 AND2_2759(.VSS(VSS),.VDD(VDD),.Y(g28110),.A(g27974),.B(g18886));
  AND2 AND2_2760(.VSS(VSS),.VDD(VDD),.Y(g21735),.A(g3057),.B(g20330));
  AND2 AND2_2761(.VSS(VSS),.VDD(VDD),.Y(g21877),.A(g6888),.B(g19801));
  AND2 AND2_2762(.VSS(VSS),.VDD(VDD),.Y(g23801),.A(g1448),.B(g19362));
  AND2 AND2_2763(.VSS(VSS),.VDD(VDD),.Y(g34858),.A(g16540),.B(g34816));
  AND2 AND2_2764(.VSS(VSS),.VDD(VDD),.Y(g30151),.A(g28607),.B(g21249));
  AND2 AND2_2765(.VSS(VSS),.VDD(VDD),.Y(g30172),.A(g28625),.B(g21286));
  AND2 AND2_2766(.VSS(VSS),.VDD(VDD),.Y(g24915),.A(g23087),.B(g20158));
  AND4 AND4_175(.VSS(VSS),.VDD(VDD),.Y(I31261),.A(g30937),.B(g31842),.C(g32831),.D(g32832));
  AND2 AND2_2767(.VSS(VSS),.VDD(VDD),.Y(g27594),.A(g26721),.B(g26694));
  AND2 AND2_2768(.VSS(VSS),.VDD(VDD),.Y(g28531),.A(g27722),.B(g15608));
  AND2 AND2_2769(.VSS(VSS),.VDD(VDD),.Y(g17391),.A(g9556),.B(g14378));
  AND2 AND2_2770(.VSS(VSS),.VDD(VDD),.Y(g22835),.A(g15803),.B(g19633));
  AND2 AND2_2771(.VSS(VSS),.VDD(VDD),.Y(g28178),.A(g27019),.B(g19397));
  AND2 AND2_2772(.VSS(VSS),.VDD(VDD),.Y(g18167),.A(g718),.B(g17433));
  AND2 AND2_2773(.VSS(VSS),.VDD(VDD),.Y(g18194),.A(g843),.B(g17821));
  AND2 AND2_2774(.VSS(VSS),.VDD(VDD),.Y(g18589),.A(g2902),.B(g16349));
  AND2 AND2_2775(.VSS(VSS),.VDD(VDD),.Y(g22014),.A(g5805),.B(g21562));
  AND2 AND2_2776(.VSS(VSS),.VDD(VDD),.Y(g34367),.A(g7404),.B(g34042));
  AND2 AND2_2777(.VSS(VSS),.VDD(VDD),.Y(g31787),.A(g21281),.B(g29385));
  AND2 AND2_2778(.VSS(VSS),.VDD(VDD),.Y(g34394),.A(g34190),.B(g21305));
  AND2 AND2_2779(.VSS(VSS),.VDD(VDD),.Y(g25071),.A(g12804),.B(g23478));
  AND2 AND2_2780(.VSS(VSS),.VDD(VDD),.Y(g33113),.A(g31964),.B(g22339));
  AND2 AND2_2781(.VSS(VSS),.VDD(VDD),.Y(g33787),.A(g33103),.B(g20595));
  AND2 AND2_2782(.VSS(VSS),.VDD(VDD),.Y(g32342),.A(g6545),.B(g31579));
  AND2 AND2_2783(.VSS(VSS),.VDD(VDD),.Y(g29574),.A(g2016),.B(g28931));
  AND2 AND2_2784(.VSS(VSS),.VDD(VDD),.Y(g31282),.A(g30130),.B(g27779));
  AND2 AND2_2785(.VSS(VSS),.VDD(VDD),.Y(g22007),.A(g5770),.B(g21562));
  AND2 AND2_2786(.VSS(VSS),.VDD(VDD),.Y(g15850),.A(g3606),.B(g14151));
  AND3 AND3_166(.VSS(VSS),.VDD(VDD),.Y(g29205),.A(g24117),.B(I27523),.C(I27524));
  AND2 AND2_2787(.VSS(VSS),.VDD(VDD),.Y(g18588),.A(g2970),.B(g16349));
  AND2 AND2_2788(.VSS(VSS),.VDD(VDD),.Y(g18524),.A(g2681),.B(g15509));
  AND2 AND2_2789(.VSS(VSS),.VDD(VDD),.Y(g28676),.A(g27570),.B(g20632));
  AND2 AND2_2790(.VSS(VSS),.VDD(VDD),.Y(g32145),.A(g31609),.B(g29977));
  AND2 AND2_2791(.VSS(VSS),.VDD(VDD),.Y(g14791),.A(g1146),.B(g10909));
  AND2 AND2_2792(.VSS(VSS),.VDD(VDD),.Y(g32031),.A(g31372),.B(g13464));
  AND2 AND2_2793(.VSS(VSS),.VDD(VDD),.Y(g24467),.A(g13761),.B(g23047));
  AND2 AND2_2794(.VSS(VSS),.VDD(VDD),.Y(g27519),.A(g26488),.B(g17710));
  AND2 AND2_2795(.VSS(VSS),.VDD(VDD),.Y(g33357),.A(g32247),.B(g20775));
  AND3 AND3_167(.VSS(VSS),.VDD(VDD),.Y(g27185),.A(g26190),.B(g8302),.C(g1917));
  AND2 AND2_2796(.VSS(VSS),.VDD(VDD),.Y(g25147),.A(g20202),.B(g23542));
  AND2 AND2_2797(.VSS(VSS),.VDD(VDD),.Y(g32199),.A(g30916),.B(g25506));
  AND2 AND2_2798(.VSS(VSS),.VDD(VDD),.Y(g18401),.A(g2036),.B(g15373));
  AND2 AND2_2799(.VSS(VSS),.VDD(VDD),.Y(g28654),.A(g1030),.B(g27108));
  AND2 AND2_2800(.VSS(VSS),.VDD(VDD),.Y(g33105),.A(g26298),.B(g32138));
  AND2 AND2_2801(.VSS(VSS),.VDD(VDD),.Y(g14168),.A(g887),.B(g10632));
  AND2 AND2_2802(.VSS(VSS),.VDD(VDD),.Y(g18477),.A(g2429),.B(g15426));
  AND2 AND2_2803(.VSS(VSS),.VDD(VDD),.Y(g26203),.A(g1632),.B(g25337));
  AND2 AND2_2804(.VSS(VSS),.VDD(VDD),.Y(g33743),.A(g33119),.B(g19574));
  AND2 AND2_2805(.VSS(VSS),.VDD(VDD),.Y(g16802),.A(g5567),.B(g14807));
  AND2 AND2_2806(.VSS(VSS),.VDD(VDD),.Y(g18119),.A(g475),.B(g17015));
  AND2 AND2_2807(.VSS(VSS),.VDD(VDD),.Y(g27518),.A(g26488),.B(g17709));
  AND2 AND2_2808(.VSS(VSS),.VDD(VDD),.Y(g27154),.A(g26055),.B(g16630));
  AND2 AND2_2809(.VSS(VSS),.VDD(VDD),.Y(g34319),.A(g9535),.B(g34156));
  AND2 AND2_2810(.VSS(VSS),.VDD(VDD),.Y(g32198),.A(g4253),.B(g31327));
  AND2 AND2_2811(.VSS(VSS),.VDD(VDD),.Y(g22116),.A(g6589),.B(g19277));
  AND2 AND2_2812(.VSS(VSS),.VDD(VDD),.Y(g16730),.A(g5212),.B(g14723));
  AND2 AND2_2813(.VSS(VSS),.VDD(VDD),.Y(g24984),.A(g22929),.B(g12818));
  AND2 AND2_2814(.VSS(VSS),.VDD(VDD),.Y(g18118),.A(g471),.B(g17015));
  AND2 AND2_2815(.VSS(VSS),.VDD(VDD),.Y(g21866),.A(g4072),.B(g19801));
  AND2 AND2_2816(.VSS(VSS),.VDD(VDD),.Y(g21917),.A(g5092),.B(g21468));
  AND2 AND2_2817(.VSS(VSS),.VDD(VDD),.Y(g30227),.A(g28708),.B(g23899));
  AND2 AND2_2818(.VSS(VSS),.VDD(VDD),.Y(g31769),.A(g30141),.B(g23986));
  AND2 AND2_2819(.VSS(VSS),.VDD(VDD),.Y(g23917),.A(g1472),.B(g19428));
  AND2 AND2_2820(.VSS(VSS),.VDD(VDD),.Y(g33640),.A(g33387),.B(g18831));
  AND4 AND4_176(.VSS(VSS),.VDD(VDD),.Y(g26281),.A(g24688),.B(g8812),.C(g8778),.D(g8757));
  AND2 AND2_2821(.VSS(VSS),.VDD(VDD),.Y(g32330),.A(g31320),.B(g20631));
  AND2 AND2_2822(.VSS(VSS),.VDD(VDD),.Y(g29592),.A(g28469),.B(g11832));
  AND2 AND2_2823(.VSS(VSS),.VDD(VDD),.Y(g30059),.A(g28106),.B(g12467));
  AND2 AND2_2824(.VSS(VSS),.VDD(VDD),.Y(g22720),.A(g9253),.B(g20619));
  AND4 AND4_177(.VSS(VSS),.VDD(VDD),.Y(I31316),.A(g29385),.B(g32911),.C(g32912),.D(g32913));
  AND2 AND2_2825(.VSS(VSS),.VDD(VDD),.Y(g30025),.A(g28492),.B(g23502));
  AND2 AND2_2826(.VSS(VSS),.VDD(VDD),.Y(g25151),.A(g17719),.B(g23549));
  AND2 AND2_2827(.VSS(VSS),.VDD(VDD),.Y(g16765),.A(g6581),.B(g15045));
  AND2 AND2_2828(.VSS(VSS),.VDD(VDD),.Y(g15716),.A(g468),.B(g13437));
  AND2 AND2_2829(.VSS(VSS),.VDD(VDD),.Y(g18749),.A(g5148),.B(g17847));
  AND2 AND2_2830(.VSS(VSS),.VDD(VDD),.Y(g22041),.A(g5957),.B(g19147));
  AND2 AND2_2831(.VSS(VSS),.VDD(VDD),.Y(g26301),.A(g2145),.B(g25244));
  AND2 AND2_2832(.VSS(VSS),.VDD(VDD),.Y(g13656),.A(g278),.B(g11144));
  AND2 AND2_2833(.VSS(VSS),.VDD(VDD),.Y(g18616),.A(g6875),.B(g17200));
  AND2 AND2_2834(.VSS(VSS),.VDD(VDD),.Y(g18313),.A(g1430),.B(g16931));
  AND2 AND2_2835(.VSS(VSS),.VDD(VDD),.Y(g33803),.A(g33231),.B(g20071));
  AND3 AND3_168(.VSS(VSS),.VDD(VDD),.Y(g24822),.A(g3010),.B(g23534),.C(I24003));
  AND2 AND2_2836(.VSS(VSS),.VDD(VDD),.Y(g26120),.A(g9809),.B(g25293));
  AND2 AND2_2837(.VSS(VSS),.VDD(VDD),.Y(g30058),.A(g29180),.B(g12950));
  AND2 AND2_2838(.VSS(VSS),.VDD(VDD),.Y(g16690),.A(g8399),.B(g13867));
  AND4 AND4_178(.VSS(VSS),.VDD(VDD),.Y(g11144),.A(g239),.B(g8136),.C(g246),.D(I14198));
  AND2 AND2_2839(.VSS(VSS),.VDD(VDD),.Y(g18748),.A(g5142),.B(g17847));
  AND2 AND2_2840(.VSS(VSS),.VDD(VDD),.Y(g8643),.A(g2927),.B(g2922));
  AND2 AND2_2841(.VSS(VSS),.VDD(VDD),.Y(g25367),.A(g6946),.B(g22407));
  AND4 AND4_179(.VSS(VSS),.VDD(VDD),.Y(I31056),.A(g30735),.B(g31805),.C(g32536),.D(g32537));
  AND2 AND2_2842(.VSS(VSS),.VDD(VDD),.Y(g21706),.A(g222),.B(g20283));
  AND2 AND2_2843(.VSS(VSS),.VDD(VDD),.Y(g18276),.A(g1351),.B(g16136));
  AND2 AND2_2844(.VSS(VSS),.VDD(VDD),.Y(g18285),.A(g1395),.B(g16164));
  AND2 AND2_2845(.VSS(VSS),.VDD(VDD),.Y(g29350),.A(g4939),.B(g28395));
  AND2 AND2_2846(.VSS(VSS),.VDD(VDD),.Y(g26146),.A(g9892),.B(g25334));
  AND2 AND2_2847(.VSS(VSS),.VDD(VDD),.Y(g30203),.A(g28668),.B(g23864));
  AND2 AND2_2848(.VSS(VSS),.VDD(VDD),.Y(g18704),.A(g4793),.B(g16782));
  AND2 AND2_2849(.VSS(VSS),.VDD(VDD),.Y(g34203),.A(g33726),.B(g24537));
  AND2 AND2_2850(.VSS(VSS),.VDD(VDD),.Y(g18305),.A(g1521),.B(g16489));
  AND2 AND2_2851(.VSS(VSS),.VDD(VDD),.Y(g33881),.A(g33292),.B(g20586));
  AND2 AND2_2852(.VSS(VSS),.VDD(VDD),.Y(g30044),.A(g29174),.B(g12944));
  AND2 AND2_2853(.VSS(VSS),.VDD(VDD),.Y(g18254),.A(g1236),.B(g16897));
  AND2 AND2_2854(.VSS(VSS),.VDD(VDD),.Y(g18809),.A(g7074),.B(g15656));
  AND2 AND2_2855(.VSS(VSS),.VDD(VDD),.Y(g21923),.A(g5029),.B(g21468));
  AND2 AND2_2856(.VSS(VSS),.VDD(VDD),.Y(g22340),.A(g19605),.B(g13522));
  AND2 AND2_2857(.VSS(VSS),.VDD(VDD),.Y(g32161),.A(g3151),.B(g31154));
  AND2 AND2_2858(.VSS(VSS),.VDD(VDD),.Y(g22035),.A(g5933),.B(g19147));
  AND2 AND2_2859(.VSS(VSS),.VDD(VDD),.Y(g28587),.A(g27487),.B(g20498));
  AND2 AND2_2860(.VSS(VSS),.VDD(VDD),.Y(g26290),.A(g2595),.B(g25498));
  AND2 AND2_2861(.VSS(VSS),.VDD(VDD),.Y(g18466),.A(g2389),.B(g15224));
  AND2 AND2_2862(.VSS(VSS),.VDD(VDD),.Y(g23280),.A(g19417),.B(g20146));
  AND2 AND2_2863(.VSS(VSS),.VDD(VDD),.Y(g27215),.A(g26055),.B(g16724));
  AND2 AND2_2864(.VSS(VSS),.VDD(VDD),.Y(g27501),.A(g26400),.B(g17673));
  AND2 AND2_2865(.VSS(VSS),.VDD(VDD),.Y(g15112),.A(g4284),.B(g14454));
  AND4 AND4_180(.VSS(VSS),.VDD(VDD),.Y(I31271),.A(g29385),.B(g32846),.C(g32847),.D(g32848));
  AND2 AND2_2866(.VSS(VSS),.VDD(VDD),.Y(g30281),.A(g28850),.B(g23992));
  AND2 AND2_2867(.VSS(VSS),.VDD(VDD),.Y(g18808),.A(g6390),.B(g15656));
  AND3 AND3_169(.VSS(VSS),.VDD(VDD),.Y(g25420),.A(g6058),.B(g22220),.C(I24555));
  AND2 AND2_2868(.VSS(VSS),.VDD(VDD),.Y(g24194),.A(g106),.B(g22722));
  AND2 AND2_2869(.VSS(VSS),.VDD(VDD),.Y(g24589),.A(g5471),.B(g23630));
  AND2 AND2_2870(.VSS(VSS),.VDD(VDD),.Y(g34281),.A(g34043),.B(g19276));
  AND2 AND2_2871(.VSS(VSS),.VDD(VDD),.Y(g29731),.A(g2089),.B(g29118));
  AND2 AND2_2872(.VSS(VSS),.VDD(VDD),.Y(g22142),.A(g7957),.B(g19140));
  AND2 AND2_2873(.VSS(VSS),.VDD(VDD),.Y(g27439),.A(g232),.B(g26831));
  AND2 AND2_2874(.VSS(VSS),.VDD(VDD),.Y(g34301),.A(g34064),.B(g19415));
  AND2 AND2_2875(.VSS(VSS),.VDD(VDD),.Y(g18177),.A(g749),.B(g17328));
  AND2 AND2_2876(.VSS(VSS),.VDD(VDD),.Y(g18560),.A(g2837),.B(g15277));
  AND2 AND2_2877(.VSS(VSS),.VDD(VDD),.Y(g30120),.A(g28576),.B(g21051));
  AND2 AND2_2878(.VSS(VSS),.VDD(VDD),.Y(g28543),.A(g27735),.B(g15628));
  AND2 AND2_2879(.VSS(VSS),.VDD(VDD),.Y(g24588),.A(g5142),.B(g23590));
  AND2 AND2_2880(.VSS(VSS),.VDD(VDD),.Y(g32087),.A(g1291),.B(g30825));
  AND2 AND2_2881(.VSS(VSS),.VDD(VDD),.Y(g34120),.A(g33930),.B(g25158));
  AND4 AND4_181(.VSS(VSS),.VDD(VDD),.Y(I31342),.A(g32949),.B(g32950),.C(g32951),.D(g32952));
  AND2 AND2_2882(.VSS(VSS),.VDD(VDD),.Y(g32258),.A(g31624),.B(g30303));
  AND2 AND2_2883(.VSS(VSS),.VDD(VDD),.Y(g28117),.A(g8075),.B(g27245));
  AND2 AND2_2884(.VSS(VSS),.VDD(VDD),.Y(g18642),.A(g15097),.B(g17096));
  AND2 AND2_2885(.VSS(VSS),.VDD(VDD),.Y(g25059),.A(g20870),.B(g23460));
  AND2 AND2_2886(.VSS(VSS),.VDD(VDD),.Y(g33890),.A(g33310),.B(g20659));
  AND2 AND2_2887(.VSS(VSS),.VDD(VDD),.Y(g19788),.A(g9983),.B(g17216));
  AND4 AND4_182(.VSS(VSS),.VDD(VDD),.Y(I31031),.A(g30614),.B(g31801),.C(g32499),.D(g32500));
  AND2 AND2_2888(.VSS(VSS),.VDD(VDD),.Y(g16128),.A(g14333),.B(g14166));
  AND2 AND2_2889(.VSS(VSS),.VDD(VDD),.Y(g34146),.A(g33788),.B(g20091));
  AND2 AND2_2890(.VSS(VSS),.VDD(VDD),.Y(g34738),.A(g34660),.B(g33442));
  AND2 AND2_2891(.VSS(VSS),.VDD(VDD),.Y(g33249),.A(g32144),.B(g20026));
  AND2 AND2_2892(.VSS(VSS),.VDD(VDD),.Y(g34562),.A(g34369),.B(g17411));
  AND2 AND2_2893(.VSS(VSS),.VDD(VDD),.Y(g28569),.A(g27453),.B(g20433));
  AND2 AND2_2894(.VSS(VSS),.VDD(VDD),.Y(g21066),.A(g10043),.B(g17625));
  AND2 AND2_2895(.VSS(VSS),.VDD(VDD),.Y(g25058),.A(g23276),.B(g20513));
  AND2 AND2_2896(.VSS(VSS),.VDD(VDD),.Y(g16245),.A(g14278),.B(g14708));
  AND2 AND2_2897(.VSS(VSS),.VDD(VDD),.Y(g32043),.A(g31482),.B(g16173));
  AND3 AND3_170(.VSS(VSS),.VDD(VDD),.Y(g33482),.A(g32614),.B(I31106),.C(I31107));
  AND2 AND2_2898(.VSS(VSS),.VDD(VDD),.Y(g32244),.A(g31609),.B(g30297));
  AND2 AND2_2899(.VSS(VSS),.VDD(VDD),.Y(g31710),.A(g29814),.B(g19128));
  AND2 AND2_2900(.VSS(VSS),.VDD(VDD),.Y(g33248),.A(g32131),.B(g19996));
  AND2 AND2_2901(.VSS(VSS),.VDD(VDD),.Y(g10676),.A(g8506),.B(g3774));
  AND4 AND4_183(.VSS(VSS),.VDD(VDD),.Y(I27514),.A(g24091),.B(g24092),.C(g24093),.D(g24094));
  AND2 AND2_2902(.VSS(VSS),.VDD(VDD),.Y(g18733),.A(g15141),.B(g16877));
  AND2 AND2_2903(.VSS(VSS),.VDD(VDD),.Y(g27083),.A(g25819),.B(g22456));
  AND2 AND2_2904(.VSS(VSS),.VDD(VDD),.Y(g27348),.A(g26488),.B(g17392));
  AND2 AND2_2905(.VSS(VSS),.VDD(VDD),.Y(g33710),.A(g14037),.B(g33246));
  AND2 AND2_2906(.VSS(VSS),.VDD(VDD),.Y(g22130),.A(g6637),.B(g19277));
  AND2 AND2_2907(.VSS(VSS),.VDD(VDD),.Y(g27284),.A(g9908),.B(g26631));
  AND2 AND2_2908(.VSS(VSS),.VDD(VDD),.Y(g24864),.A(g11201),.B(g22305));
  AND2 AND2_2909(.VSS(VSS),.VDD(VDD),.Y(g22193),.A(g19880),.B(g20682));
  AND2 AND2_2910(.VSS(VSS),.VDD(VDD),.Y(g28242),.A(g27769),.B(g23626));
  AND2 AND2_2911(.VSS(VSS),.VDD(VDD),.Y(g21876),.A(g4119),.B(g19801));
  AND2 AND2_2912(.VSS(VSS),.VDD(VDD),.Y(g21885),.A(g4122),.B(g19801));
  AND2 AND2_2913(.VSS(VSS),.VDD(VDD),.Y(g26547),.A(g13283),.B(g25027));
  AND2 AND2_2914(.VSS(VSS),.VDD(VDD),.Y(g10654),.A(g3085),.B(g8434));
  AND2 AND2_2915(.VSS(VSS),.VDD(VDD),.Y(g11023),.A(g9669),.B(g5084));
  AND2 AND2_2916(.VSS(VSS),.VDD(VDD),.Y(g15857),.A(g3199),.B(g14038));
  AND2 AND2_2917(.VSS(VSS),.VDD(VDD),.Y(g23885),.A(g4132),.B(g19513));
  AND2 AND2_2918(.VSS(VSS),.VDD(VDD),.Y(g27304),.A(g2273),.B(g26682));
  AND2 AND2_2919(.VSS(VSS),.VDD(VDD),.Y(g24749),.A(g17511),.B(g22432));
  AND2 AND2_2920(.VSS(VSS),.VDD(VDD),.Y(g32069),.A(g10878),.B(g30735));
  AND2 AND2_2921(.VSS(VSS),.VDD(VDD),.Y(g12284),.A(g1532),.B(g7557));
  AND2 AND2_2922(.VSS(VSS),.VDD(VDD),.Y(g14654),.A(g7178),.B(g10476));
  AND2 AND2_2923(.VSS(VSS),.VDD(VDD),.Y(g24313),.A(g4504),.B(g22228));
  AND2 AND2_2924(.VSS(VSS),.VDD(VDD),.Y(g22165),.A(g15594),.B(g18903));
  AND2 AND2_2925(.VSS(VSS),.VDD(VDD),.Y(g18630),.A(g3689),.B(g17226));
  AND2 AND2_2926(.VSS(VSS),.VDD(VDD),.Y(g21854),.A(g3921),.B(g21070));
  AND2 AND2_2927(.VSS(VSS),.VDD(VDD),.Y(g15793),.A(g3219),.B(g13873));
  AND2 AND2_2928(.VSS(VSS),.VDD(VDD),.Y(g18693),.A(g4717),.B(g16053));
  AND2 AND2_2929(.VSS(VSS),.VDD(VDD),.Y(g23854),.A(g4093),.B(g19506));
  AND2 AND2_2930(.VSS(VSS),.VDD(VDD),.Y(g31778),.A(g21369),.B(g29385));
  AND2 AND2_2931(.VSS(VSS),.VDD(VDD),.Y(g24748),.A(g17656),.B(g22457));
  AND4 AND4_184(.VSS(VSS),.VDD(VDD),.Y(g26226),.A(g24688),.B(g8812),.C(g10658),.D(g10627));
  AND2 AND2_2932(.VSS(VSS),.VDD(VDD),.Y(g32068),.A(g31515),.B(g10862));
  AND2 AND2_2933(.VSS(VSS),.VDD(VDD),.Y(g33081),.A(g32388),.B(g18875));
  AND2 AND2_2934(.VSS(VSS),.VDD(VDD),.Y(g17193),.A(g2504),.B(g13023));
  AND2 AND2_2935(.VSS(VSS),.VDD(VDD),.Y(g21763),.A(g3223),.B(g20785));
  AND2 AND2_2936(.VSS(VSS),.VDD(VDD),.Y(g18166),.A(g655),.B(g17433));
  AND2 AND2_2937(.VSS(VSS),.VDD(VDD),.Y(g24285),.A(g4388),.B(g22550));
  AND2 AND2_2938(.VSS(VSS),.VDD(VDD),.Y(g25902),.A(g24398),.B(g19373));
  AND2 AND2_2939(.VSS(VSS),.VDD(VDD),.Y(g18665),.A(g4584),.B(g17367));
  AND4 AND4_185(.VSS(VSS),.VDD(VDD),.Y(I31132),.A(g32645),.B(g32646),.C(g32647),.D(g32648));
  AND2 AND2_2940(.VSS(VSS),.VDD(VDD),.Y(g31786),.A(g30189),.B(g24010));
  AND2 AND2_2941(.VSS(VSS),.VDD(VDD),.Y(g25957),.A(g17190),.B(g24960));
  AND2 AND2_2942(.VSS(VSS),.VDD(VDD),.Y(g24704),.A(g17593),.B(g22384));
  AND3 AND3_171(.VSS(VSS),.VDD(VDD),.Y(g25377),.A(g5712),.B(g22210),.C(I24530));
  AND2 AND2_2943(.VSS(VSS),.VDD(VDD),.Y(g33786),.A(g33130),.B(g20572));
  AND2 AND2_2944(.VSS(VSS),.VDD(VDD),.Y(g24305),.A(g4477),.B(g22228));
  AND2 AND2_2945(.VSS(VSS),.VDD(VDD),.Y(g16737),.A(g6645),.B(g15042));
  AND2 AND2_2946(.VSS(VSS),.VDD(VDD),.Y(g26572),.A(g7443),.B(g24439));
  AND2 AND2_2947(.VSS(VSS),.VDD(VDD),.Y(g22006),.A(g5767),.B(g21562));
  AND2 AND2_2948(.VSS(VSS),.VDD(VDD),.Y(g28639),.A(g27767),.B(g20597));
  AND3 AND3_172(.VSS(VSS),.VDD(VDD),.Y(g24900),.A(g3752),.B(g23582),.C(I24067));
  AND2 AND2_2949(.VSS(VSS),.VDD(VDD),.Y(g33647),.A(g33390),.B(g18878));
  AND2 AND2_2950(.VSS(VSS),.VDD(VDD),.Y(g32337),.A(g31465),.B(g20663));
  AND2 AND2_2951(.VSS(VSS),.VDD(VDD),.Y(g27139),.A(g26055),.B(g16608));
  AND3 AND3_173(.VSS(VSS),.VDD(VDD),.Y(g28293),.A(g7424),.B(g2495),.C(g27474));
  AND2 AND2_2952(.VSS(VSS),.VDD(VDD),.Y(g33356),.A(g32245),.B(g20772));
  AND2 AND2_2953(.VSS(VSS),.VDD(VDD),.Y(g22863),.A(g9547),.B(g20388));
  AND2 AND2_2954(.VSS(VSS),.VDD(VDD),.Y(g27653),.A(g26549),.B(g15562));
  AND2 AND2_2955(.VSS(VSS),.VDD(VDD),.Y(g28638),.A(g27551),.B(g20583));
  AND2 AND2_2956(.VSS(VSS),.VDD(VDD),.Y(g32171),.A(g31706),.B(g27800));
  AND4 AND4_186(.VSS(VSS),.VDD(VDD),.Y(I31161),.A(g30614),.B(g31824),.C(g32687),.D(g32688));
  AND2 AND2_2957(.VSS(VSS),.VDD(VDD),.Y(g18476),.A(g2433),.B(g15426));
  AND2 AND2_2958(.VSS(VSS),.VDD(VDD),.Y(g18485),.A(g2465),.B(g15426));
  AND2 AND2_2959(.VSS(VSS),.VDD(VDD),.Y(g29787),.A(g28334),.B(g23249));
  AND2 AND2_2960(.VSS(VSS),.VDD(VDD),.Y(g26127),.A(g2236),.B(g25119));
  AND2 AND2_2961(.VSS(VSS),.VDD(VDD),.Y(g27138),.A(g26055),.B(g16607));
  AND2 AND2_2962(.VSS(VSS),.VDD(VDD),.Y(g28265),.A(g11367),.B(g27989));
  AND2 AND2_2963(.VSS(VSS),.VDD(VDD),.Y(g34661),.A(g34575),.B(g18907));
  AND2 AND2_2964(.VSS(VSS),.VDD(VDD),.Y(g18555),.A(g2834),.B(g15277));
  AND2 AND2_2965(.VSS(VSS),.VDD(VDD),.Y(g18454),.A(g2303),.B(g15224));
  AND3 AND3_174(.VSS(VSS),.VDD(VDD),.Y(g25290),.A(g5022),.B(g22173),.C(I24482));
  AND2 AND2_2966(.VSS(VSS),.VDD(VDD),.Y(g14216),.A(g7631),.B(g10608));
  AND2 AND2_2967(.VSS(VSS),.VDD(VDD),.Y(g21916),.A(g5084),.B(g21468));
  AND2 AND2_2968(.VSS(VSS),.VDD(VDD),.Y(g30226),.A(g28707),.B(g23898));
  AND2 AND2_2969(.VSS(VSS),.VDD(VDD),.Y(g18570),.A(g2848),.B(g16349));
  AND2 AND2_2970(.VSS(VSS),.VDD(VDD),.Y(g18712),.A(g4843),.B(g15915));
  AND2 AND2_2971(.VSS(VSS),.VDD(VDD),.Y(g33233),.A(g32094),.B(g23005));
  AND2 AND2_2972(.VSS(VSS),.VDD(VDD),.Y(g31182),.A(g30240),.B(g20682));
  AND2 AND2_2973(.VSS(VSS),.VDD(VDD),.Y(g31672),.A(g29814),.B(g19050));
  AND2 AND2_2974(.VSS(VSS),.VDD(VDD),.Y(g27333),.A(g10180),.B(g26765));
  AND2 AND2_2975(.VSS(VSS),.VDD(VDD),.Y(g24642),.A(g8290),.B(g22898));
  AND2 AND2_2976(.VSS(VSS),.VDD(VDD),.Y(g34226),.A(g33914),.B(g21467));
  AND2 AND2_2977(.VSS(VSS),.VDD(VDD),.Y(g14587),.A(g10584),.B(g10567));
  AND2 AND2_2978(.VSS(VSS),.VDD(VDD),.Y(g29743),.A(g28206),.B(g10233));
  AND4 AND4_187(.VSS(VSS),.VDD(VDD),.Y(I31087),.A(g32580),.B(g32581),.C(g32582),.D(g32583));
  AND2 AND2_2979(.VSS(VSS),.VDD(VDD),.Y(g34715),.A(g34570),.B(g33375));
  AND2 AND2_2980(.VSS(VSS),.VDD(VDD),.Y(g34481),.A(g34404),.B(g18916));
  AND2 AND2_2981(.VSS(VSS),.VDD(VDD),.Y(g23314),.A(g9104),.B(g19200));
  AND2 AND2_2982(.VSS(VSS),.VDD(VDD),.Y(g32425),.A(g31668),.B(g21604));
  AND2 AND2_2983(.VSS(VSS),.VDD(VDD),.Y(g26103),.A(g2185),.B(g25100));
  AND2 AND2_2984(.VSS(VSS),.VDD(VDD),.Y(g34572),.A(g34387),.B(g33326));
  AND2 AND2_2985(.VSS(VSS),.VDD(VDD),.Y(g10543),.A(g8238),.B(g437));
  AND2 AND2_2986(.VSS(VSS),.VDD(VDD),.Y(g26095),.A(g11923),.B(g25090));
  AND2 AND2_2987(.VSS(VSS),.VDD(VDD),.Y(g27963),.A(g25952),.B(g16047));
  AND2 AND2_2988(.VSS(VSS),.VDD(VDD),.Y(g23076),.A(g19128),.B(g9104));
  AND2 AND2_2989(.VSS(VSS),.VDD(VDD),.Y(g29640),.A(g28498),.B(g8125));
  AND2 AND2_2990(.VSS(VSS),.VDD(VDD),.Y(g25366),.A(g7733),.B(g22406));
  AND2 AND2_2991(.VSS(VSS),.VDD(VDD),.Y(g29769),.A(g28319),.B(g23237));
  AND2 AND2_2992(.VSS(VSS),.VDD(VDD),.Y(g18239),.A(g1135),.B(g16326));
  AND2 AND2_2993(.VSS(VSS),.VDD(VDD),.Y(g21721),.A(g385),.B(g21037));
  AND2 AND2_2994(.VSS(VSS),.VDD(VDD),.Y(g33331),.A(g32216),.B(g20607));
  AND2 AND2_2995(.VSS(VSS),.VDD(VDD),.Y(g27664),.A(g1024),.B(g25911));
  AND2 AND2_2996(.VSS(VSS),.VDD(VDD),.Y(g18567),.A(g2894),.B(g16349));
  AND2 AND2_2997(.VSS(VSS),.VDD(VDD),.Y(g18594),.A(g12858),.B(g16349));
  AND2 AND2_2998(.VSS(VSS),.VDD(VDD),.Y(g31513),.A(g2606),.B(g29318));
  AND2 AND2_2999(.VSS(VSS),.VDD(VDD),.Y(g32010),.A(g31785),.B(g22303));
  AND3 AND3_175(.VSS(VSS),.VDD(VDD),.Y(g33513),.A(g32837),.B(I31261),.C(I31262));
  AND2 AND2_3000(.VSS(VSS),.VDD(VDD),.Y(g29803),.A(g28414),.B(g26836));
  AND2 AND2_3001(.VSS(VSS),.VDD(VDD),.Y(g18238),.A(g1152),.B(g16326));
  AND2 AND2_3002(.VSS(VSS),.VDD(VDD),.Y(g26181),.A(g2652),.B(g25157));
  AND2 AND2_3003(.VSS(VSS),.VDD(VDD),.Y(g26671),.A(g316),.B(g24429));
  AND2 AND2_3004(.VSS(VSS),.VDD(VDD),.Y(g28586),.A(g27484),.B(g20497));
  AND2 AND2_3005(.VSS(VSS),.VDD(VDD),.Y(g24630),.A(g23255),.B(g14149));
  AND2 AND2_3006(.VSS(VSS),.VDD(VDD),.Y(g31961),.A(g31751),.B(g22154));
  AND2 AND2_3007(.VSS(VSS),.VDD(VDD),.Y(g33897),.A(g33315),.B(g20777));
  AND4 AND4_188(.VSS(VSS),.VDD(VDD),.Y(g17781),.A(g6772),.B(g11592),.C(g6789),.D(I18785));
  AND2 AND2_3008(.VSS(VSS),.VDD(VDD),.Y(g31505),.A(g30195),.B(g24379));
  AND2 AND2_3009(.VSS(VSS),.VDD(VDD),.Y(g28442),.A(g27278),.B(g20072));
  AND3 AND3_176(.VSS(VSS),.VDD(VDD),.Y(g33505),.A(g32779),.B(I31221),.C(I31222));
  AND2 AND2_3010(.VSS(VSS),.VDD(VDD),.Y(g18382),.A(g1936),.B(g15171));
  AND2 AND2_3011(.VSS(VSS),.VDD(VDD),.Y(g24009),.A(g19671),.B(g10971));
  AND2 AND2_3012(.VSS(VSS),.VDD(VDD),.Y(g33404),.A(g32353),.B(g21397));
  AND2 AND2_3013(.VSS(VSS),.VDD(VDD),.Y(g29881),.A(g2040),.B(g29150));
  AND2 AND2_3014(.VSS(VSS),.VDD(VDD),.Y(g21773),.A(g3263),.B(g20785));
  AND2 AND2_3015(.VSS(VSS),.VDD(VDD),.Y(g18519),.A(g2648),.B(g15509));
  AND2 AND2_3016(.VSS(VSS),.VDD(VDD),.Y(g11016),.A(g4888),.B(g8984));
  AND2 AND2_3017(.VSS(VSS),.VDD(VDD),.Y(g21942),.A(g5236),.B(g18997));
  AND2 AND2_3018(.VSS(VSS),.VDD(VDD),.Y(g13525),.A(g10019),.B(g11911));
  AND2 AND2_3019(.VSS(VSS),.VDD(VDD),.Y(g18176),.A(g732),.B(g17328));
  AND2 AND2_3020(.VSS(VSS),.VDD(VDD),.Y(g18185),.A(g790),.B(g17328));
  AND2 AND2_3021(.VSS(VSS),.VDD(VDD),.Y(g22063),.A(g6109),.B(g21611));
  AND2 AND2_3022(.VSS(VSS),.VDD(VDD),.Y(g18675),.A(g4349),.B(g15758));
  AND2 AND2_3023(.VSS(VSS),.VDD(VDD),.Y(g34385),.A(g34168),.B(g20642));
  AND2 AND2_3024(.VSS(VSS),.VDD(VDD),.Y(g33717),.A(g14092),.B(g33306));
  AND2 AND2_3025(.VSS(VSS),.VDD(VDD),.Y(g24008),.A(g7909),.B(g19502));
  AND2 AND2_3026(.VSS(VSS),.VDD(VDD),.Y(g32086),.A(g7597),.B(g30735));
  AND2 AND2_3027(.VSS(VSS),.VDD(VDD),.Y(g30095),.A(g28545),.B(g20768));
  AND2 AND2_3028(.VSS(VSS),.VDD(VDD),.Y(g31212),.A(g20028),.B(g29669));
  AND2 AND2_3029(.VSS(VSS),.VDD(VDD),.Y(g28116),.A(g27366),.B(g26183));
  AND2 AND2_3030(.VSS(VSS),.VDD(VDD),.Y(g18518),.A(g2657),.B(g15509));
  AND2 AND2_3031(.VSS(VSS),.VDD(VDD),.Y(g18154),.A(g622),.B(g17533));
  AND2 AND2_3032(.VSS(VSS),.VDD(VDD),.Y(g27312),.A(g12019),.B(g26700));
  AND2 AND2_3033(.VSS(VSS),.VDD(VDD),.Y(g24892),.A(g11559),.B(g23264));
  AND4 AND4_189(.VSS(VSS),.VDD(VDD),.Y(g26190),.A(g25357),.B(g11724),.C(g7586),.D(g11686));
  AND2 AND2_3034(.VSS(VSS),.VDD(VDD),.Y(g24485),.A(g10710),.B(g22319));
  AND2 AND2_3035(.VSS(VSS),.VDD(VDD),.Y(g24476),.A(g18879),.B(g22330));
  AND4 AND4_190(.VSS(VSS),.VDD(VDD),.Y(I31337),.A(g32942),.B(g32943),.C(g32944),.D(g32945));
  AND2 AND2_3036(.VSS(VSS),.VDD(VDD),.Y(g16611),.A(g5583),.B(g14727));
  AND2 AND2_3037(.VSS(VSS),.VDD(VDD),.Y(g27115),.A(g26026),.B(g16526));
  AND2 AND2_3038(.VSS(VSS),.VDD(VDD),.Y(g11893),.A(g1668),.B(g7268));
  AND4 AND4_191(.VSS(VSS),.VDD(VDD),.Y(g13830),.A(g11543),.B(g11424),.C(g11395),.D(I16143));
  AND2 AND2_3039(.VSS(VSS),.VDD(VDD),.Y(g22873),.A(g19854),.B(g19683));
  AND2 AND2_3040(.VSS(VSS),.VDD(VDD),.Y(g25551),.A(g23822),.B(g21511));
  AND2 AND2_3041(.VSS(VSS),.VDD(VDD),.Y(g18637),.A(g3821),.B(g17096));
  AND2 AND2_3042(.VSS(VSS),.VDD(VDD),.Y(g25572),.A(I24699),.B(I24700));
  AND4 AND4_192(.VSS(VSS),.VDD(VDD),.Y(I31171),.A(g31528),.B(g31826),.C(g32701),.D(g32702));
  AND2 AND2_3043(.VSS(VSS),.VDD(VDD),.Y(g30181),.A(g28636),.B(g23821));
  AND2 AND2_3044(.VSS(VSS),.VDD(VDD),.Y(g30671),.A(g29319),.B(g22317));
  AND2 AND2_3045(.VSS(VSS),.VDD(VDD),.Y(g18935),.A(g4322),.B(g15574));
  AND2 AND2_3046(.VSS(VSS),.VDD(VDD),.Y(g32322),.A(g31308),.B(g20605));
  AND2 AND2_3047(.VSS(VSS),.VDD(VDD),.Y(g24555),.A(g23184),.B(g21024));
  AND2 AND2_3048(.VSS(VSS),.VDD(VDD),.Y(g29662),.A(g1848),.B(g29049));
  AND2 AND2_3049(.VSS(VSS),.VDD(VDD),.Y(g9217),.A(g632),.B(g626));
  AND2 AND2_3050(.VSS(VSS),.VDD(VDD),.Y(g21734),.A(g3040),.B(g20330));
  AND2 AND2_3051(.VSS(VSS),.VDD(VDD),.Y(g32159),.A(g31658),.B(g30040));
  AND2 AND2_3052(.VSS(VSS),.VDD(VDD),.Y(g24712),.A(g19592),.B(g23001));
  AND2 AND2_3053(.VSS(VSS),.VDD(VDD),.Y(g29890),.A(g28419),.B(g23355));
  AND2 AND2_3054(.VSS(VSS),.VDD(VDD),.Y(g24914),.A(g8721),.B(g23301));
  AND2 AND2_3055(.VSS(VSS),.VDD(VDD),.Y(g21839),.A(g3763),.B(g20453));
  AND2 AND2_3056(.VSS(VSS),.VDD(VDD),.Y(g21930),.A(g5180),.B(g18997));
  AND2 AND2_3057(.VSS(VSS),.VDD(VDD),.Y(g25127),.A(g13997),.B(g23524));
  AND2 AND2_3058(.VSS(VSS),.VDD(VDD),.Y(g21993),.A(g5603),.B(g19074));
  AND2 AND2_3059(.VSS(VSS),.VDD(VDD),.Y(g32158),.A(g31658),.B(g30022));
  AND2 AND2_3060(.VSS(VSS),.VDD(VDD),.Y(g22209),.A(g19907),.B(g20751));
  AND2 AND2_3061(.VSS(VSS),.VDD(VDD),.Y(g15856),.A(g9056),.B(g14223));
  AND3 AND3_177(.VSS(VSS),.VDD(VDD),.Y(g15995),.A(g13314),.B(g1157),.C(g10666));
  AND2 AND2_3062(.VSS(VSS),.VDD(VDD),.Y(g33723),.A(g14091),.B(g33299));
  AND2 AND2_3063(.VSS(VSS),.VDD(VDD),.Y(g28237),.A(g9492),.B(g27597));
  AND2 AND2_3064(.VSS(VSS),.VDD(VDD),.Y(g21838),.A(g3747),.B(g20453));
  AND2 AND2_3065(.VSS(VSS),.VDD(VDD),.Y(g22834),.A(g102),.B(g19630));
  AND2 AND2_3066(.VSS(VSS),.VDD(VDD),.Y(g15880),.A(g3211),.B(g13980));
  AND2 AND2_3067(.VSS(VSS),.VDD(VDD),.Y(g31149),.A(g29508),.B(g23021));
  AND2 AND2_3068(.VSS(VSS),.VDD(VDD),.Y(g21965),.A(g15149),.B(g21514));
  AND2 AND2_3069(.VSS(VSS),.VDD(VDD),.Y(g26088),.A(g6545),.B(g25080));
  AND2 AND2_3070(.VSS(VSS),.VDD(VDD),.Y(g26024),.A(g2619),.B(g25039));
  AND2 AND2_3071(.VSS(VSS),.VDD(VDD),.Y(g22208),.A(g19906),.B(g20739));
  AND2 AND2_3072(.VSS(VSS),.VDD(VDD),.Y(g29710),.A(g2380),.B(g29094));
  AND3 AND3_178(.VSS(VSS),.VDD(VDD),.Y(g28035),.A(g24103),.B(I26530),.C(I26531));
  AND2 AND2_3073(.VSS(VSS),.VDD(VDD),.Y(g29552),.A(g2223),.B(g28579));
  AND2 AND2_3074(.VSS(VSS),.VDD(VDD),.Y(g33433),.A(g32238),.B(g29694));
  AND2 AND2_3075(.VSS(VSS),.VDD(VDD),.Y(g23131),.A(g13919),.B(g19930));
  AND2 AND2_3076(.VSS(VSS),.VDD(VDD),.Y(g32295),.A(g27931),.B(g31376));
  AND2 AND2_3077(.VSS(VSS),.VDD(VDD),.Y(g10841),.A(g8509),.B(g8567));
  AND3 AND3_179(.VSS(VSS),.VDD(VDD),.Y(g29204),.A(g24110),.B(I27518),.C(I27519));
  AND2 AND2_3078(.VSS(VSS),.VDD(VDD),.Y(g31148),.A(g2661),.B(g30055));
  AND2 AND2_3079(.VSS(VSS),.VDD(VDD),.Y(g30190),.A(g28646),.B(g23842));
  AND2 AND2_3080(.VSS(VSS),.VDD(VDD),.Y(g13042),.A(g433),.B(g11048));
  AND2 AND2_3081(.VSS(VSS),.VDD(VDD),.Y(g16199),.A(g3614),.B(g14051));
  AND2 AND2_3082(.VSS(VSS),.VDD(VDD),.Y(g18215),.A(g943),.B(g15979));
  AND2 AND2_3083(.VSS(VSS),.VDD(VDD),.Y(g25103),.A(g4927),.B(g22908));
  AND2 AND2_3084(.VSS(VSS),.VDD(VDD),.Y(g27184),.A(g26628),.B(g13756));
  AND2 AND2_3085(.VSS(VSS),.VDD(VDD),.Y(g16736),.A(g6303),.B(g15036));
  AND2 AND2_3086(.VSS(VSS),.VDD(VDD),.Y(g18501),.A(g12854),.B(g15509));
  AND2 AND2_3087(.VSS(VSS),.VDD(VDD),.Y(g18729),.A(g15139),.B(g16821));
  AND2 AND2_3088(.VSS(VSS),.VDD(VDD),.Y(g22021),.A(g5869),.B(g19147));
  AND2 AND2_3089(.VSS(VSS),.VDD(VDD),.Y(g27674),.A(g26873),.B(g23543));
  AND2 AND2_3090(.VSS(VSS),.VDD(VDD),.Y(g25980),.A(g1926),.B(g25006));
  AND2 AND2_3091(.VSS(VSS),.VDD(VDD),.Y(g18577),.A(g2988),.B(g16349));
  AND2 AND2_3092(.VSS(VSS),.VDD(VDD),.Y(g33104),.A(g26296),.B(g32137));
  AND2 AND2_3093(.VSS(VSS),.VDD(VDD),.Y(g25095),.A(g23319),.B(g20556));
  AND2 AND2_3094(.VSS(VSS),.VDD(VDD),.Y(g33811),.A(g33439),.B(g17573));
  AND2 AND2_3095(.VSS(VSS),.VDD(VDD),.Y(g33646),.A(g33389),.B(g18876));
  AND2 AND2_3096(.VSS(VSS),.VDD(VDD),.Y(g19767),.A(g16810),.B(g14203));
  AND2 AND2_3097(.VSS(VSS),.VDD(VDD),.Y(g32336),.A(g31596),.B(g11842));
  AND2 AND2_3098(.VSS(VSS),.VDD(VDD),.Y(g34520),.A(g34294),.B(g19505));
  AND2 AND2_3099(.VSS(VSS),.VDD(VDD),.Y(g23619),.A(g19453),.B(g13045));
  AND2 AND2_3100(.VSS(VSS),.VDD(VDD),.Y(g33343),.A(g32227),.B(g20665));
  AND2 AND2_3101(.VSS(VSS),.VDD(VDD),.Y(g21557),.A(g12980),.B(g15674));
  AND2 AND2_3102(.VSS(VSS),.VDD(VDD),.Y(g18728),.A(g4939),.B(g16821));
  AND2 AND2_3103(.VSS(VSS),.VDD(VDD),.Y(g18439),.A(g2250),.B(g18008));
  AND2 AND2_3104(.VSS(VSS),.VDD(VDD),.Y(g30089),.A(g28538),.B(g20709));
  AND2 AND2_3105(.VSS(VSS),.VDD(VDD),.Y(g24941),.A(g23171),.B(g20190));
  AND2 AND2_3106(.VSS(VSS),.VDD(VDD),.Y(g26126),.A(g1959),.B(g25118));
  AND2 AND2_3107(.VSS(VSS),.VDD(VDD),.Y(g30211),.A(g28685),.B(g23878));
  AND2 AND2_3108(.VSS(VSS),.VDD(VDD),.Y(g11939),.A(g2361),.B(g7380));
  AND2 AND2_3109(.VSS(VSS),.VDD(VDD),.Y(g23618),.A(g19388),.B(g11917));
  AND2 AND2_3110(.VSS(VSS),.VDD(VDD),.Y(g25181),.A(g23405),.B(g20696));
  AND3 AND3_180(.VSS(VSS),.VDD(VDD),.Y(g34089),.A(g22957),.B(g9104),.C(g33744));
  AND2 AND2_3111(.VSS(VSS),.VDD(VDD),.Y(g16843),.A(g6251),.B(g14864));
  AND2 AND2_3112(.VSS(VSS),.VDD(VDD),.Y(g18438),.A(g2236),.B(g18008));
  AND2 AND2_3113(.VSS(VSS),.VDD(VDD),.Y(g34211),.A(g33891),.B(g21349));
  AND2 AND2_3114(.VSS(VSS),.VDD(VDD),.Y(g26250),.A(g1902),.B(g25429));
  AND2 AND2_3115(.VSS(VSS),.VDD(VDD),.Y(g13383),.A(g4765),.B(g11797));
  AND2 AND2_3116(.VSS(VSS),.VDD(VDD),.Y(g24675),.A(g17568),.B(g22342));
  AND2 AND2_3117(.VSS(VSS),.VDD(VDD),.Y(g29647),.A(g28934),.B(g22457));
  AND2 AND2_3118(.VSS(VSS),.VDD(VDD),.Y(g30024),.A(g28497),.B(g23501));
  AND2 AND2_3119(.VSS(VSS),.VDD(VDD),.Y(g33369),.A(g32277),.B(g21060));
  AND3 AND3_181(.VSS(VSS),.VDD(VDD),.Y(I24048),.A(g3034),.B(g3040),.C(g8426));
  AND2 AND2_3120(.VSS(VSS),.VDD(VDD),.Y(g17726),.A(g1467),.B(g13315));
  AND2 AND2_3121(.VSS(VSS),.VDD(VDD),.Y(g16764),.A(g6307),.B(g14776));
  AND3 AND3_182(.VSS(VSS),.VDD(VDD),.Y(g34088),.A(g33736),.B(g9104),.C(g18957));
  AND2 AND2_3122(.VSS(VSS),.VDD(VDD),.Y(g13030),.A(g429),.B(g11048));
  AND2 AND2_3123(.VSS(VSS),.VDD(VDD),.Y(g22073),.A(g6235),.B(g19210));
  AND2 AND2_3124(.VSS(VSS),.VDD(VDD),.Y(g18349),.A(g1768),.B(g17955));
  AND2 AND2_3125(.VSS(VSS),.VDD(VDD),.Y(g14586),.A(g11953),.B(g11970));
  AND2 AND2_3126(.VSS(VSS),.VDD(VDD),.Y(g13294),.A(g1564),.B(g11513));
  AND4 AND4_193(.VSS(VSS),.VDD(VDD),.Y(I31086),.A(g31554),.B(g31811),.C(g32578),.D(g32579));
  AND2 AND2_3127(.VSS(VSS),.VDD(VDD),.Y(g29380),.A(g28134),.B(g19396));
  AND2 AND2_3128(.VSS(VSS),.VDD(VDD),.Y(g33368),.A(g32275),.B(g21057));
  AND2 AND2_3129(.VSS(VSS),.VDD(VDD),.Y(g34860),.A(g16540),.B(g34823));
  AND2 AND2_3130(.VSS(VSS),.VDD(VDD),.Y(g16869),.A(g6259),.B(g14902));
  AND2 AND2_3131(.VSS(VSS),.VDD(VDD),.Y(g27692),.A(g26392),.B(g20697));
  AND2 AND2_3132(.VSS(VSS),.VDD(VDD),.Y(g28130),.A(g27353),.B(g23063));
  AND2 AND2_3133(.VSS(VSS),.VDD(VDD),.Y(g28193),.A(g8851),.B(g27629));
  AND2 AND2_3134(.VSS(VSS),.VDD(VDD),.Y(g26339),.A(g225),.B(g24836));
  AND2 AND2_3135(.VSS(VSS),.VDD(VDD),.Y(g25931),.A(g24574),.B(g19477));
  AND2 AND2_3136(.VSS(VSS),.VDD(VDD),.Y(g18906),.A(g13568),.B(g16264));
  AND2 AND2_3137(.VSS(VSS),.VDD(VDD),.Y(g18348),.A(g1744),.B(g17955));
  AND2 AND2_3138(.VSS(VSS),.VDD(VDD),.Y(g24637),.A(g16586),.B(g22884));
  AND2 AND2_3139(.VSS(VSS),.VDD(VDD),.Y(g19521),.A(g513),.B(g16739));
  AND2 AND2_3140(.VSS(VSS),.VDD(VDD),.Y(g22122),.A(g6601),.B(g19277));
  AND3 AND3_183(.VSS(VSS),.VDD(VDD),.Y(g12692),.A(g10323),.B(g3522),.C(g3530));
  AND2 AND2_3141(.VSS(VSS),.VDD(VDD),.Y(g12761),.A(g969),.B(g7567));
  AND2 AND2_3142(.VSS(VSS),.VDD(VDD),.Y(g18284),.A(g15071),.B(g16164));
  AND2 AND2_3143(.VSS(VSS),.VDD(VDD),.Y(g16868),.A(g5813),.B(g14297));
  AND2 AND2_3144(.VSS(VSS),.VDD(VDD),.Y(g34497),.A(g34275),.B(g33072));
  AND2 AND2_3145(.VSS(VSS),.VDD(VDD),.Y(g28165),.A(g27018),.B(g22455));
  AND2 AND2_3146(.VSS(VSS),.VDD(VDD),.Y(g28523),.A(g27704),.B(g15585));
  AND2 AND2_3147(.VSS(VSS),.VDD(VDD),.Y(g18304),.A(g1542),.B(g16489));
  AND2 AND2_3148(.VSS(VSS),.VDD(VDD),.Y(g29182),.A(g27163),.B(g12730));
  AND2 AND2_3149(.VSS(VSS),.VDD(VDD),.Y(g29651),.A(g2537),.B(g29134));
  AND2 AND2_3150(.VSS(VSS),.VDD(VDD),.Y(g33412),.A(g32362),.B(g21411));
  AND4 AND4_194(.VSS(VSS),.VDD(VDD),.Y(I31322),.A(g32921),.B(g32922),.C(g32923),.D(g32924));
  AND2 AND2_3151(.VSS(VSS),.VDD(VDD),.Y(g16161),.A(g5841),.B(g14297));
  AND2 AND2_3152(.VSS(VSS),.VDD(VDD),.Y(g15611),.A(g471),.B(g13437));
  AND2 AND2_3153(.VSS(VSS),.VDD(VDD),.Y(g15722),.A(g464),.B(g13437));
  AND2 AND2_3154(.VSS(VSS),.VDD(VDD),.Y(g18622),.A(g3480),.B(g17062));
  AND2 AND2_3155(.VSS(VSS),.VDD(VDD),.Y(g22034),.A(g5929),.B(g19147));
  AND2 AND2_3156(.VSS(VSS),.VDD(VDD),.Y(g15080),.A(g12855),.B(g12983));
  AND2 AND2_3157(.VSS(VSS),.VDD(VDD),.Y(g18566),.A(g2860),.B(g16349));
  AND2 AND2_3158(.VSS(VSS),.VDD(VDD),.Y(g30126),.A(g28582),.B(g21058));
  AND2 AND2_3159(.VSS(VSS),.VDD(VDD),.Y(g14615),.A(g10604),.B(g10587));
  AND2 AND2_3160(.VSS(VSS),.VDD(VDD),.Y(g27214),.A(g26026),.B(g13901));
  AND2 AND2_3161(.VSS(VSS),.VDD(VDD),.Y(g34700),.A(g34535),.B(g20129));
  AND2 AND2_3162(.VSS(VSS),.VDD(VDD),.Y(g31229),.A(g30288),.B(g23949));
  AND3 AND3_184(.VSS(VSS),.VDD(VDD),.Y(g10720),.A(g2704),.B(g10219),.C(g2689));
  AND2 AND2_3163(.VSS(VSS),.VDD(VDD),.Y(g21815),.A(g3598),.B(g20924));
  AND2 AND2_3164(.VSS(VSS),.VDD(VDD),.Y(g30250),.A(g28744),.B(g23939));
  AND2 AND2_3165(.VSS(VSS),.VDD(VDD),.Y(g27329),.A(g12052),.B(g26743));
  AND2 AND2_3166(.VSS(VSS),.VDD(VDD),.Y(g32309),.A(g5160),.B(g31528));
  AND2 AND2_3167(.VSS(VSS),.VDD(VDD),.Y(g27207),.A(g26055),.B(g16692));
  AND2 AND2_3168(.VSS(VSS),.VDD(VDD),.Y(g33896),.A(g33314),.B(g20771));
  AND2 AND2_3169(.VSS(VSS),.VDD(VDD),.Y(g31228),.A(g20028),.B(g29713));
  AND2 AND2_3170(.VSS(VSS),.VDD(VDD),.Y(g27539),.A(g26576),.B(g17745));
  AND2 AND2_3171(.VSS(VSS),.VDD(VDD),.Y(g29331),.A(g29143),.B(g22169));
  AND2 AND2_3172(.VSS(VSS),.VDD(VDD),.Y(g32224),.A(g4300),.B(g31327));
  AND2 AND2_3173(.VSS(VSS),.VDD(VDD),.Y(g34658),.A(g34574),.B(g18896));
  AND2 AND2_3174(.VSS(VSS),.VDD(VDD),.Y(g23187),.A(g13989),.B(g20010));
  AND2 AND2_3175(.VSS(VSS),.VDD(VDD),.Y(g26855),.A(g2960),.B(g24535));
  AND2 AND2_3176(.VSS(VSS),.VDD(VDD),.Y(g21975),.A(g5523),.B(g19074));
  AND2 AND2_3177(.VSS(VSS),.VDD(VDD),.Y(g27328),.A(g12482),.B(g26736));
  AND2 AND2_3178(.VSS(VSS),.VDD(VDD),.Y(g25089),.A(g23317),.B(g20553));
  AND2 AND2_3179(.VSS(VSS),.VDD(VDD),.Y(g32308),.A(g31293),.B(g23503));
  AND2 AND2_3180(.VSS(VSS),.VDD(VDD),.Y(g20215),.A(g16479),.B(g10476));
  AND2 AND2_3181(.VSS(VSS),.VDD(VDD),.Y(g29513),.A(g28448),.B(g14095));
  AND2 AND2_3182(.VSS(VSS),.VDD(VDD),.Y(g18139),.A(g542),.B(g17249));
  AND2 AND2_3183(.VSS(VSS),.VDD(VDD),.Y(g27538),.A(g26549),.B(g14744));
  AND2 AND2_3184(.VSS(VSS),.VDD(VDD),.Y(g18653),.A(g4176),.B(g16249));
  AND2 AND2_3185(.VSS(VSS),.VDD(VDD),.Y(g24501),.A(g14000),.B(g23182));
  AND2 AND2_3186(.VSS(VSS),.VDD(VDD),.Y(g24729),.A(g22719),.B(g23018));
  AND2 AND2_3187(.VSS(VSS),.VDD(VDD),.Y(g25088),.A(g17601),.B(g23491));
  AND2 AND2_3188(.VSS(VSS),.VDD(VDD),.Y(g17292),.A(g1075),.B(g13093));
  AND4 AND4_195(.VSS(VSS),.VDD(VDD),.Y(g11160),.A(g6336),.B(g7074),.C(g6322),.D(g10003));
  AND2 AND2_3189(.VSS(VSS),.VDD(VDD),.Y(g17153),.A(g6311),.B(g14943));
  AND3 AND3_185(.VSS(VSS),.VDD(VDD),.Y(I24033),.A(g8219),.B(g8443),.C(g3747));
  AND2 AND2_3190(.VSS(VSS),.VDD(VDD),.Y(g18138),.A(g546),.B(g17249));
  AND4 AND4_196(.VSS(VSS),.VDD(VDD),.Y(I26531),.A(g24099),.B(g24100),.C(g24101),.D(g24102));
  AND2 AND2_3191(.VSS(VSS),.VDD(VDD),.Y(g21937),.A(g5208),.B(g18997));
  AND3 AND3_186(.VSS(VSS),.VDD(VDD),.Y(I17552),.A(g13156),.B(g11450),.C(g11498));
  AND2 AND2_3192(.VSS(VSS),.VDD(VDD),.Y(g34338),.A(g34099),.B(g19905));
  AND2 AND2_3193(.VSS(VSS),.VDD(VDD),.Y(g24728),.A(g16513),.B(g23017));
  AND4 AND4_197(.VSS(VSS),.VDD(VDD),.Y(g16244),.A(g11547),.B(g11592),.C(g6789),.D(I17585));
  AND4 AND4_198(.VSS(VSS),.VDD(VDD),.Y(I31336),.A(g31672),.B(g31855),.C(g32940),.D(g32941));
  AND2 AND2_3194(.VSS(VSS),.VDD(VDD),.Y(g14035),.A(g699),.B(g11048));
  AND2 AND2_3195(.VSS(VSS),.VDD(VDD),.Y(g15650),.A(g8362),.B(g13413));
  AND2 AND2_3196(.VSS(VSS),.VDD(VDD),.Y(g34969),.A(g34960),.B(g19570));
  AND2 AND2_3197(.VSS(VSS),.VDD(VDD),.Y(g10684),.A(g7998),.B(g411));
  AND2 AND2_3198(.VSS(VSS),.VDD(VDD),.Y(g28703),.A(g27925),.B(g20680));
  AND2 AND2_3199(.VSS(VSS),.VDD(VDD),.Y(g18636),.A(g3817),.B(g17096));
  AND2 AND2_3200(.VSS(VSS),.VDD(VDD),.Y(g18415),.A(g2108),.B(g15373));
  AND2 AND2_3201(.VSS(VSS),.VDD(VDD),.Y(g31310),.A(g30157),.B(g27886));
  AND2 AND2_3202(.VSS(VSS),.VDD(VDD),.Y(g18333),.A(g1691),.B(g17873));
  AND2 AND2_3203(.VSS(VSS),.VDD(VDD),.Y(g30060),.A(g29146),.B(g10581));
  AND2 AND2_3204(.VSS(VSS),.VDD(VDD),.Y(g21791),.A(g3368),.B(g20391));
  AND2 AND2_3205(.VSS(VSS),.VDD(VDD),.Y(g28253),.A(g23719),.B(g27700));
  AND2 AND2_3206(.VSS(VSS),.VDD(VDD),.Y(g21884),.A(g4104),.B(g19801));
  AND2 AND2_3207(.VSS(VSS),.VDD(VDD),.Y(g11915),.A(g1802),.B(g7315));
  AND2 AND2_3208(.VSS(VSS),.VDD(VDD),.Y(g34968),.A(g34952),.B(g23203));
  AND2 AND2_3209(.VSS(VSS),.VDD(VDD),.Y(g23884),.A(g4119),.B(g19510));
  AND2 AND2_3210(.VSS(VSS),.VDD(VDD),.Y(g30197),.A(g28661),.B(g23859));
  AND2 AND2_3211(.VSS(VSS),.VDD(VDD),.Y(g31959),.A(g4907),.B(g30673));
  AND2 AND2_3212(.VSS(VSS),.VDD(VDD),.Y(g33379),.A(g30984),.B(g32364));
  AND4 AND4_199(.VSS(VSS),.VDD(VDD),.Y(g19462),.A(g7850),.B(g14182),.C(g14177),.D(g16646));
  AND2 AND2_3213(.VSS(VSS),.VDD(VDD),.Y(g25126),.A(g16839),.B(g23523));
  AND2 AND2_3214(.VSS(VSS),.VDD(VDD),.Y(g25987),.A(g9501),.B(g25015));
  AND4 AND4_200(.VSS(VSS),.VDD(VDD),.Y(I31017),.A(g32480),.B(g32481),.C(g32482),.D(g32483));
  AND2 AND2_3215(.VSS(VSS),.VDD(VDD),.Y(g13277),.A(g3195),.B(g11432));
  AND2 AND2_3216(.VSS(VSS),.VDD(VDD),.Y(g28236),.A(g8515),.B(g27971));
  AND2 AND2_3217(.VSS(VSS),.VDD(VDD),.Y(g34870),.A(g34820),.B(g19882));
  AND2 AND2_3218(.VSS(VSS),.VDD(VDD),.Y(g34527),.A(g34303),.B(g19603));
  AND2 AND2_3219(.VSS(VSS),.VDD(VDD),.Y(g24284),.A(g4375),.B(g22550));
  AND2 AND2_3220(.VSS(VSS),.VDD(VDD),.Y(g18664),.A(g4332),.B(g17367));
  AND2 AND2_3221(.VSS(VSS),.VDD(VDD),.Y(g27235),.A(g25910),.B(g19579));
  AND2 AND2_3222(.VSS(VSS),.VDD(VDD),.Y(g24304),.A(g12875),.B(g22228));
  AND2 AND2_3223(.VSS(VSS),.VDD(VDD),.Y(g26819),.A(g106),.B(g24490));
  AND2 AND2_3224(.VSS(VSS),.VDD(VDD),.Y(g27683),.A(g25770),.B(g23567));
  AND2 AND2_3225(.VSS(VSS),.VDD(VDD),.Y(g24622),.A(g19856),.B(g22866));
  AND3 AND3_187(.VSS(VSS),.VDD(VDD),.Y(g33742),.A(g7828),.B(g33142),.C(I31600));
  AND2 AND2_3226(.VSS(VSS),.VDD(VDD),.Y(g26257),.A(g4253),.B(g25197));
  AND2 AND2_3227(.VSS(VSS),.VDD(VDD),.Y(g31944),.A(g31745),.B(g22146));
  AND2 AND2_3228(.VSS(VSS),.VDD(VDD),.Y(g11037),.A(g6128),.B(g9184));
  AND2 AND2_3229(.VSS(VSS),.VDD(VDD),.Y(g18576),.A(g2868),.B(g16349));
  AND2 AND2_3230(.VSS(VSS),.VDD(VDD),.Y(g18585),.A(g2960),.B(g16349));
  AND2 AND2_3231(.VSS(VSS),.VDD(VDD),.Y(g14193),.A(g7178),.B(g10590));
  AND2 AND2_3232(.VSS(VSS),.VDD(VDD),.Y(g18484),.A(g2491),.B(g15426));
  AND2 AND2_3233(.VSS(VSS),.VDD(VDD),.Y(g22109),.A(g6455),.B(g18833));
  AND2 AND2_3234(.VSS(VSS),.VDD(VDD),.Y(g32260),.A(g31250),.B(g20385));
  AND3 AND3_188(.VSS(VSS),.VDD(VDD),.Y(g28264),.A(g7315),.B(g1802),.C(g27416));
  AND2 AND2_3235(.VSS(VSS),.VDD(VDD),.Y(g34503),.A(g34278),.B(g19437));
  AND2 AND2_3236(.VSS(VSS),.VDD(VDD),.Y(g34867),.A(g34826),.B(g20145));
  AND2 AND2_3237(.VSS(VSS),.VDD(VDD),.Y(g25969),.A(g9310),.B(g24987));
  AND2 AND2_3238(.VSS(VSS),.VDD(VDD),.Y(g18554),.A(g2831),.B(g15277));
  AND2 AND2_3239(.VSS(VSS),.VDD(VDD),.Y(g29620),.A(g2399),.B(g29097));
  AND2 AND2_3240(.VSS(VSS),.VDD(VDD),.Y(g33681),.A(g33129),.B(g7991));
  AND2 AND2_3241(.VSS(VSS),.VDD(VDD),.Y(g22108),.A(g6439),.B(g18833));
  AND2 AND2_3242(.VSS(VSS),.VDD(VDD),.Y(g18609),.A(g3147),.B(g16987));
  AND2 AND2_3243(.VSS(VSS),.VDD(VDD),.Y(g27414),.A(g255),.B(g26827));
  AND2 AND2_3244(.VSS(VSS),.VDD(VDD),.Y(g32195),.A(g30734),.B(g25451));
  AND2 AND2_3245(.VSS(VSS),.VDD(VDD),.Y(g24139),.A(g17619),.B(g21653));
  AND2 AND2_3246(.VSS(VSS),.VDD(VDD),.Y(g25968),.A(g25215),.B(g20739));
  AND2 AND2_3247(.VSS(VSS),.VDD(VDD),.Y(g18312),.A(g1579),.B(g16931));
  AND2 AND2_3248(.VSS(VSS),.VDD(VDD),.Y(g33802),.A(g33097),.B(g14545));
  AND2 AND2_3249(.VSS(VSS),.VDD(VDD),.Y(g33429),.A(g32231),.B(g29676));
  AND2 AND2_3250(.VSS(VSS),.VDD(VDD),.Y(g33857),.A(g33267),.B(g20445));
  AND2 AND2_3251(.VSS(VSS),.VDD(VDD),.Y(g29646),.A(g1816),.B(g28675));
  AND3 AND3_189(.VSS(VSS),.VDD(VDD),.Y(g30315),.A(g29182),.B(g7028),.C(g5644));
  AND2 AND2_3252(.VSS(VSS),.VDD(VDD),.Y(g34581),.A(g22864),.B(g34312));
  AND2 AND2_3253(.VSS(VSS),.VDD(VDD),.Y(g18608),.A(g15087),.B(g16987));
  AND2 AND2_3254(.VSS(VSS),.VDD(VDD),.Y(g27407),.A(g26488),.B(g17522));
  AND2 AND2_3255(.VSS(VSS),.VDD(VDD),.Y(g18115),.A(g460),.B(g17015));
  AND4 AND4_201(.VSS(VSS),.VDD(VDD),.Y(I27534),.A(g28039),.B(g24128),.C(g24129),.D(g24130));
  AND4 AND4_202(.VSS(VSS),.VDD(VDD),.Y(g33730),.A(g7202),.B(g4621),.C(g33127),.D(g4633));
  AND2 AND2_3256(.VSS(VSS),.VDD(VDD),.Y(g32016),.A(g8522),.B(g31138));
  AND2 AND2_3257(.VSS(VSS),.VDD(VDD),.Y(g33428),.A(g32230),.B(g29672));
  AND2 AND2_3258(.VSS(VSS),.VDD(VDD),.Y(g34707),.A(g34544),.B(g20579));
  AND2 AND2_3259(.VSS(VSS),.VDD(VDD),.Y(g30202),.A(g28667),.B(g23863));
  AND2 AND2_3260(.VSS(VSS),.VDD(VDD),.Y(g25870),.A(g24840),.B(g16182));
  AND2 AND2_3261(.VSS(VSS),.VDD(VDD),.Y(g30257),.A(g28750),.B(g23952));
  AND3 AND3_190(.VSS(VSS),.VDD(VDD),.Y(g25411),.A(g5062),.B(g23764),.C(I24546));
  AND2 AND2_3262(.VSS(VSS),.VDD(VDD),.Y(g26094),.A(g24936),.B(g9664));
  AND2 AND2_3263(.VSS(VSS),.VDD(VDD),.Y(g31765),.A(g30128),.B(g23968));
  AND2 AND2_3264(.VSS(VSS),.VDD(VDD),.Y(g24415),.A(g4760),.B(g22869));
  AND2 AND2_3265(.VSS(VSS),.VDD(VDD),.Y(g7763),.A(g2965),.B(g2960));
  AND2 AND2_3266(.VSS(VSS),.VDD(VDD),.Y(g24333),.A(g4512),.B(g22228));
  AND2 AND2_3267(.VSS(VSS),.VDD(VDD),.Y(g29369),.A(g28209),.B(g22341));
  AND2 AND2_3268(.VSS(VSS),.VDD(VDD),.Y(g14222),.A(g8655),.B(g11826));
  AND2 AND2_3269(.VSS(VSS),.VDD(VDD),.Y(g21922),.A(g5112),.B(g21468));
  AND2 AND2_3270(.VSS(VSS),.VDD(VDD),.Y(g22982),.A(g19535),.B(g19747));
  AND2 AND2_3271(.VSS(VSS),.VDD(VDD),.Y(g30111),.A(g28565),.B(g20917));
  AND2 AND2_3272(.VSS(VSS),.VDD(VDD),.Y(g18745),.A(g5128),.B(g17847));
  AND2 AND2_3273(.VSS(VSS),.VDD(VDD),.Y(g33690),.A(g33146),.B(g16280));
  AND2 AND2_3274(.VSS(VSS),.VDD(VDD),.Y(g30070),.A(g29167),.B(g9529));
  AND2 AND2_3275(.VSS(VSS),.VDD(VDD),.Y(g34111),.A(g33733),.B(g22936));
  AND2 AND2_3276(.VSS(VSS),.VDD(VDD),.Y(g18799),.A(g6181),.B(g15348));
  AND2 AND2_3277(.VSS(VSS),.VDD(VDD),.Y(g22091),.A(g6415),.B(g18833));
  AND2 AND2_3278(.VSS(VSS),.VDD(VDD),.Y(g23531),.A(g10760),.B(g18930));
  AND2 AND2_3279(.VSS(VSS),.VDD(VDD),.Y(g13853),.A(g4549),.B(g10620));
  AND2 AND2_3280(.VSS(VSS),.VDD(VDD),.Y(g18813),.A(g6513),.B(g15483));
  AND2 AND2_3281(.VSS(VSS),.VDD(VDD),.Y(g30590),.A(g18911),.B(g29812));
  AND2 AND2_3282(.VSS(VSS),.VDD(VDD),.Y(g21740),.A(g3085),.B(g20330));
  AND2 AND2_3283(.VSS(VSS),.VDD(VDD),.Y(g16599),.A(g6601),.B(g15030));
  AND2 AND2_3284(.VSS(VSS),.VDD(VDD),.Y(g26019),.A(g5507),.B(g25032));
  AND2 AND2_3285(.VSS(VSS),.VDD(VDD),.Y(g25503),.A(g6888),.B(g22529));
  AND2 AND2_3286(.VSS(VSS),.VDD(VDD),.Y(g18798),.A(g6177),.B(g15348));
  AND2 AND2_3287(.VSS(VSS),.VDD(VDD),.Y(g28542),.A(g27405),.B(g20275));
  AND2 AND2_3288(.VSS(VSS),.VDD(VDD),.Y(g31504),.A(g29370),.B(g10553));
  AND2 AND2_3289(.VSS(VSS),.VDD(VDD),.Y(g28453),.A(g27582),.B(g10233));
  AND2 AND2_3290(.VSS(VSS),.VDD(VDD),.Y(g27206),.A(g26055),.B(g16691));
  AND3 AND3_191(.VSS(VSS),.VDD(VDD),.Y(g33504),.A(g32772),.B(I31216),.C(I31217));
  AND2 AND2_3291(.VSS(VSS),.VDD(VDD),.Y(g24664),.A(g22652),.B(g19741));
  AND2 AND2_3292(.VSS(VSS),.VDD(VDD),.Y(g29850),.A(g28340),.B(g24893));
  AND2 AND2_3293(.VSS(VSS),.VDD(VDD),.Y(g19911),.A(g14707),.B(g17748));
  AND2 AND2_3294(.VSS(VSS),.VDD(VDD),.Y(g34741),.A(g8899),.B(g34697));
  AND2 AND2_3295(.VSS(VSS),.VDD(VDD),.Y(g16598),.A(g6283),.B(g14899));
  AND2 AND2_3296(.VSS(VSS),.VDD(VDD),.Y(g15810),.A(g3937),.B(g14055));
  AND2 AND2_3297(.VSS(VSS),.VDD(VDD),.Y(g13524),.A(g9995),.B(g11910));
  AND2 AND2_3298(.VSS(VSS),.VDD(VDD),.Y(g17091),.A(g8659),.B(g12940));
  AND2 AND2_3299(.VSS(VSS),.VDD(VDD),.Y(g18184),.A(g785),.B(g17328));
  AND2 AND2_3300(.VSS(VSS),.VDD(VDD),.Y(g21953),.A(g5377),.B(g21514));
  AND2 AND2_3301(.VSS(VSS),.VDD(VDD),.Y(g18805),.A(g6377),.B(g15656));
  AND2 AND2_3302(.VSS(VSS),.VDD(VDD),.Y(g18674),.A(g4340),.B(g15758));
  AND2 AND2_3303(.VSS(VSS),.VDD(VDD),.Y(g23373),.A(g13699),.B(g20195));
  AND2 AND2_3304(.VSS(VSS),.VDD(VDD),.Y(g30094),.A(g28544),.B(g20767));
  AND4 AND4_203(.VSS(VSS),.VDD(VDD),.Y(g27759),.A(g22457),.B(g25224),.C(g26424),.D(g26213));
  AND2 AND2_3305(.VSS(VSS),.VDD(VDD),.Y(g25581),.A(g19338),.B(g24150));
  AND2 AND2_3306(.VSS(VSS),.VDD(VDD),.Y(g25450),.A(g6888),.B(g22497));
  AND2 AND2_3307(.VSS(VSS),.VDD(VDD),.Y(g32042),.A(g27244),.B(g31070));
  AND2 AND2_3308(.VSS(VSS),.VDD(VDD),.Y(g21800),.A(g3546),.B(g20924));
  AND2 AND2_3309(.VSS(VSS),.VDD(VDD),.Y(g24484),.A(g16288),.B(g23208));
  AND2 AND2_3310(.VSS(VSS),.VDD(VDD),.Y(g29896),.A(g2599),.B(g29171));
  AND2 AND2_3311(.VSS(VSS),.VDD(VDD),.Y(g27114),.A(g25997),.B(g16523));
  AND2 AND2_3312(.VSS(VSS),.VDD(VDD),.Y(g32255),.A(g31248),.B(g20381));
  AND2 AND2_3313(.VSS(VSS),.VDD(VDD),.Y(g31129),.A(g1968),.B(g30017));
  AND2 AND2_3314(.VSS(VSS),.VDD(VDD),.Y(g32189),.A(g30824),.B(g25369));
  AND2 AND2_3315(.VSS(VSS),.VDD(VDD),.Y(g21936),.A(g5200),.B(g18997));
  AND2 AND2_3316(.VSS(VSS),.VDD(VDD),.Y(g18732),.A(g4961),.B(g16877));
  AND2 AND2_3317(.VSS(VSS),.VDD(VDD),.Y(g27435),.A(g26549),.B(g17585));
  AND2 AND2_3318(.VSS(VSS),.VDD(VDD),.Y(g18934),.A(g3133),.B(g16096));
  AND2 AND2_3319(.VSS(VSS),.VDD(VDD),.Y(g30735),.A(g29814),.B(g22319));
  AND2 AND2_3320(.VSS(VSS),.VDD(VDD),.Y(g24554),.A(g22490),.B(g19541));
  AND2 AND2_3321(.VSS(VSS),.VDD(VDD),.Y(g27107),.A(g26055),.B(g16514));
  AND2 AND2_3322(.VSS(VSS),.VDD(VDD),.Y(g32270),.A(g31254),.B(g20444));
  AND2 AND2_3323(.VSS(VSS),.VDD(VDD),.Y(g16125),.A(g5152),.B(g14238));
  AND2 AND2_3324(.VSS(VSS),.VDD(VDD),.Y(g16532),.A(g5252),.B(g14841));
  AND2 AND2_3325(.VSS(VSS),.VDD(VDD),.Y(g25818),.A(g8124),.B(g24605));
  AND2 AND2_3326(.VSS(VSS),.VDD(VDD),.Y(g28530),.A(g27383),.B(g20240));
  AND2 AND2_3327(.VSS(VSS),.VDD(VDD),.Y(g31128),.A(g12187),.B(g30016));
  AND2 AND2_3328(.VSS(VSS),.VDD(VDD),.Y(g32188),.A(g27586),.B(g31376));
  AND2 AND2_3329(.VSS(VSS),.VDD(VDD),.Y(g25979),.A(g24517),.B(g19650));
  AND2 AND2_3330(.VSS(VSS),.VDD(VDD),.Y(g28346),.A(g27243),.B(g19800));
  AND2 AND2_3331(.VSS(VSS),.VDD(VDD),.Y(g7251),.A(g452),.B(g392));
  AND2 AND2_3332(.VSS(VSS),.VDD(VDD),.Y(g24312),.A(g4501),.B(g22228));
  AND2 AND2_3333(.VSS(VSS),.VDD(VDD),.Y(g18692),.A(g4732),.B(g16053));
  AND2 AND2_3334(.VSS(VSS),.VDD(VDD),.Y(g18761),.A(g5471),.B(g17929));
  AND2 AND2_3335(.VSS(VSS),.VDD(VDD),.Y(g33245),.A(g32125),.B(g19961));
  AND2 AND2_3336(.VSS(VSS),.VDD(VDD),.Y(g24608),.A(g6500),.B(g23425));
  AND2 AND2_3337(.VSS(VSS),.VDD(VDD),.Y(g25978),.A(g9391),.B(g25001));
  AND2 AND2_3338(.VSS(VSS),.VDD(VDD),.Y(g13313),.A(g475),.B(g11048));
  AND2 AND2_3339(.VSS(VSS),.VDD(VDD),.Y(g15967),.A(g3913),.B(g14058));
  AND2 AND2_3340(.VSS(VSS),.VDD(VDD),.Y(g30196),.A(g28659),.B(g23858));
  AND2 AND2_3341(.VSS(VSS),.VDD(VDD),.Y(g31323),.A(g30150),.B(g27907));
  AND2 AND2_3342(.VSS(VSS),.VDD(VDD),.Y(g29582),.A(g27766),.B(g28608));
  AND2 AND2_3343(.VSS(VSS),.VDD(VDD),.Y(g31299),.A(g30123),.B(g27800));
  AND2 AND2_3344(.VSS(VSS),.VDD(VDD),.Y(g17192),.A(g1677),.B(g13022));
  AND2 AND2_3345(.VSS(VSS),.VDD(VDD),.Y(g34196),.A(g33682),.B(g24485));
  AND2 AND2_3346(.VSS(VSS),.VDD(VDD),.Y(g21762),.A(g3219),.B(g20785));
  AND2 AND2_3347(.VSS(VSS),.VDD(VDD),.Y(g21964),.A(g5441),.B(g21514));
  AND2 AND2_3348(.VSS(VSS),.VDD(VDD),.Y(g25986),.A(g5160),.B(g25013));
  AND2 AND2_3349(.VSS(VSS),.VDD(VDD),.Y(g32030),.A(g4172),.B(g30937));
  AND2 AND2_3350(.VSS(VSS),.VDD(VDD),.Y(g24921),.A(g23721),.B(g20739));
  AND4 AND4_204(.VSS(VSS),.VDD(VDD),.Y(I31016),.A(g30825),.B(g31798),.C(g32478),.D(g32479));
  AND2 AND2_3351(.VSS(VSS),.VDD(VDD),.Y(g31298),.A(g30169),.B(g27886));
  AND2 AND2_3352(.VSS(VSS),.VDD(VDD),.Y(g34526),.A(g34300),.B(g19569));
  AND2 AND2_3353(.VSS(VSS),.VDD(VDD),.Y(g18400),.A(g2012),.B(g15373));
  AND2 AND2_3354(.VSS(VSS),.VDD(VDD),.Y(g10873),.A(g3004),.B(g9015));
  AND2 AND2_3355(.VSS(VSS),.VDD(VDD),.Y(g26077),.A(g9607),.B(g25233));
  AND2 AND2_3356(.VSS(VSS),.VDD(VDD),.Y(g24745),.A(g650),.B(g23550));
  AND2 AND2_3357(.VSS(VSS),.VDD(VDD),.Y(g29627),.A(g28493),.B(g11884));
  AND2 AND2_3358(.VSS(VSS),.VDD(VDD),.Y(g18214),.A(g939),.B(g15979));
  AND2 AND2_3359(.VSS(VSS),.VDD(VDD),.Y(g28292),.A(g23781),.B(g27762));
  AND2 AND2_3360(.VSS(VSS),.VDD(VDD),.Y(g29959),.A(g28953),.B(g12823));
  AND2 AND2_3361(.VSS(VSS),.VDD(VDD),.Y(g22862),.A(g1570),.B(g19673));
  AND3 AND3_192(.VSS(VSS),.VDD(VDD),.Y(g28153),.A(g26424),.B(g22763),.C(g27031));
  AND2 AND2_3362(.VSS(VSS),.VDD(VDD),.Y(g18329),.A(g1612),.B(g17873));
  AND2 AND2_3363(.VSS(VSS),.VDD(VDD),.Y(g25067),.A(g4722),.B(g22885));
  AND2 AND2_3364(.VSS(VSS),.VDD(VDD),.Y(g25094),.A(g23318),.B(g20554));
  AND2 AND2_3365(.VSS(VSS),.VDD(VDD),.Y(g18207),.A(g925),.B(g15938));
  AND2 AND2_3366(.VSS(VSS),.VDD(VDD),.Y(g26689),.A(g15754),.B(g24431));
  AND2 AND2_3367(.VSS(VSS),.VDD(VDD),.Y(g29378),.A(g28137),.B(g22493));
  AND2 AND2_3368(.VSS(VSS),.VDD(VDD),.Y(g13808),.A(g4543),.B(g10607));
  AND2 AND2_3369(.VSS(VSS),.VDD(VDD),.Y(g18539),.A(g2763),.B(g15277));
  AND2 AND2_3370(.VSS(VSS),.VDD(VDD),.Y(g11036),.A(g9806),.B(g5774));
  AND2 AND2_3371(.VSS(VSS),.VDD(VDD),.Y(g26280),.A(g13051),.B(g25248));
  AND2 AND2_3372(.VSS(VSS),.VDD(VDD),.Y(g18328),.A(g1657),.B(g17873));
  AND2 AND2_3373(.VSS(VSS),.VDD(VDD),.Y(g27263),.A(g25940),.B(g19713));
  AND2 AND2_3374(.VSS(VSS),.VDD(VDD),.Y(g21909),.A(g5041),.B(g21468));
  AND2 AND2_3375(.VSS(VSS),.VDD(VDD),.Y(g31232),.A(g30294),.B(g23972));
  AND2 AND2_3376(.VSS(VSS),.VDD(VDD),.Y(g25150),.A(g17480),.B(g23547));
  AND2 AND2_3377(.VSS(VSS),.VDD(VDD),.Y(g22040),.A(g5953),.B(g19147));
  AND2 AND2_3378(.VSS(VSS),.VDD(VDD),.Y(g25801),.A(g8097),.B(g24585));
  AND2 AND2_3379(.VSS(VSS),.VDD(VDD),.Y(g26300),.A(g1968),.B(g25341));
  AND2 AND2_3380(.VSS(VSS),.VDD(VDD),.Y(g34866),.A(g34819),.B(g20106));
  AND2 AND2_3381(.VSS(VSS),.VDD(VDD),.Y(g28136),.A(g27382),.B(g23135));
  AND2 AND2_3382(.VSS(VSS),.VDD(VDD),.Y(g18538),.A(g2759),.B(g15277));
  AND2 AND2_3383(.VSS(VSS),.VDD(VDD),.Y(g15079),.A(g2151),.B(g12955));
  AND2 AND2_3384(.VSS(VSS),.VDD(VDD),.Y(g27332),.A(g12538),.B(g26758));
  AND2 AND2_3385(.VSS(VSS),.VDD(VDD),.Y(g29603),.A(g2265),.B(g29060));
  AND2 AND2_3386(.VSS(VSS),.VDD(VDD),.Y(g24674),.A(g446),.B(g23496));
  AND2 AND2_3387(.VSS(VSS),.VDD(VDD),.Y(g29742),.A(g28288),.B(g10233));
  AND2 AND2_3388(.VSS(VSS),.VDD(VDD),.Y(g21908),.A(g5037),.B(g21468));
  AND2 AND2_3389(.VSS(VSS),.VDD(VDD),.Y(g15078),.A(g10361),.B(g12955));
  AND2 AND2_3390(.VSS(VSS),.VDD(VDD),.Y(g33697),.A(g33160),.B(g13330));
  AND2 AND2_3391(.VSS(VSS),.VDD(VDD),.Y(g30001),.A(g28490),.B(g23486));
  AND2 AND2_3392(.VSS(VSS),.VDD(VDD),.Y(g31995),.A(g28274),.B(g30569));
  AND2 AND2_3393(.VSS(VSS),.VDD(VDD),.Y(g33856),.A(g33266),.B(g20442));
  AND2 AND2_3394(.VSS(VSS),.VDD(VDD),.Y(g26102),.A(g1825),.B(g25099));
  AND2 AND2_3395(.VSS(VSS),.VDD(VDD),.Y(g12135),.A(g9684),.B(g9959));
  AND2 AND2_3396(.VSS(VSS),.VDD(VDD),.Y(g31261),.A(g14754),.B(g30259));
  AND2 AND2_3397(.VSS(VSS),.VDD(VDD),.Y(g26157),.A(g2093),.B(g25136));
  AND2 AND2_3398(.VSS(VSS),.VDD(VDD),.Y(g27406),.A(g26488),.B(g17521));
  AND3 AND3_193(.VSS(VSS),.VDD(VDD),.Y(g34077),.A(g22957),.B(g9104),.C(g33736));
  AND2 AND2_3399(.VSS(VSS),.VDD(VDD),.Y(g27962),.A(g25954),.B(g19597));
  AND2 AND2_3400(.VSS(VSS),.VDD(VDD),.Y(g27361),.A(g26519),.B(g17419));
  AND2 AND2_3401(.VSS(VSS),.VDD(VDD),.Y(g33880),.A(g33290),.B(g20568));
  AND4 AND4_205(.VSS(VSS),.VDD(VDD),.Y(I31042),.A(g32515),.B(g32516),.C(g32517),.D(g32518));
  AND2 AND2_3402(.VSS(VSS),.VDD(VDD),.Y(g18241),.A(g1183),.B(g16431));
  AND2 AND2_3403(.VSS(VSS),.VDD(VDD),.Y(g34706),.A(g34496),.B(g10570));
  AND2 AND2_3404(.VSS(VSS),.VDD(VDD),.Y(g21747),.A(g3061),.B(g20330));
  AND2 AND2_3405(.VSS(VSS),.VDD(VDD),.Y(g32160),.A(g31001),.B(g22995));
  AND2 AND2_3406(.VSS(VSS),.VDD(VDD),.Y(g30256),.A(g28749),.B(g23947));
  AND2 AND2_3407(.VSS(VSS),.VDD(VDD),.Y(g25526),.A(g23720),.B(g21400));
  AND2 AND2_3408(.VSS(VSS),.VDD(VDD),.Y(g28164),.A(g8651),.B(g27528));
  AND2 AND2_3409(.VSS(VSS),.VDD(VDD),.Y(g26231),.A(g1854),.B(g25300));
  AND3 AND3_194(.VSS(VSS),.VDD(VDD),.Y(g33512),.A(g32830),.B(I31256),.C(I31257));
  AND2 AND2_3410(.VSS(VSS),.VDD(VDD),.Y(g14913),.A(g1442),.B(g10939));
  AND2 AND2_3411(.VSS(VSS),.VDD(VDD),.Y(g27500),.A(g26400),.B(g17672));
  AND2 AND2_3412(.VSS(VSS),.VDD(VDD),.Y(g29857),.A(g28386),.B(g23304));
  AND2 AND2_3413(.VSS(VSS),.VDD(VDD),.Y(g15817),.A(g3921),.B(g13929));
  AND2 AND2_3414(.VSS(VSS),.VDD(VDD),.Y(g14614),.A(g11975),.B(g11997));
  AND2 AND2_3415(.VSS(VSS),.VDD(VDD),.Y(g24761),.A(g22751),.B(g19852));
  AND2 AND2_3416(.VSS(VSS),.VDD(VDD),.Y(g19540),.A(g1124),.B(g15904));
  AND2 AND2_3417(.VSS(VSS),.VDD(VDD),.Y(g21814),.A(g3594),.B(g20924));
  AND2 AND2_3418(.VSS(VSS),.VDD(VDD),.Y(g18771),.A(g5685),.B(g15615));
  AND2 AND2_3419(.VSS(VSS),.VDD(VDD),.Y(g16023),.A(g3813),.B(g13584));
  AND2 AND2_3420(.VSS(VSS),.VDD(VDD),.Y(g16224),.A(g14583),.B(g14232));
  AND4 AND4_206(.VSS(VSS),.VDD(VDD),.Y(g11166),.A(g8363),.B(g269),.C(g8296),.D(I14225));
  AND2 AND2_3421(.VSS(VSS),.VDD(VDD),.Y(g18235),.A(g1141),.B(g16326));
  AND2 AND2_3422(.VSS(VSS),.VDD(VDD),.Y(g21751),.A(g3167),.B(g20785));
  AND2 AND2_3423(.VSS(VSS),.VDD(VDD),.Y(g21807),.A(g3566),.B(g20924));
  AND2 AND2_3424(.VSS(VSS),.VDD(VDD),.Y(g21772),.A(g3259),.B(g20785));
  AND2 AND2_3425(.VSS(VSS),.VDD(VDD),.Y(g26854),.A(g2868),.B(g24534));
  AND2 AND2_3426(.VSS(VSS),.VDD(VDD),.Y(g15783),.A(g3215),.B(g14098));
  AND2 AND2_3427(.VSS(VSS),.VDD(VDD),.Y(g21974),.A(g5517),.B(g19074));
  AND2 AND2_3428(.VSS(VSS),.VDD(VDD),.Y(g22062),.A(g6093),.B(g21611));
  AND2 AND2_3429(.VSS(VSS),.VDD(VDD),.Y(g18683),.A(g4674),.B(g15885));
  AND2 AND2_3430(.VSS(VSS),.VDD(VDD),.Y(g25866),.A(g3853),.B(g24648));
  AND2 AND2_3431(.VSS(VSS),.VDD(VDD),.Y(g24400),.A(g3466),.B(g23112));
  AND2 AND2_3432(.VSS(VSS),.VDD(VDD),.Y(g27221),.A(g26055),.B(g16747));
  AND3 AND3_195(.VSS(VSS),.VDD(VDD),.Y(g33831),.A(g23088),.B(g33149),.C(g9104));
  AND2 AND2_3433(.VSS(VSS),.VDD(VDD),.Y(g28327),.A(g27365),.B(g19785));
  AND2 AND2_3434(.VSS(VSS),.VDD(VDD),.Y(g29549),.A(g2012),.B(g28900));
  AND2 AND2_3435(.VSS(VSS),.VDD(VDD),.Y(g34102),.A(g33912),.B(g23599));
  AND2 AND2_3436(.VSS(VSS),.VDD(VDD),.Y(g26511),.A(g19265),.B(g24364));
  AND2 AND2_3437(.VSS(VSS),.VDD(VDD),.Y(g34157),.A(g33794),.B(g20159));
  AND2 AND2_3438(.VSS(VSS),.VDD(VDD),.Y(g23639),.A(g19050),.B(g9104));
  AND4 AND4_207(.VSS(VSS),.VDD(VDD),.Y(I31267),.A(g32840),.B(g32841),.C(g32842),.D(g32843));
  AND2 AND2_3439(.VSS(VSS),.VDD(VDD),.Y(g10565),.A(g8182),.B(g424));
  AND2 AND2_3440(.VSS(VSS),.VDD(VDD),.Y(g28537),.A(g6832),.B(g27089));
  AND2 AND2_3441(.VSS(VSS),.VDD(VDD),.Y(g31499),.A(g29801),.B(g23446));
  AND3 AND3_196(.VSS(VSS),.VDD(VDD),.Y(g33499),.A(g32737),.B(I31191),.C(I31192));
  AND2 AND2_3442(.VSS(VSS),.VDD(VDD),.Y(g14565),.A(g11934),.B(g11952));
  AND2 AND2_3443(.VSS(VSS),.VDD(VDD),.Y(g29548),.A(g1798),.B(g28575));
  AND2 AND2_3444(.VSS(VSS),.VDD(VDD),.Y(g23293),.A(g9104),.B(g19200));
  AND2 AND2_3445(.VSS(VSS),.VDD(VDD),.Y(g24329),.A(g4462),.B(g22228));
  AND2 AND2_3446(.VSS(VSS),.VDD(VDD),.Y(g30066),.A(g28518),.B(g20636));
  AND2 AND2_3447(.VSS(VSS),.VDD(VDD),.Y(g22851),.A(g496),.B(g19654));
  AND2 AND2_3448(.VSS(VSS),.VDD(VDD),.Y(g28108),.A(g7975),.B(g27237));
  AND2 AND2_3449(.VSS(VSS),.VDD(VDD),.Y(g30231),.A(g28718),.B(g23907));
  AND2 AND2_3450(.VSS(VSS),.VDD(VDD),.Y(g15823),.A(g3945),.B(g14116));
  AND2 AND2_3451(.VSS(VSS),.VDD(VDD),.Y(g34066),.A(g33730),.B(g19352));
  AND2 AND2_3452(.VSS(VSS),.VDD(VDD),.Y(g10034),.A(g1521),.B(g1500));
  AND2 AND2_3453(.VSS(VSS),.VDD(VDD),.Y(g25077),.A(g23297),.B(g20536));
  AND3 AND3_197(.VSS(VSS),.VDD(VDD),.Y(g33498),.A(g32730),.B(I31186),.C(I31187));
  AND2 AND2_3454(.VSS(VSS),.VDD(VDD),.Y(g23265),.A(g20069),.B(g20132));
  AND2 AND2_3455(.VSS(VSS),.VDD(VDD),.Y(g24328),.A(g4567),.B(g22228));
  AND3 AND3_198(.VSS(VSS),.VDD(VDD),.Y(g28283),.A(g7380),.B(g2361),.C(g27445));
  AND2 AND2_3456(.VSS(VSS),.VDD(VDD),.Y(g18515),.A(g2643),.B(g15509));
  AND2 AND2_3457(.VSS(VSS),.VDD(VDD),.Y(g23416),.A(g20082),.B(g20321));
  AND2 AND2_3458(.VSS(VSS),.VDD(VDD),.Y(g18414),.A(g2102),.B(g15373));
  AND2 AND2_3459(.VSS(VSS),.VDD(VDD),.Y(g31989),.A(g31770),.B(g22200));
  AND2 AND2_3460(.VSS(VSS),.VDD(VDD),.Y(g14641),.A(g11994),.B(g12020));
  AND3 AND3_199(.VSS(VSS),.VDD(VDD),.Y(g28303),.A(g7462),.B(g2629),.C(g27494));
  AND2 AND2_3461(.VSS(VSS),.VDD(VDD),.Y(g27106),.A(g26026),.B(g16512));
  AND2 AND2_3462(.VSS(VSS),.VDD(VDD),.Y(g21841),.A(g3857),.B(g21070));
  AND2 AND2_3463(.VSS(VSS),.VDD(VDD),.Y(g21992),.A(g5599),.B(g19074));
  AND2 AND2_3464(.VSS(VSS),.VDD(VDD),.Y(g34876),.A(g34844),.B(g20534));
  AND2 AND2_3465(.VSS(VSS),.VDD(VDD),.Y(g18407),.A(g2016),.B(g15373));
  AND2 AND2_3466(.VSS(VSS),.VDD(VDD),.Y(g25923),.A(g24443),.B(g19443));
  AND2 AND2_3467(.VSS(VSS),.VDD(VDD),.Y(g31988),.A(g31768),.B(g22199));
  AND2 AND2_3468(.VSS(VSS),.VDD(VDD),.Y(g33722),.A(g33175),.B(g19445));
  AND2 AND2_3469(.VSS(VSS),.VDD(VDD),.Y(g33924),.A(g33335),.B(g33346));
  AND2 AND2_3470(.VSS(VSS),.VDD(VDD),.Y(g32419),.A(g4955),.B(g31000));
  AND2 AND2_3471(.VSS(VSS),.VDD(VDD),.Y(g15966),.A(g3462),.B(g13555));
  AND4 AND4_208(.VSS(VSS),.VDD(VDD),.Y(g28982),.A(g27163),.B(g12687),.C(g20682),.D(I27349));
  AND2 AND2_3472(.VSS(VSS),.VDD(VDD),.Y(g31271),.A(g29706),.B(g23300));
  AND2 AND2_3473(.VSS(VSS),.VDD(VDD),.Y(g12812),.A(g518),.B(g9158));
  AND2 AND2_3474(.VSS(VSS),.VDD(VDD),.Y(g34763),.A(g34689),.B(g19915));
  AND2 AND2_3475(.VSS(VSS),.VDD(VDD),.Y(g15631),.A(g168),.B(g13437));
  AND2 AND2_3476(.VSS(VSS),.VDD(VDD),.Y(g27033),.A(g25767),.B(g19273));
  AND2 AND2_3477(.VSS(VSS),.VDD(VDD),.Y(g27371),.A(g26400),.B(g17473));
  AND2 AND2_3478(.VSS(VSS),.VDD(VDD),.Y(g32418),.A(g31126),.B(g16239));
  AND2 AND2_3479(.VSS(VSS),.VDD(VDD),.Y(g26287),.A(g2138),.B(g25225));
  AND2 AND2_3480(.VSS(VSS),.VDD(VDD),.Y(g27234),.A(g26055),.B(g16814));
  AND2 AND2_3481(.VSS(VSS),.VDD(VDD),.Y(g25102),.A(g4727),.B(g22885));
  AND2 AND2_3482(.VSS(VSS),.VDD(VDD),.Y(g21835),.A(g3802),.B(g20453));
  AND2 AND2_3483(.VSS(VSS),.VDD(VDD),.Y(g32170),.A(g31671),.B(g27779));
  AND2 AND2_3484(.VSS(VSS),.VDD(VDD),.Y(g13567),.A(g10102),.B(g11948));
  AND2 AND2_3485(.VSS(VSS),.VDD(VDD),.Y(g22047),.A(g6077),.B(g21611));
  AND2 AND2_3486(.VSS(VSS),.VDD(VDD),.Y(g26307),.A(g13070),.B(g25288));
  AND2 AND2_3487(.VSS(VSS),.VDD(VDD),.Y(g26085),.A(g11906),.B(g25070));
  AND2 AND2_3488(.VSS(VSS),.VDD(VDD),.Y(g29626),.A(g28584),.B(g11415));
  AND3 AND3_200(.VSS(VSS),.VDD(VDD),.Y(g33461),.A(g32463),.B(I31001),.C(I31002));
  AND2 AND2_3489(.VSS(VSS),.VDD(VDD),.Y(g16669),.A(g5611),.B(g14993));
  AND2 AND2_3490(.VSS(VSS),.VDD(VDD),.Y(g33342),.A(g32226),.B(g20660));
  AND3 AND3_201(.VSS(VSS),.VDD(VDD),.Y(g29323),.A(g28539),.B(g6905),.C(g3639));
  AND2 AND2_3491(.VSS(VSS),.VDD(VDD),.Y(g23007),.A(g681),.B(g20248));
  AND2 AND2_3492(.VSS(VSS),.VDD(VDD),.Y(g31145),.A(g9970),.B(g30052));
  AND2 AND2_3493(.VSS(VSS),.VDD(VDD),.Y(g18441),.A(g2246),.B(g18008));
  AND2 AND2_3494(.VSS(VSS),.VDD(VDD),.Y(g18584),.A(g2950),.B(g16349));
  AND2 AND2_3495(.VSS(VSS),.VDD(VDD),.Y(g24771),.A(g7028),.B(g23605));
  AND2 AND2_3496(.VSS(VSS),.VDD(VDD),.Y(g18206),.A(g918),.B(g15938));
  AND2 AND2_3497(.VSS(VSS),.VDD(VDD),.Y(g29533),.A(g28958),.B(g22417));
  AND2 AND2_3498(.VSS(VSS),.VDD(VDD),.Y(g12795),.A(g1312),.B(g7601));
  AND2 AND2_3499(.VSS(VSS),.VDD(VDD),.Y(g16668),.A(g5543),.B(g14962));
  AND2 AND2_3500(.VSS(VSS),.VDD(VDD),.Y(g16842),.A(g6279),.B(g14861));
  AND2 AND2_3501(.VSS(VSS),.VDD(VDD),.Y(g17574),.A(g9554),.B(g14546));
  AND2 AND2_3502(.VSS(VSS),.VDD(VDD),.Y(g33887),.A(g33298),.B(g20615));
  AND2 AND2_3503(.VSS(VSS),.VDD(VDD),.Y(g18759),.A(g5467),.B(g17929));
  AND2 AND2_3504(.VSS(VSS),.VDD(VDD),.Y(g22051),.A(g6105),.B(g21611));
  AND2 AND2_3505(.VSS(VSS),.VDD(VDD),.Y(g22072),.A(g6259),.B(g19210));
  AND2 AND2_3506(.VSS(VSS),.VDD(VDD),.Y(g18725),.A(g4912),.B(g16077));
  AND2 AND2_3507(.VSS(VSS),.VDD(VDD),.Y(g32167),.A(g3853),.B(g31194));
  AND2 AND2_3508(.VSS(VSS),.VDD(VDD),.Y(g32194),.A(g30601),.B(g28436));
  AND2 AND2_3509(.VSS(VSS),.VDD(VDD),.Y(g25876),.A(g3470),.B(g24667));
  AND3 AND3_202(.VSS(VSS),.VDD(VDD),.Y(g33529),.A(g32953),.B(I31341),.C(I31342));
  AND4 AND4_209(.VSS(VSS),.VDD(VDD),.Y(I31201),.A(g31672),.B(g31831),.C(g32745),.D(g32746));
  AND2 AND2_3510(.VSS(VSS),.VDD(VDD),.Y(g27507),.A(g26549),.B(g17683));
  AND4 AND4_210(.VSS(VSS),.VDD(VDD),.Y(I31277),.A(g32856),.B(g32857),.C(g32858),.D(g32859));
  AND2 AND2_3511(.VSS(VSS),.VDD(VDD),.Y(g18114),.A(g452),.B(g17015));
  AND2 AND2_3512(.VSS(VSS),.VDD(VDD),.Y(g28192),.A(g8891),.B(g27415));
  AND2 AND2_3513(.VSS(VSS),.VDD(VDD),.Y(g18758),.A(g7004),.B(g15595));
  AND2 AND2_3514(.VSS(VSS),.VDD(VDD),.Y(g31528),.A(g19050),.B(g29814));
  AND2 AND2_3515(.VSS(VSS),.VDD(VDD),.Y(g26341),.A(g24746),.B(g20105));
  AND2 AND2_3516(.VSS(VSS),.VDD(VDD),.Y(g18435),.A(g2173),.B(g18008));
  AND3 AND3_203(.VSS(VSS),.VDD(VDD),.Y(g33528),.A(g32946),.B(I31336),.C(I31337));
  AND2 AND2_3517(.VSS(VSS),.VDD(VDD),.Y(g34287),.A(g11370),.B(g34124));
  AND2 AND2_3518(.VSS(VSS),.VDD(VDD),.Y(g19661),.A(g5489),.B(g16969));
  AND2 AND2_3519(.VSS(VSS),.VDD(VDD),.Y(g33843),.A(g33256),.B(g20325));
  AND2 AND2_3520(.VSS(VSS),.VDD(VDD),.Y(g21720),.A(g376),.B(g21037));
  AND2 AND2_3521(.VSS(VSS),.VDD(VDD),.Y(g33330),.A(g32211),.B(g20588));
  AND2 AND2_3522(.VSS(VSS),.VDD(VDD),.Y(g26156),.A(g2028),.B(g25135));
  AND2 AND2_3523(.VSS(VSS),.VDD(VDD),.Y(g18107),.A(g429),.B(g17015));
  AND4 AND4_211(.VSS(VSS),.VDD(VDD),.Y(g27421),.A(g8038),.B(g26314),.C(g9187),.D(g9077));
  AND3 AND3_204(.VSS(VSS),.VDD(VDD),.Y(g34085),.A(g33761),.B(g9104),.C(g18957));
  AND2 AND2_3524(.VSS(VSS),.VDD(VDD),.Y(g28663),.A(g27566),.B(g20624));
  AND2 AND2_3525(.VSS(VSS),.VDD(VDD),.Y(g32401),.A(g31116),.B(g13432));
  AND2 AND2_3526(.VSS(VSS),.VDD(VDD),.Y(g34076),.A(g33694),.B(g19519));
  AND2 AND2_3527(.VSS(VSS),.VDD(VDD),.Y(g30596),.A(g30279),.B(g18947));
  AND2 AND2_3528(.VSS(VSS),.VDD(VDD),.Y(g26180),.A(g2587),.B(g25156));
  AND2 AND2_3529(.VSS(VSS),.VDD(VDD),.Y(g26670),.A(g13385),.B(g24428));
  AND2 AND2_3530(.VSS(VSS),.VDD(VDD),.Y(g21746),.A(g3045),.B(g20330));
  AND2 AND2_3531(.VSS(VSS),.VDD(VDD),.Y(g33365),.A(g32267),.B(g20994));
  AND2 AND2_3532(.VSS(VSS),.VDD(VDD),.Y(g32119),.A(g31609),.B(g29939));
  AND2 AND2_3533(.VSS(VSS),.VDD(VDD),.Y(g30243),.A(g28731),.B(g23929));
  AND2 AND2_3534(.VSS(VSS),.VDD(VDD),.Y(g31132),.A(g29504),.B(g22987));
  AND2 AND2_3535(.VSS(VSS),.VDD(VDD),.Y(g18744),.A(g5124),.B(g17847));
  AND2 AND2_3536(.VSS(VSS),.VDD(VDD),.Y(g34054),.A(g33778),.B(g22942));
  AND2 AND2_3537(.VSS(VSS),.VDD(VDD),.Y(g31960),.A(g31749),.B(g22153));
  AND2 AND2_3538(.VSS(VSS),.VDD(VDD),.Y(g33869),.A(g33279),.B(g20543));
  AND2 AND2_3539(.VSS(VSS),.VDD(VDD),.Y(g14537),.A(g10550),.B(g10529));
  AND2 AND2_3540(.VSS(VSS),.VDD(VDD),.Y(g18345),.A(g1736),.B(g17955));
  AND2 AND2_3541(.VSS(VSS),.VDD(VDD),.Y(g19715),.A(g9679),.B(g17120));
  AND4 AND4_212(.VSS(VSS),.VDD(VDD),.Y(I31037),.A(g32508),.B(g32509),.C(g32510),.D(g32511));
  AND2 AND2_3542(.VSS(VSS),.VDD(VDD),.Y(g29856),.A(g28385),.B(g23303));
  AND4 AND4_213(.VSS(VSS),.VDD(VDD),.Y(g17780),.A(g6772),.B(g11592),.C(g11640),.D(I18782));
  AND2 AND2_3543(.VSS(VSS),.VDD(VDD),.Y(g21465),.A(g16155),.B(g13663));
  AND2 AND2_3544(.VSS(VSS),.VDD(VDD),.Y(g18399),.A(g2024),.B(g15373));
  AND2 AND2_3545(.VSS(VSS),.VDD(VDD),.Y(g29880),.A(g1936),.B(g29149));
  AND2 AND2_3546(.VSS(VSS),.VDD(VDD),.Y(g33868),.A(g33278),.B(g20542));
  AND2 AND2_3547(.VSS(VSS),.VDD(VDD),.Y(g26839),.A(g2988),.B(g24516));
  AND2 AND2_3548(.VSS(VSS),.VDD(VDD),.Y(g27541),.A(g26278),.B(g23334));
  AND2 AND2_3549(.VSS(VSS),.VDD(VDD),.Y(g30269),.A(g28778),.B(g23970));
  AND2 AND2_3550(.VSS(VSS),.VDD(VDD),.Y(g22846),.A(g9386),.B(g20676));
  AND2 AND2_3551(.VSS(VSS),.VDD(VDD),.Y(g21983),.A(g5555),.B(g19074));
  AND2 AND2_3552(.VSS(VSS),.VDD(VDD),.Y(g28553),.A(g27187),.B(g10290));
  AND3 AND3_205(.VSS(VSS),.VDD(VDD),.Y(g25456),.A(g5752),.B(g22210),.C(I24579));
  AND2 AND2_3553(.VSS(VSS),.VDD(VDD),.Y(g18398),.A(g2020),.B(g15373));
  AND2 AND2_3554(.VSS(VSS),.VDD(VDD),.Y(g29512),.A(g2161),.B(g28793));
  AND2 AND2_3555(.VSS(VSS),.VDD(VDD),.Y(g32313),.A(g31303),.B(g23515));
  AND4 AND4_214(.VSS(VSS),.VDD(VDD),.Y(I31352),.A(g32963),.B(g32964),.C(g32965),.D(g32966));
  AND2 AND2_3556(.VSS(VSS),.VDD(VDD),.Y(g21806),.A(g3558),.B(g20924));
  AND2 AND2_3557(.VSS(VSS),.VDD(VDD),.Y(g26838),.A(g2860),.B(g24515));
  AND2 AND2_3558(.VSS(VSS),.VDD(VDD),.Y(g18141),.A(g568),.B(g17533));
  AND2 AND2_3559(.VSS(VSS),.VDD(VDD),.Y(g30268),.A(g28777),.B(g23969));
  AND2 AND2_3560(.VSS(VSS),.VDD(VDD),.Y(g18652),.A(g4172),.B(g16249));
  AND2 AND2_3561(.VSS(VSS),.VDD(VDD),.Y(g18804),.A(g15163),.B(g15656));
  AND2 AND2_3562(.VSS(VSS),.VDD(VDD),.Y(g34341),.A(g34101),.B(g19952));
  AND2 AND2_3563(.VSS(VSS),.VDD(VDD),.Y(g25916),.A(g24432),.B(g19434));
  AND2 AND2_3564(.VSS(VSS),.VDD(VDD),.Y(g16610),.A(g5260),.B(g14918));
  AND2 AND2_3565(.VSS(VSS),.VDD(VDD),.Y(g16705),.A(g6299),.B(g15024));
  AND2 AND2_3566(.VSS(VSS),.VDD(VDD),.Y(g17152),.A(g8635),.B(g12997));
  AND2 AND2_3567(.VSS(VSS),.VDD(VDD),.Y(g31225),.A(g30276),.B(g21012));
  AND2 AND2_3568(.VSS(VSS),.VDD(VDD),.Y(g32276),.A(g31646),.B(g30313));
  AND4 AND4_215(.VSS(VSS),.VDD(VDD),.Y(g27724),.A(g22417),.B(g25208),.C(g26424),.D(g26190));
  AND2 AND2_3569(.VSS(VSS),.VDD(VDD),.Y(g34655),.A(g34573),.B(g18885));
  AND4 AND4_216(.VSS(VSS),.VDD(VDD),.Y(I31266),.A(g31327),.B(g31843),.C(g32838),.D(g32839));
  AND2 AND2_3570(.VSS(VSS),.VDD(VDD),.Y(g27359),.A(g26488),.B(g17416));
  AND2 AND2_3571(.VSS(VSS),.VDD(VDD),.Y(g30180),.A(g28635),.B(g23820));
  AND2 AND2_3572(.VSS(VSS),.VDD(VDD),.Y(g27325),.A(g12478),.B(g26724));
  AND2 AND2_3573(.VSS(VSS),.VDD(VDD),.Y(g30670),.A(g11330),.B(g29359));
  AND2 AND2_3574(.VSS(VSS),.VDD(VDD),.Y(g31471),.A(g29754),.B(g23399));
  AND2 AND2_3575(.VSS(VSS),.VDD(VDD),.Y(g32305),.A(g31287),.B(g20567));
  AND2 AND2_3576(.VSS(VSS),.VDD(VDD),.Y(g32053),.A(g14176),.B(g31509));
  AND3 AND3_206(.VSS(VSS),.VDD(VDD),.Y(g33471),.A(g32535),.B(I31051),.C(I31052));
  AND2 AND2_3577(.VSS(VSS),.VDD(VDD),.Y(g34180),.A(g33716),.B(g24373));
  AND2 AND2_3578(.VSS(VSS),.VDD(VDD),.Y(g33087),.A(g32391),.B(g18888));
  AND2 AND2_3579(.VSS(VSS),.VDD(VDD),.Y(g18263),.A(g1249),.B(g16000));
  AND2 AND2_3580(.VSS(VSS),.VDD(VDD),.Y(g32254),.A(g31247),.B(g20379));
  AND2 AND2_3581(.VSS(VSS),.VDD(VDD),.Y(g27535),.A(g26519),.B(g17737));
  AND2 AND2_3582(.VSS(VSS),.VDD(VDD),.Y(g26487),.A(g15702),.B(g24359));
  AND2 AND2_3583(.VSS(VSS),.VDD(VDD),.Y(g27434),.A(g26549),.B(g17584));
  AND2 AND2_3584(.VSS(VSS),.VDD(VDD),.Y(g27358),.A(g26400),.B(g17415));
  AND2 AND2_3585(.VSS(VSS),.VDD(VDD),.Y(g25076),.A(g12805),.B(g23479));
  AND2 AND2_3586(.VSS(VSS),.VDD(VDD),.Y(g25085),.A(g4912),.B(g22908));
  AND2 AND2_3587(.VSS(VSS),.VDD(VDD),.Y(g18332),.A(g1677),.B(g17873));
  AND2 AND2_3588(.VSS(VSS),.VDD(VDD),.Y(g19784),.A(g2775),.B(g15877));
  AND2 AND2_3589(.VSS(VSS),.VDD(VDD),.Y(g28252),.A(g27159),.B(g19682));
  AND2 AND2_3590(.VSS(VSS),.VDD(VDD),.Y(g12920),.A(g1227),.B(g10960));
  AND2 AND2_3591(.VSS(VSS),.VDD(VDD),.Y(g18135),.A(g136),.B(g17249));
  AND2 AND2_3592(.VSS(VSS),.VDD(VDD),.Y(g34335),.A(g8461),.B(g34197));
  AND2 AND2_3593(.VSS(VSS),.VDD(VDD),.Y(g25054),.A(g12778),.B(g23452));
  AND2 AND2_3594(.VSS(VSS),.VDD(VDD),.Y(g24725),.A(g19587),.B(g23012));
  AND2 AND2_3595(.VSS(VSS),.VDD(VDD),.Y(g30930),.A(g29915),.B(g23342));
  AND2 AND2_3596(.VSS(VSS),.VDD(VDD),.Y(g32036),.A(g31469),.B(g13486));
  AND2 AND2_3597(.VSS(VSS),.VDD(VDD),.Y(g27121),.A(g136),.B(g26326));
  AND3 AND3_207(.VSS(VSS),.VDD(VDD),.Y(g29316),.A(g28528),.B(g6875),.C(g3288));
  AND2 AND2_3598(.VSS(VSS),.VDD(VDD),.Y(g19354),.A(g471),.B(g16235));
  AND2 AND2_3599(.VSS(VSS),.VDD(VDD),.Y(g33244),.A(g32190),.B(g23152));
  AND2 AND2_3600(.VSS(VSS),.VDD(VDD),.Y(g32177),.A(g30608),.B(g25214));
  AND2 AND2_3601(.VSS(VSS),.VDD(VDD),.Y(g18406),.A(g2060),.B(g15373));
  AND2 AND2_3602(.VSS(VSS),.VDD(VDD),.Y(g13349),.A(g4933),.B(g11780));
  AND4 AND4_217(.VSS(VSS),.VDD(VDD),.Y(I31167),.A(g32696),.B(g32697),.C(g32698),.D(g32699));
  AND3 AND3_208(.VSS(VSS),.VDD(VDD),.Y(I18785),.A(g13156),.B(g6767),.C(g11498));
  AND2 AND2_3603(.VSS(VSS),.VDD(VDD),.Y(g26279),.A(g4249),.B(g25213));
  AND2 AND2_3604(.VSS(VSS),.VDD(VDD),.Y(g18361),.A(g1821),.B(g17955));
  AND2 AND2_3605(.VSS(VSS),.VDD(VDD),.Y(g24758),.A(g6523),.B(g23733));
  AND2 AND2_3606(.VSS(VSS),.VDD(VDD),.Y(g23130),.A(g728),.B(g20248));
  AND2 AND2_3607(.VSS(VSS),.VDD(VDD),.Y(g34667),.A(g34471),.B(g33424));
  AND2 AND2_3608(.VSS(VSS),.VDD(VDD),.Y(g34694),.A(g34530),.B(g19885));
  AND2 AND2_3609(.VSS(VSS),.VDD(VDD),.Y(g17405),.A(g1422),.B(g13137));
  AND2 AND2_3610(.VSS(VSS),.VDD(VDD),.Y(g11083),.A(g8836),.B(g802));
  AND2 AND2_3611(.VSS(VSS),.VDD(VDD),.Y(g34965),.A(g34949),.B(g23084));
  AND2 AND2_3612(.VSS(VSS),.VDD(VDD),.Y(g30131),.A(g28589),.B(g21178));
  AND2 AND2_3613(.VSS(VSS),.VDD(VDD),.Y(g31069),.A(g29793),.B(g14150));
  AND2 AND2_3614(.VSS(VSS),.VDD(VDD),.Y(g19671),.A(g1454),.B(g16155));
  AND2 AND2_3615(.VSS(VSS),.VDD(VDD),.Y(g29989),.A(g29006),.B(g10489));
  AND2 AND2_3616(.VSS(VSS),.VDD(VDD),.Y(g18500),.A(g2421),.B(g15426));
  AND2 AND2_3617(.VSS(VSS),.VDD(VDD),.Y(g22020),.A(g5863),.B(g19147));
  AND2 AND2_3618(.VSS(VSS),.VDD(VDD),.Y(g27682),.A(g25777),.B(g23565));
  AND2 AND2_3619(.VSS(VSS),.VDD(VDD),.Y(g23165),.A(g13954),.B(g19964));
  AND2 AND2_3620(.VSS(VSS),.VDD(VDD),.Y(g28183),.A(g27024),.B(g19421));
  AND2 AND2_3621(.VSS(VSS),.VDD(VDD),.Y(g28673),.A(g1373),.B(g27122));
  AND2 AND2_3622(.VSS(VSS),.VDD(VDD),.Y(g33810),.A(g33427),.B(g12768));
  AND2 AND2_3623(.VSS(VSS),.VDD(VDD),.Y(g27291),.A(g11969),.B(g26653));
  AND2 AND2_3624(.VSS(VSS),.VDD(VDD),.Y(g29611),.A(g28540),.B(g14209));
  AND2 AND2_3625(.VSS(VSS),.VDD(VDD),.Y(g33657),.A(g30991),.B(g33443));
  AND2 AND2_3626(.VSS(VSS),.VDD(VDD),.Y(g26286),.A(g2126),.B(g25389));
  AND2 AND2_3627(.VSS(VSS),.VDD(VDD),.Y(g29988),.A(g29187),.B(g12235));
  AND2 AND2_3628(.VSS(VSS),.VDD(VDD),.Y(g29924),.A(g13031),.B(g29190));
  AND2 AND2_3629(.VSS(VSS),.VDD(VDD),.Y(g34487),.A(g34416),.B(g18983));
  AND2 AND2_3630(.VSS(VSS),.VDD(VDD),.Y(g13566),.A(g7092),.B(g12358));
  AND2 AND2_3631(.VSS(VSS),.VDD(VDD),.Y(g22046),.A(g6073),.B(g21611));
  AND2 AND2_3632(.VSS(VSS),.VDD(VDD),.Y(g26306),.A(g13087),.B(g25286));
  AND2 AND2_3633(.VSS(VSS),.VDD(VDD),.Y(g24849),.A(g4165),.B(g22227));
  AND2 AND2_3634(.VSS(VSS),.VDD(VDD),.Y(g33879),.A(g33289),.B(g20566));
  AND2 AND2_3635(.VSS(VSS),.VDD(VDD),.Y(g24940),.A(g5011),.B(g23971));
  AND2 AND2_3636(.VSS(VSS),.VDD(VDD),.Y(g24399),.A(g3133),.B(g23067));
  AND2 AND2_3637(.VSS(VSS),.VDD(VDD),.Y(g34502),.A(g26363),.B(g34343));
  AND2 AND2_3638(.VSS(VSS),.VDD(VDD),.Y(g30210),.A(g28684),.B(g23877));
  AND2 AND2_3639(.VSS(VSS),.VDD(VDD),.Y(g34557),.A(g34352),.B(g20555));
  AND2 AND2_3640(.VSS(VSS),.VDD(VDD),.Y(g23006),.A(g19575),.B(g19776));
  AND2 AND2_3641(.VSS(VSS),.VDD(VDD),.Y(g23475),.A(g19070),.B(g8971));
  AND2 AND2_3642(.VSS(VSS),.VDD(VDD),.Y(g33878),.A(g33288),.B(g20565));
  AND4 AND4_218(.VSS(VSS),.VDD(VDD),.Y(I31022),.A(g32487),.B(g32488),.C(g32489),.D(g32490));
  AND2 AND2_3643(.VSS(VSS),.VDD(VDD),.Y(g18221),.A(g1018),.B(g16100));
  AND2 AND2_3644(.VSS(VSS),.VDD(VDD),.Y(g22113),.A(g6561),.B(g19277));
  AND2 AND2_3645(.VSS(VSS),.VDD(VDD),.Y(g21863),.A(g3957),.B(g21070));
  AND2 AND2_3646(.VSS(VSS),.VDD(VDD),.Y(g26815),.A(g4108),.B(g24528));
  AND2 AND2_3647(.VSS(VSS),.VDD(VDD),.Y(g24141),.A(g17657),.B(g21656));
  AND2 AND2_3648(.VSS(VSS),.VDD(VDD),.Y(g34279),.A(g34231),.B(g19208));
  AND4 AND4_219(.VSS(VSS),.VDD(VDD),.Y(g11139),.A(g5990),.B(g7051),.C(g5976),.D(g9935));
  AND2 AND2_3649(.VSS(VSS),.VDD(VDD),.Y(g33886),.A(g33297),.B(g20614));
  AND2 AND2_3650(.VSS(VSS),.VDD(VDD),.Y(g27134),.A(g25997),.B(g16602));
  AND2 AND2_3651(.VSS(VSS),.VDD(VDD),.Y(g30278),.A(g28818),.B(g23988));
  AND2 AND2_3652(.VSS(VSS),.VDD(VDD),.Y(g27029),.A(g26327),.B(g11031));
  AND2 AND2_3653(.VSS(VSS),.VDD(VDD),.Y(g18613),.A(g3338),.B(g17200));
  AND2 AND2_3654(.VSS(VSS),.VDD(VDD),.Y(g31792),.A(g30214),.B(g24017));
  AND2 AND2_3655(.VSS(VSS),.VDD(VDD),.Y(g32166),.A(g31007),.B(g23029));
  AND2 AND2_3656(.VSS(VSS),.VDD(VDD),.Y(g32009),.A(g31782),.B(g22224));
  AND2 AND2_3657(.VSS(VSS),.VDD(VDD),.Y(g25993),.A(g2610),.B(g25025));
  AND2 AND2_3658(.VSS(VSS),.VDD(VDD),.Y(g31967),.A(g31755),.B(g22167));
  AND2 AND2_3659(.VSS(VSS),.VDD(VDD),.Y(g31994),.A(g31775),.B(g22215));
  AND2 AND2_3660(.VSS(VSS),.VDD(VDD),.Y(g22105),.A(g6494),.B(g18833));
  AND4 AND4_220(.VSS(VSS),.VDD(VDD),.Y(I31276),.A(g31376),.B(g31844),.C(g32854),.D(g32855));
  AND2 AND2_3661(.VSS(VSS),.VDD(VDD),.Y(g27028),.A(g26342),.B(g1157));
  AND2 AND2_3662(.VSS(VSS),.VDD(VDD),.Y(g29199),.A(g27187),.B(g12687));
  AND2 AND2_3663(.VSS(VSS),.VDD(VDD),.Y(g32008),.A(g31781),.B(g22223));
  AND2 AND2_3664(.VSS(VSS),.VDD(VDD),.Y(g25965),.A(g2208),.B(g24980));
  AND2 AND2_3665(.VSS(VSS),.VDD(VDD),.Y(g29650),.A(g28949),.B(g22472));
  AND2 AND2_3666(.VSS(VSS),.VDD(VDD),.Y(g29736),.A(g28522),.B(g10233));
  AND2 AND2_3667(.VSS(VSS),.VDD(VDD),.Y(g16160),.A(g5499),.B(g14262));
  AND2 AND2_3668(.VSS(VSS),.VDD(VDD),.Y(g29887),.A(g28417),.B(g23351));
  AND2 AND2_3669(.VSS(VSS),.VDD(VDD),.Y(g21703),.A(g146),.B(g20283));
  AND2 AND2_3670(.VSS(VSS),.VDD(VDD),.Y(g18273),.A(g1287),.B(g16031));
  AND2 AND2_3671(.VSS(VSS),.VDD(VDD),.Y(g24332),.A(g4459),.B(g22228));
  AND2 AND2_3672(.VSS(VSS),.VDD(VDD),.Y(g18106),.A(g411),.B(g17015));
  AND2 AND2_3673(.VSS(VSS),.VDD(VDD),.Y(g20135),.A(g16258),.B(g16695));
  AND2 AND2_3674(.VSS(VSS),.VDD(VDD),.Y(g18605),.A(g3129),.B(g16987));
  AND2 AND2_3675(.VSS(VSS),.VDD(VDD),.Y(g13415),.A(g837),.B(g11048));
  AND2 AND2_3676(.VSS(VSS),.VDD(VDD),.Y(g21347),.A(g1339),.B(g15750));
  AND2 AND2_3677(.VSS(VSS),.VDD(VDD),.Y(g13333),.A(g4743),.B(g11755));
  AND2 AND2_3678(.VSS(VSS),.VDD(VDD),.Y(g33425),.A(g32380),.B(g21466));
  AND2 AND2_3679(.VSS(VSS),.VDD(VDD),.Y(g28213),.A(g27720),.B(g23380));
  AND2 AND2_3680(.VSS(VSS),.VDD(VDD),.Y(g15679),.A(g3470),.B(g13555));
  AND2 AND2_3681(.VSS(VSS),.VDD(VDD),.Y(g18812),.A(g6509),.B(g15483));
  AND2 AND2_3682(.VSS(VSS),.VDD(VDD),.Y(g10948),.A(g7880),.B(g1478));
  AND2 AND2_3683(.VSS(VSS),.VDD(VDD),.Y(g18463),.A(g2375),.B(g15224));
  AND2 AND2_3684(.VSS(VSS),.VDD(VDD),.Y(g33919),.A(g33438),.B(g10795));
  AND2 AND2_3685(.VSS(VSS),.VDD(VDD),.Y(g24406),.A(g13623),.B(g22860));
  AND2 AND2_3686(.VSS(VSS),.VDD(VDD),.Y(g29528),.A(g2429),.B(g28874));
  AND4 AND4_221(.VSS(VSS),.VDD(VDD),.Y(I31036),.A(g30673),.B(g31802),.C(g32506),.D(g32507));
  AND2 AND2_3687(.VSS(VSS),.VDD(VDD),.Y(g24962),.A(g23194),.B(g20210));
  AND2 AND2_3688(.VSS(VSS),.VDD(VDD),.Y(g29843),.A(g28373),.B(g23289));
  AND2 AND2_3689(.VSS(VSS),.VDD(VDD),.Y(g21781),.A(g3408),.B(g20391));
  AND2 AND2_3690(.VSS(VSS),.VDD(VDD),.Y(g29330),.A(g29114),.B(g18894));
  AND2 AND2_3691(.VSS(VSS),.VDD(VDD),.Y(g16617),.A(g6287),.B(g14940));
  AND2 AND2_3692(.VSS(VSS),.VDD(VDD),.Y(g25502),.A(g6946),.B(g22527));
  AND2 AND2_3693(.VSS(VSS),.VDD(VDD),.Y(g15678),.A(g1094),.B(g13846));
  AND4 AND4_222(.VSS(VSS),.VDD(VDD),.Y(I31101),.A(g30735),.B(g31813),.C(g32601),.D(g32602));
  AND4 AND4_223(.VSS(VSS),.VDD(VDD),.Y(I31177),.A(g32710),.B(g32711),.C(g32712),.D(g32713));
  AND2 AND2_3694(.VSS(VSS),.VDD(VDD),.Y(g18951),.A(g3484),.B(g16124));
  AND2 AND2_3695(.VSS(VSS),.VDD(VDD),.Y(g30187),.A(g28643),.B(g23840));
  AND2 AND2_3696(.VSS(VSS),.VDD(VDD),.Y(g18371),.A(g1870),.B(g15171));
  AND3 AND3_209(.VSS(VSS),.VDD(VDD),.Y(g8721),.A(g385),.B(g376),.C(g365));
  AND2 AND2_3697(.VSS(VSS),.VDD(VDD),.Y(g28205),.A(g27516),.B(g16746));
  AND2 AND2_3698(.VSS(VSS),.VDD(VDD),.Y(g18234),.A(g1129),.B(g16326));
  AND2 AND2_3699(.VSS(VSS),.VDD(VDD),.Y(g34187),.A(g33708),.B(g24397));
  AND2 AND2_3700(.VSS(VSS),.VDD(VDD),.Y(g17769),.A(g1146),.B(g13188));
  AND2 AND2_3701(.VSS(VSS),.VDD(VDD),.Y(g21952),.A(g5366),.B(g21514));
  AND2 AND2_3702(.VSS(VSS),.VDD(VDD),.Y(g28311),.A(g9792),.B(g27679));
  AND2 AND2_3703(.VSS(VSS),.VDD(VDD),.Y(g23372),.A(g16448),.B(g20194));
  AND2 AND2_3704(.VSS(VSS),.VDD(VDD),.Y(g29869),.A(g2331),.B(g29129));
  AND2 AND2_3705(.VSS(VSS),.VDD(VDD),.Y(g21821),.A(g3723),.B(g20453));
  AND2 AND2_3706(.VSS(VSS),.VDD(VDD),.Y(g17768),.A(g13325),.B(g10741));
  AND4 AND4_224(.VSS(VSS),.VDD(VDD),.Y(I26530),.A(g26365),.B(g24096),.C(g24097),.D(g24098));
  AND2 AND2_3707(.VSS(VSS),.VDD(VDD),.Y(g18795),.A(g6163),.B(g15348));
  AND2 AND2_3708(.VSS(VSS),.VDD(VDD),.Y(g30937),.A(g22626),.B(g29814));
  AND2 AND2_3709(.VSS(VSS),.VDD(VDD),.Y(g29868),.A(g2227),.B(g29128));
  AND2 AND2_3710(.VSS(VSS),.VDD(VDD),.Y(g27649),.A(g10820),.B(g25820));
  AND2 AND2_3711(.VSS(VSS),.VDD(VDD),.Y(g34143),.A(g33934),.B(g23828));
  AND2 AND2_3712(.VSS(VSS),.VDD(VDD),.Y(g16595),.A(g5921),.B(g14697));
  AND2 AND2_3713(.VSS(VSS),.VDD(VDD),.Y(g21790),.A(g3454),.B(g20391));
  AND2 AND2_3714(.VSS(VSS),.VDD(VDD),.Y(g24004),.A(g37),.B(g21225));
  AND2 AND2_3715(.VSS(VSS),.VDD(VDD),.Y(g33086),.A(g32390),.B(g18887));
  AND2 AND2_3716(.VSS(VSS),.VDD(VDD),.Y(g27648),.A(g25882),.B(g8974));
  AND2 AND2_3717(.VSS(VSS),.VDD(VDD),.Y(g24221),.A(g232),.B(g22594));
  AND2 AND2_3718(.VSS(VSS),.VDD(VDD),.Y(g27491),.A(g26576),.B(g17652));
  AND2 AND2_3719(.VSS(VSS),.VDD(VDD),.Y(g26486),.A(g4423),.B(g24358));
  AND2 AND2_3720(.VSS(VSS),.VDD(VDD),.Y(g18514),.A(g2629),.B(g15509));
  AND2 AND2_3721(.VSS(VSS),.VDD(VDD),.Y(g29709),.A(g2116),.B(g29121));
  AND2 AND2_3722(.VSS(VSS),.VDD(VDD),.Y(g34169),.A(g33804),.B(g31227));
  AND2 AND2_3723(.VSS(VSS),.VDD(VDD),.Y(g21873),.A(g6946),.B(g19801));
  AND2 AND2_3724(.VSS(VSS),.VDD(VDD),.Y(g18507),.A(g2595),.B(g15509));
  AND2 AND2_3725(.VSS(VSS),.VDD(VDD),.Y(g22027),.A(g5889),.B(g19147));
  AND2 AND2_3726(.VSS(VSS),.VDD(VDD),.Y(g23873),.A(g21222),.B(g10815));
  AND2 AND2_3727(.VSS(VSS),.VDD(VDD),.Y(g15875),.A(g3961),.B(g13963));
  AND2 AND2_3728(.VSS(VSS),.VDD(VDD),.Y(g30168),.A(g28623),.B(g23794));
  AND2 AND2_3729(.VSS(VSS),.VDD(VDD),.Y(g29708),.A(g1955),.B(g29082));
  AND2 AND2_3730(.VSS(VSS),.VDD(VDD),.Y(g33817),.A(g33235),.B(g20102));
  AND2 AND2_3731(.VSS(VSS),.VDD(VDD),.Y(g11115),.A(g6133),.B(g9954));
  AND2 AND2_3732(.VSS(VSS),.VDD(VDD),.Y(g33322),.A(g32202),.B(g20450));
  AND2 AND2_3733(.VSS(VSS),.VDD(VDD),.Y(g34410),.A(g34204),.B(g21427));
  AND2 AND2_3734(.VSS(VSS),.VDD(VDD),.Y(g27981),.A(g26751),.B(g23924));
  AND2 AND2_3735(.VSS(VSS),.VDD(VDD),.Y(g25815),.A(g8155),.B(g24603));
  AND2 AND2_3736(.VSS(VSS),.VDD(VDD),.Y(g31125),.A(g29502),.B(g22973));
  AND2 AND2_3737(.VSS(VSS),.VDD(VDD),.Y(g32176),.A(g2779),.B(g31623));
  AND4 AND4_225(.VSS(VSS),.VDD(VDD),.Y(I31166),.A(g30673),.B(g31825),.C(g32694),.D(g32695));
  AND4 AND4_226(.VSS(VSS),.VDD(VDD),.Y(g26223),.A(g24688),.B(g10678),.C(g10658),.D(g8757));
  AND2 AND2_3738(.VSS(VSS),.VDD(VDD),.Y(g31977),.A(g31764),.B(g22179));
  AND3 AND3_210(.VSS(VSS),.VDD(VDD),.Y(g33532),.A(g32974),.B(I31356),.C(I31357));
  AND2 AND2_3739(.VSS(VSS),.VDD(VDD),.Y(g33901),.A(g33317),.B(g20920));
  AND2 AND2_3740(.VSS(VSS),.VDD(VDD),.Y(g34479),.A(g34403),.B(g18905));
  AND2 AND2_3741(.VSS(VSS),.VDD(VDD),.Y(g34666),.A(g34587),.B(g19144));
  AND2 AND2_3742(.VSS(VSS),.VDD(VDD),.Y(g25187),.A(g12296),.B(g23629));
  AND2 AND2_3743(.VSS(VSS),.VDD(VDD),.Y(g18163),.A(g79),.B(g17433));
  AND2 AND2_3744(.VSS(VSS),.VDD(VDD),.Y(g15837),.A(g3255),.B(g14127));
  AND2 AND2_3745(.VSS(VSS),.VDD(VDD),.Y(g32154),.A(g31277),.B(g14184));
  AND2 AND2_3746(.VSS(VSS),.VDD(VDD),.Y(g34363),.A(g34148),.B(g20389));
  AND2 AND2_3747(.VSS(VSS),.VDD(VDD),.Y(g25975),.A(g9434),.B(g24999));
  AND2 AND2_3748(.VSS(VSS),.VDD(VDD),.Y(g34217),.A(g33736),.B(g22876));
  AND2 AND2_3749(.VSS(VSS),.VDD(VDD),.Y(g22710),.A(g19358),.B(g19600));
  AND2 AND2_3750(.VSS(VSS),.VDD(VDD),.Y(g30015),.A(g29040),.B(g10519));
  AND2 AND2_3751(.VSS(VSS),.VDD(VDD),.Y(g21834),.A(g3752),.B(g20453));
  AND2 AND2_3752(.VSS(VSS),.VDD(VDD),.Y(g22003),.A(g5736),.B(g21562));
  AND2 AND2_3753(.VSS(VSS),.VDD(VDD),.Y(g34478),.A(g34402),.B(g18904));
  AND2 AND2_3754(.VSS(VSS),.VDD(VDD),.Y(g28152),.A(g26297),.B(g27279));
  AND2 AND2_3755(.VSS(VSS),.VDD(VDD),.Y(g26084),.A(g24926),.B(g9602));
  AND4 AND4_227(.VSS(VSS),.VDD(VDD),.Y(g28846),.A(g21434),.B(g26424),.C(g25399),.D(g27474));
  AND2 AND2_3756(.VSS(VSS),.VDD(VDD),.Y(g24812),.A(g19662),.B(g22192));
  AND2 AND2_3757(.VSS(VSS),.VDD(VDD),.Y(g19855),.A(g2787),.B(g15962));
  AND2 AND2_3758(.VSS(VSS),.VDD(VDD),.Y(g33353),.A(g32240),.B(g20732));
  AND2 AND2_3759(.VSS(VSS),.VDD(VDD),.Y(g25143),.A(g4922),.B(g22908));
  AND2 AND2_3760(.VSS(VSS),.VDD(VDD),.Y(g34486),.A(g34412),.B(g18953));
  AND2 AND2_3761(.VSS(VSS),.VDD(VDD),.Y(g18541),.A(g2767),.B(g15277));
  AND4 AND4_228(.VSS(VSS),.VDD(VDD),.Y(g27395),.A(g8046),.B(g26314),.C(g9187),.D(g9077));
  AND2 AND2_3762(.VSS(VSS),.VDD(VDD),.Y(g33680),.A(g33128),.B(g4688));
  AND2 AND2_3763(.VSS(VSS),.VDD(VDD),.Y(g18473),.A(g2342),.B(g15224));
  AND2 AND2_3764(.VSS(VSS),.VDD(VDD),.Y(g27262),.A(g25997),.B(g17092));
  AND2 AND2_3765(.VSS(VSS),.VDD(VDD),.Y(g26179),.A(g2504),.B(g25155));
  AND2 AND2_3766(.VSS(VSS),.VDD(VDD),.Y(g12794),.A(g1008),.B(g7567));
  AND3 AND3_211(.VSS(VSS),.VDD(VDD),.Y(I17529),.A(g13156),.B(g11450),.C(g6756));
  AND2 AND2_3767(.VSS(VSS),.VDD(VDD),.Y(g34556),.A(g34350),.B(g20537));
  AND2 AND2_3768(.VSS(VSS),.VDD(VDD),.Y(g18789),.A(g6035),.B(g15634));
  AND2 AND2_3769(.VSS(VSS),.VDD(VDD),.Y(g21453),.A(g16713),.B(g13625));
  AND2 AND2_3770(.VSS(VSS),.VDD(VDD),.Y(g22081),.A(g6279),.B(g19210));
  AND2 AND2_3771(.VSS(VSS),.VDD(VDD),.Y(g29602),.A(g2020),.B(g28962));
  AND2 AND2_3772(.VSS(VSS),.VDD(VDD),.Y(g29810),.A(g28259),.B(g11317));
  AND2 AND2_3773(.VSS(VSS),.VDD(VDD),.Y(g29774),.A(g28287),.B(g10233));
  AND2 AND2_3774(.VSS(VSS),.VDD(VDD),.Y(g34580),.A(g29539),.B(g34311));
  AND2 AND2_3775(.VSS(VSS),.VDD(VDD),.Y(g26178),.A(g2389),.B(g25473));
  AND4 AND4_229(.VSS(VSS),.VDD(VDD),.Y(g16194),.A(g11547),.B(g6782),.C(g11640),.D(I17529));
  AND2 AND2_3776(.VSS(VSS),.VDD(VDD),.Y(g27633),.A(g13076),.B(g25766));
  AND2 AND2_3777(.VSS(VSS),.VDD(VDD),.Y(g21913),.A(g5069),.B(g21468));
  AND2 AND2_3778(.VSS(VSS),.VDD(VDD),.Y(g29375),.A(g13946),.B(g28370));
  AND2 AND2_3779(.VSS(VSS),.VDD(VDD),.Y(g30223),.A(g28702),.B(g23895));
  AND4 AND4_230(.VSS(VSS),.VDD(VDD),.Y(g13805),.A(g11489),.B(g11394),.C(g11356),.D(I16129));
  AND2 AND2_3780(.VSS(VSS),.VDD(VDD),.Y(g18788),.A(g6031),.B(g15634));
  AND2 AND2_3781(.VSS(VSS),.VDD(VDD),.Y(g18724),.A(g4907),.B(g16077));
  AND2 AND2_3782(.VSS(VSS),.VDD(VDD),.Y(g25884),.A(g11153),.B(g24711));
  AND2 AND2_3783(.VSS(VSS),.VDD(VDD),.Y(g18359),.A(g1825),.B(g17955));
  AND2 AND2_3784(.VSS(VSS),.VDD(VDD),.Y(g34223),.A(g33744),.B(g22876));
  AND2 AND2_3785(.VSS(VSS),.VDD(VDD),.Y(g18325),.A(g1624),.B(g17873));
  AND2 AND2_3786(.VSS(VSS),.VDD(VDD),.Y(g26186),.A(g24580),.B(g23031));
  AND2 AND2_3787(.VSS(VSS),.VDD(VDD),.Y(g23436),.A(g676),.B(g20375));
  AND2 AND2_3788(.VSS(VSS),.VDD(VDD),.Y(g18535),.A(g2741),.B(g15277));
  AND2 AND2_3789(.VSS(VSS),.VDD(VDD),.Y(g18434),.A(g2217),.B(g18008));
  AND2 AND2_3790(.VSS(VSS),.VDD(VDD),.Y(g18358),.A(g1811),.B(g17955));
  AND2 AND2_3791(.VSS(VSS),.VDD(VDD),.Y(g31966),.A(g31754),.B(g22166));
  AND2 AND2_3792(.VSS(VSS),.VDD(VDD),.Y(g30084),.A(g28534),.B(g20700));
  AND2 AND2_3793(.VSS(VSS),.VDD(VDD),.Y(g27521),.A(g26519),.B(g14700));
  AND2 AND2_3794(.VSS(VSS),.VDD(VDD),.Y(g29337),.A(g29166),.B(g22180));
  AND2 AND2_3795(.VSS(VSS),.VDD(VDD),.Y(g17786),.A(g1489),.B(g13216));
  AND2 AND2_3796(.VSS(VSS),.VDD(VDD),.Y(g30110),.A(g28564),.B(g20916));
  AND2 AND2_3797(.VSS(VSS),.VDD(VDD),.Y(g25479),.A(g22646),.B(g9917));
  AND2 AND2_3798(.VSS(VSS),.VDD(VDD),.Y(g34084),.A(g9214),.B(g33851));
  AND2 AND2_3799(.VSS(VSS),.VDD(VDD),.Y(g15075),.A(g12850),.B(g12955));
  AND2 AND2_3800(.VSS(VSS),.VDD(VDD),.Y(g31017),.A(g29479),.B(g22841));
  AND2 AND2_3801(.VSS(VSS),.VDD(VDD),.Y(g34110),.A(g33732),.B(g22935));
  AND2 AND2_3802(.VSS(VSS),.VDD(VDD),.Y(g25217),.A(g12418),.B(g23698));
  AND2 AND2_3803(.VSS(VSS),.VDD(VDD),.Y(g33364),.A(g32264),.B(g20921));
  AND2 AND2_3804(.VSS(VSS),.VDD(VDD),.Y(g18121),.A(g424),.B(g17015));
  AND2 AND2_3805(.VSS(VSS),.VDD(VDD),.Y(g22090),.A(g6404),.B(g18833));
  AND2 AND2_3806(.VSS(VSS),.VDD(VDD),.Y(g30179),.A(g28634),.B(g23819));
  AND2 AND2_3807(.VSS(VSS),.VDD(VDD),.Y(g24507),.A(g22304),.B(g19429));
  AND2 AND2_3808(.VSS(VSS),.VDD(VDD),.Y(g18344),.A(g1740),.B(g17955));
  AND3 AND3_212(.VSS(VSS),.VDD(VDD),.Y(g19581),.A(g15843),.B(g1500),.C(g10918));
  AND2 AND2_3809(.VSS(VSS),.VDD(VDD),.Y(g34179),.A(g33686),.B(g24372));
  AND4 AND4_231(.VSS(VSS),.VDD(VDD),.Y(g27440),.A(g8046),.B(g26314),.C(g518),.D(g504));
  AND2 AND2_3810(.VSS(VSS),.VDD(VDD),.Y(g21464),.A(g16181),.B(g10872));
  AND4 AND4_232(.VSS(VSS),.VDD(VDD),.Y(g28020),.A(g23032),.B(g26241),.C(g26424),.D(g25542));
  AND2 AND2_3811(.VSS(VSS),.VDD(VDD),.Y(g28583),.A(g12009),.B(g27112));
  AND2 AND2_3812(.VSS(VSS),.VDD(VDD),.Y(g30178),.A(g28632),.B(g23815));
  AND2 AND2_3813(.VSS(VSS),.VDD(VDD),.Y(g9479),.A(g305),.B(g324));
  AND2 AND2_3814(.VSS(VSS),.VDD(VDD),.Y(g24421),.A(g3835),.B(g23139));
  AND2 AND2_3815(.VSS(VSS),.VDD(VDD),.Y(g34178),.A(g33712),.B(g24361));
  AND2 AND2_3816(.VSS(VSS),.VDD(VDD),.Y(g34740),.A(g34664),.B(g19414));
  AND2 AND2_3817(.VSS(VSS),.VDD(VDD),.Y(g16616),.A(g6267),.B(g14741));
  AND4 AND4_233(.VSS(VSS),.VDD(VDD),.Y(g10756),.A(g3990),.B(g6928),.C(g3976),.D(g8595));
  AND2 AND2_3818(.VSS(VSS),.VDD(VDD),.Y(g18682),.A(g4646),.B(g15885));
  AND4 AND4_234(.VSS(VSS),.VDD(VDD),.Y(I31176),.A(g31579),.B(g31827),.C(g32708),.D(g32709));
  AND2 AND2_3819(.VSS(VSS),.VDD(VDD),.Y(g30186),.A(g28641),.B(g23839));
  AND2 AND2_3820(.VSS(VSS),.VDD(VDD),.Y(g27247),.A(g2759),.B(g26745));
  AND4 AND4_235(.VSS(VSS),.VDD(VDD),.Y(I31092),.A(g32589),.B(g32590),.C(g32591),.D(g32592));
  AND2 AND2_3821(.VSS(VSS),.VDD(VDD),.Y(g18291),.A(g1437),.B(g16449));
  AND2 AND2_3822(.VSS(VSS),.VDD(VDD),.Y(g24012),.A(g14496),.B(g21561));
  AND2 AND2_3823(.VSS(VSS),.VDD(VDD),.Y(g17182),.A(g8579),.B(g13016));
  AND2 AND2_3824(.VSS(VSS),.VDD(VDD),.Y(g21797),.A(g3518),.B(g20924));
  AND2 AND2_3825(.VSS(VSS),.VDD(VDD),.Y(g34186),.A(g33705),.B(g24396));
  AND2 AND2_3826(.VSS(VSS),.VDD(VDD),.Y(g34685),.A(g14164),.B(g34550));
  AND2 AND2_3827(.VSS(VSS),.VDD(VDD),.Y(g25580),.A(g19268),.B(g24149));
  AND2 AND2_3828(.VSS(VSS),.VDD(VDD),.Y(g18173),.A(g736),.B(g17328));
  AND2 AND2_3829(.VSS(VSS),.VDD(VDD),.Y(g27389),.A(g26519),.B(g17503));
  AND2 AND2_3830(.VSS(VSS),.VDD(VDD),.Y(g34953),.A(g34935),.B(g19957));
  AND4 AND4_236(.VSS(VSS),.VDD(VDD),.Y(g27045),.A(g10295),.B(g3171),.C(g3179),.D(g26244));
  AND2 AND2_3831(.VSS(VSS),.VDD(VDD),.Y(g31309),.A(g30132),.B(g27837));
  AND4 AND4_237(.VSS(VSS),.VDD(VDD),.Y(I24699),.A(g21127),.B(g24054),.C(g24055),.D(g24056));
  AND2 AND2_3832(.VSS(VSS),.VDD(VDD),.Y(g32083),.A(g947),.B(g30735));
  AND2 AND2_3833(.VSS(VSS),.VDD(VDD),.Y(g32348),.A(g2145),.B(g31672));
  AND2 AND2_3834(.VSS(VSS),.VDD(VDD),.Y(g23292),.A(g19879),.B(g16726));
  AND2 AND2_3835(.VSS(VSS),.VDD(VDD),.Y(g25223),.A(g22523),.B(g10652));
  AND2 AND2_3836(.VSS(VSS),.VDD(VDD),.Y(g16704),.A(g5957),.B(g15018));
  AND2 AND2_3837(.VSS(VSS),.VDD(VDD),.Y(g27612),.A(g25887),.B(g8844));
  AND2 AND2_3838(.VSS(VSS),.VDD(VDD),.Y(g31224),.A(g30280),.B(g23932));
  AND2 AND2_3839(.VSS(VSS),.VDD(VDD),.Y(g32284),.A(g31260),.B(g20507));
  AND2 AND2_3840(.VSS(VSS),.VDD(VDD),.Y(g28113),.A(g8016),.B(g27242));
  AND2 AND2_3841(.VSS(VSS),.VDD(VDD),.Y(g26423),.A(g19488),.B(g24356));
  AND2 AND2_3842(.VSS(VSS),.VDD(VDD),.Y(g27099),.A(g14094),.B(g26352));
  AND2 AND2_3843(.VSS(VSS),.VDD(VDD),.Y(g15822),.A(g3925),.B(g13960));
  AND2 AND2_3844(.VSS(VSS),.VDD(VDD),.Y(g27388),.A(g26519),.B(g17502));
  AND2 AND2_3845(.VSS(VSS),.VDD(VDD),.Y(g27324),.A(g10150),.B(g26720));
  AND2 AND2_3846(.VSS(VSS),.VDD(VDD),.Y(g24541),.A(g22626),.B(g10851));
  AND2 AND2_3847(.VSS(VSS),.VDD(VDD),.Y(g32304),.A(g31284),.B(g20564));
  AND2 AND2_3848(.VSS(VSS),.VDD(VDD),.Y(g30936),.A(g8830),.B(g29916));
  AND2 AND2_3849(.VSS(VSS),.VDD(VDD),.Y(g28282),.A(g23762),.B(g27727));
  AND2 AND2_3850(.VSS(VSS),.VDD(VDD),.Y(g12099),.A(g9619),.B(g9888));
  AND2 AND2_3851(.VSS(VSS),.VDD(VDD),.Y(g27534),.A(g26488),.B(g17735));
  AND2 AND2_3852(.VSS(VSS),.VDD(VDD),.Y(g27098),.A(g25868),.B(g22528));
  AND2 AND2_3853(.VSS(VSS),.VDD(VDD),.Y(g28302),.A(g23809),.B(g27817));
  AND2 AND2_3854(.VSS(VSS),.VDD(VDD),.Y(g25084),.A(g4737),.B(g22885));
  AND2 AND2_3855(.VSS(VSS),.VDD(VDD),.Y(g27251),.A(g26721),.B(g26694));
  AND2 AND2_3856(.VSS(VSS),.VDD(VDD),.Y(g27272),.A(g26055),.B(g17144));
  AND2 AND2_3857(.VSS(VSS),.VDD(VDD),.Y(g25110),.A(g10427),.B(g23509));
  AND2 AND2_3858(.VSS(VSS),.VDD(VDD),.Y(g16808),.A(g6653),.B(g14825));
  AND2 AND2_3859(.VSS(VSS),.VDD(VDD),.Y(g19384),.A(g667),.B(g16310));
  AND2 AND2_3860(.VSS(VSS),.VDD(VDD),.Y(g18760),.A(g5462),.B(g17929));
  AND2 AND2_3861(.VSS(VSS),.VDD(VDD),.Y(g18134),.A(g534),.B(g17249));
  AND2 AND2_3862(.VSS(VSS),.VDD(VDD),.Y(g25922),.A(g24959),.B(g20065));
  AND2 AND2_3863(.VSS(VSS),.VDD(VDD),.Y(g34334),.A(g34090),.B(g19865));
  AND2 AND2_3864(.VSS(VSS),.VDD(VDD),.Y(g24788),.A(g11384),.B(g23111));
  AND2 AND2_3865(.VSS(VSS),.VDD(VDD),.Y(g31495),.A(g1913),.B(g30309));
  AND2 AND2_3866(.VSS(VSS),.VDD(VDD),.Y(g24724),.A(g17624),.B(g22432));
  AND2 AND2_3867(.VSS(VSS),.VDD(VDD),.Y(g29599),.A(g1710),.B(g29018));
  AND3 AND3_213(.VSS(VSS),.VDD(VDD),.Y(g33495),.A(g32707),.B(I31171),.C(I31172));
  AND2 AND2_3868(.VSS(VSS),.VDD(VDD),.Y(g22717),.A(g9291),.B(g20212));
  AND2 AND2_3869(.VSS(VSS),.VDD(VDD),.Y(g16177),.A(g5128),.B(g14238));
  AND2 AND2_3870(.VSS(VSS),.VDD(VDD),.Y(g24325),.A(g4543),.B(g22228));
  AND2 AND2_3871(.VSS(VSS),.VDD(VDD),.Y(g25179),.A(g16928),.B(g23611));
  AND2 AND2_3872(.VSS(VSS),.VDD(VDD),.Y(g26543),.A(g12910),.B(g24377));
  AND4 AND4_238(.VSS(VSS),.VDD(VDD),.Y(I27503),.A(g19890),.B(g24075),.C(g24076),.D(g28032));
  AND2 AND2_3873(.VSS(VSS),.VDD(VDD),.Y(g18506),.A(g2571),.B(g15509));
  AND2 AND2_3874(.VSS(VSS),.VDD(VDD),.Y(g22026),.A(g5913),.B(g19147));
  AND2 AND2_3875(.VSS(VSS),.VDD(VDD),.Y(g27462),.A(g26576),.B(g17612));
  AND2 AND2_3876(.VSS(VSS),.VDD(VDD),.Y(g33816),.A(g33234),.B(g20096));
  AND2 AND2_3877(.VSS(VSS),.VDD(VDD),.Y(g29598),.A(g28823),.B(g22342));
  AND2 AND2_3878(.VSS(VSS),.VDD(VDD),.Y(g16642),.A(g6633),.B(g14981));
  AND2 AND2_3879(.VSS(VSS),.VDD(VDD),.Y(g25178),.A(g20241),.B(g23608));
  AND2 AND2_3880(.VSS(VSS),.VDD(VDD),.Y(g15589),.A(g411),.B(g13334));
  AND2 AND2_3881(.VSS(VSS),.VDD(VDD),.Y(g32139),.A(g31601),.B(g29960));
  AND4 AND4_239(.VSS(VSS),.VDD(VDD),.Y(g27032),.A(g7704),.B(g5180),.C(g5188),.D(g26200));
  AND2 AND2_3882(.VSS(VSS),.VDD(VDD),.Y(g34964),.A(g34947),.B(g23060));
  AND2 AND2_3883(.VSS(VSS),.VDD(VDD),.Y(g33687),.A(g33132),.B(g4878));
  AND2 AND2_3884(.VSS(VSS),.VDD(VDD),.Y(g31976),.A(g31762),.B(g22178));
  AND2 AND2_3885(.VSS(VSS),.VDD(VDD),.Y(g31985),.A(g4722),.B(g30614));
  AND2 AND2_3886(.VSS(VSS),.VDD(VDD),.Y(g19735),.A(g9740),.B(g17135));
  AND2 AND2_3887(.VSS(VSS),.VDD(VDD),.Y(g27140),.A(g25885),.B(g22593));
  AND2 AND2_3888(.VSS(VSS),.VDD(VDD),.Y(g30216),.A(g28691),.B(g23882));
  AND2 AND2_3889(.VSS(VSS),.VDD(VDD),.Y(g27997),.A(g26813),.B(g23995));
  AND4 AND4_240(.VSS(VSS),.VDD(VDD),.Y(g28768),.A(g21434),.B(g26424),.C(g25308),.D(g27421));
  AND2 AND2_3890(.VSS(VSS),.VDD(VDD),.Y(g15836),.A(g3187),.B(g14104));
  AND2 AND2_3891(.VSS(VSS),.VDD(VDD),.Y(g31752),.A(g30104),.B(g23928));
  AND2 AND2_3892(.VSS(VSS),.VDD(VDD),.Y(g34216),.A(g33778),.B(g22689));
  AND2 AND2_3893(.VSS(VSS),.VDD(VDD),.Y(g31374),.A(g29748),.B(g23390));
  AND3 AND3_214(.VSS(VSS),.VDD(VDD),.Y(g29322),.A(g29192),.B(g7074),.C(g6336));
  AND2 AND2_3894(.VSS(VSS),.VDD(VDD),.Y(g33374),.A(g32289),.B(g21221));
  AND2 AND2_3895(.VSS(VSS),.VDD(VDD),.Y(g16733),.A(g5893),.B(g14889));
  AND3 AND3_215(.VSS(VSS),.VDD(VDD),.Y(I18671),.A(g13156),.B(g11450),.C(g6756));
  AND2 AND2_3896(.VSS(VSS),.VDD(VDD),.Y(g29532),.A(g1878),.B(g28861));
  AND2 AND2_3897(.VSS(VSS),.VDD(VDD),.Y(g29901),.A(g28429),.B(g23376));
  AND2 AND2_3898(.VSS(VSS),.VDD(VDD),.Y(g32333),.A(g31326),.B(g23559));
  AND2 AND2_3899(.VSS(VSS),.VDD(VDD),.Y(g15119),.A(g4249),.B(g14454));
  AND2 AND2_3900(.VSS(VSS),.VDD(VDD),.Y(g20682),.A(g16238),.B(g4646));
  AND4 AND4_241(.VSS(VSS),.VDD(VDD),.Y(g13771),.A(g11441),.B(g11355),.C(g11302),.D(I16111));
  AND3 AND3_216(.VSS(VSS),.VDD(VDD),.Y(g25417),.A(g5712),.B(g23816),.C(I24552));
  AND2 AND2_3901(.VSS(VSS),.VDD(VDD),.Y(g23474),.A(g13830),.B(g20533));
  AND2 AND2_3902(.VSS(VSS),.VDD(VDD),.Y(g24682),.A(g22662),.B(g19754));
  AND2 AND2_3903(.VSS(VSS),.VDD(VDD),.Y(g22149),.A(g14581),.B(g18880));
  AND2 AND2_3904(.VSS(VSS),.VDD(VDD),.Y(g29783),.A(g28329),.B(g23246));
  AND2 AND2_3905(.VSS(VSS),.VDD(VDD),.Y(g21711),.A(g291),.B(g20283));
  AND2 AND2_3906(.VSS(VSS),.VDD(VDD),.Y(g26123),.A(g1696),.B(g25382));
  AND2 AND2_3907(.VSS(VSS),.VDD(VDD),.Y(g15118),.A(g4253),.B(g14454));
  AND2 AND2_3908(.VSS(VSS),.VDD(VDD),.Y(g34909),.A(g34856),.B(g20130));
  AND2 AND2_3909(.VSS(VSS),.VDD(VDD),.Y(g24291),.A(g18660),.B(g22550));
  AND2 AND2_3910(.VSS(VSS),.VDD(VDD),.Y(g30000),.A(g23685),.B(g29029));
  AND2 AND2_3911(.VSS(VSS),.VDD(VDD),.Y(g29656),.A(g28515),.B(g11666));
  AND2 AND2_3912(.VSS(VSS),.VDD(VDD),.Y(g34117),.A(g33742),.B(g19755));
  AND2 AND2_3913(.VSS(VSS),.VDD(VDD),.Y(g15749),.A(g1454),.B(g13273));
  AND2 AND2_3914(.VSS(VSS),.VDD(VDD),.Y(g18649),.A(g4049),.B(g17271));
  AND2 AND2_3915(.VSS(VSS),.VDD(VDD),.Y(g22097),.A(g6451),.B(g18833));
  AND2 AND2_3916(.VSS(VSS),.VDD(VDD),.Y(g27360),.A(g26488),.B(g17417));
  AND2 AND2_3917(.VSS(VSS),.VDD(VDD),.Y(g33842),.A(g33255),.B(g20322));
  AND2 AND2_3918(.VSS(VSS),.VDD(VDD),.Y(g18240),.A(g15066),.B(g16431));
  AND2 AND2_3919(.VSS(VSS),.VDD(VDD),.Y(g22104),.A(g6444),.B(g18833));
  AND2 AND2_3920(.VSS(VSS),.VDD(VDD),.Y(g17149),.A(g232),.B(g13255));
  AND2 AND2_3921(.VSS(VSS),.VDD(VDD),.Y(g33392),.A(g32344),.B(g21362));
  AND2 AND2_3922(.VSS(VSS),.VDD(VDD),.Y(g18648),.A(g4045),.B(g17271));
  AND2 AND2_3923(.VSS(VSS),.VDD(VDD),.Y(g18491),.A(g2518),.B(g15426));
  AND2 AND2_3924(.VSS(VSS),.VDD(VDD),.Y(g31489),.A(g2204),.B(g30305));
  AND2 AND2_3925(.VSS(VSS),.VDD(VDD),.Y(g26230),.A(g1768),.B(g25385));
  AND2 AND2_3926(.VSS(VSS),.VDD(VDD),.Y(g25964),.A(g1783),.B(g24979));
  AND3 AND3_217(.VSS(VSS),.VDD(VDD),.Y(g33489),.A(g32665),.B(I31141),.C(I31142));
  AND2 AND2_3927(.VSS(VSS),.VDD(VDD),.Y(g21606),.A(g15959),.B(g13763));
  AND3 AND3_218(.VSS(VSS),.VDD(VDD),.Y(g27162),.A(g26171),.B(g8259),.C(g2208));
  AND2 AND2_3928(.VSS(VSS),.VDD(VDD),.Y(g34568),.A(g34379),.B(g17512));
  AND2 AND2_3929(.VSS(VSS),.VDD(VDD),.Y(g34747),.A(g34671),.B(g19527));
  AND2 AND2_3930(.VSS(VSS),.VDD(VDD),.Y(g23606),.A(g16927),.B(g20679));
  AND2 AND2_3931(.VSS(VSS),.VDD(VDD),.Y(g29336),.A(g4704),.B(g28363));
  AND2 AND2_3932(.VSS(VSS),.VDD(VDD),.Y(g15704),.A(g3440),.B(g13504));
  AND2 AND2_3933(.VSS(VSS),.VDD(VDD),.Y(g30242),.A(g28730),.B(g23927));
  AND2 AND2_3934(.VSS(VSS),.VDD(VDD),.Y(g18604),.A(g3125),.B(g16987));
  AND2 AND2_3935(.VSS(VSS),.VDD(VDD),.Y(g21303),.A(g10120),.B(g17625));
  AND2 AND2_3936(.VSS(VSS),.VDD(VDD),.Y(g16485),.A(g5563),.B(g14924));
  AND2 AND2_3937(.VSS(VSS),.VDD(VDD),.Y(g18755),.A(g5343),.B(g15595));
  AND2 AND2_3938(.VSS(VSS),.VDD(VDD),.Y(g31525),.A(g29892),.B(g23526));
  AND2 AND2_3939(.VSS(VSS),.VDD(VDD),.Y(g31488),.A(g1779),.B(g30302));
  AND2 AND2_3940(.VSS(VSS),.VDD(VDD),.Y(g31016),.A(g29478),.B(g22840));
  AND3 AND3_219(.VSS(VSS),.VDD(VDD),.Y(g33525),.A(g32925),.B(I31321),.C(I31322));
  AND3 AND3_220(.VSS(VSS),.VDD(VDD),.Y(g33488),.A(g32658),.B(I31136),.C(I31137));
  AND2 AND2_3941(.VSS(VSS),.VDD(VDD),.Y(g28249),.A(g27152),.B(g19677));
  AND2 AND2_3942(.VSS(VSS),.VDD(VDD),.Y(g15809),.A(g3917),.B(g14154));
  AND2 AND2_3943(.VSS(VSS),.VDD(VDD),.Y(g18770),.A(g15153),.B(g15615));
  AND3 AND3_221(.VSS(VSS),.VDD(VDD),.Y(g22369),.A(g9354),.B(g7717),.C(g20783));
  AND2 AND2_3944(.VSS(VSS),.VDD(VDD),.Y(g18563),.A(g2890),.B(g16349));
  AND2 AND2_3945(.VSS(VSS),.VDD(VDD),.Y(g18981),.A(g11206),.B(g16158));
  AND2 AND2_3946(.VSS(VSS),.VDD(VDD),.Y(g21750),.A(g3161),.B(g20785));
  AND2 AND2_3947(.VSS(VSS),.VDD(VDD),.Y(g28248),.A(g27150),.B(g19676));
  AND2 AND2_3948(.VSS(VSS),.VDD(VDD),.Y(g29966),.A(g23617),.B(g28970));
  AND2 AND2_3949(.VSS(VSS),.VDD(VDD),.Y(g28710),.A(g27589),.B(g20703));
  AND2 AND2_3950(.VSS(VSS),.VDD(VDD),.Y(g15808),.A(g3590),.B(g14048));
  AND2 AND2_3951(.VSS(VSS),.VDD(VDD),.Y(g21982),.A(g5547),.B(g19074));
  AND2 AND2_3952(.VSS(VSS),.VDD(VDD),.Y(g27451),.A(g26400),.B(g17599));
  AND2 AND2_3953(.VSS(VSS),.VDD(VDD),.Y(g26391),.A(g19593),.B(g25555));
  AND3 AND3_222(.VSS(VSS),.VDD(VDD),.Y(I26948),.A(g24981),.B(g26424),.C(g22698));
  AND2 AND2_3954(.VSS(VSS),.VDD(VDD),.Y(g23381),.A(g7239),.B(g21413));
  AND2 AND2_3955(.VSS(VSS),.VDD(VDD),.Y(g27220),.A(g26026),.B(g16743));
  AND2 AND2_3956(.VSS(VSS),.VDD(VDD),.Y(g33830),.A(g33382),.B(g20166));
  AND2 AND2_3957(.VSS(VSS),.VDD(VDD),.Y(g29631),.A(g1682),.B(g28656));
  AND2 AND2_3958(.VSS(VSS),.VDD(VDD),.Y(g32312),.A(g31302),.B(g20591));
  AND2 AND2_3959(.VSS(VSS),.VDD(VDD),.Y(g32200),.A(g27468),.B(g31376));
  AND2 AND2_3960(.VSS(VSS),.VDD(VDD),.Y(g33893),.A(g33313),.B(g20706));
  AND2 AND2_3961(.VSS(VSS),.VDD(VDD),.Y(g28204),.A(g26098),.B(g27654));
  AND2 AND2_3962(.VSS(VSS),.VDD(VDD),.Y(g27628),.A(g26400),.B(g18061));
  AND2 AND2_3963(.VSS(VSS),.VDD(VDD),.Y(g34751),.A(g34674),.B(g19543));
  AND2 AND2_3964(.VSS(VSS),.VDD(VDD),.Y(g29364),.A(g27400),.B(g28321));
  AND2 AND2_3965(.VSS(VSS),.VDD(VDD),.Y(g10827),.A(g8914),.B(g4258));
  AND2 AND2_3966(.VSS(VSS),.VDD(VDD),.Y(g25909),.A(g8745),.B(g24875));
  AND2 AND2_3967(.VSS(VSS),.VDD(VDD),.Y(g32115),.A(g31631),.B(g29928));
  AND2 AND2_3968(.VSS(VSS),.VDD(VDD),.Y(g25543),.A(g23795),.B(g21461));
  AND2 AND2_3969(.VSS(VSS),.VDD(VDD),.Y(g12220),.A(g1521),.B(g7535));
  AND2 AND2_3970(.VSS(VSS),.VDD(VDD),.Y(g27246),.A(g26690),.B(g26673));
  AND2 AND2_3971(.VSS(VSS),.VDD(VDD),.Y(g33865),.A(g33275),.B(g20526));
  AND2 AND2_3972(.VSS(VSS),.VDD(VDD),.Y(g21796),.A(g3512),.B(g20924));
  AND2 AND2_3973(.VSS(VSS),.VDD(VDD),.Y(g30230),.A(g28717),.B(g23906));
  AND2 AND2_3974(.VSS(VSS),.VDD(VDD),.Y(g25908),.A(g24782),.B(g22520));
  AND2 AND2_3975(.VSS(VSS),.VDD(VDD),.Y(g18767),.A(g15150),.B(g17929));
  AND2 AND2_3976(.VSS(VSS),.VDD(VDD),.Y(g18794),.A(g6154),.B(g15348));
  AND2 AND2_3977(.VSS(VSS),.VDD(VDD),.Y(g34230),.A(g33761),.B(g22942));
  AND2 AND2_3978(.VSS(VSS),.VDD(VDD),.Y(g18395),.A(g12849),.B(g15373));
  AND2 AND2_3979(.VSS(VSS),.VDD(VDD),.Y(g32052),.A(g31507),.B(g13885));
  AND2 AND2_3980(.VSS(VSS),.VDD(VDD),.Y(g18262),.A(g1259),.B(g16000));
  AND2 AND2_3981(.VSS(VSS),.VDD(VDD),.Y(g22133),.A(g6649),.B(g19277));
  AND2 AND2_3982(.VSS(VSS),.VDD(VDD),.Y(g25569),.A(I24684),.B(I24685));
  AND2 AND2_3983(.VSS(VSS),.VDD(VDD),.Y(g21840),.A(g15099),.B(g21070));
  AND2 AND2_3984(.VSS(VSS),.VDD(VDD),.Y(g25568),.A(I24679),.B(I24680));
  AND2 AND2_3985(.VSS(VSS),.VDD(VDD),.Y(g18633),.A(g6905),.B(g17226));
  AND2 AND2_3986(.VSS(VSS),.VDD(VDD),.Y(g17133),.A(g10683),.B(g13222));
  AND2 AND2_3987(.VSS(VSS),.VDD(VDD),.Y(g34841),.A(g34761),.B(g20080));
  AND2 AND2_3988(.VSS(VSS),.VDD(VDD),.Y(g18191),.A(g827),.B(g17821));
  AND2 AND2_3989(.VSS(VSS),.VDD(VDD),.Y(g18719),.A(g4894),.B(g16795));
  AND2 AND2_3990(.VSS(VSS),.VDD(VDD),.Y(g22011),.A(g15154),.B(g21562));
  AND2 AND2_3991(.VSS(VSS),.VDD(VDD),.Y(g15874),.A(g3893),.B(g14079));
  AND2 AND2_3992(.VSS(VSS),.VDD(VDD),.Y(g24649),.A(g6527),.B(g23733));
  AND2 AND2_3993(.VSS(VSS),.VDD(VDD),.Y(g29571),.A(g28452),.B(g11762));
  AND2 AND2_3994(.VSS(VSS),.VDD(VDD),.Y(g11114),.A(g5689),.B(g10160));
  AND2 AND2_3995(.VSS(VSS),.VDD(VDD),.Y(g31270),.A(g29692),.B(g23282));
  AND2 AND2_3996(.VSS(VSS),.VDD(VDD),.Y(g16519),.A(g5591),.B(g14804));
  AND2 AND2_3997(.VSS(VSS),.VDD(VDD),.Y(g16176),.A(g14596),.B(g11779));
  AND2 AND2_3998(.VSS(VSS),.VDD(VDD),.Y(g16185),.A(g3263),.B(g14011));
  AND2 AND2_3999(.VSS(VSS),.VDD(VDD),.Y(g25123),.A(g4732),.B(g22885));
  AND2 AND2_4000(.VSS(VSS),.VDD(VDD),.Y(g18718),.A(g4854),.B(g15915));
  AND2 AND2_4001(.VSS(VSS),.VDD(VDD),.Y(g15693),.A(g269),.B(g13474));
  AND2 AND2_4002(.VSS(VSS),.VDD(VDD),.Y(g18521),.A(g2667),.B(g15509));
  AND2 AND2_4003(.VSS(VSS),.VDD(VDD),.Y(g31188),.A(g20028),.B(g29653));
  AND2 AND2_4004(.VSS(VSS),.VDD(VDD),.Y(g25814),.A(g24760),.B(g13323));
  AND2 AND2_4005(.VSS(VSS),.VDD(VDD),.Y(g27370),.A(g26400),.B(g17472));
  AND2 AND2_4006(.VSS(VSS),.VDD(VDD),.Y(g31124),.A(g2259),.B(g29997));
  AND2 AND2_4007(.VSS(VSS),.VDD(VDD),.Y(g32184),.A(g30611),.B(g25249));
  AND4 AND4_242(.VSS(VSS),.VDD(VDD),.Y(g28998),.A(g17424),.B(g25212),.C(g26424),.D(g27474));
  AND2 AND2_4008(.VSS(VSS),.VDD(VDD),.Y(g33124),.A(g8945),.B(g32296));
  AND3 AND3_223(.VSS(VSS),.VDD(VDD),.Y(g33678),.A(g33149),.B(g10710),.C(g22319));
  AND2 AND2_4009(.VSS(VSS),.VDD(VDD),.Y(g24491),.A(g10727),.B(g22332));
  AND2 AND2_4010(.VSS(VSS),.VDD(VDD),.Y(g24903),.A(g128),.B(g23889));
  AND2 AND2_4011(.VSS(VSS),.VDD(VDD),.Y(g28233),.A(g27827),.B(g23411));
  AND2 AND2_4012(.VSS(VSS),.VDD(VDD),.Y(g16518),.A(g5571),.B(g14956));
  AND2 AND2_4013(.VSS(VSS),.VDD(VDD),.Y(g28182),.A(g8770),.B(g27349));
  AND2 AND2_4014(.VSS(VSS),.VDD(VDD),.Y(g25772),.A(g24944),.B(g24934));
  AND2 AND2_4015(.VSS(VSS),.VDD(VDD),.Y(g28672),.A(g7577),.B(g27017));
  AND2 AND2_4016(.VSS(VSS),.VDD(VDD),.Y(g24755),.A(g16022),.B(g23030));
  AND2 AND2_4017(.VSS(VSS),.VDD(VDD),.Y(g27151),.A(g26026),.B(g16626));
  AND2 AND2_4018(.VSS(VSS),.VDD(VDD),.Y(g34578),.A(g24578),.B(g34308));
  AND2 AND2_4019(.VSS(VSS),.VDD(VDD),.Y(g16637),.A(g5949),.B(g14968));
  AND2 AND2_4020(.VSS(VSS),.VDD(VDD),.Y(g22310),.A(g19662),.B(g20235));
  AND2 AND2_4021(.VSS(VSS),.VDD(VDD),.Y(g18440),.A(g2255),.B(g18008));
  AND2 AND2_4022(.VSS(VSS),.VDD(VDD),.Y(g13345),.A(g4754),.B(g11773));
  AND2 AND2_4023(.VSS(VSS),.VDD(VDD),.Y(g26275),.A(g2417),.B(g25349));
  AND2 AND2_4024(.VSS(VSS),.VDD(VDD),.Y(g30007),.A(g29141),.B(g12929));
  AND3 AND3_224(.VSS(VSS),.VDD(VDD),.Y(I24546),.A(g5046),.B(g5052),.C(g9716));
  AND2 AND2_4025(.VSS(VSS),.VDD(VDD),.Y(g34586),.A(g11025),.B(g34317));
  AND2 AND2_4026(.VSS(VSS),.VDD(VDD),.Y(g18573),.A(g2898),.B(g16349));
  AND2 AND2_4027(.VSS(VSS),.VDD(VDD),.Y(g29687),.A(g2407),.B(g29097));
  AND2 AND2_4028(.VSS(VSS),.VDD(VDD),.Y(g22112),.A(g6555),.B(g19277));
  AND2 AND2_4029(.VSS(VSS),.VDD(VDD),.Y(g18247),.A(g1178),.B(g16431));
  AND2 AND2_4030(.VSS(VSS),.VDD(VDD),.Y(g29985),.A(g28127),.B(g20532));
  AND2 AND2_4031(.VSS(VSS),.VDD(VDD),.Y(g10890),.A(g7858),.B(g1105));
  AND2 AND2_4032(.VSS(VSS),.VDD(VDD),.Y(g21862),.A(g3953),.B(g21070));
  AND2 AND2_4033(.VSS(VSS),.VDD(VDD),.Y(g22050),.A(g6088),.B(g21611));
  AND2 AND2_4034(.VSS(VSS),.VDD(VDD),.Y(g23553),.A(g19413),.B(g11875));
  AND2 AND2_4035(.VSS(VSS),.VDD(VDD),.Y(g18389),.A(g1974),.B(g15171));
  AND2 AND2_4036(.VSS(VSS),.VDD(VDD),.Y(g29752),.A(g28516),.B(g10233));
  AND4 AND4_243(.VSS(VSS),.VDD(VDD),.Y(I31312),.A(g32905),.B(g32906),.C(g32907),.D(g32908));
  AND2 AND2_4037(.VSS(VSS),.VDD(VDD),.Y(g29954),.A(g2299),.B(g28796));
  AND2 AND2_4038(.VSS(VSS),.VDD(VDD),.Y(g21949),.A(g5264),.B(g18997));
  AND2 AND2_4039(.VSS(VSS),.VDD(VDD),.Y(g15712),.A(g3791),.B(g13521));
  AND2 AND2_4040(.VSS(VSS),.VDD(VDD),.Y(g18612),.A(g3329),.B(g17200));
  AND2 AND2_4041(.VSS(VSS),.VDD(VDD),.Y(g15914),.A(g3905),.B(g14024));
  AND2 AND2_4042(.VSS(VSS),.VDD(VDD),.Y(g25992),.A(g2485),.B(g25024));
  AND2 AND2_4043(.VSS(VSS),.VDD(VDD),.Y(g18388),.A(g1968),.B(g15171));
  AND2 AND2_4044(.VSS(VSS),.VDD(VDD),.Y(g19660),.A(g12001),.B(g16968));
  AND2 AND2_4045(.VSS(VSS),.VDD(VDD),.Y(g18324),.A(g1644),.B(g17873));
  AND2 AND2_4046(.VSS(VSS),.VDD(VDD),.Y(g24794),.A(g11414),.B(g23138));
  AND2 AND2_4047(.VSS(VSS),.VDD(VDD),.Y(g31219),.A(g30265),.B(g20875));
  AND2 AND2_4048(.VSS(VSS),.VDD(VDD),.Y(g34116),.A(g33933),.B(g25140));
  AND2 AND2_4049(.VSS(VSS),.VDD(VDD),.Y(g24395),.A(g4704),.B(g22845));
  AND3 AND3_225(.VSS(VSS),.VDD(VDD),.Y(g25510),.A(g6444),.B(g22300),.C(I24619));
  AND2 AND2_4050(.VSS(VSS),.VDD(VDD),.Y(g18701),.A(g4771),.B(g16856));
  AND2 AND2_4051(.VSS(VSS),.VDD(VDD),.Y(g26684),.A(g25407),.B(g20673));
  AND2 AND2_4052(.VSS(VSS),.VDD(VDD),.Y(g21948),.A(g5260),.B(g18997));
  AND2 AND2_4053(.VSS(VSS),.VDD(VDD),.Y(g22096),.A(g6434),.B(g18833));
  AND2 AND2_4054(.VSS(VSS),.VDD(VDD),.Y(g32400),.A(g4743),.B(g30989));
  AND2 AND2_4055(.VSS(VSS),.VDD(VDD),.Y(g18777),.A(g5808),.B(g18065));
  AND2 AND2_4056(.VSS(VSS),.VDD(VDD),.Y(g18534),.A(g2735),.B(g15277));
  AND4 AND4_244(.VSS(VSS),.VDD(VDD),.Y(I14198),.A(g225),.B(g8237),.C(g232),.D(g8180));
  AND2 AND2_4057(.VSS(VSS),.VDD(VDD),.Y(g32013),.A(g8673),.B(g30614));
  AND2 AND2_4058(.VSS(VSS),.VDD(VDD),.Y(g30041),.A(g28511),.B(g23518));
  AND4 AND4_245(.VSS(VSS),.VDD(VDD),.Y(I31052),.A(g32531),.B(g32532),.C(g32533),.D(g32534));
  AND2 AND2_4059(.VSS(VSS),.VDD(VDD),.Y(g18251),.A(g996),.B(g16897));
  AND2 AND2_4060(.VSS(VSS),.VDD(VDD),.Y(g21702),.A(g157),.B(g20283));
  AND2 AND2_4061(.VSS(VSS),.VDD(VDD),.Y(g31218),.A(g30271),.B(g23909));
  AND2 AND2_4062(.VSS(VSS),.VDD(VDD),.Y(g16729),.A(g5240),.B(g14720));
  AND2 AND2_4063(.VSS(VSS),.VDD(VDD),.Y(g18272),.A(g1283),.B(g16031));
  AND2 AND2_4064(.VSS(VSS),.VDD(VDD),.Y(g21757),.A(g3187),.B(g20785));
  AND2 AND2_4065(.VSS(VSS),.VDD(VDD),.Y(g25579),.A(g19422),.B(g24147));
  AND2 AND2_4066(.VSS(VSS),.VDD(VDD),.Y(g30275),.A(g28816),.B(g23984));
  AND4 AND4_246(.VSS(VSS),.VDD(VDD),.Y(I24700),.A(g24057),.B(g24058),.C(g24059),.D(g24060));
  AND2 AND2_4067(.VSS(VSS),.VDD(VDD),.Y(g27227),.A(g26026),.B(g16771));
  AND2 AND2_4068(.VSS(VSS),.VDD(VDD),.Y(g33837),.A(g33251),.B(g20233));
  AND3 AND3_226(.VSS(VSS),.VDD(VDD),.Y(I24625),.A(g6428),.B(g6434),.C(g10014));
  AND2 AND2_4069(.VSS(VSS),.VDD(VDD),.Y(g32207),.A(g31221),.B(g23323));
  AND2 AND2_4070(.VSS(VSS),.VDD(VDD),.Y(g26517),.A(g15708),.B(g24367));
  AND2 AND2_4071(.VSS(VSS),.VDD(VDD),.Y(g34746),.A(g34670),.B(g19526));
  AND2 AND2_4072(.VSS(VSS),.VDD(VDD),.Y(g34493),.A(g34273),.B(g19360));
  AND2 AND2_4073(.VSS(VSS),.VDD(VDD),.Y(g25578),.A(g19402),.B(g24146));
  AND2 AND2_4074(.VSS(VSS),.VDD(VDD),.Y(g15567),.A(g392),.B(g13312));
  AND2 AND2_4075(.VSS(VSS),.VDD(VDD),.Y(g27025),.A(g26334),.B(g7917));
  AND2 AND2_4076(.VSS(VSS),.VDD(VDD),.Y(g24191),.A(g319),.B(g22722));
  AND2 AND2_4077(.VSS(VSS),.VDD(VDD),.Y(g24719),.A(g681),.B(g23530));
  AND2 AND2_4078(.VSS(VSS),.VDD(VDD),.Y(g18462),.A(g2361),.B(g15224));
  AND2 AND2_4079(.VSS(VSS),.VDD(VDD),.Y(g25014),.A(g17474),.B(g23420));
  AND2 AND2_4080(.VSS(VSS),.VDD(VDD),.Y(g32328),.A(g5853),.B(g31554));
  AND2 AND2_4081(.VSS(VSS),.VDD(VDD),.Y(g29668),.A(g28527),.B(g14255));
  AND2 AND2_4082(.VSS(VSS),.VDD(VDD),.Y(g29842),.A(g28372),.B(g23284));
  AND2 AND2_4083(.VSS(VSS),.VDD(VDD),.Y(g27540),.A(g26576),.B(g17746));
  AND2 AND2_4084(.VSS(VSS),.VDD(VDD),.Y(g23564),.A(g16882),.B(g20648));
  AND4 AND4_247(.VSS(VSS),.VDD(VDD),.Y(g27058),.A(g10323),.B(g3522),.C(g3530),.D(g26264));
  AND2 AND2_4085(.VSS(VSS),.VDD(VDD),.Y(g30035),.A(g22539),.B(g28120));
  AND2 AND2_4086(.VSS(VSS),.VDD(VDD),.Y(g18140),.A(g559),.B(g17533));
  AND2 AND2_4087(.VSS(VSS),.VDD(VDD),.Y(g34340),.A(g34100),.B(g19950));
  AND2 AND2_4088(.VSS(VSS),.VDD(VDD),.Y(g27203),.A(g26026),.B(g16688));
  AND2 AND2_4089(.VSS(VSS),.VDD(VDD),.Y(g19596),.A(g1094),.B(g16681));
  AND2 AND2_4090(.VSS(VSS),.VDD(VDD),.Y(g26130),.A(g24890),.B(g19772));
  AND2 AND2_4091(.VSS(VSS),.VDD(VDD),.Y(g29525),.A(g2169),.B(g28837));
  AND2 AND2_4092(.VSS(VSS),.VDD(VDD),.Y(g21847),.A(g3905),.B(g21070));
  AND2 AND2_4093(.VSS(VSS),.VDD(VDD),.Y(g34684),.A(g14178),.B(g34545));
  AND2 AND2_4094(.VSS(VSS),.VDD(VDD),.Y(g10999),.A(g7880),.B(g1472));
  AND2 AND2_4095(.VSS(VSS),.VDD(VDD),.Y(g13833),.A(g4546),.B(g10613));
  AND3 AND3_227(.VSS(VSS),.VDD(VDD),.Y(I18819),.A(g13156),.B(g11450),.C(g11498));
  AND2 AND2_4096(.VSS(VSS),.VDD(VDD),.Y(g26362),.A(g19557),.B(g25538));
  AND4 AND4_248(.VSS(VSS),.VDD(VDD),.Y(g27044),.A(g7766),.B(g5873),.C(g5881),.D(g26241));
  AND2 AND2_4097(.VSS(VSS),.VDD(VDD),.Y(g31470),.A(g29753),.B(g23398));
  AND2 AND2_4098(.VSS(VSS),.VDD(VDD),.Y(g23397),.A(g11154),.B(g20239));
  AND3 AND3_228(.VSS(VSS),.VDD(VDD),.Y(g33470),.A(g32528),.B(I31046),.C(I31047));
  AND2 AND2_4099(.VSS(VSS),.VDD(VDD),.Y(g33915),.A(g33140),.B(g7846));
  AND2 AND2_4100(.VSS(VSS),.VDD(VDD),.Y(g32241),.A(g31244),.B(g20323));
  AND2 AND2_4101(.VSS(VSS),.VDD(VDD),.Y(g26165),.A(g11980),.B(g25153));
  AND4 AND4_249(.VSS(VSS),.VDD(VDD),.Y(g17793),.A(g6772),.B(g11592),.C(g6789),.D(I18803));
  AND4 AND4_250(.VSS(VSS),.VDD(VDD),.Y(g10998),.A(g8567),.B(g8509),.C(g8451),.D(g7650));
  AND2 AND2_4102(.VSS(VSS),.VDD(VDD),.Y(g18766),.A(g5495),.B(g17929));
  AND2 AND2_4103(.VSS(VSS),.VDD(VDD),.Y(g13048),.A(g8558),.B(g11043));
  AND2 AND2_4104(.VSS(VSS),.VDD(VDD),.Y(g23062),.A(g718),.B(g20248));
  AND2 AND2_4105(.VSS(VSS),.VDD(VDD),.Y(g27281),.A(g9830),.B(g26615));
  AND3 AND3_229(.VSS(VSS),.VDD(VDD),.Y(g24861),.A(g3712),.B(g23582),.C(I24033));
  AND2 AND2_4106(.VSS(VSS),.VDD(VDD),.Y(g24573),.A(g17198),.B(g23716));
  AND2 AND2_4107(.VSS(VSS),.VDD(VDD),.Y(g34517),.A(g34290),.B(g19493));
  AND2 AND2_4108(.VSS(VSS),.VDD(VDD),.Y(g28148),.A(g27355),.B(g26093));
  AND2 AND2_4109(.VSS(VSS),.VDD(VDD),.Y(g14233),.A(g8639),.B(g11855));
  AND2 AND2_4110(.VSS(VSS),.VDD(VDD),.Y(g21933),.A(g5212),.B(g18997));
  AND2 AND2_4111(.VSS(VSS),.VDD(VDD),.Y(g27301),.A(g11992),.B(g26679));
  AND4 AND4_251(.VSS(VSS),.VDD(VDD),.Y(I14225),.A(g8457),.B(g255),.C(g8406),.D(g262));
  AND2 AND2_4112(.VSS(VSS),.VDD(VDD),.Y(g27957),.A(g25947),.B(g15995));
  AND2 AND2_4113(.VSS(VSS),.VDD(VDD),.Y(g7804),.A(g2975),.B(g2970));
  AND2 AND2_4114(.VSS(VSS),.VDD(VDD),.Y(g25041),.A(g23261),.B(g20494));
  AND2 AND2_4115(.VSS(VSS),.VDD(VDD),.Y(g13221),.A(g6946),.B(g11425));
  AND2 AND2_4116(.VSS(VSS),.VDD(VDD),.Y(g27120),.A(g25878),.B(g22543));
  AND4 AND4_252(.VSS(VSS),.VDD(VDD),.Y(g17690),.A(g11547),.B(g11592),.C(g11640),.D(I18671));
  AND2 AND2_4117(.VSS(VSS),.VDD(VDD),.Y(g29865),.A(g1802),.B(g29115));
  AND2 AND2_4118(.VSS(VSS),.VDD(VDD),.Y(g21851),.A(g3901),.B(g21070));
  AND2 AND2_4119(.VSS(VSS),.VDD(VDD),.Y(g21872),.A(g4098),.B(g19801));
  AND2 AND2_4120(.VSS(VSS),.VDD(VDD),.Y(g23872),.A(g19389),.B(g4157));
  AND2 AND2_4121(.VSS(VSS),.VDD(VDD),.Y(g15883),.A(g9180),.B(g14258));
  AND2 AND2_4122(.VSS(VSS),.VDD(VDD),.Y(g18360),.A(g1830),.B(g17955));
  AND2 AND2_4123(.VSS(VSS),.VDD(VDD),.Y(g31467),.A(g30162),.B(g27937));
  AND2 AND2_4124(.VSS(VSS),.VDD(VDD),.Y(g31494),.A(g29792),.B(g23435));
  AND2 AND2_4125(.VSS(VSS),.VDD(VDD),.Y(g28343),.A(g27380),.B(g19799));
  AND3 AND3_230(.VSS(VSS),.VDD(VDD),.Y(I24527),.A(g9672),.B(g9264),.C(g5401));
  AND2 AND2_4126(.VSS(VSS),.VDD(VDD),.Y(g19655),.A(g2729),.B(g16966));
  AND3 AND3_231(.VSS(VSS),.VDD(VDD),.Y(g33467),.A(g32505),.B(I31031),.C(I31032));
  AND3 AND3_232(.VSS(VSS),.VDD(VDD),.Y(g33494),.A(g32700),.B(I31166),.C(I31167));
  AND2 AND2_4127(.VSS(VSS),.VDD(VDD),.Y(g24324),.A(g4540),.B(g22228));
  AND3 AND3_233(.VSS(VSS),.VDD(VDD),.Y(g27146),.A(g26148),.B(g8187),.C(g1648));
  AND2 AND2_4128(.VSS(VSS),.VDD(VDD),.Y(g27645),.A(g26488),.B(g15344));
  AND2 AND2_4129(.VSS(VSS),.VDD(VDD),.Y(g26863),.A(g24974),.B(g24957));
  AND2 AND2_4130(.VSS(VSS),.VDD(VDD),.Y(g18447),.A(g2208),.B(g18008));
  AND2 AND2_4131(.VSS(VSS),.VDD(VDD),.Y(g30193),.A(g28650),.B(g23848));
  AND2 AND2_4132(.VSS(VSS),.VDD(VDD),.Y(g24777),.A(g11345),.B(g23066));
  AND2 AND2_4133(.VSS(VSS),.VDD(VDD),.Y(g27699),.A(g26396),.B(g20766));
  AND2 AND2_4134(.VSS(VSS),.VDD(VDD),.Y(g16653),.A(g8343),.B(g13850));
  AND2 AND2_4135(.VSS(VSS),.VDD(VDD),.Y(g18162),.A(g686),.B(g17433));
  AND2 AND2_4136(.VSS(VSS),.VDD(VDD),.Y(g25983),.A(g2476),.B(g25009));
  AND2 AND2_4137(.VSS(VSS),.VDD(VDD),.Y(g29610),.A(g28483),.B(g8026));
  AND2 AND2_4138(.VSS(VSS),.VDD(VDD),.Y(g30165),.A(g28619),.B(g23788));
  AND2 AND2_4139(.VSS(VSS),.VDD(VDD),.Y(g22129),.A(g6633),.B(g19277));
  AND2 AND2_4140(.VSS(VSS),.VDD(VDD),.Y(g34523),.A(g9162),.B(g34351));
  AND2 AND2_4141(.VSS(VSS),.VDD(VDD),.Y(g22002),.A(g5706),.B(g21562));
  AND2 AND2_4142(.VSS(VSS),.VDD(VDD),.Y(g22057),.A(g15159),.B(g21611));
  AND2 AND2_4143(.VSS(VSS),.VDD(VDD),.Y(g17317),.A(g1079),.B(g13124));
  AND2 AND2_4144(.VSS(VSS),.VDD(VDD),.Y(g22128),.A(g6629),.B(g19277));
  AND2 AND2_4145(.VSS(VSS),.VDD(VDD),.Y(g33352),.A(g32237),.B(g20712));
  AND4 AND4_253(.VSS(VSS),.VDD(VDD),.Y(I31207),.A(g32754),.B(g32755),.C(g32756),.D(g32757));
  AND2 AND2_4146(.VSS(VSS),.VDD(VDD),.Y(g16636),.A(g5929),.B(g14768));
  AND2 AND2_4147(.VSS(VSS),.VDD(VDD),.Y(g18629),.A(g3680),.B(g17226));
  AND2 AND2_4148(.VSS(VSS),.VDD(VDD),.Y(g25142),.A(g4717),.B(g22885));
  AND2 AND2_4149(.VSS(VSS),.VDD(VDD),.Y(g18451),.A(g2295),.B(g15224));
  AND2 AND2_4150(.VSS(VSS),.VDD(VDD),.Y(g26347),.A(g262),.B(g24850));
  AND2 AND2_4151(.VSS(VSS),.VDD(VDD),.Y(g18472),.A(g2413),.B(g15224));
  AND2 AND2_4152(.VSS(VSS),.VDD(VDD),.Y(g32414),.A(g4944),.B(g30999));
  AND2 AND2_4153(.VSS(VSS),.VDD(VDD),.Y(g29188),.A(g27163),.B(g12762));
  AND2 AND2_4154(.VSS(VSS),.VDD(VDD),.Y(g33418),.A(g32372),.B(g21425));
  AND2 AND2_4155(.VSS(VSS),.VDD(VDD),.Y(g33822),.A(g33385),.B(g20157));
  AND2 AND2_4156(.VSS(VSS),.VDD(VDD),.Y(g18220),.A(g1002),.B(g16100));
  AND2 AND2_4157(.VSS(VSS),.VDD(VDD),.Y(g26253),.A(g2327),.B(g25435));
  AND2 AND2_4158(.VSS(VSS),.VDD(VDD),.Y(g30006),.A(g29032),.B(g9259));
  AND2 AND2_4159(.VSS(VSS),.VDD(VDD),.Y(g31266),.A(g30129),.B(g27742));
  AND2 AND2_4160(.VSS(VSS),.VDD(VDD),.Y(g31170),.A(g19128),.B(g29814));
  AND2 AND2_4161(.VSS(VSS),.VDD(VDD),.Y(g21452),.A(g16119),.B(g13624));
  AND2 AND2_4162(.VSS(VSS),.VDD(VDD),.Y(g18628),.A(g15095),.B(g17226));
  AND2 AND2_4163(.VSS(VSS),.VDD(VDD),.Y(g27427),.A(g26400),.B(g17575));
  AND2 AND2_4164(.VSS(VSS),.VDD(VDD),.Y(g34475),.A(g27450),.B(g34327));
  AND2 AND2_4165(.VSS(VSS),.VDD(VDD),.Y(g17057),.A(g446),.B(g13173));
  AND2 AND2_4166(.VSS(VSS),.VDD(VDD),.Y(g24140),.A(g17663),.B(g21654));
  AND2 AND2_4167(.VSS(VSS),.VDD(VDD),.Y(g22299),.A(g19999),.B(g21024));
  AND2 AND2_4168(.VSS(VSS),.VDD(VDD),.Y(g29686),.A(g2246),.B(g29057));
  AND2 AND2_4169(.VSS(VSS),.VDD(VDD),.Y(g24997),.A(g22929),.B(g10419));
  AND2 AND2_4170(.VSS(VSS),.VDD(VDD),.Y(g18246),.A(g1199),.B(g16431));
  AND2 AND2_4171(.VSS(VSS),.VDD(VDD),.Y(g21912),.A(g5052),.B(g21468));
  AND2 AND2_4172(.VSS(VSS),.VDD(VDD),.Y(g29383),.A(g28138),.B(g19412));
  AND2 AND2_4173(.VSS(VSS),.VDD(VDD),.Y(g30222),.A(g28701),.B(g23894));
  AND2 AND2_4174(.VSS(VSS),.VDD(VDD),.Y(g34863),.A(g16540),.B(g34833));
  AND2 AND2_4175(.VSS(VSS),.VDD(VDD),.Y(g28133),.A(g27367),.B(g23108));
  AND2 AND2_4176(.VSS(VSS),.VDD(VDD),.Y(g22298),.A(g19997),.B(g21012));
  AND4 AND4_254(.VSS(VSS),.VDD(VDD),.Y(g26236),.A(g25357),.B(g6856),.C(g7586),.D(g7558));
  AND2 AND2_4177(.VSS(VSS),.VDD(VDD),.Y(g28229),.A(g27345),.B(g17213));
  AND2 AND2_4178(.VSS(VSS),.VDD(VDD),.Y(g19487),.A(g499),.B(g16680));
  AND2 AND2_4179(.VSS(VSS),.VDD(VDD),.Y(g29938),.A(g23552),.B(g28889));
  AND2 AND2_4180(.VSS(VSS),.VDD(VDD),.Y(g26351),.A(g239),.B(g24869));
  AND2 AND2_4181(.VSS(VSS),.VDD(VDD),.Y(g28228),.A(g27126),.B(g19636));
  AND2 AND2_4182(.VSS(VSS),.VDD(VDD),.Y(g25130),.A(g23358),.B(g20600));
  AND2 AND2_4183(.VSS(VSS),.VDD(VDD),.Y(g26821),.A(g24821),.B(g13103));
  AND2 AND2_4184(.VSS(VSS),.VDD(VDD),.Y(g27661),.A(g26576),.B(g15568));
  AND4 AND4_255(.VSS(VSS),.VDD(VDD),.Y(I31241),.A(g30825),.B(g31838),.C(g32803),.D(g32804));
  AND2 AND2_4185(.VSS(VSS),.VDD(VDD),.Y(g27547),.A(g26549),.B(g17759));
  AND2 AND2_4186(.VSS(VSS),.VDD(VDD),.Y(g18591),.A(g2965),.B(g16349));
  AND2 AND2_4187(.VSS(VSS),.VDD(VDD),.Y(g31194),.A(g19128),.B(g29814));
  AND2 AND2_4188(.VSS(VSS),.VDD(VDD),.Y(g31167),.A(g10080),.B(g30076));
  AND2 AND2_4189(.VSS(VSS),.VDD(VDD),.Y(g18776),.A(g5813),.B(g18065));
  AND2 AND2_4190(.VSS(VSS),.VDD(VDD),.Y(g18785),.A(g5849),.B(g18065));
  AND2 AND2_4191(.VSS(VSS),.VDD(VDD),.Y(g15083),.A(g10362),.B(g12983));
  AND2 AND2_4192(.VSS(VSS),.VDD(VDD),.Y(g21756),.A(g3211),.B(g20785));
  AND2 AND2_4193(.VSS(VSS),.VDD(VDD),.Y(g18147),.A(g599),.B(g17533));
  AND2 AND2_4194(.VSS(VSS),.VDD(VDD),.Y(g25165),.A(g14062),.B(g23570));
  AND2 AND2_4195(.VSS(VSS),.VDD(VDD),.Y(g30253),.A(g28746),.B(g23943));
  AND2 AND2_4196(.VSS(VSS),.VDD(VDD),.Y(g16484),.A(g5244),.B(g14755));
  AND2 AND2_4197(.VSS(VSS),.VDD(VDD),.Y(g18754),.A(g5339),.B(g15595));
  AND2 AND2_4198(.VSS(VSS),.VDD(VDD),.Y(g31524),.A(g29897),.B(g20593));
  AND3 AND3_234(.VSS(VSS),.VDD(VDD),.Y(g33524),.A(g32918),.B(I31316),.C(I31317));
  AND2 AND2_4199(.VSS(VSS),.VDD(VDD),.Y(g18355),.A(g1748),.B(g17955));
  AND4 AND4_256(.VSS(VSS),.VDD(VDD),.Y(g26264),.A(g24688),.B(g8812),.C(g8778),.D(g10627));
  AND2 AND2_4200(.VSS(VSS),.VDD(VDD),.Y(g33836),.A(g33096),.B(g27020));
  AND2 AND2_4201(.VSS(VSS),.VDD(VDD),.Y(g21780),.A(g3391),.B(g20391));
  AND2 AND2_4202(.VSS(VSS),.VDD(VDD),.Y(g29875),.A(g28403),.B(g23337));
  AND2 AND2_4203(.VSS(VSS),.VDD(VDD),.Y(g32206),.A(g30609),.B(g25524));
  AND2 AND2_4204(.VSS(VSS),.VDD(VDD),.Y(g26516),.A(g24968),.B(g8876));
  AND2 AND2_4205(.VSS(VSS),.VDD(VDD),.Y(g13507),.A(g7023),.B(g12198));
  AND2 AND2_4206(.VSS(VSS),.VDD(VDD),.Y(g27481),.A(g26400),.B(g14630));
  AND2 AND2_4207(.VSS(VSS),.VDD(VDD),.Y(g30600),.A(g30287),.B(g18975));
  AND2 AND2_4208(.VSS(VSS),.VDD(VDD),.Y(g18825),.A(g6736),.B(g15680));
  AND2 AND2_4209(.VSS(VSS),.VDD(VDD),.Y(g18950),.A(g11193),.B(g16123));
  AND2 AND2_4210(.VSS(VSS),.VDD(VDD),.Y(g18370),.A(g1874),.B(g15171));
  AND2 AND2_4211(.VSS(VSS),.VDD(VDD),.Y(g31477),.A(g29763),.B(g23409));
  AND2 AND2_4212(.VSS(VSS),.VDD(VDD),.Y(g33401),.A(g32349),.B(g21381));
  AND3 AND3_235(.VSS(VSS),.VDD(VDD),.Y(g33477),.A(g32577),.B(I31081),.C(I31082));
  AND2 AND2_4213(.VSS(VSS),.VDD(VDD),.Y(g20162),.A(g8737),.B(g16750));
  AND2 AND2_4214(.VSS(VSS),.VDD(VDD),.Y(g30236),.A(g28724),.B(g23916));
  AND2 AND2_4215(.VSS(VSS),.VDD(VDD),.Y(g14148),.A(g884),.B(g10632));
  AND2 AND2_4216(.VSS(VSS),.VDD(VDD),.Y(g29837),.A(g28369),.B(g20144));
  AND2 AND2_4217(.VSS(VSS),.VDD(VDD),.Y(g14097),.A(g878),.B(g10632));
  AND2 AND2_4218(.VSS(VSS),.VDD(VDD),.Y(g21820),.A(g3712),.B(g20453));
  AND2 AND2_4219(.VSS(VSS),.VDD(VDD),.Y(g11163),.A(g6727),.B(g10224));
  AND3 AND3_236(.VSS(VSS),.VDD(VDD),.Y(I24067),.A(g3731),.B(g3736),.C(g8553));
  AND2 AND2_4220(.VSS(VSS),.VDD(VDD),.Y(g9906),.A(g996),.B(g1157));
  AND2 AND2_4221(.VSS(VSS),.VDD(VDD),.Y(g18151),.A(g617),.B(g17533));
  AND2 AND2_4222(.VSS(VSS),.VDD(VDD),.Y(g31118),.A(g29490),.B(g22906));
  AND2 AND2_4223(.VSS(VSS),.VDD(VDD),.Y(g18172),.A(g15058),.B(g17328));
  AND2 AND2_4224(.VSS(VSS),.VDD(VDD),.Y(g28627),.A(g27543),.B(g20574));
  AND2 AND2_4225(.VSS(VSS),.VDD(VDD),.Y(g32114),.A(g31624),.B(g29927));
  AND4 AND4_257(.VSS(VSS),.VDD(VDD),.Y(g28959),.A(g17401),.B(g25194),.C(g26424),.D(g27440));
  AND2 AND2_4226(.VSS(VSS),.VDD(VDD),.Y(g30175),.A(g28629),.B(g23813));
  AND2 AND2_4227(.VSS(VSS),.VDD(VDD),.Y(g32082),.A(g4917),.B(g30673));
  AND2 AND2_4228(.VSS(VSS),.VDD(VDD),.Y(g33864),.A(g33274),.B(g20524));
  AND2 AND2_4229(.VSS(VSS),.VDD(VDD),.Y(g27127),.A(g25997),.B(g16582));
  AND2 AND2_4230(.VSS(VSS),.VDD(VDD),.Y(g21846),.A(g3897),.B(g21070));
  AND2 AND2_4231(.VSS(VSS),.VDD(VDD),.Y(g28112),.A(g27352),.B(g26162));
  AND2 AND2_4232(.VSS(VSS),.VDD(VDD),.Y(g32107),.A(g31624),.B(g29912));
  AND2 AND2_4233(.VSS(VSS),.VDD(VDD),.Y(g15653),.A(g3119),.B(g13530));
  AND2 AND2_4234(.VSS(VSS),.VDD(VDD),.Y(g24629),.A(g6163),.B(g23699));
  AND2 AND2_4235(.VSS(VSS),.VDD(VDD),.Y(g23396),.A(g20051),.B(g20229));
  AND2 AND2_4236(.VSS(VSS),.VDD(VDD),.Y(g18367),.A(g1783),.B(g17955));
  AND2 AND2_4237(.VSS(VSS),.VDD(VDD),.Y(g18394),.A(g1862),.B(g15171));
  AND2 AND2_4238(.VSS(VSS),.VDD(VDD),.Y(g31313),.A(g30160),.B(g27907));
  AND2 AND2_4239(.VSS(VSS),.VDD(VDD),.Y(g24451),.A(g3476),.B(g23112));
  AND2 AND2_4240(.VSS(VSS),.VDD(VDD),.Y(g21731),.A(g3029),.B(g20330));
  AND2 AND2_4241(.VSS(VSS),.VDD(VDD),.Y(g24220),.A(g255),.B(g22594));
  AND2 AND2_4242(.VSS(VSS),.VDD(VDD),.Y(g20628),.A(g1046),.B(g15789));
  AND2 AND2_4243(.VSS(VSS),.VDD(VDD),.Y(g27490),.A(g26576),.B(g17651));
  AND2 AND2_4244(.VSS(VSS),.VDD(VDD),.Y(g13541),.A(g7069),.B(g12308));
  AND2 AND2_4245(.VSS(VSS),.VDD(VDD),.Y(g30264),.A(g28774),.B(g23963));
  AND2 AND2_4246(.VSS(VSS),.VDD(VDD),.Y(g34063),.A(g33806),.B(g23121));
  AND2 AND2_4247(.VSS(VSS),.VDD(VDD),.Y(g13473),.A(g9797),.B(g11841));
  AND2 AND2_4248(.VSS(VSS),.VDD(VDD),.Y(g30137),.A(g28594),.B(g21181));
  AND2 AND2_4249(.VSS(VSS),.VDD(VDD),.Y(g19601),.A(g16198),.B(g11149));
  AND2 AND2_4250(.VSS(VSS),.VDD(VDD),.Y(g24628),.A(g5835),.B(g23666));
  AND2 AND2_4251(.VSS(VSS),.VDD(VDD),.Y(g32345),.A(g2138),.B(g31672));
  AND2 AND2_4252(.VSS(VSS),.VDD(VDD),.Y(g34137),.A(g33928),.B(g23802));
  AND2 AND2_4253(.VSS(VSS),.VDD(VDD),.Y(g31285),.A(g30134),.B(g27800));
  AND2 AND2_4254(.VSS(VSS),.VDD(VDD),.Y(g34516),.A(g34289),.B(g19492));
  AND2 AND2_4255(.VSS(VSS),.VDD(VDD),.Y(g27376),.A(g26549),.B(g17481));
  AND2 AND2_4256(.VSS(VSS),.VDD(VDD),.Y(g27385),.A(g26400),.B(g17497));
  AND3 AND3_237(.VSS(VSS),.VDD(VDD),.Y(g33704),.A(g33176),.B(g10710),.C(g22319));
  AND2 AND2_4257(.VSS(VSS),.VDD(VDD),.Y(g29617),.A(g2024),.B(g28987));
  AND2 AND2_4258(.VSS(VSS),.VDD(VDD),.Y(g31305),.A(g29741),.B(g23354));
  AND4 AND4_258(.VSS(VSS),.VDD(VDD),.Y(I24695),.A(g24050),.B(g24051),.C(g24052),.D(g24053));
  AND3 AND3_238(.VSS(VSS),.VDD(VDD),.Y(I24018),.A(g8155),.B(g8390),.C(g3396));
  AND2 AND2_4259(.VSS(VSS),.VDD(VDD),.Y(g27103),.A(g25997),.B(g16509));
  AND2 AND2_4260(.VSS(VSS),.VDD(VDD),.Y(g33305),.A(g31935),.B(g17811));
  AND2 AND2_4261(.VSS(VSS),.VDD(VDD),.Y(g22831),.A(g19441),.B(g19629));
  AND2 AND2_4262(.VSS(VSS),.VDD(VDD),.Y(g23691),.A(g14731),.B(g20993));
  AND2 AND2_4263(.VSS(VSS),.VDD(VDD),.Y(g26542),.A(g13102),.B(g24376));
  AND2 AND2_4264(.VSS(VSS),.VDD(VDD),.Y(g34873),.A(g34830),.B(g20046));
  AND2 AND2_4265(.VSS(VSS),.VDD(VDD),.Y(g26021),.A(g9568),.B(g25035));
  AND2 AND2_4266(.VSS(VSS),.VDD(VDD),.Y(g18420),.A(g1996),.B(g15373));
  AND2 AND2_4267(.VSS(VSS),.VDD(VDD),.Y(g15852),.A(g13820),.B(g13223));
  AND2 AND2_4268(.VSS(VSS),.VDD(VDD),.Y(g27095),.A(g25997),.B(g16473));
  AND2 AND2_4269(.VSS(VSS),.VDD(VDD),.Y(g18319),.A(g1600),.B(g17873));
  AND2 AND2_4270(.VSS(VSS),.VDD(VDD),.Y(g33809),.A(g33432),.B(g30184));
  AND2 AND2_4271(.VSS(VSS),.VDD(VDD),.Y(g33900),.A(g33316),.B(g20913));
  AND3 AND3_239(.VSS(VSS),.VDD(VDD),.Y(g33466),.A(g32498),.B(I31026),.C(I31027));
  AND2 AND2_4272(.VSS(VSS),.VDD(VDD),.Y(g16184),.A(g9285),.B(g14183));
  AND2 AND2_4273(.VSS(VSS),.VDD(VDD),.Y(g16805),.A(g7187),.B(g12972));
  AND2 AND2_4274(.VSS(VSS),.VDD(VDD),.Y(g21405),.A(g13377),.B(g15811));
  AND2 AND2_4275(.VSS(VSS),.VDD(VDD),.Y(g16674),.A(g6637),.B(g15014));
  AND3 AND3_240(.VSS(VSS),.VDD(VDD),.Y(g29201),.A(g24081),.B(I27503),.C(I27504));
  AND2 AND2_4276(.VSS(VSS),.VDD(VDD),.Y(g32141),.A(g31639),.B(g29963));
  AND2 AND2_4277(.VSS(VSS),.VDD(VDD),.Y(g22316),.A(g2837),.B(g20270));
  AND2 AND2_4278(.VSS(VSS),.VDD(VDD),.Y(g18318),.A(g1604),.B(g17873));
  AND2 AND2_4279(.VSS(VSS),.VDD(VDD),.Y(g18446),.A(g2279),.B(g18008));
  AND2 AND2_4280(.VSS(VSS),.VDD(VDD),.Y(g33808),.A(g33109),.B(g22161));
  AND2 AND2_4281(.VSS(VSS),.VDD(VDD),.Y(g24785),.A(g7051),.B(g23645));
  AND2 AND2_4282(.VSS(VSS),.VDD(VDD),.Y(g18227),.A(g1052),.B(g16129));
  AND3 AND3_241(.VSS(VSS),.VDD(VDD),.Y(g7777),.A(g723),.B(g822),.C(g817));
  AND2 AND2_4283(.VSS(VSS),.VDD(VDD),.Y(g27181),.A(g26026),.B(g16655));
  AND2 AND2_4284(.VSS(VSS),.VDD(VDD),.Y(g30209),.A(g28682),.B(g23876));
  AND3 AND3_242(.VSS(VSS),.VDD(VDD),.Y(g22498),.A(g7753),.B(g7717),.C(g21334));
  AND2 AND2_4285(.VSS(VSS),.VDD(VDD),.Y(g33101),.A(g32398),.B(g18976));
  AND2 AND2_4286(.VSS(VSS),.VDD(VDD),.Y(g19791),.A(g14253),.B(g17189));
  AND2 AND2_4287(.VSS(VSS),.VDD(VDD),.Y(g24754),.A(g19604),.B(g23027));
  AND2 AND2_4288(.VSS(VSS),.VDD(VDD),.Y(g29595),.A(g28475),.B(g11833));
  AND2 AND2_4289(.VSS(VSS),.VDD(VDD),.Y(g29494),.A(g9073),.B(g28479));
  AND2 AND2_4290(.VSS(VSS),.VDD(VDD),.Y(g30208),.A(g28681),.B(g23875));
  AND2 AND2_4291(.VSS(VSS),.VDD(VDD),.Y(g16732),.A(g5555),.B(g14882));
  AND2 AND2_4292(.VSS(VSS),.VDD(VDD),.Y(g21929),.A(g5176),.B(g18997));
  AND2 AND2_4293(.VSS(VSS),.VDD(VDD),.Y(g32263),.A(g31631),.B(g30306));
  AND2 AND2_4294(.VSS(VSS),.VDD(VDD),.Y(g18540),.A(g2775),.B(g15277));
  AND2 AND2_4295(.VSS(VSS),.VDD(VDD),.Y(g10896),.A(g1205),.B(g8654));
  AND2 AND2_4296(.VSS(VSS),.VDD(VDD),.Y(g22056),.A(g6133),.B(g21611));
  AND2 AND2_4297(.VSS(VSS),.VDD(VDD),.Y(g26274),.A(g2130),.B(g25210));
  AND2 AND2_4298(.VSS(VSS),.VDD(VDD),.Y(g29623),.A(g28496),.B(g11563));
  AND2 AND2_4299(.VSS(VSS),.VDD(VDD),.Y(g32332),.A(g31325),.B(g23558));
  AND4 AND4_259(.VSS(VSS),.VDD(VDD),.Y(I31206),.A(g31710),.B(g31832),.C(g32752),.D(g32753));
  AND2 AND2_4300(.VSS(VSS),.VDD(VDD),.Y(g21928),.A(g5170),.B(g18997));
  AND2 AND2_4301(.VSS(VSS),.VDD(VDD),.Y(g22080),.A(g6275),.B(g19210));
  AND2 AND2_4302(.VSS(VSS),.VDD(VDD),.Y(g25063),.A(g13078),.B(g22325));
  AND3 AND3_243(.VSS(VSS),.VDD(VDD),.Y(g24858),.A(g3361),.B(g23223),.C(I24030));
  AND2 AND2_4303(.VSS(VSS),.VDD(VDD),.Y(g29782),.A(g28328),.B(g23245));
  AND2 AND2_4304(.VSS(VSS),.VDD(VDD),.Y(g18203),.A(g911),.B(g15938));
  AND2 AND2_4305(.VSS(VSS),.VDD(VDD),.Y(g26122),.A(g24557),.B(g19762));
  AND2 AND2_4306(.VSS(VSS),.VDD(VDD),.Y(g16761),.A(g7170),.B(g12947));
  AND2 AND2_4307(.VSS(VSS),.VDD(VDD),.Y(g29984),.A(g2567),.B(g28877));
  AND2 AND2_4308(.VSS(VSS),.VDD(VDD),.Y(g34542),.A(g34332),.B(g20089));
  AND3 AND3_244(.VSS(VSS),.VDD(VDD),.Y(g22432),.A(g9354),.B(g7717),.C(g21187));
  AND2 AND2_4309(.VSS(VSS),.VDD(VDD),.Y(g12931),.A(g392),.B(g11048));
  AND2 AND2_4310(.VSS(VSS),.VDD(VDD),.Y(g29352),.A(g4950),.B(g28410));
  AND2 AND2_4311(.VSS(VSS),.VDD(VDD),.Y(g25873),.A(g24854),.B(g16197));
  AND2 AND2_4312(.VSS(VSS),.VDD(VDD),.Y(g30614),.A(g20154),.B(g29814));
  AND3 AND3_245(.VSS(VSS),.VDD(VDD),.Y(I24597),.A(g5736),.B(g5742),.C(g9875));
  AND4 AND4_260(.VSS(VSS),.VDD(VDD),.Y(I31082),.A(g32573),.B(g32574),.C(g32575),.D(g32576));
  AND2 AND2_4313(.VSS(VSS),.VDD(VDD),.Y(g18281),.A(g1373),.B(g16136));
  AND2 AND2_4314(.VSS(VSS),.VDD(VDD),.Y(g27520),.A(g26519),.B(g17714));
  AND2 AND2_4315(.VSS(VSS),.VDD(VDD),.Y(g21787),.A(g15091),.B(g20391));
  AND2 AND2_4316(.VSS(VSS),.VDD(VDD),.Y(g15115),.A(g2946),.B(g14454));
  AND4 AND4_261(.VSS(VSS),.VDD(VDD),.Y(I31107),.A(g32610),.B(g32611),.C(g32612),.D(g32613));
  AND3 AND3_246(.VSS(VSS),.VDD(VDD),.Y(g22342),.A(g9354),.B(g9285),.C(g21287));
  AND2 AND2_4317(.VSS(VSS),.VDD(VDD),.Y(g18301),.A(g1532),.B(g16489));
  AND2 AND2_4318(.VSS(VSS),.VDD(VDD),.Y(g30607),.A(g30291),.B(g18989));
  AND2 AND2_4319(.VSS(VSS),.VDD(VDD),.Y(g32049),.A(g10902),.B(g30735));
  AND4 AND4_262(.VSS(VSS),.VDD(VDD),.Y(I24689),.A(g20841),.B(g24040),.C(g24041),.D(g24042));
  AND2 AND2_4320(.VSS(VSS),.VDD(VDD),.Y(g26292),.A(g2689),.B(g25228));
  AND2 AND2_4321(.VSS(VSS),.VDD(VDD),.Y(g33693),.A(g33145),.B(g13594));
  AND2 AND2_4322(.VSS(VSS),.VDD(VDD),.Y(g18377),.A(g1894),.B(g15171));
  AND2 AND2_4323(.VSS(VSS),.VDD(VDD),.Y(g19556),.A(g11932),.B(g16809));
  AND2 AND2_4324(.VSS(VSS),.VDD(VDD),.Y(g30073),.A(g1379),.B(g28194));
  AND2 AND2_4325(.VSS(VSS),.VDD(VDD),.Y(g22145),.A(g14555),.B(g18832));
  AND2 AND2_4326(.VSS(VSS),.VDD(VDD),.Y(g18120),.A(g457),.B(g17015));
  AND2 AND2_4327(.VSS(VSS),.VDD(VDD),.Y(g26153),.A(g24565),.B(g19780));
  AND2 AND2_4328(.VSS(VSS),.VDD(VDD),.Y(g18739),.A(g5008),.B(g16826));
  AND2 AND2_4329(.VSS(VSS),.VDD(VDD),.Y(g21302),.A(g956),.B(g15731));
  AND2 AND2_4330(.VSS(VSS),.VDD(VDD),.Y(g22031),.A(g5917),.B(g19147));
  AND2 AND2_4331(.VSS(VSS),.VDD(VDD),.Y(g27546),.A(g26549),.B(g17758));
  AND2 AND2_4332(.VSS(VSS),.VDD(VDD),.Y(g30274),.A(g28815),.B(g23983));
  AND2 AND2_4333(.VSS(VSS),.VDD(VDD),.Y(g31166),.A(g1816),.B(g30074));
  AND2 AND2_4334(.VSS(VSS),.VDD(VDD),.Y(g34073),.A(g8948),.B(g33823));
  AND2 AND2_4335(.VSS(VSS),.VDD(VDD),.Y(g10925),.A(g7858),.B(g956));
  AND2 AND2_4336(.VSS(VSS),.VDD(VDD),.Y(g16207),.A(g9839),.B(g14204));
  AND2 AND2_4337(.VSS(VSS),.VDD(VDD),.Y(g27211),.A(g25997),.B(g16716));
  AND2 AND2_4338(.VSS(VSS),.VDD(VDD),.Y(g32048),.A(g31498),.B(g13869));
  AND4 AND4_263(.VSS(VSS),.VDD(VDD),.Y(g16539),.A(g11547),.B(g6782),.C(g6789),.D(I17741));
  AND2 AND2_4339(.VSS(VSS),.VDD(VDD),.Y(g21743),.A(g3100),.B(g20330));
  AND2 AND2_4340(.VSS(VSS),.VDD(VDD),.Y(g21827),.A(g3759),.B(g20453));
  AND2 AND2_4341(.VSS(VSS),.VDD(VDD),.Y(g11029),.A(g5782),.B(g9103));
  AND2 AND2_4342(.VSS(VSS),.VDD(VDD),.Y(g17753),.A(g13281),.B(g13175));
  AND2 AND2_4343(.VSS(VSS),.VDD(VDD),.Y(g18146),.A(g595),.B(g17533));
  AND2 AND2_4344(.VSS(VSS),.VDD(VDD),.Y(g18738),.A(g15142),.B(g16826));
  AND2 AND2_4345(.VSS(VSS),.VDD(VDD),.Y(g13029),.A(g8359),.B(g11030));
  AND2 AND2_4346(.VSS(VSS),.VDD(VDD),.Y(g15745),.A(g686),.B(g13223));
  AND2 AND2_4347(.VSS(VSS),.VDD(VDD),.Y(g18645),.A(g15100),.B(g17271));
  AND2 AND2_4348(.VSS(VSS),.VDD(VDD),.Y(g30122),.A(g28578),.B(g21054));
  AND2 AND2_4349(.VSS(VSS),.VDD(VDD),.Y(g24420),.A(g23997),.B(g18980));
  AND2 AND2_4350(.VSS(VSS),.VDD(VDD),.Y(g24319),.A(g4561),.B(g22228));
  AND2 AND2_4351(.VSS(VSS),.VDD(VDD),.Y(g29853),.A(g1862),.B(g29081));
  AND2 AND2_4352(.VSS(VSS),.VDD(VDD),.Y(g16538),.A(g6255),.B(g15005));
  AND2 AND2_4353(.VSS(VSS),.VDD(VDD),.Y(g17145),.A(g7469),.B(g13249));
  AND2 AND2_4354(.VSS(VSS),.VDD(VDD),.Y(g26635),.A(g25321),.B(g20617));
  AND2 AND2_4355(.VSS(VSS),.VDD(VDD),.Y(g11028),.A(g9730),.B(g5428));
  AND2 AND2_4356(.VSS(VSS),.VDD(VDD),.Y(g18699),.A(g4760),.B(g16816));
  AND2 AND2_4357(.VSS(VSS),.VDD(VDD),.Y(g34565),.A(g34374),.B(g17471));
  AND2 AND2_4358(.VSS(VSS),.VDD(VDD),.Y(g15813),.A(g3247),.B(g14069));
  AND2 AND2_4359(.VSS(VSS),.VDD(VDD),.Y(g31485),.A(g29776),.B(g23421));
  AND2 AND2_4360(.VSS(VSS),.VDD(VDD),.Y(g29589),.A(g2575),.B(g28977));
  AND2 AND2_4361(.VSS(VSS),.VDD(VDD),.Y(g33892),.A(g33312),.B(g20701));
  AND2 AND2_4362(.VSS(VSS),.VDD(VDD),.Y(g18290),.A(g1467),.B(g16449));
  AND2 AND2_4363(.VSS(VSS),.VDD(VDD),.Y(g17199),.A(g2236),.B(g13034));
  AND2 AND2_4364(.VSS(VSS),.VDD(VDD),.Y(g24318),.A(g4555),.B(g22228));
  AND3 AND3_247(.VSS(VSS),.VDD(VDD),.Y(g33476),.A(g32570),.B(I31076),.C(I31077));
  AND3 AND3_248(.VSS(VSS),.VDD(VDD),.Y(g33485),.A(g32635),.B(I31121),.C(I31122));
  AND2 AND2_4365(.VSS(VSS),.VDD(VDD),.Y(g21769),.A(g3247),.B(g20785));
  AND2 AND2_4366(.VSS(VSS),.VDD(VDD),.Y(g30034),.A(g29077),.B(g10541));
  AND2 AND2_4367(.VSS(VSS),.VDD(VDD),.Y(g22843),.A(g9429),.B(g20272));
  AND2 AND2_4368(.VSS(VSS),.VDD(VDD),.Y(g24227),.A(g890),.B(g22594));
  AND2 AND2_4369(.VSS(VSS),.VDD(VDD),.Y(g18698),.A(g15131),.B(g16777));
  AND4 AND4_264(.VSS(VSS),.VDD(VDD),.Y(I31141),.A(g31376),.B(g31820),.C(g32659),.D(g32660));
  AND3 AND3_249(.VSS(VSS),.VDD(VDD),.Y(g25453),.A(g5406),.B(g23789),.C(I24576));
  AND2 AND2_4370(.VSS(VSS),.VDD(VDD),.Y(g29588),.A(g2311),.B(g28942));
  AND2 AND2_4371(.VSS(VSS),.VDD(VDD),.Y(g29524),.A(g2004),.B(g28864));
  AND2 AND2_4372(.VSS(VSS),.VDD(VDD),.Y(g29836),.A(g28425),.B(g26841));
  AND2 AND2_4373(.VSS(VSS),.VDD(VDD),.Y(g21768),.A(g3243),.B(g20785));
  AND2 AND2_4374(.VSS(VSS),.VDD(VDD),.Y(g21803),.A(g3538),.B(g20924));
  AND2 AND2_4375(.VSS(VSS),.VDD(VDD),.Y(g28245),.A(g11367),.B(g27975));
  AND2 AND2_4376(.VSS(VSS),.VDD(VDD),.Y(g15805),.A(g3243),.B(g14041));
  AND2 AND2_4377(.VSS(VSS),.VDD(VDD),.Y(g28626),.A(g27542),.B(g20573));
  AND2 AND2_4378(.VSS(VSS),.VDD(VDD),.Y(g30153),.A(g28610),.B(g23768));
  AND2 AND2_4379(.VSS(VSS),.VDD(VDD),.Y(g28299),.A(g9716),.B(g27670));
  AND4 AND4_265(.VSS(VSS),.VDD(VDD),.Y(g27700),.A(g22342),.B(g25182),.C(g26424),.D(g26148));
  AND2 AND2_4380(.VSS(VSS),.VDD(VDD),.Y(g22132),.A(g6645),.B(g19277));
  AND2 AND2_4381(.VSS(VSS),.VDD(VDD),.Y(g29477),.A(g14090),.B(g28441));
  AND2 AND2_4382(.VSS(VSS),.VDD(VDD),.Y(g32273),.A(g31255),.B(g20446));
  AND2 AND2_4383(.VSS(VSS),.VDD(VDD),.Y(g32106),.A(g31601),.B(g29911));
  AND2 AND2_4384(.VSS(VSS),.VDD(VDD),.Y(g18427),.A(g2181),.B(g18008));
  AND2 AND2_4385(.VSS(VSS),.VDD(VDD),.Y(g14681),.A(g4392),.B(g10476));
  AND2 AND2_4386(.VSS(VSS),.VDD(VDD),.Y(g19740),.A(g2783),.B(g15907));
  AND2 AND2_4387(.VSS(VSS),.VDD(VDD),.Y(g20203),.A(g6195),.B(g17789));
  AND3 AND3_250(.VSS(VSS),.VDD(VDD),.Y(g33907),.A(g23088),.B(g33219),.C(g9104));
  AND2 AND2_4388(.VSS(VSS),.VDD(VDD),.Y(g18366),.A(g1854),.B(g17955));
  AND4 AND4_266(.VSS(VSS),.VDD(VDD),.Y(I31332),.A(g32935),.B(g32936),.C(g32937),.D(g32938));
  AND2 AND2_4389(.VSS(VSS),.VDD(VDD),.Y(g21881),.A(g4064),.B(g19801));
  AND2 AND2_4390(.VSS(VSS),.VDD(VDD),.Y(g27658),.A(g22491),.B(g25786));
  AND2 AND2_4391(.VSS(VSS),.VDD(VDD),.Y(g18632),.A(g3698),.B(g17226));
  AND2 AND2_4392(.VSS(VSS),.VDD(VDD),.Y(g25905),.A(g24879),.B(g16311));
  AND2 AND2_4393(.VSS(VSS),.VDD(VDD),.Y(g17365),.A(g7650),.B(g13036));
  AND2 AND2_4394(.VSS(VSS),.VDD(VDD),.Y(g22161),.A(g13202),.B(g19071));
  AND2 AND2_4395(.VSS(VSS),.VDD(VDD),.Y(g33074),.A(g32387),.B(g18830));
  AND2 AND2_4396(.VSS(VSS),.VDD(VDD),.Y(g34136),.A(g33850),.B(g23293));
  AND2 AND2_4397(.VSS(VSS),.VDD(VDD),.Y(g33239),.A(g32117),.B(g19902));
  AND2 AND2_4398(.VSS(VSS),.VDD(VDD),.Y(g25530),.A(g23750),.B(g21414));
  AND2 AND2_4399(.VSS(VSS),.VDD(VDD),.Y(g27339),.A(g26400),.B(g17308));
  AND2 AND2_4400(.VSS(VSS),.VDD(VDD),.Y(g29749),.A(g28295),.B(g23214));
  AND2 AND2_4401(.VSS(VSS),.VDD(VDD),.Y(g29616),.A(g1974),.B(g29085));
  AND3 AND3_251(.VSS(VSS),.VDD(VDD),.Y(g7511),.A(g2145),.B(g2138),.C(g2130));
  AND2 AND2_4402(.VSS(VSS),.VDD(VDD),.Y(g26711),.A(g25446),.B(g20713));
  AND2 AND2_4403(.VSS(VSS),.VDD(VDD),.Y(g31238),.A(g29583),.B(g20053));
  AND2 AND2_4404(.VSS(VSS),.VDD(VDD),.Y(g32234),.A(g31601),.B(g30292));
  AND2 AND2_4405(.VSS(VSS),.VDD(VDD),.Y(g25122),.A(g23374),.B(g20592));
  AND2 AND2_4406(.VSS(VSS),.VDD(VDD),.Y(g18403),.A(g2028),.B(g15373));
  AND2 AND2_4407(.VSS(VSS),.VDD(VDD),.Y(g18547),.A(g121),.B(g15277));
  AND2 AND2_4408(.VSS(VSS),.VDD(VDD),.Y(g25565),.A(g13013),.B(g22660));
  AND2 AND2_4409(.VSS(VSS),.VDD(VDD),.Y(g24301),.A(g6961),.B(g22228));
  AND2 AND2_4410(.VSS(VSS),.VDD(VDD),.Y(g28232),.A(g27732),.B(g23586));
  AND2 AND2_4411(.VSS(VSS),.VDD(VDD),.Y(g20739),.A(g16259),.B(g4674));
  AND2 AND2_4412(.VSS(VSS),.VDD(VDD),.Y(g13491),.A(g6999),.B(g12160));
  AND2 AND2_4413(.VSS(VSS),.VDD(VDD),.Y(g22087),.A(g6303),.B(g19210));
  AND2 AND2_4414(.VSS(VSS),.VDD(VDD),.Y(g30164),.A(g28618),.B(g23787));
  AND2 AND2_4415(.VSS(VSS),.VDD(VDD),.Y(g31941),.A(g1283),.B(g30825));
  AND2 AND2_4416(.VSS(VSS),.VDD(VDD),.Y(g33941),.A(g33380),.B(g21560));
  AND2 AND2_4417(.VSS(VSS),.VDD(VDD),.Y(g18226),.A(g15064),.B(g16129));
  AND2 AND2_4418(.VSS(VSS),.VDD(VDD),.Y(g21890),.A(g4125),.B(g19801));
  AND2 AND2_4419(.VSS(VSS),.VDD(VDD),.Y(g13604),.A(g4495),.B(g10487));
  AND2 AND2_4420(.VSS(VSS),.VDD(VDD),.Y(g31519),.A(g29864),.B(g23490));
  AND2 AND2_4421(.VSS(VSS),.VDD(VDD),.Y(g18715),.A(g4871),.B(g15915));
  AND2 AND2_4422(.VSS(VSS),.VDD(VDD),.Y(g27968),.A(g25958),.B(g19614));
  AND2 AND2_4423(.VSS(VSS),.VDD(VDD),.Y(g28697),.A(g27581),.B(g20669));
  AND2 AND2_4424(.VSS(VSS),.VDD(VDD),.Y(g31185),.A(g10114),.B(g30087));
  AND2 AND2_4425(.VSS(VSS),.VDD(VDD),.Y(g18481),.A(g2461),.B(g15426));
  AND3 AND3_252(.VSS(VSS),.VDD(VDD),.Y(g33519),.A(g32881),.B(I31291),.C(I31292));
  AND2 AND2_4426(.VSS(VSS),.VDD(VDD),.Y(g29809),.A(g28362),.B(g23274));
  AND3 AND3_253(.VSS(VSS),.VDD(VDD),.Y(g33675),.A(g33164),.B(g10727),.C(g22332));
  AND2 AND2_4427(.VSS(VSS),.VDD(VDD),.Y(g24645),.A(g22639),.B(g19709));
  AND2 AND2_4428(.VSS(VSS),.VDD(VDD),.Y(g28261),.A(g27878),.B(g23695));
  AND2 AND2_4429(.VSS(VSS),.VDD(VDD),.Y(g26606),.A(g1018),.B(g24510));
  AND4 AND4_267(.VSS(VSS),.VDD(VDD),.Y(g28880),.A(g21434),.B(g26424),.C(g25438),.D(g27494));
  AND2 AND2_4430(.VSS(VSS),.VDD(VDD),.Y(g18551),.A(g2811),.B(g15277));
  AND2 AND2_4431(.VSS(VSS),.VDD(VDD),.Y(g22043),.A(g5965),.B(g19147));
  AND2 AND2_4432(.VSS(VSS),.VDD(VDD),.Y(g26303),.A(g2685),.B(g25439));
  AND2 AND2_4433(.VSS(VSS),.VDD(VDD),.Y(g31518),.A(g20041),.B(g29970));
  AND2 AND2_4434(.VSS(VSS),.VDD(VDD),.Y(g31154),.A(g19128),.B(g29814));
  AND2 AND2_4435(.VSS(VSS),.VDD(VDD),.Y(g18572),.A(g2864),.B(g16349));
  AND3 AND3_254(.VSS(VSS),.VDD(VDD),.Y(g33518),.A(g32874),.B(I31286),.C(I31287));
  AND2 AND2_4436(.VSS(VSS),.VDD(VDD),.Y(g29808),.A(g28361),.B(g23273));
  AND2 AND2_4437(.VSS(VSS),.VDD(VDD),.Y(g21710),.A(g287),.B(g20283));
  AND4 AND4_268(.VSS(VSS),.VDD(VDD),.Y(I31221),.A(g31327),.B(g31835),.C(g32773),.D(g32774));
  AND2 AND2_4438(.VSS(VSS),.VDD(VDD),.Y(g24290),.A(g4430),.B(g22550));
  AND4 AND4_269(.VSS(VSS),.VDD(VDD),.Y(g29036),.A(g27163),.B(g12762),.C(g20875),.D(I27381));
  AND2 AND2_4439(.VSS(VSS),.VDD(VDD),.Y(g27411),.A(g26549),.B(g17528));
  AND2 AND2_4440(.VSS(VSS),.VDD(VDD),.Y(g34474),.A(g20083),.B(g34326));
  AND2 AND2_4441(.VSS(VSS),.VDD(VDD),.Y(g24698),.A(g22664),.B(g19761));
  AND2 AND2_4442(.VSS(VSS),.VDD(VDD),.Y(g21779),.A(g3385),.B(g20391));
  AND2 AND2_4443(.VSS(VSS),.VDD(VDD),.Y(g26750),.A(g24514),.B(g24474));
  AND2 AND2_4444(.VSS(VSS),.VDD(VDD),.Y(g12527),.A(g8680),.B(g667));
  AND2 AND2_4445(.VSS(VSS),.VDD(VDD),.Y(g23779),.A(g1105),.B(g19355));
  AND2 AND2_4446(.VSS(VSS),.VDD(VDD),.Y(g18127),.A(g499),.B(g16971));
  AND2 AND2_4447(.VSS(VSS),.VDD(VDD),.Y(g22069),.A(g6227),.B(g19210));
  AND2 AND2_4448(.VSS(VSS),.VDD(VDD),.Y(g25408),.A(g22682),.B(g9772));
  AND2 AND2_4449(.VSS(VSS),.VDD(VDD),.Y(g30109),.A(g28562),.B(g20912));
  AND2 AND2_4450(.VSS(VSS),.VDD(VDD),.Y(g26381),.A(g4456),.B(g25548));
  AND2 AND2_4451(.VSS(VSS),.VDD(VDD),.Y(g34109),.A(g33918),.B(g23708));
  AND2 AND2_4452(.VSS(VSS),.VDD(VDD),.Y(g29642),.A(g27954),.B(g28669));
  AND2 AND2_4453(.VSS(VSS),.VDD(VDD),.Y(g33883),.A(g33294),.B(g20589));
  AND2 AND2_4454(.VSS(VSS),.VDD(VDD),.Y(g21778),.A(g3355),.B(g20391));
  AND2 AND2_4455(.VSS(VSS),.VDD(VDD),.Y(g22068),.A(g6219),.B(g19210));
  AND2 AND2_4456(.VSS(VSS),.VDD(VDD),.Y(g26091),.A(g1691),.B(g25082));
  AND2 AND2_4457(.VSS(VSS),.VDD(VDD),.Y(g18490),.A(g2504),.B(g15426));
  AND2 AND2_4458(.VSS(VSS),.VDD(VDD),.Y(g30108),.A(g28561),.B(g20910));
  AND2 AND2_4459(.VSS(VSS),.VDD(VDD),.Y(g32163),.A(g3502),.B(g31170));
  AND2 AND2_4460(.VSS(VSS),.VDD(VDD),.Y(g32012),.A(g8297),.B(g31233));
  AND3 AND3_255(.VSS(VSS),.VDD(VDD),.Y(g34108),.A(g22957),.B(g9104),.C(g33766));
  AND2 AND2_4461(.VSS(VSS),.VDD(VDD),.Y(g24427),.A(g4961),.B(g22919));
  AND2 AND2_4462(.VSS(VSS),.VDD(VDD),.Y(g21786),.A(g3436),.B(g20391));
  AND2 AND2_4463(.VSS(VSS),.VDD(VDD),.Y(g27503),.A(g26488),.B(g14668));
  AND3 AND3_256(.VSS(VSS),.VDD(VDD),.Y(I24054),.A(g8443),.B(g8075),.C(g3747));
  AND2 AND2_4464(.VSS(VSS),.VDD(VDD),.Y(g30283),.A(g28851),.B(g23993));
  AND4 AND4_270(.VSS(VSS),.VDD(VDD),.Y(I31106),.A(g30825),.B(g31814),.C(g32608),.D(g32609));
  AND2 AND2_4465(.VSS(VSS),.VDD(VDD),.Y(g18784),.A(g15155),.B(g18065));
  AND2 AND2_4466(.VSS(VSS),.VDD(VDD),.Y(g18376),.A(g1913),.B(g15171));
  AND2 AND2_4467(.VSS(VSS),.VDD(VDD),.Y(g18385),.A(g1959),.B(g15171));
  AND2 AND2_4468(.VSS(VSS),.VDD(VDD),.Y(g29733),.A(g2675),.B(g29157));
  AND2 AND2_4469(.VSS(VSS),.VDD(VDD),.Y(g18297),.A(g1478),.B(g16449));
  AND2 AND2_4470(.VSS(VSS),.VDD(VDD),.Y(g17810),.A(g1495),.B(g13246));
  AND2 AND2_4471(.VSS(VSS),.VDD(VDD),.Y(g18103),.A(g401),.B(g17015));
  AND2 AND2_4472(.VSS(VSS),.VDD(VDD),.Y(g10626),.A(g4057),.B(g7927));
  AND2 AND2_4473(.VSS(VSS),.VDD(VDD),.Y(g34492),.A(g34272),.B(g33430));
  AND2 AND2_4474(.VSS(VSS),.VDD(VDD),.Y(g13633),.A(g4567),.B(g10509));
  AND2 AND2_4475(.VSS(VSS),.VDD(VDD),.Y(g25164),.A(g16883),.B(g23569));
  AND2 AND2_4476(.VSS(VSS),.VDD(VDD),.Y(g21945),.A(g5248),.B(g18997));
  AND2 AND2_4477(.VSS(VSS),.VDD(VDD),.Y(g28499),.A(g27982),.B(g17762));
  AND2 AND2_4478(.VSS(VSS),.VDD(VDD),.Y(g18354),.A(g1792),.B(g17955));
  AND2 AND2_4479(.VSS(VSS),.VDD(VDD),.Y(g29874),.A(g28402),.B(g23336));
  AND4 AND4_271(.VSS(VSS),.VDD(VDD),.Y(g27714),.A(g22384),.B(g25195),.C(g26424),.D(g26171));
  AND2 AND2_4480(.VSS(VSS),.VDD(VDD),.Y(g21826),.A(g3742),.B(g20453));
  AND2 AND2_4481(.VSS(VSS),.VDD(VDD),.Y(g21999),.A(g5723),.B(g21562));
  AND2 AND2_4482(.VSS(VSS),.VDD(VDD),.Y(g26390),.A(g4423),.B(g25554));
  AND2 AND2_4483(.VSS(VSS),.VDD(VDD),.Y(g31501),.A(g2047),.B(g29310));
  AND2 AND2_4484(.VSS(VSS),.VDD(VDD),.Y(g18824),.A(g6732),.B(g15680));
  AND2 AND2_4485(.VSS(VSS),.VDD(VDD),.Y(g27315),.A(g12022),.B(g26709));
  AND3 AND3_257(.VSS(VSS),.VDD(VDD),.Y(g33501),.A(g32751),.B(I31201),.C(I31202));
  AND2 AND2_4486(.VSS(VSS),.VDD(VDD),.Y(g29630),.A(g28212),.B(g19781));
  AND2 AND2_4487(.VSS(VSS),.VDD(VDD),.Y(g24403),.A(g4894),.B(g22858));
  AND2 AND2_4488(.VSS(VSS),.VDD(VDD),.Y(g29693),.A(g28207),.B(g10233));
  AND2 AND2_4489(.VSS(VSS),.VDD(VDD),.Y(g30982),.A(g8895),.B(g29933));
  AND2 AND2_4490(.VSS(VSS),.VDD(VDD),.Y(g34750),.A(g34673),.B(g19542));
  AND2 AND2_4491(.VSS(VSS),.VDD(VDD),.Y(g16759),.A(g5587),.B(g14761));
  AND2 AND2_4492(.VSS(VSS),.VDD(VDD),.Y(g18181),.A(g772),.B(g17328));
  AND2 AND2_4493(.VSS(VSS),.VDD(VDD),.Y(g21998),.A(g5712),.B(g21562));
  AND2 AND2_4494(.VSS(VSS),.VDD(VDD),.Y(g18671),.A(g4628),.B(g15758));
  AND2 AND2_4495(.VSS(VSS),.VDD(VDD),.Y(g34381),.A(g34166),.B(g20594));
  AND2 AND2_4496(.VSS(VSS),.VDD(VDD),.Y(g23998),.A(g19631),.B(g10971));
  AND3 AND3_258(.VSS(VSS),.VDD(VDD),.Y(g33728),.A(g22626),.B(g10851),.C(g33187));
  AND2 AND2_4497(.VSS(VSS),.VDD(VDD),.Y(g27202),.A(g25997),.B(g13876));
  AND2 AND2_4498(.VSS(VSS),.VDD(VDD),.Y(g19568),.A(g1467),.B(g15959));
  AND2 AND2_4499(.VSS(VSS),.VDD(VDD),.Y(g30091),.A(g28127),.B(g20716));
  AND2 AND2_4500(.VSS(VSS),.VDD(VDD),.Y(g32325),.A(g31316),.B(g23538));
  AND2 AND2_4501(.VSS(VSS),.VDD(VDD),.Y(g29665),.A(g2375),.B(g28696));
  AND2 AND2_4502(.VSS(VSS),.VDD(VDD),.Y(g16758),.A(g5220),.B(g14758));
  AND3 AND3_259(.VSS(VSS),.VDD(VDD),.Y(g34091),.A(g22957),.B(g9104),.C(g33761));
  AND2 AND2_4503(.VSS(VSS),.VDD(VDD),.Y(g24226),.A(g446),.B(g22594));
  AND2 AND2_4504(.VSS(VSS),.VDD(VDD),.Y(g13832),.A(g8880),.B(g10612));
  AND2 AND2_4505(.VSS(VSS),.VDD(VDD),.Y(g28722),.A(g27955),.B(g20738));
  AND4 AND4_272(.VSS(VSS),.VDD(VDD),.Y(g28924),.A(g17317),.B(g25183),.C(g26424),.D(g27416));
  AND2 AND2_4506(.VSS(VSS),.VDD(VDD),.Y(g30174),.A(g28628),.B(g23812));
  AND4 AND4_273(.VSS(VSS),.VDD(VDD),.Y(g29008),.A(g27163),.B(g12730),.C(g20739),.D(I27364));
  AND2 AND2_4507(.VSS(VSS),.VDD(VDD),.Y(g12979),.A(g424),.B(g11048));
  AND2 AND2_4508(.VSS(VSS),.VDD(VDD),.Y(g24551),.A(g17148),.B(g23331));
  AND2 AND2_4509(.VSS(VSS),.VDD(VDD),.Y(g24572),.A(g5462),.B(g23393));
  AND2 AND2_4510(.VSS(VSS),.VDD(VDD),.Y(g33349),.A(g32233),.B(g20699));
  AND2 AND2_4511(.VSS(VSS),.VDD(VDD),.Y(g25108),.A(g23345),.B(g20576));
  AND2 AND2_4512(.VSS(VSS),.VDD(VDD),.Y(g21932),.A(g5204),.B(g18997));
  AND2 AND2_4513(.VSS(VSS),.VDD(VDD),.Y(g32121),.A(g31616),.B(g29942));
  AND2 AND2_4514(.VSS(VSS),.VDD(VDD),.Y(g18426),.A(g2177),.B(g18008));
  AND2 AND2_4515(.VSS(VSS),.VDD(VDD),.Y(g33906),.A(g33084),.B(g22311));
  AND2 AND2_4516(.VSS(VSS),.VDD(VDD),.Y(g13247),.A(g8964),.B(g11316));
  AND2 AND2_4517(.VSS(VSS),.VDD(VDD),.Y(g29555),.A(g29004),.B(g22498));
  AND2 AND2_4518(.VSS(VSS),.VDD(VDD),.Y(g21513),.A(g16196),.B(g10882));
  AND2 AND2_4519(.VSS(VSS),.VDD(VDD),.Y(g18190),.A(g822),.B(g17821));
  AND2 AND2_4520(.VSS(VSS),.VDD(VDD),.Y(g22010),.A(g5787),.B(g21562));
  AND2 AND2_4521(.VSS(VSS),.VDD(VDD),.Y(g23513),.A(g19430),.B(g13007));
  AND2 AND2_4522(.VSS(VSS),.VDD(VDD),.Y(g34390),.A(g34172),.B(g21069));
  AND2 AND2_4523(.VSS(VSS),.VDD(VDD),.Y(g10856),.A(g4269),.B(g8967));
  AND2 AND2_4524(.VSS(VSS),.VDD(VDD),.Y(g11045),.A(g5787),.B(g9883));
  AND2 AND2_4525(.VSS(VSS),.VDD(VDD),.Y(g15882),.A(g3554),.B(g13986));
  AND2 AND2_4526(.VSS(VSS),.VDD(VDD),.Y(g27384),.A(g26400),.B(g17496));
  AND2 AND2_4527(.VSS(VSS),.VDD(VDD),.Y(g29570),.A(g2763),.B(g28598));
  AND2 AND2_4528(.VSS(VSS),.VDD(VDD),.Y(g29712),.A(g2643),.B(g28726));
  AND4 AND4_274(.VSS(VSS),.VDD(VDD),.Y(I24694),.A(g20982),.B(g24047),.C(g24048),.D(g24049));
  AND2 AND2_4529(.VSS(VSS),.VDD(VDD),.Y(g33304),.A(g32427),.B(g31971));
  AND2 AND2_4530(.VSS(VSS),.VDD(VDD),.Y(g14261),.A(g4507),.B(g10738));
  AND2 AND2_4531(.VSS(VSS),.VDD(VDD),.Y(g18520),.A(g2661),.B(g15509));
  AND2 AND2_4532(.VSS(VSS),.VDD(VDD),.Y(g21961),.A(g5424),.B(g21514));
  AND2 AND2_4533(.VSS(VSS),.VDD(VDD),.Y(g22079),.A(g6271),.B(g19210));
  AND2 AND2_4534(.VSS(VSS),.VDD(VDD),.Y(g27094),.A(g25997),.B(g16472));
  AND2 AND2_4535(.VSS(VSS),.VDD(VDD),.Y(g30192),.A(g28649),.B(g23847));
  AND2 AND2_4536(.VSS(VSS),.VDD(VDD),.Y(g31566),.A(g19050),.B(g29814));
  AND2 AND2_4537(.VSS(VSS),.VDD(VDD),.Y(g13324),.A(g854),.B(g11326));
  AND2 AND2_4538(.VSS(VSS),.VDD(VDD),.Y(g29907),.A(g2629),.B(g29177));
  AND2 AND2_4539(.VSS(VSS),.VDD(VDD),.Y(g32291),.A(g31268),.B(g20527));
  AND2 AND2_4540(.VSS(VSS),.VDD(VDD),.Y(g16804),.A(g5905),.B(g14813));
  AND2 AND2_4541(.VSS(VSS),.VDD(VDD),.Y(g21404),.A(g16069),.B(g13569));
  AND2 AND2_4542(.VSS(VSS),.VDD(VDD),.Y(g28199),.A(g27479),.B(g16684));
  AND2 AND2_4543(.VSS(VSS),.VDD(VDD),.Y(g22078),.A(g6267),.B(g19210));
  AND2 AND2_4544(.VSS(VSS),.VDD(VDD),.Y(g23404),.A(g20063),.B(g20247));
  AND2 AND2_4545(.VSS(VSS),.VDD(VDD),.Y(g32173),.A(g160),.B(g31134));
  AND2 AND2_4546(.VSS(VSS),.VDD(VDD),.Y(g18546),.A(g2795),.B(g15277));
  AND2 AND2_4547(.VSS(VSS),.VDD(VDD),.Y(g25982),.A(g2351),.B(g25008));
  AND4 AND4_275(.VSS(VSS),.VDD(VDD),.Y(I31012),.A(g32473),.B(g32474),.C(g32475),.D(g32476));
  AND2 AND2_4548(.VSS(VSS),.VDD(VDD),.Y(g18211),.A(g15062),.B(g15979));
  AND2 AND2_4549(.VSS(VSS),.VDD(VDD),.Y(g21717),.A(g15051),.B(g21037));
  AND2 AND2_4550(.VSS(VSS),.VDD(VDD),.Y(g28198),.A(g26649),.B(g27492));
  AND2 AND2_4551(.VSS(VSS),.VDD(VDD),.Y(g24297),.A(g4455),.B(g22550));
  AND2 AND2_4552(.VSS(VSS),.VDD(VDD),.Y(g22086),.A(g6299),.B(g19210));
  AND2 AND2_4553(.VSS(VSS),.VDD(VDD),.Y(g25091),.A(g12830),.B(g23492));
  AND2 AND2_4554(.VSS(VSS),.VDD(VDD),.Y(g20095),.A(g8873),.B(g16632));
  AND3 AND3_260(.VSS(VSS),.VDD(VDD),.Y(I24619),.A(g6423),.B(g6428),.C(g10014));
  AND2 AND2_4555(.VSS(VSS),.VDD(VDD),.Y(g29567),.A(g2357),.B(g28593));
  AND2 AND2_4556(.VSS(VSS),.VDD(VDD),.Y(g29594),.A(g28529),.B(g14192));
  AND3 AND3_261(.VSS(VSS),.VDD(VDD),.Y(g12735),.A(g7121),.B(g3873),.C(g3881));
  AND2 AND2_4557(.VSS(VSS),.VDD(VDD),.Y(g31139),.A(g12221),.B(g30036));
  AND2 AND2_4558(.VSS(VSS),.VDD(VDD),.Y(g28528),.A(g27187),.B(g12730));
  AND2 AND2_4559(.VSS(VSS),.VDD(VDD),.Y(g28330),.A(g27238),.B(g19786));
  AND2 AND2_4560(.VSS(VSS),.VDD(VDD),.Y(g26252),.A(g2283),.B(g25309));
  AND2 AND2_4561(.VSS(VSS),.VDD(VDD),.Y(g11032),.A(g9354),.B(g7717));
  AND2 AND2_4562(.VSS(VSS),.VDD(VDD),.Y(g34483),.A(g34406),.B(g18938));
  AND2 AND2_4563(.VSS(VSS),.VDD(VDD),.Y(g18497),.A(g2541),.B(g15426));
  AND2 AND2_4564(.VSS(VSS),.VDD(VDD),.Y(g32029),.A(g31318),.B(g16482));
  AND2 AND2_4565(.VSS(VSS),.VDD(VDD),.Y(g24671),.A(g5481),.B(g23630));
  AND2 AND2_4566(.VSS(VSS),.VDD(VDD),.Y(g14831),.A(g1152),.B(g10909));
  AND2 AND2_4567(.VSS(VSS),.VDD(VDD),.Y(g22125),.A(g6617),.B(g19277));
  AND3 AND3_262(.VSS(VSS),.VDD(VDD),.Y(g29382),.A(g26424),.B(g22763),.C(g28172));
  AND2 AND2_4568(.VSS(VSS),.VDD(VDD),.Y(g27526),.A(g26576),.B(g17721));
  AND2 AND2_4569(.VSS(VSS),.VDD(VDD),.Y(g34862),.A(g16540),.B(g34830));
  AND2 AND2_4570(.VSS(VSS),.VDD(VDD),.Y(g29519),.A(g2295),.B(g28840));
  AND2 AND2_4571(.VSS(VSS),.VDD(VDD),.Y(g32028),.A(g30569),.B(g29339));
  AND2 AND2_4572(.VSS(VSS),.VDD(VDD),.Y(g19578),.A(g16183),.B(g11130));
  AND2 AND2_4573(.VSS(VSS),.VDD(VDD),.Y(g33415),.A(g32368),.B(g21422));
  AND2 AND2_4574(.VSS(VSS),.VDD(VDD),.Y(g22158),.A(g13698),.B(g19609));
  AND2 AND2_4575(.VSS(VSS),.VDD(VDD),.Y(g14316),.A(g2370),.B(g11920));
  AND2 AND2_4576(.VSS(VSS),.VDD(VDD),.Y(g33333),.A(g32218),.B(g20612));
  AND2 AND2_4577(.VSS(VSS),.VDD(VDD),.Y(g18700),.A(g15132),.B(g16816));
  AND4 AND4_276(.VSS(VSS),.VDD(VDD),.Y(g17817),.A(g11547),.B(g6782),.C(g11640),.D(I18819));
  AND2 AND2_4578(.VSS(VSS),.VDD(VDD),.Y(g18126),.A(g15054),.B(g16971));
  AND2 AND2_4579(.VSS(VSS),.VDD(VDD),.Y(g18659),.A(g4366),.B(g17183));
  AND2 AND2_4580(.VSS(VSS),.VDD(VDD),.Y(g18625),.A(g15092),.B(g17062));
  AND2 AND2_4581(.VSS(VSS),.VDD(VDD),.Y(g18987),.A(g182),.B(g16162));
  AND2 AND2_4582(.VSS(VSS),.VDD(VDD),.Y(g29518),.A(g28906),.B(g22384));
  AND2 AND2_4583(.VSS(VSS),.VDD(VDD),.Y(g18250),.A(g6821),.B(g16897));
  AND2 AND2_4584(.VSS(VSS),.VDD(VDD),.Y(g24931),.A(g23153),.B(g20178));
  AND2 AND2_4585(.VSS(VSS),.VDD(VDD),.Y(g15114),.A(g4239),.B(g14454));
  AND2 AND2_4586(.VSS(VSS),.VDD(VDD),.Y(g25192),.A(g20276),.B(g23648));
  AND2 AND2_4587(.VSS(VSS),.VDD(VDD),.Y(g26847),.A(g2873),.B(g24525));
  AND2 AND2_4588(.VSS(VSS),.VDD(VDD),.Y(g34948),.A(g16540),.B(g34935));
  AND2 AND2_4589(.VSS(VSS),.VDD(VDD),.Y(g18658),.A(g15121),.B(g17183));
  AND2 AND2_4590(.VSS(VSS),.VDD(VDD),.Y(g27457),.A(g26519),.B(g17606));
  AND2 AND2_4591(.VSS(VSS),.VDD(VDD),.Y(g26397),.A(g19475),.B(g25563));
  AND2 AND2_4592(.VSS(VSS),.VDD(VDD),.Y(g15082),.A(g2697),.B(g12983));
  AND2 AND2_4593(.VSS(VSS),.VDD(VDD),.Y(g23387),.A(g16506),.B(g20211));
  AND2 AND2_4594(.VSS(VSS),.VDD(VDD),.Y(g31963),.A(g30731),.B(g18895));
  AND2 AND2_4595(.VSS(VSS),.VDD(VDD),.Y(g29637),.A(g2533),.B(g29134));
  AND2 AND2_4596(.VSS(VSS),.VDD(VDD),.Y(g22680),.A(g19530),.B(g7781));
  AND2 AND2_4597(.VSS(VSS),.VDD(VDD),.Y(g34702),.A(g34537),.B(g20208));
  AND2 AND2_4598(.VSS(VSS),.VDD(VDD),.Y(g15107),.A(g4258),.B(g14454));
  AND2 AND2_4599(.VSS(VSS),.VDD(VDD),.Y(g23148),.A(g19128),.B(g9104));
  AND2 AND2_4600(.VSS(VSS),.VDD(VDD),.Y(g34757),.A(g34682),.B(g19635));
  AND2 AND2_4601(.VSS(VSS),.VDD(VDD),.Y(g17783),.A(g7851),.B(g13110));
  AND2 AND2_4602(.VSS(VSS),.VDD(VDD),.Y(g25522),.A(g6888),.B(g22544));
  AND4 AND4_277(.VSS(VSS),.VDD(VDD),.Y(I31121),.A(g30614),.B(g31817),.C(g32629),.D(g32630));
  AND2 AND2_4603(.VSS(VSS),.VDD(VDD),.Y(g24190),.A(g329),.B(g22722));
  AND2 AND2_4604(.VSS(VSS),.VDD(VDD),.Y(g18339),.A(g1714),.B(g17873));
  AND2 AND2_4605(.VSS(VSS),.VDD(VDD),.Y(g18943),.A(g269),.B(g16099));
  AND2 AND2_4606(.VSS(VSS),.VDD(VDD),.Y(g29883),.A(g2465),.B(g29152));
  AND2 AND2_4607(.VSS(VSS),.VDD(VDD),.Y(g18296),.A(g1495),.B(g16449));
  AND2 AND2_4608(.VSS(VSS),.VDD(VDD),.Y(g21811),.A(g3582),.B(g20924));
  AND2 AND2_4609(.VSS(VSS),.VDD(VDD),.Y(g28225),.A(g27770),.B(g23400));
  AND2 AND2_4610(.VSS(VSS),.VDD(VDD),.Y(g23104),.A(g661),.B(g20248));
  AND2 AND2_4611(.VSS(VSS),.VDD(VDD),.Y(g23811),.A(g4087),.B(g19364));
  AND2 AND2_4612(.VSS(VSS),.VDD(VDD),.Y(g23646),.A(g16959),.B(g20737));
  AND2 AND2_4613(.VSS(VSS),.VDD(VDD),.Y(g18644),.A(g15098),.B(g17125));
  AND4 AND4_278(.VSS(VSS),.VDD(VDD),.Y(g28471),.A(g27187),.B(g12762),.C(g21024),.D(I26960));
  AND2 AND2_4614(.VSS(VSS),.VDD(VDD),.Y(g16221),.A(g5791),.B(g14231));
  AND2 AND2_4615(.VSS(VSS),.VDD(VDD),.Y(g18338),.A(g1710),.B(g17873));
  AND2 AND2_4616(.VSS(VSS),.VDD(VDD),.Y(g30564),.A(g21358),.B(g29385));
  AND2 AND2_4617(.VSS(VSS),.VDD(VDD),.Y(g9967),.A(g1178),.B(g1157));
  AND2 AND2_4618(.VSS(VSS),.VDD(VDD),.Y(g28258),.A(g27182),.B(g19687));
  AND2 AND2_4619(.VSS(VSS),.VDD(VDD),.Y(g21971),.A(g5417),.B(g21514));
  AND2 AND2_4620(.VSS(VSS),.VDD(VDD),.Y(g34564),.A(g34373),.B(g17466));
  AND2 AND2_4621(.VSS(VSS),.VDD(VDD),.Y(g15849),.A(g3538),.B(g14136));
  AND2 AND2_4622(.VSS(VSS),.VDD(VDD),.Y(g31484),.A(g29775),.B(g23418));
  AND2 AND2_4623(.VSS(VSS),.VDD(VDD),.Y(g24546),.A(g22447),.B(g19523));
  AND3 AND3_263(.VSS(VSS),.VDD(VDD),.Y(g33484),.A(g32628),.B(I31116),.C(I31117));
  AND2 AND2_4624(.VSS(VSS),.VDD(VDD),.Y(g16613),.A(g5925),.B(g14732));
  AND4 AND4_279(.VSS(VSS),.VDD(VDD),.Y(I31291),.A(g31021),.B(g31847),.C(g32875),.D(g32876));
  AND2 AND2_4625(.VSS(VSS),.VDD(VDD),.Y(g15848),.A(g3259),.B(g13892));
  AND2 AND2_4626(.VSS(VSS),.VDD(VDD),.Y(g19275),.A(g7823),.B(g16044));
  AND2 AND2_4627(.VSS(VSS),.VDD(VDD),.Y(g31554),.A(g19050),.B(g29814));
  AND2 AND2_4628(.VSS(VSS),.VDD(VDD),.Y(g30673),.A(g20175),.B(g29814));
  AND2 AND2_4629(.VSS(VSS),.VDD(VDD),.Y(g27256),.A(g25937),.B(g19698));
  AND2 AND2_4630(.VSS(VSS),.VDD(VDD),.Y(g19746),.A(g9816),.B(g17147));
  AND2 AND2_4631(.VSS(VSS),.VDD(VDD),.Y(g28244),.A(g27926),.B(g26715));
  AND2 AND2_4632(.VSS(VSS),.VDD(VDD),.Y(g34183),.A(g33695),.B(g24385));
  AND2 AND2_4633(.VSS(VSS),.VDD(VDD),.Y(g18197),.A(g854),.B(g17821));
  AND2 AND2_4634(.VSS(VSS),.VDD(VDD),.Y(g22017),.A(g5763),.B(g21562));
  AND2 AND2_4635(.VSS(VSS),.VDD(VDD),.Y(g15652),.A(g174),.B(g13437));
  AND2 AND2_4636(.VSS(VSS),.VDD(VDD),.Y(g15804),.A(g3223),.B(g13889));
  AND2 AND2_4637(.VSS(VSS),.VDD(VDD),.Y(g34397),.A(g7673),.B(g34068));
  AND2 AND2_4638(.VSS(VSS),.VDD(VDD),.Y(g25949),.A(g24701),.B(g19559));
  AND2 AND2_4639(.VSS(VSS),.VDD(VDD),.Y(g27280),.A(g9825),.B(g26614));
  AND2 AND2_4640(.VSS(VSS),.VDD(VDD),.Y(g31312),.A(g30136),.B(g27858));
  AND2 AND2_4641(.VSS(VSS),.VDD(VDD),.Y(g29577),.A(g2441),.B(g28946));
  AND2 AND2_4642(.VSS(VSS),.VDD(VDD),.Y(g30062),.A(g13129),.B(g28174));
  AND2 AND2_4643(.VSS(VSS),.VDD(VDD),.Y(g27300),.A(g12370),.B(g26672));
  AND2 AND2_4644(.VSS(VSS),.VDD(VDD),.Y(g10736),.A(g4040),.B(g8751));
  AND3 AND3_264(.VSS(VSS),.VDD(VDD),.Y(g10887),.A(g7812),.B(g6565),.C(g6573));
  AND2 AND2_4645(.VSS(VSS),.VDD(VDD),.Y(g31115),.A(g29487),.B(g22882));
  AND2 AND2_4646(.VSS(VSS),.VDD(VDD),.Y(g18411),.A(g2093),.B(g15373));
  AND2 AND2_4647(.VSS(VSS),.VDD(VDD),.Y(g25536),.A(g23770),.B(g21431));
  AND2 AND2_4648(.VSS(VSS),.VDD(VDD),.Y(g25040),.A(g12738),.B(g23443));
  AND4 AND4_280(.VSS(VSS),.VDD(VDD),.Y(g26213),.A(g25357),.B(g11724),.C(g7586),.D(g7558));
  AND2 AND2_4649(.VSS(VSS),.VDD(VDD),.Y(g34509),.A(g34283),.B(g19473));
  AND2 AND2_4650(.VSS(VSS),.VDD(VDD),.Y(g21850),.A(g3893),.B(g21070));
  AND2 AND2_4651(.VSS(VSS),.VDD(VDD),.Y(g28602),.A(g27509),.B(g20515));
  AND2 AND2_4652(.VSS(VSS),.VDD(VDD),.Y(g23412),.A(g7297),.B(g21510));
  AND2 AND2_4653(.VSS(VSS),.VDD(VDD),.Y(g28657),.A(g27562),.B(g20606));
  AND2 AND2_4654(.VSS(VSS),.VDD(VDD),.Y(g25904),.A(g14001),.B(g24791));
  AND3 AND3_265(.VSS(VSS),.VDD(VDD),.Y(g33921),.A(g33187),.B(g9104),.C(g19200));
  AND2 AND2_4655(.VSS(VSS),.VDD(VDD),.Y(g19684),.A(g2735),.B(g17297));
  AND2 AND2_4656(.VSS(VSS),.VDD(VDD),.Y(g34508),.A(g34282),.B(g19472));
  AND2 AND2_4657(.VSS(VSS),.VDD(VDD),.Y(g10528),.A(g1576),.B(g9051));
  AND2 AND2_4658(.VSS(VSS),.VDD(VDD),.Y(g34872),.A(g34827),.B(g19954));
  AND3 AND3_266(.VSS(VSS),.VDD(VDD),.Y(I18740),.A(g13156),.B(g11450),.C(g11498));
  AND2 AND2_4659(.VSS(VSS),.VDD(VDD),.Y(g24700),.A(g645),.B(g23512));
  AND4 AND4_281(.VSS(VSS),.VDD(VDD),.Y(g28970),.A(g17405),.B(g25196),.C(g26424),.D(g27445));
  AND2 AND2_4660(.VSS(VSS),.VDD(VDD),.Y(g24659),.A(g5134),.B(g23590));
  AND4 AND4_282(.VSS(VSS),.VDD(VDD),.Y(g14528),.A(g12459),.B(g12306),.C(g12245),.D(I16646));
  AND2 AND2_4661(.VSS(VSS),.VDD(VDD),.Y(g26205),.A(g2098),.B(g25492));
  AND2 AND2_4662(.VSS(VSS),.VDD(VDD),.Y(g23229),.A(g18994),.B(g4521));
  AND4 AND4_283(.VSS(VSS),.VDD(VDD),.Y(g16234),.A(g6772),.B(g6782),.C(g11640),.D(I17575));
  AND2 AND2_4663(.VSS(VSS),.VDD(VDD),.Y(g29349),.A(g4760),.B(g28391));
  AND2 AND2_4664(.VSS(VSS),.VDD(VDD),.Y(g22309),.A(g1478),.B(g19751));
  AND2 AND2_4665(.VSS(VSS),.VDD(VDD),.Y(g20658),.A(g1389),.B(g15800));
  AND2 AND2_4666(.VSS(VSS),.VDD(VDD),.Y(g18503),.A(g2563),.B(g15509));
  AND2 AND2_4667(.VSS(VSS),.VDD(VDD),.Y(g22023),.A(g5881),.B(g19147));
  AND2 AND2_4668(.VSS(VSS),.VDD(VDD),.Y(g26311),.A(g2527),.B(g25400));
  AND2 AND2_4669(.VSS(VSS),.VDD(VDD),.Y(g24658),.A(g22645),.B(g19732));
  AND3 AND3_267(.VSS(VSS),.VDD(VDD),.Y(I24015),.A(g8334),.B(g7975),.C(g3045));
  AND3 AND3_268(.VSS(VSS),.VDD(VDD),.Y(g10869),.A(g7766),.B(g5873),.C(g5881));
  AND2 AND2_4670(.VSS(VSS),.VDD(VDD),.Y(g22308),.A(g1135),.B(g19738));
  AND2 AND2_4671(.VSS(VSS),.VDD(VDD),.Y(g28171),.A(g27016),.B(g19385));
  AND2 AND2_4672(.VSS(VSS),.VDD(VDD),.Y(g33798),.A(g33227),.B(g20058));
  AND2 AND2_4673(.VSS(VSS),.VDD(VDD),.Y(g21716),.A(g301),.B(g20283));
  AND2 AND2_4674(.VSS(VSS),.VDD(VDD),.Y(g30213),.A(g28688),.B(g23880));
  AND2 AND2_4675(.VSS(VSS),.VDD(VDD),.Y(g24296),.A(g4382),.B(g22550));
  AND2 AND2_4676(.VSS(VSS),.VDD(VDD),.Y(g18581),.A(g2912),.B(g16349));
  AND2 AND2_4677(.VSS(VSS),.VDD(VDD),.Y(g18714),.A(g4864),.B(g15915));
  AND2 AND2_4678(.VSS(VSS),.VDD(VDD),.Y(g26051),.A(g24896),.B(g14169));
  AND2 AND2_4679(.VSS(VSS),.VDD(VDD),.Y(g18450),.A(g2299),.B(g15224));
  AND2 AND2_4680(.VSS(VSS),.VDD(VDD),.Y(g31184),.A(g1950),.B(g30085));
  AND2 AND2_4681(.VSS(VSS),.VDD(VDD),.Y(g34213),.A(g33766),.B(g22689));
  AND2 AND2_4682(.VSS(VSS),.VDD(VDD),.Y(g18315),.A(g1548),.B(g16931));
  AND2 AND2_4683(.VSS(VSS),.VDD(VDD),.Y(g33805),.A(g33232),.B(g20079));
  AND3 AND3_269(.VSS(VSS),.VDD(VDD),.Y(g33674),.A(g33164),.B(g10710),.C(g22319));
  AND2 AND2_4684(.VSS(VSS),.VDD(VDD),.Y(g24644),.A(g11714),.B(g22903));
  AND2 AND2_4685(.VSS(VSS),.VDD(VDD),.Y(g29622),.A(g2579),.B(g29001));
  AND2 AND2_4686(.VSS(VSS),.VDD(VDD),.Y(g29566),.A(g2307),.B(g28907));
  AND2 AND2_4687(.VSS(VSS),.VDD(VDD),.Y(g18707),.A(g15134),.B(g16782));
  AND2 AND2_4688(.VSS(VSS),.VDD(VDD),.Y(g18819),.A(g6541),.B(g15483));
  AND2 AND2_4689(.VSS(VSS),.VDD(VDD),.Y(g18910),.A(g16227),.B(g16075));
  AND2 AND2_4690(.VSS(VSS),.VDD(VDD),.Y(g18202),.A(g907),.B(g15938));
  AND2 AND2_4691(.VSS(VSS),.VDD(VDD),.Y(g30047),.A(g29109),.B(g9407));
  AND2 AND2_4692(.VSS(VSS),.VDD(VDD),.Y(g18257),.A(g1205),.B(g16897));
  AND2 AND2_4693(.VSS(VSS),.VDD(VDD),.Y(g26780),.A(g4098),.B(g24437));
  AND2 AND2_4694(.VSS(VSS),.VDD(VDD),.Y(g30205),.A(g28671),.B(g23869));
  AND2 AND2_4695(.VSS(VSS),.VDD(VDD),.Y(g32191),.A(g27593),.B(g31376));
  AND2 AND2_4696(.VSS(VSS),.VDD(VDD),.Y(g18818),.A(g15165),.B(g15483));
  AND2 AND2_4697(.VSS(VSS),.VDD(VDD),.Y(g18496),.A(g2537),.B(g15426));
  AND2 AND2_4698(.VSS(VSS),.VDD(VDD),.Y(g34205),.A(g33729),.B(g24541));
  AND2 AND2_4699(.VSS(VSS),.VDD(VDD),.Y(g31934),.A(g31670),.B(g18827));
  AND2 AND2_4700(.VSS(VSS),.VDD(VDD),.Y(g18111),.A(g174),.B(g17015));
  AND2 AND2_4701(.VSS(VSS),.VDD(VDD),.Y(g21959),.A(g5413),.B(g21514));
  AND2 AND2_4702(.VSS(VSS),.VDD(VDD),.Y(g21925),.A(g5073),.B(g21468));
  AND2 AND2_4703(.VSS(VSS),.VDD(VDD),.Y(g26350),.A(g13087),.B(g25517));
  AND2 AND2_4704(.VSS(VSS),.VDD(VDD),.Y(g25872),.A(g3119),.B(g24655));
  AND2 AND2_4705(.VSS(VSS),.VDD(VDD),.Y(g28919),.A(g27663),.B(g21295));
  AND2 AND2_4706(.VSS(VSS),.VDD(VDD),.Y(g14708),.A(g74),.B(g12369));
  AND3 AND3_270(.VSS(VSS),.VDD(VDD),.Y(I18762),.A(g13156),.B(g6767),.C(g11498));
  AND4 AND4_284(.VSS(VSS),.VDD(VDD),.Y(g28458),.A(g27187),.B(g12730),.C(g20887),.D(I26948));
  AND2 AND2_4707(.VSS(VSS),.VDD(VDD),.Y(g24197),.A(g347),.B(g22722));
  AND3 AND3_271(.VSS(VSS),.VDD(VDD),.Y(g24855),.A(g3050),.B(g23534),.C(I24027));
  AND3 AND3_272(.VSS(VSS),.VDD(VDD),.Y(g27660),.A(g24688),.B(g26424),.C(g22763));
  AND2 AND2_4708(.VSS(VSS),.VDD(VDD),.Y(g16163),.A(g14254),.B(g14179));
  AND2 AND2_4709(.VSS(VSS),.VDD(VDD),.Y(g22752),.A(g15792),.B(g19612));
  AND2 AND2_4710(.VSS(VSS),.VDD(VDD),.Y(g15613),.A(g3490),.B(g13555));
  AND2 AND2_4711(.VSS(VSS),.VDD(VDD),.Y(g18590),.A(g2917),.B(g16349));
  AND2 AND2_4712(.VSS(VSS),.VDD(VDD),.Y(g21958),.A(g5396),.B(g21514));
  AND2 AND2_4713(.VSS(VSS),.VDD(VDD),.Y(g21378),.A(g7887),.B(g16090));
  AND2 AND2_4714(.VSS(VSS),.VDD(VDD),.Y(g23050),.A(g655),.B(g20248));
  AND4 AND4_285(.VSS(VSS),.VDD(VDD),.Y(g28010),.A(g23032),.B(g26223),.C(g26424),.D(g25535));
  AND2 AND2_4715(.VSS(VSS),.VDD(VDD),.Y(g23958),.A(g9104),.B(g19200));
  AND2 AND2_4716(.VSS(VSS),.VDD(VDD),.Y(g24411),.A(g4584),.B(g22161));
  AND2 AND2_4717(.VSS(VSS),.VDD(VDD),.Y(g30051),.A(g28513),.B(g20604));
  AND2 AND2_4718(.VSS(VSS),.VDD(VDD),.Y(g26846),.A(g37),.B(g24524));
  AND2 AND2_4719(.VSS(VSS),.VDD(VDD),.Y(g18741),.A(g15143),.B(g17384));
  AND2 AND2_4720(.VSS(VSS),.VDD(VDD),.Y(g34072),.A(g33839),.B(g24872));
  AND2 AND2_4721(.VSS(VSS),.VDD(VDD),.Y(g23386),.A(g20034),.B(g20207));
  AND2 AND2_4722(.VSS(VSS),.VDD(VDD),.Y(g30592),.A(g30270),.B(g18929));
  AND2 AND2_4723(.VSS(VSS),.VDD(VDD),.Y(g18384),.A(g1945),.B(g15171));
  AND2 AND2_4724(.VSS(VSS),.VDD(VDD),.Y(g29636),.A(g2403),.B(g29097));
  AND2 AND2_4725(.VSS(VSS),.VDD(VDD),.Y(g21742),.A(g3050),.B(g20330));
  AND2 AND2_4726(.VSS(VSS),.VDD(VDD),.Y(g17752),.A(g7841),.B(g13174));
  AND2 AND2_4727(.VSS(VSS),.VDD(VDD),.Y(g27480),.A(g26400),.B(g17638));
  AND2 AND2_4728(.VSS(VSS),.VDD(VDD),.Y(g34756),.A(g34680),.B(g19618));
  AND2 AND2_4729(.VSS(VSS),.VDD(VDD),.Y(g23742),.A(g19128),.B(g9104));
  AND2 AND2_4730(.VSS(VSS),.VDD(VDD),.Y(g28599),.A(g27027),.B(g8922));
  AND2 AND2_4731(.VSS(VSS),.VDD(VDD),.Y(g21944),.A(g5244),.B(g18997));
  AND2 AND2_4732(.VSS(VSS),.VDD(VDD),.Y(g33400),.A(g32347),.B(g21380));
  AND2 AND2_4733(.VSS(VSS),.VDD(VDD),.Y(g29852),.A(g1772),.B(g29080));
  AND2 AND2_4734(.VSS(VSS),.VDD(VDD),.Y(g17643),.A(g9681),.B(g14599));
  AND2 AND2_4735(.VSS(VSS),.VDD(VDD),.Y(g15812),.A(g3227),.B(g13915));
  AND4 AND4_286(.VSS(VSS),.VDD(VDD),.Y(g13319),.A(g4076),.B(g8812),.C(g10658),.D(g8757));
  AND2 AND2_4736(.VSS(VSS),.VDD(VDD),.Y(g27314),.A(g12436),.B(g26702));
  AND2 AND2_4737(.VSS(VSS),.VDD(VDD),.Y(g24503),.A(g22225),.B(g19409));
  AND2 AND2_4738(.VSS(VSS),.VDD(VDD),.Y(g27287),.A(g26545),.B(g23011));
  AND2 AND2_4739(.VSS(VSS),.VDD(VDD),.Y(g32045),.A(g31491),.B(g16187));
  AND4 AND4_287(.VSS(VSS),.VDD(VDD),.Y(I24685),.A(g24036),.B(g24037),.C(g24038),.D(g24039));
  AND2 AND2_4740(.VSS(VSS),.VDD(VDD),.Y(g33329),.A(g32210),.B(g20585));
  AND2 AND2_4741(.VSS(VSS),.VDD(VDD),.Y(g31207),.A(g30252),.B(g20739));
  AND2 AND2_4742(.VSS(VSS),.VDD(VDD),.Y(g18150),.A(g604),.B(g17533));
  AND2 AND2_4743(.VSS(VSS),.VDD(VDD),.Y(g10657),.A(g8451),.B(g4064));
  AND2 AND2_4744(.VSS(VSS),.VDD(VDD),.Y(g18801),.A(g15160),.B(g15348));
  AND2 AND2_4745(.VSS(VSS),.VDD(VDD),.Y(g18735),.A(g4983),.B(g16826));
  AND2 AND2_4746(.VSS(VSS),.VDD(VDD),.Y(g25574),.A(I24709),.B(I24710));
  AND2 AND2_4747(.VSS(VSS),.VDD(VDD),.Y(g27085),.A(g25835),.B(g22494));
  AND2 AND2_4748(.VSS(VSS),.VDD(VDD),.Y(g32324),.A(g31315),.B(g23537));
  AND2 AND2_4749(.VSS(VSS),.VDD(VDD),.Y(g29664),.A(g2273),.B(g29060));
  AND2 AND2_4750(.VSS(VSS),.VDD(VDD),.Y(g33328),.A(g32209),.B(g20584));
  AND2 AND2_4751(.VSS(VSS),.VDD(VDD),.Y(g21802),.A(g3562),.B(g20924));
  AND2 AND2_4752(.VSS(VSS),.VDD(VDD),.Y(g22489),.A(g12954),.B(g19386));
  AND2 AND2_4753(.VSS(VSS),.VDD(VDD),.Y(g21857),.A(g3933),.B(g21070));
  AND2 AND2_4754(.VSS(VSS),.VDD(VDD),.Y(g23802),.A(g9104),.B(g19050));
  AND2 AND2_4755(.VSS(VSS),.VDD(VDD),.Y(g16535),.A(g5595),.B(g14848));
  AND2 AND2_4756(.VSS(VSS),.VDD(VDD),.Y(g20581),.A(g10801),.B(g15571));
  AND2 AND2_4757(.VSS(VSS),.VDD(VDD),.Y(g10970),.A(g854),.B(g9582));
  AND2 AND2_4758(.VSS(VSS),.VDD(VDD),.Y(g23857),.A(g19626),.B(g7908));
  AND2 AND2_4759(.VSS(VSS),.VDD(VDD),.Y(g13059),.A(g6900),.B(g11303));
  AND2 AND2_4760(.VSS(VSS),.VDD(VDD),.Y(g13025),.A(g8431),.B(g11026));
  AND2 AND2_4761(.VSS(VSS),.VDD(VDD),.Y(g30152),.A(g28609),.B(g23767));
  AND2 AND2_4762(.VSS(VSS),.VDD(VDD),.Y(g24581),.A(g5124),.B(g23590));
  AND2 AND2_4763(.VSS(VSS),.VDD(VDD),.Y(g24714),.A(g6173),.B(g23699));
  AND2 AND2_4764(.VSS(VSS),.VDD(VDD),.Y(g32098),.A(g4732),.B(g30614));
  AND2 AND2_4765(.VSS(VSS),.VDD(VDD),.Y(g24450),.A(g3129),.B(g23067));
  AND2 AND2_4766(.VSS(VSS),.VDD(VDD),.Y(g21730),.A(g3025),.B(g20330));
  AND2 AND2_4767(.VSS(VSS),.VDD(VDD),.Y(g24315),.A(g4521),.B(g22228));
  AND2 AND2_4768(.VSS(VSS),.VDD(VDD),.Y(g21793),.A(g3412),.B(g20391));
  AND2 AND2_4769(.VSS(VSS),.VDD(VDD),.Y(g32272),.A(g31639),.B(g30310));
  AND2 AND2_4770(.VSS(VSS),.VDD(VDD),.Y(g22525),.A(g13006),.B(g19411));
  AND2 AND2_4771(.VSS(VSS),.VDD(VDD),.Y(g28159),.A(g8553),.B(g27317));
  AND4 AND4_288(.VSS(VSS),.VDD(VDD),.Y(I31262),.A(g32833),.B(g32834),.C(g32835),.D(g32836));
  AND2 AND2_4772(.VSS(VSS),.VDD(VDD),.Y(g10878),.A(g7858),.B(g1135));
  AND2 AND2_4773(.VSS(VSS),.VDD(VDD),.Y(g18196),.A(g703),.B(g17821));
  AND2 AND2_4774(.VSS(VSS),.VDD(VDD),.Y(g22016),.A(g5747),.B(g21562));
  AND2 AND2_4775(.VSS(VSS),.VDD(VDD),.Y(g28125),.A(g27381),.B(g26209));
  AND2 AND2_4776(.VSS(VSS),.VDD(VDD),.Y(g15795),.A(g3566),.B(g14130));
  AND2 AND2_4777(.VSS(VSS),.VDD(VDD),.Y(g18695),.A(g4737),.B(g16053));
  AND2 AND2_4778(.VSS(VSS),.VDD(VDD),.Y(g28532),.A(g27394),.B(g20265));
  AND2 AND2_4779(.VSS(VSS),.VDD(VDD),.Y(g34396),.A(g34194),.B(g21337));
  AND3 AND3_273(.VSS(VSS),.VDD(VDD),.Y(I18568),.A(g13156),.B(g11450),.C(g11498));
  AND2 AND2_4780(.VSS(VSS),.VDD(VDD),.Y(g24707),.A(g13295),.B(g22997));
  AND2 AND2_4781(.VSS(VSS),.VDD(VDD),.Y(g30731),.A(g11374),.B(g29361));
  AND2 AND2_4782(.VSS(VSS),.VDD(VDD),.Y(g29576),.A(g2177),.B(g28903));
  AND2 AND2_4783(.VSS(VSS),.VDD(VDD),.Y(g29585),.A(g1756),.B(g28920));
  AND2 AND2_4784(.VSS(VSS),.VDD(VDD),.Y(g21765),.A(g3231),.B(g20785));
  AND3 AND3_274(.VSS(VSS),.VDD(VDD),.Y(g28158),.A(g26424),.B(g22763),.C(g27037));
  AND4 AND4_289(.VSS(VSS),.VDD(VDD),.Y(I27523),.A(g20857),.B(g24111),.C(g24112),.D(g24113));
  AND2 AND2_4785(.VSS(VSS),.VDD(VDD),.Y(g18526),.A(g2555),.B(g15509));
  AND2 AND2_4786(.VSS(VSS),.VDD(VDD),.Y(g27269),.A(g25943),.B(g19734));
  AND2 AND2_4787(.VSS(VSS),.VDD(VDD),.Y(g29554),.A(g28997),.B(g22472));
  AND2 AND2_4788(.VSS(VSS),.VDD(VDD),.Y(g23690),.A(g14726),.B(g20978));
  AND2 AND2_4789(.VSS(VSS),.VDD(VDD),.Y(g19372),.A(g686),.B(g16289));
  AND2 AND2_4790(.VSS(VSS),.VDD(VDD),.Y(g26020),.A(g9559),.B(g25034));
  AND2 AND2_4791(.VSS(VSS),.VDD(VDD),.Y(g33241),.A(g32173),.B(g23128));
  AND2 AND2_4792(.VSS(VSS),.VDD(VDD),.Y(g34413),.A(g34094),.B(g22670));
  AND2 AND2_4793(.VSS(VSS),.VDD(VDD),.Y(g17424),.A(g1426),.B(g13176));
  AND2 AND2_4794(.VSS(VSS),.VDD(VDD),.Y(g11044),.A(g5343),.B(g10124));
  AND4 AND4_290(.VSS(VSS),.VDD(VDD),.Y(I31191),.A(g30735),.B(g31829),.C(g32731),.D(g32732));
  AND2 AND2_4795(.VSS(VSS),.VDD(VDD),.Y(g27341),.A(g10203),.B(g26788));
  AND2 AND2_4796(.VSS(VSS),.VDD(VDD),.Y(g10967),.A(g7880),.B(g1448));
  AND2 AND2_4797(.VSS(VSS),.VDD(VDD),.Y(g29609),.A(g28482),.B(g11861));
  AND2 AND2_4798(.VSS(VSS),.VDD(VDD),.Y(g27268),.A(g25942),.B(g19733));
  AND2 AND2_4799(.VSS(VSS),.VDD(VDD),.Y(g32032),.A(g31373),.B(g16515));
  AND2 AND2_4800(.VSS(VSS),.VDD(VDD),.Y(g25780),.A(g25532),.B(g25527));
  AND2 AND2_4801(.VSS(VSS),.VDD(VDD),.Y(g15507),.A(g10970),.B(g13305));
  AND2 AND2_4802(.VSS(VSS),.VDD(VDD),.Y(g32140),.A(g31609),.B(g29961));
  AND2 AND2_4803(.VSS(VSS),.VDD(VDD),.Y(g28144),.A(g4608),.B(g27020));
  AND2 AND2_4804(.VSS(VSS),.VDD(VDD),.Y(g18402),.A(g2047),.B(g15373));
  AND2 AND2_4805(.VSS(VSS),.VDD(VDD),.Y(g18457),.A(g2319),.B(g15224));
  AND2 AND2_4806(.VSS(VSS),.VDD(VDD),.Y(g24590),.A(g6154),.B(g23413));
  AND2 AND2_4807(.VSS(VSS),.VDD(VDD),.Y(g29608),.A(g28568),.B(g11385));
  AND2 AND2_4808(.VSS(VSS),.VDD(VDD),.Y(g27180),.A(g26026),.B(g16654));
  AND2 AND2_4809(.VSS(VSS),.VDD(VDD),.Y(g19516),.A(g7824),.B(g16097));
  AND2 AND2_4810(.VSS(VSS),.VDD(VDD),.Y(g20094),.A(g8872),.B(g16631));
  AND2 AND2_4811(.VSS(VSS),.VDD(VDD),.Y(g27335),.A(g12087),.B(g26776));
  AND3 AND3_275(.VSS(VSS),.VDD(VDD),.Y(g33683),.A(g33149),.B(g10727),.C(g22332));
  AND2 AND2_4812(.VSS(VSS),.VDD(VDD),.Y(g13738),.A(g8880),.B(g10572));
  AND2 AND2_4813(.VSS(VSS),.VDD(VDD),.Y(g25152),.A(g23383),.B(g20626));
  AND2 AND2_4814(.VSS(VSS),.VDD(VDD),.Y(g22042),.A(g5961),.B(g19147));
  AND2 AND2_4815(.VSS(VSS),.VDD(VDD),.Y(g26302),.A(g2393),.B(g25349));
  AND2 AND2_4816(.VSS(VSS),.VDD(VDD),.Y(g26357),.A(g22547),.B(g25525));
  AND2 AND2_4817(.VSS(VSS),.VDD(VDD),.Y(g29799),.A(g28271),.B(g10233));
  AND2 AND2_4818(.VSS(VSS),.VDD(VDD),.Y(g30583),.A(g19666),.B(g29355));
  AND2 AND2_4819(.VSS(VSS),.VDD(VDD),.Y(g16760),.A(g5559),.B(g14764));
  AND2 AND2_4820(.VSS(VSS),.VDD(VDD),.Y(g27667),.A(g26361),.B(g20601));
  AND4 AND4_291(.VSS(VSS),.VDD(VDD),.Y(I31247),.A(g32812),.B(g32813),.C(g32814),.D(g32815));
  AND2 AND2_4821(.VSS(VSS),.VDD(VDD),.Y(g18706),.A(g4785),.B(g16782));
  AND2 AND2_4822(.VSS(VSS),.VDD(VDD),.Y(g18597),.A(g2975),.B(g16349));
  AND2 AND2_4823(.VSS(VSS),.VDD(VDD),.Y(g27965),.A(g25834),.B(g13117));
  AND2 AND2_4824(.VSS(VSS),.VDD(VDD),.Y(g13290),.A(g3897),.B(g11534));
  AND2 AND2_4825(.VSS(VSS),.VDD(VDD),.Y(g29798),.A(g28348),.B(g23260));
  AND2 AND2_4826(.VSS(VSS),.VDD(VDD),.Y(g22124),.A(g6613),.B(g19277));
  AND2 AND2_4827(.VSS(VSS),.VDD(VDD),.Y(g27131),.A(g26055),.B(g16588));
  AND2 AND2_4828(.VSS(VSS),.VDD(VDD),.Y(g30046),.A(g29108),.B(g10564));
  AND2 AND2_4829(.VSS(VSS),.VDD(VDD),.Y(g18256),.A(g1242),.B(g16897));
  AND2 AND2_4830(.VSS(VSS),.VDD(VDD),.Y(g29973),.A(g28981),.B(g9206));
  AND2 AND2_4831(.VSS(VSS),.VDD(VDD),.Y(g18689),.A(g15129),.B(g16752));
  AND2 AND2_4832(.VSS(VSS),.VDD(VDD),.Y(g31991),.A(g4912),.B(g30673));
  AND3 AND3_276(.VSS(VSS),.VDD(VDD),.Y(g33515),.A(g32853),.B(I31271),.C(I31272));
  AND2 AND2_4833(.VSS(VSS),.VDD(VDD),.Y(g33882),.A(g33293),.B(g20587));
  AND2 AND2_4834(.VSS(VSS),.VDD(VDD),.Y(g18280),.A(g1367),.B(g16136));
  AND2 AND2_4835(.VSS(VSS),.VDD(VDD),.Y(g29805),.A(g28357),.B(g23270));
  AND2 AND2_4836(.VSS(VSS),.VDD(VDD),.Y(g33414),.A(g32367),.B(g21421));
  AND2 AND2_4837(.VSS(VSS),.VDD(VDD),.Y(g22686),.A(g19335),.B(g19577));
  AND2 AND2_4838(.VSS(VSS),.VDD(VDD),.Y(g22939),.A(g9708),.B(g21062));
  AND2 AND2_4839(.VSS(VSS),.VDD(VDD),.Y(g18688),.A(g4704),.B(g16752));
  AND2 AND2_4840(.VSS(VSS),.VDD(VDD),.Y(g18624),.A(g3490),.B(g17062));
  AND2 AND2_4841(.VSS(VSS),.VDD(VDD),.Y(g32162),.A(g31002),.B(g23014));
  AND2 AND2_4842(.VSS(VSS),.VDD(VDD),.Y(g18300),.A(g1306),.B(g16489));
  AND2 AND2_4843(.VSS(VSS),.VDD(VDD),.Y(g24196),.A(g333),.B(g22722));
  AND2 AND2_4844(.VSS(VSS),.VDD(VDD),.Y(g33407),.A(g32357),.B(g21406));
  AND2 AND2_4845(.VSS(VSS),.VDD(VDD),.Y(g34113),.A(g33734),.B(g19744));
  AND2 AND2_4846(.VSS(VSS),.VDD(VDD),.Y(g27502),.A(g26488),.B(g17677));
  AND4 AND4_292(.VSS(VSS),.VDD(VDD),.Y(I31251),.A(g31710),.B(g31840),.C(g32817),.D(g32818));
  AND2 AND2_4847(.VSS(VSS),.VDD(VDD),.Y(g11427),.A(g5706),.B(g7158));
  AND2 AND2_4848(.VSS(VSS),.VDD(VDD),.Y(g22030),.A(g5909),.B(g19147));
  AND4 AND4_293(.VSS(VSS),.VDD(VDD),.Y(I31272),.A(g32849),.B(g32850),.C(g32851),.D(g32852));
  AND2 AND2_4849(.VSS(VSS),.VDD(VDD),.Y(g22938),.A(g19782),.B(g19739));
  AND2 AND2_4850(.VSS(VSS),.VDD(VDD),.Y(g27557),.A(g26549),.B(g17774));
  AND2 AND2_4851(.VSS(VSS),.VDD(VDD),.Y(g22093),.A(g6423),.B(g18833));
  AND2 AND2_4852(.VSS(VSS),.VDD(VDD),.Y(g23533),.A(g19436),.B(g13015));
  AND2 AND2_4853(.VSS(VSS),.VDD(VDD),.Y(g11366),.A(g5016),.B(g10338));
  AND3 AND3_277(.VSS(VSS),.VDD(VDD),.Y(g27210),.A(g26218),.B(g8373),.C(g2476));
  AND2 AND2_4854(.VSS(VSS),.VDD(VDD),.Y(g21298),.A(g7697),.B(g15825));
  AND2 AND2_4855(.VSS(VSS),.VDD(VDD),.Y(g29732),.A(g2514),.B(g29131));
  AND2 AND2_4856(.VSS(VSS),.VDD(VDD),.Y(g28289),.A(g27734),.B(g26575));
  AND2 AND2_4857(.VSS(VSS),.VDD(VDD),.Y(g21775),.A(g3372),.B(g20391));
  AND3 AND3_278(.VSS(VSS),.VDD(VDD),.Y(I16671),.A(g10185),.B(g12461),.C(g12415));
  AND2 AND2_4858(.VSS(VSS),.VDD(VDD),.Y(g13632),.A(g10232),.B(g12228));
  AND2 AND2_4859(.VSS(VSS),.VDD(VDD),.Y(g18157),.A(g15057),.B(g17433));
  AND2 AND2_4860(.VSS(VSS),.VDD(VDD),.Y(g23775),.A(g14872),.B(g21267));
  AND2 AND2_4861(.VSS(VSS),.VDD(VDD),.Y(g22065),.A(g6203),.B(g19210));
  AND3 AND3_279(.VSS(VSS),.VDD(VDD),.Y(g34105),.A(g33778),.B(g9104),.C(g18957));
  AND3 AND3_280(.VSS(VSS),.VDD(VDD),.Y(g28224),.A(g27163),.B(g22763),.C(g27064));
  AND2 AND2_4862(.VSS(VSS),.VDD(VDD),.Y(g34743),.A(g8951),.B(g34703));
  AND3 AND3_281(.VSS(VSS),.VDD(VDD),.Y(I17585),.A(g14988),.B(g11450),.C(g11498));
  AND2 AND2_4863(.VSS(VSS),.VDD(VDD),.Y(g28571),.A(g27458),.B(g20435));
  AND2 AND2_4864(.VSS(VSS),.VDD(VDD),.Y(g24402),.A(g4749),.B(g22857));
  AND2 AND2_4865(.VSS(VSS),.VDD(VDD),.Y(g29761),.A(g28310),.B(g23228));
  AND4 AND4_294(.VSS(VSS),.VDD(VDD),.Y(I31032),.A(g32501),.B(g32502),.C(g32503),.D(g32504));
  AND2 AND2_4866(.VSS(VSS),.VDD(VDD),.Y(g18231),.A(g1105),.B(g16326));
  AND2 AND2_4867(.VSS(VSS),.VDD(VDD),.Y(g21737),.A(g3068),.B(g20330));
  AND2 AND2_4868(.VSS(VSS),.VDD(VDD),.Y(g32246),.A(g31246),.B(g20326));
  AND4 AND4_295(.VSS(VSS),.VDD(VDD),.Y(g27469),.A(g8046),.B(g26314),.C(g518),.D(g9077));
  AND2 AND2_4869(.VSS(VSS),.VDD(VDD),.Y(g22219),.A(g19953),.B(g20887));
  AND2 AND2_4870(.VSS(VSS),.VDD(VDD),.Y(g25928),.A(g25022),.B(g23436));
  AND2 AND2_4871(.VSS(VSS),.VDD(VDD),.Y(g8583),.A(g2917),.B(g2912));
  AND2 AND2_4872(.VSS(VSS),.VDD(VDD),.Y(g27286),.A(g6856),.B(g26634));
  AND2 AND2_4873(.VSS(VSS),.VDD(VDD),.Y(g33441),.A(g32251),.B(g29722));
  AND2 AND2_4874(.VSS(VSS),.VDD(VDD),.Y(g31206),.A(g30260),.B(g23890));
  AND2 AND2_4875(.VSS(VSS),.VDD(VDD),.Y(g10656),.A(g3782),.B(g7952));
  AND4 AND4_296(.VSS(VSS),.VDD(VDD),.Y(g27039),.A(g7738),.B(g5527),.C(g5535),.D(g26223));
  AND2 AND2_4876(.VSS(VSS),.VDD(VDD),.Y(g22218),.A(g19951),.B(g20875));
  AND2 AND2_4877(.VSS(VSS),.VDD(VDD),.Y(g28495),.A(g27012),.B(g12465));
  AND2 AND2_4878(.VSS(VSS),.VDD(VDD),.Y(g32071),.A(g27236),.B(g31070));
  AND4 AND4_297(.VSS(VSS),.VDD(VDD),.Y(I31061),.A(g30825),.B(g31806),.C(g32543),.D(g32544));
  AND2 AND2_4879(.VSS(VSS),.VDD(VDD),.Y(g21856),.A(g3929),.B(g21070));
  AND3 AND3_282(.VSS(VSS),.VDD(VDD),.Y(g10823),.A(g7704),.B(g5180),.C(g5188));
  AND2 AND2_4880(.VSS(VSS),.VDD(VDD),.Y(g14295),.A(g1811),.B(g11894));
  AND2 AND2_4881(.VSS(VSS),.VDD(VDD),.Y(g21995),.A(g5611),.B(g19074));
  AND2 AND2_4882(.VSS(VSS),.VDD(VDD),.Y(g31759),.A(g21291),.B(g29385));
  AND2 AND2_4883(.VSS(VSS),.VDD(VDD),.Y(g23856),.A(g4116),.B(g19483));
  AND2 AND2_4884(.VSS(VSS),.VDD(VDD),.Y(g14680),.A(g12024),.B(g12053));
  AND2 AND2_4885(.VSS(VSS),.VDD(VDD),.Y(g33759),.A(g33123),.B(g22847));
  AND3 AND3_283(.VSS(VSS),.VDD(VDD),.Y(g33725),.A(g22626),.B(g10851),.C(g33176));
  AND2 AND2_4886(.VSS(VSS),.VDD(VDD),.Y(g24001),.A(g19651),.B(g10951));
  AND2 AND2_4887(.VSS(VSS),.VDD(VDD),.Y(g21880),.A(g4135),.B(g19801));
  AND2 AND2_4888(.VSS(VSS),.VDD(VDD),.Y(g29329),.A(g7995),.B(g28353));
  AND2 AND2_4889(.VSS(VSS),.VDD(VDD),.Y(g25113),.A(g23346),.B(g20577));
  AND2 AND2_4890(.VSS(VSS),.VDD(VDD),.Y(g18511),.A(g2599),.B(g15509));
  AND3 AND3_284(.VSS(VSS),.VDD(VDD),.Y(g29207),.A(g24131),.B(I27533),.C(I27534));
  AND2 AND2_4891(.VSS(VSS),.VDD(VDD),.Y(g25787),.A(g24792),.B(g20887));
  AND2 AND2_4892(.VSS(VSS),.VDD(VDD),.Y(g32147),.A(g31616),.B(g29980));
  AND2 AND2_4893(.VSS(VSS),.VDD(VDD),.Y(g18763),.A(g5481),.B(g17929));
  AND2 AND2_4894(.VSS(VSS),.VDD(VDD),.Y(g31758),.A(g30115),.B(g23945));
  AND2 AND2_4895(.VSS(VSS),.VDD(VDD),.Y(g33114),.A(g22139),.B(g31945));
  AND2 AND2_4896(.VSS(VSS),.VDD(VDD),.Y(g24706),.A(g15910),.B(g22996));
  AND2 AND2_4897(.VSS(VSS),.VDD(VDD),.Y(g26249),.A(g1858),.B(g25300));
  AND2 AND2_4898(.VSS(VSS),.VDD(VDD),.Y(g33758),.A(g33133),.B(g20269));
  AND2 AND2_4899(.VSS(VSS),.VDD(VDD),.Y(g22160),.A(g8005),.B(g19795));
  AND2 AND2_4900(.VSS(VSS),.VDD(VDD),.Y(g27601),.A(g26766),.B(g26737));
  AND2 AND2_4901(.VSS(VSS),.VDD(VDD),.Y(g33082),.A(g32389),.B(g18877));
  AND2 AND2_4902(.VSS(VSS),.VDD(VDD),.Y(g21512),.A(g16225),.B(g10881));
  AND3 AND3_285(.VSS(VSS),.VDD(VDD),.Y(g29328),.A(g28553),.B(g6928),.C(g3990));
  AND2 AND2_4903(.VSS(VSS),.VDD(VDD),.Y(g27677),.A(g13021),.B(g25888));
  AND2 AND2_4904(.VSS(VSS),.VDD(VDD),.Y(g25357),.A(g23810),.B(g23786));
  AND2 AND2_4905(.VSS(VSS),.VDD(VDD),.Y(g29538),.A(g2563),.B(g28914));
  AND2 AND2_4906(.VSS(VSS),.VDD(VDD),.Y(g11127),.A(g6479),.B(g10022));
  AND2 AND2_4907(.VSS(VSS),.VDD(VDD),.Y(g24923),.A(g23129),.B(g20167));
  AND2 AND2_4908(.VSS(VSS),.VDD(VDD),.Y(g25105),.A(g13973),.B(g23505));
  AND2 AND2_4909(.VSS(VSS),.VDD(VDD),.Y(g10966),.A(g9226),.B(g7948));
  AND2 AND2_4910(.VSS(VSS),.VDD(VDD),.Y(g31744),.A(g30092),.B(g23902));
  AND2 AND2_4911(.VSS(VSS),.VDD(VDD),.Y(g24688),.A(g22681),.B(g22663));
  AND2 AND2_4912(.VSS(VSS),.VDD(VDD),.Y(g26204),.A(g1720),.B(g25275));
  AND2 AND2_4913(.VSS(VSS),.VDD(VDD),.Y(g24624),.A(g16524),.B(g22867));
  AND2 AND2_4914(.VSS(VSS),.VDD(VDD),.Y(g24300),.A(g15123),.B(g22228));
  AND3 AND3_286(.VSS(VSS),.VDD(VDD),.Y(I24579),.A(g5731),.B(g5736),.C(g9875));
  AND2 AND2_4915(.VSS(VSS),.VDD(VDD),.Y(g26779),.A(g24497),.B(g23620));
  AND2 AND2_4916(.VSS(VSS),.VDD(VDD),.Y(g33345),.A(g32229),.B(g20671));
  AND2 AND2_4917(.VSS(VSS),.VDD(VDD),.Y(g32151),.A(g31639),.B(g29996));
  AND2 AND2_4918(.VSS(VSS),.VDD(VDD),.Y(g32172),.A(g2767),.B(g31608));
  AND4 AND4_298(.VSS(VSS),.VDD(VDD),.Y(I31162),.A(g32689),.B(g32690),.C(g32691),.D(g32692));
  AND2 AND2_4919(.VSS(VSS),.VDD(VDD),.Y(g31940),.A(g943),.B(g30735));
  AND2 AND2_4920(.VSS(VSS),.VDD(VDD),.Y(g18456),.A(g2338),.B(g15224));
  AND2 AND2_4921(.VSS(VSS),.VDD(VDD),.Y(g33849),.A(g33262),.B(g20387));
  AND2 AND2_4922(.VSS(VSS),.VDD(VDD),.Y(g30027),.A(g29104),.B(g12550));
  AND2 AND2_4923(.VSS(VSS),.VDD(VDD),.Y(g33399),.A(g32346),.B(g21379));
  AND2 AND2_4924(.VSS(VSS),.VDD(VDD),.Y(g21831),.A(g3782),.B(g20453));
  AND2 AND2_4925(.VSS(VSS),.VDD(VDD),.Y(g26778),.A(g25501),.B(g20923));
  AND2 AND2_4926(.VSS(VSS),.VDD(VDD),.Y(g34662),.A(g34576),.B(g18931));
  AND2 AND2_4927(.VSS(VSS),.VDD(VDD),.Y(g16845),.A(g6593),.B(g15011));
  AND2 AND2_4928(.VSS(VSS),.VDD(VDD),.Y(g11956),.A(g2070),.B(g7411));
  AND2 AND2_4929(.VSS(VSS),.VDD(VDD),.Y(g18480),.A(g2437),.B(g15426));
//
  OR2 OR2_0(.VSS(VSS),.VDD(VDD),.Y(g32367),.A(g29880),.B(g31309));
  OR2 OR2_1(.VSS(VSS),.VDD(VDD),.Y(g34890),.A(g34863),.B(g21674));
  OR2 OR2_2(.VSS(VSS),.VDD(VDD),.Y(g28668),.A(g27411),.B(g16617));
  OR2 OR2_3(.VSS(VSS),.VDD(VDD),.Y(g34249),.A(g34110),.B(g21702));
  OR2 OR2_4(.VSS(VSS),.VDD(VDD),.Y(g13095),.A(g11374),.B(g1287));
  OR2 OR2_5(.VSS(VSS),.VDD(VDD),.Y(g30482),.A(g30230),.B(g21978));
  OR2 OR2_6(.VSS(VSS),.VDD(VDD),.Y(g24231),.A(g22589),.B(g18201));
  OR2 OR2_7(.VSS(VSS),.VDD(VDD),.Y(g13888),.A(g2941),.B(g11691));
  OR2 OR2_8(.VSS(VSS),.VDD(VDD),.Y(g26945),.A(g26379),.B(g24283));
  OR2 OR2_9(.VSS(VSS),.VDD(VDD),.Y(g30552),.A(g30283),.B(g22123));
  OR2 OR2_10(.VSS(VSS),.VDD(VDD),.Y(g34003),.A(g33866),.B(g18452));
  OR2 OR2_11(.VSS(VSS),.VDD(VDD),.Y(g23989),.A(g20581),.B(g17179));
  OR2 OR2_12(.VSS(VSS),.VDD(VDD),.Y(g29235),.A(g28110),.B(g18260));
  OR2 OR2_13(.VSS(VSS),.VDD(VDD),.Y(g28525),.A(g27284),.B(g26176));
  OR2 OR2_14(.VSS(VSS),.VDD(VDD),.Y(g34204),.A(g33832),.B(g33833));
  OR4 OR4_0(.VSS(VSS),.VDD(VDD),.Y(I28566),.A(g29201),.B(g29202),.C(g29203),.D(g28035));
  OR2 OR2_15(.VSS(VSS),.VDD(VDD),.Y(g14309),.A(g10320),.B(g11048));
  OR4 OR4_1(.VSS(VSS),.VDD(VDD),.Y(I30330),.A(g29385),.B(g31376),.C(g30735),.D(g30825));
  OR2 OR2_16(.VSS(VSS),.VDD(VDD),.Y(g24854),.A(g21453),.B(g24002));
  OR2 OR2_17(.VSS(VSS),.VDD(VDD),.Y(g30081),.A(g28454),.B(g11366));
  OR2 OR2_18(.VSS(VSS),.VDD(VDD),.Y(g32227),.A(g31146),.B(g29648));
  OR2 OR2_19(.VSS(VSS),.VDD(VDD),.Y(g33962),.A(g33822),.B(g18123));
  OR2 OR2_20(.VSS(VSS),.VDD(VDD),.Y(g19575),.A(g15693),.B(g13042));
  OR2 OR2_21(.VSS(VSS),.VDD(VDD),.Y(g27556),.A(g26097),.B(g24687));
  OR2 OR2_22(.VSS(VSS),.VDD(VDD),.Y(g25662),.A(g24656),.B(g21787));
  OR2 OR2_23(.VSS(VSS),.VDD(VDD),.Y(g28544),.A(g27300),.B(g26229));
  OR2 OR2_24(.VSS(VSS),.VDD(VDD),.Y(g30356),.A(g30096),.B(g18365));
  OR2 OR2_25(.VSS(VSS),.VDD(VDD),.Y(g27580),.A(g26159),.B(g24749));
  OR2 OR2_26(.VSS(VSS),.VDD(VDD),.Y(g34647),.A(g34558),.B(g18820));
  OR2 OR2_27(.VSS(VSS),.VDD(VDD),.Y(g26932),.A(g26684),.B(g18549));
  OR4 OR4_2(.VSS(VSS),.VDD(VDD),.Y(I31859),.A(g33501),.B(g33502),.C(g33503),.D(g33504));
  OR2 OR2_28(.VSS(VSS),.VDD(VDD),.Y(g33049),.A(g31966),.B(g21929));
  OR2 OR2_29(.VSS(VSS),.VDD(VDD),.Y(g30380),.A(g30161),.B(g18492));
  OR2 OR2_30(.VSS(VSS),.VDD(VDD),.Y(g34826),.A(g34742),.B(g34685));
  OR3 OR3_0(.VSS(VSS),.VDD(VDD),.Y(g16926),.A(g14061),.B(g11804),.C(g11780));
  OR3 OR3_1(.VSS(VSS),.VDD(VDD),.Y(I25736),.A(g12),.B(g22150),.C(g20277));
  OR4 OR4_3(.VSS(VSS),.VDD(VDD),.Y(I31858),.A(g33497),.B(g33498),.C(g33499),.D(g33500));
  OR2 OR2_31(.VSS(VSS),.VDD(VDD),.Y(g33048),.A(g31960),.B(g21928));
  OR2 OR2_32(.VSS(VSS),.VDD(VDD),.Y(g7684),.A(g4072),.B(g4176));
  OR2 OR2_33(.VSS(VSS),.VDD(VDD),.Y(g25710),.A(g25031),.B(g21961));
  OR2 OR2_34(.VSS(VSS),.VDD(VDD),.Y(g28610),.A(g27347),.B(g16484));
  OR2 OR2_35(.VSS(VSS),.VDD(VDD),.Y(g26897),.A(g26611),.B(g18176));
  OR2 OR2_36(.VSS(VSS),.VDD(VDD),.Y(g34090),.A(g33676),.B(g33680));
  OR2 OR2_37(.VSS(VSS),.VDD(VDD),.Y(g26961),.A(g26280),.B(g24306));
  OR2 OR2_38(.VSS(VSS),.VDD(VDD),.Y(g28705),.A(g27460),.B(g16672));
  OR2 OR2_39(.VSS(VSS),.VDD(VDD),.Y(g28042),.A(g24148),.B(g26879));
  OR2 OR2_40(.VSS(VSS),.VDD(VDD),.Y(g30672),.A(g13737),.B(g29752));
  OR2 OR2_41(.VSS(VSS),.VDD(VDD),.Y(g34233),.A(g32455),.B(g33951));
  OR2 OR2_42(.VSS(VSS),.VDD(VDD),.Y(g13211),.A(g11294),.B(g7567));
  OR2 OR2_43(.VSS(VSS),.VDD(VDD),.Y(g33004),.A(g32246),.B(g18431));
  OR2 OR2_44(.VSS(VSS),.VDD(VDD),.Y(g31221),.A(g29494),.B(g28204));
  OR3 OR3_2(.VSS(VSS),.VDD(VDD),.Y(g23198),.A(g20214),.B(g20199),.C(I22298));
  OR4 OR4_4(.VSS(VSS),.VDD(VDD),.Y(I31844),.A(g33474),.B(g33475),.C(g33476),.D(g33477));
  OR2 OR2_45(.VSS(VSS),.VDD(VDD),.Y(g27179),.A(g25816),.B(g24409));
  OR2 OR2_46(.VSS(VSS),.VDD(VDD),.Y(g28188),.A(g22535),.B(g27108));
  OR2 OR2_47(.VSS(VSS),.VDD(VDD),.Y(g33613),.A(g33248),.B(g18649));
  OR2 OR2_48(.VSS(VSS),.VDD(VDD),.Y(g34331),.A(g27121),.B(g34072));
  OR2 OR2_49(.VSS(VSS),.VDD(VDD),.Y(g30513),.A(g30200),.B(g22034));
  OR2 OR2_50(.VSS(VSS),.VDD(VDD),.Y(g30449),.A(g29845),.B(g21858));
  OR2 OR2_51(.VSS(VSS),.VDD(VDD),.Y(g33947),.A(g32438),.B(g33457));
  OR2 OR2_52(.VSS(VSS),.VDD(VDD),.Y(g34449),.A(g34279),.B(g18662));
  OR2 OR2_53(.VSS(VSS),.VDD(VDD),.Y(g25647),.A(g24725),.B(g21740));
  OR2 OR2_54(.VSS(VSS),.VDD(VDD),.Y(g24243),.A(g22992),.B(g18254));
  OR2 OR2_55(.VSS(VSS),.VDD(VDD),.Y(g33273),.A(g32122),.B(g29553));
  OR2 OR2_56(.VSS(VSS),.VDD(VDD),.Y(g28030),.A(g24018),.B(g26874));
  OR2 OR2_57(.VSS(VSS),.VDD(VDD),.Y(g33605),.A(g33352),.B(g18521));
  OR2 OR2_58(.VSS(VSS),.VDD(VDD),.Y(g25945),.A(g24427),.B(g22307));
  OR2 OR2_59(.VSS(VSS),.VDD(VDD),.Y(g28093),.A(g27981),.B(g21951));
  OR2 OR2_60(.VSS(VSS),.VDD(VDD),.Y(g30448),.A(g29809),.B(g21857));
  OR2 OR2_61(.VSS(VSS),.VDD(VDD),.Y(g34897),.A(g34861),.B(g21682));
  OR2 OR2_62(.VSS(VSS),.VDD(VDD),.Y(g34448),.A(g34365),.B(g18553));
  OR2 OR2_63(.VSS(VSS),.VDD(VDD),.Y(g30505),.A(g30168),.B(g22026));
  OR2 OR2_64(.VSS(VSS),.VDD(VDD),.Y(g29114),.A(g27646),.B(g26602));
  OR2 OR2_65(.VSS(VSS),.VDD(VDD),.Y(g30404),.A(g29758),.B(g21763));
  OR2 OR2_66(.VSS(VSS),.VDD(VDD),.Y(g28065),.A(g27299),.B(g21792));
  OR2 OR2_67(.VSS(VSS),.VDD(VDD),.Y(g27800),.A(g17321),.B(g26703));
  OR2 OR2_68(.VSS(VSS),.VDD(VDD),.Y(g24269),.A(g23131),.B(g18613));
  OR2 OR2_69(.VSS(VSS),.VDD(VDD),.Y(g34404),.A(g34182),.B(g25102));
  OR3 OR3_3(.VSS(VSS),.VDD(VDD),.Y(g33951),.A(g33469),.B(I31838),.C(I31839));
  OR2 OR2_70(.VSS(VSS),.VDD(VDD),.Y(g33972),.A(g33941),.B(g18335));
  OR2 OR2_71(.VSS(VSS),.VDD(VDD),.Y(g24341),.A(g23564),.B(g18771));
  OR2 OR2_72(.VSS(VSS),.VDD(VDD),.Y(g33033),.A(g32333),.B(g21843));
  OR2 OR2_73(.VSS(VSS),.VDD(VDD),.Y(g24268),.A(g23025),.B(g18612));
  OR2 OR2_74(.VSS(VSS),.VDD(VDD),.Y(g25651),.A(g24680),.B(g21744));
  OR2 OR2_75(.VSS(VSS),.VDD(VDD),.Y(g25672),.A(g24647),.B(g21829));
  OR2 OR2_76(.VSS(VSS),.VDD(VDD),.Y(g33234),.A(g32039),.B(g32043));
  OR2 OR2_77(.VSS(VSS),.VDD(VDD),.Y(g34026),.A(g33715),.B(g18682));
  OR2 OR2_78(.VSS(VSS),.VDD(VDD),.Y(g32427),.A(g8928),.B(g30583));
  OR2 OR2_79(.VSS(VSS),.VDD(VDD),.Y(g13296),.A(g10626),.B(g10657));
  OR2 OR2_80(.VSS(VSS),.VDD(VDD),.Y(g23087),.A(g19487),.B(g15852));
  OR2 OR2_81(.VSS(VSS),.VDD(VDD),.Y(g29849),.A(g26049),.B(g28273));
  OR2 OR2_82(.VSS(VSS),.VDD(VDD),.Y(g13969),.A(g11448),.B(g8913));
  OR2 OR2_83(.VSS(VSS),.VDD(VDD),.Y(g26343),.A(g1514),.B(g24609));
  OR2 OR2_84(.VSS(VSS),.VDD(VDD),.Y(g19522),.A(g17057),.B(g14180));
  OR2 OR2_85(.VSS(VSS),.VDD(VDD),.Y(g29848),.A(g28260),.B(g26077));
  OR2 OR2_86(.VSS(VSS),.VDD(VDD),.Y(g24335),.A(g22165),.B(g18678));
  OR2 OR2_87(.VSS(VSS),.VDD(VDD),.Y(g26971),.A(g26325),.B(g24333));
  OR2 OR2_88(.VSS(VSS),.VDD(VDD),.Y(g34723),.A(g34710),.B(g18139));
  OR2 OR2_89(.VSS(VSS),.VDD(VDD),.Y(g30433),.A(g29899),.B(g21817));
  OR2 OR2_90(.VSS(VSS),.VDD(VDD),.Y(g34149),.A(g33760),.B(g19674));
  OR2 OR2_91(.VSS(VSS),.VDD(VDD),.Y(g30387),.A(g30151),.B(g18524));
  OR2 OR2_92(.VSS(VSS),.VDD(VDD),.Y(g24965),.A(g22667),.B(g23825));
  OR2 OR2_93(.VSS(VSS),.VDD(VDD),.Y(g32226),.A(g31145),.B(g29645));
  OR2 OR2_94(.VSS(VSS),.VDD(VDD),.Y(g29263),.A(g28239),.B(g18617));
  OR2 OR2_95(.VSS(VSS),.VDD(VDD),.Y(g34620),.A(g34529),.B(g18582));
  OR2 OR2_96(.VSS(VSS),.VDD(VDD),.Y(g34148),.A(g33758),.B(g19656));
  OR2 OR2_97(.VSS(VSS),.VDD(VDD),.Y(g25717),.A(g25106),.B(g21968));
  OR2 OR2_98(.VSS(VSS),.VDD(VDD),.Y(g27543),.A(g26085),.B(g24670));
  OR2 OR2_99(.VSS(VSS),.VDD(VDD),.Y(g30104),.A(g28478),.B(g11427));
  OR2 OR2_100(.VSS(VSS),.VDD(VDD),.Y(g33012),.A(g32274),.B(g18483));
  OR2 OR2_101(.VSS(VSS),.VDD(VDD),.Y(g19949),.A(g17671),.B(g14681));
  OR2 OR2_102(.VSS(VSS),.VDD(VDD),.Y(g30343),.A(g29344),.B(g18278));
  OR2 OR2_103(.VSS(VSS),.VDD(VDD),.Y(g34646),.A(g34557),.B(g18803));
  OR2 OR2_104(.VSS(VSS),.VDD(VDD),.Y(g24557),.A(g22308),.B(g19207));
  OR2 OR2_105(.VSS(VSS),.VDD(VDD),.Y(g24210),.A(g22900),.B(g18125));
  OR2 OR2_106(.VSS(VSS),.VDD(VDD),.Y(g27569),.A(g26124),.B(g24721));
  OR2 OR2_107(.VSS(VSS),.VDD(VDD),.Y(g34971),.A(g34869),.B(g34962));
  OR2 OR2_108(.VSS(VSS),.VDD(VDD),.Y(g33541),.A(g33101),.B(g18223));
  OR2 OR2_109(.VSS(VSS),.VDD(VDD),.Y(g31473),.A(g26180),.B(g29666));
  OR2 OR2_110(.VSS(VSS),.VDD(VDD),.Y(g28075),.A(g27083),.B(g21877));
  OR2 OR2_111(.VSS(VSS),.VDD(VDD),.Y(g30369),.A(g30066),.B(g18439));
  OR2 OR2_112(.VSS(VSS),.VDD(VDD),.Y(g24443),.A(g23917),.B(g21378));
  OR2 OR2_113(.VSS(VSS),.VDD(VDD),.Y(g19904),.A(g17636),.B(g14654));
  OR2 OR2_114(.VSS(VSS),.VDD(VDD),.Y(g23171),.A(g19536),.B(g15903));
  OR2 OR2_115(.VSS(VSS),.VDD(VDD),.Y(g24279),.A(g23218),.B(g15105));
  OR2 OR2_116(.VSS(VSS),.VDD(VDD),.Y(g26896),.A(g26341),.B(g18171));
  OR2 OR2_117(.VSS(VSS),.VDD(VDD),.Y(g34369),.A(g26279),.B(g34136));
  OR2 OR2_118(.VSS(VSS),.VDD(VDD),.Y(g28595),.A(g27335),.B(g26290));
  OR2 OR2_119(.VSS(VSS),.VDD(VDD),.Y(g14030),.A(g11037),.B(g11046));
  OR2 OR2_120(.VSS(VSS),.VDD(VDD),.Y(g30368),.A(g30098),.B(g18435));
  OR2 OR2_121(.VSS(VSS),.VDD(VDD),.Y(g24278),.A(g23201),.B(g18648));
  OR2 OR2_122(.VSS(VSS),.VDD(VDD),.Y(g25723),.A(g25033),.B(g22006));
  OR2 OR2_123(.VSS(VSS),.VDD(VDD),.Y(g28623),.A(g27361),.B(g16520));
  OR2 OR2_124(.VSS(VSS),.VDD(VDD),.Y(g34368),.A(g26274),.B(g34135));
  OR2 OR2_125(.VSS(VSS),.VDD(VDD),.Y(g33788),.A(g33122),.B(g32041));
  OR2 OR2_126(.VSS(VSS),.VDD(VDD),.Y(g31325),.A(g29625),.B(g29639));
  OR2 OR2_127(.VSS(VSS),.VDD(VDD),.Y(g32385),.A(g31480),.B(g29938));
  OR2 OR2_128(.VSS(VSS),.VDD(VDD),.Y(g31920),.A(g31493),.B(g22045));
  OR2 OR2_129(.VSS(VSS),.VDD(VDD),.Y(g32980),.A(g32254),.B(g18198));
  OR2 OR2_130(.VSS(VSS),.VDD(VDD),.Y(g30412),.A(g29885),.B(g21771));
  OR2 OR2_131(.VSS(VSS),.VDD(VDD),.Y(g33535),.A(g33233),.B(g21711));
  OR2 OR2_132(.VSS(VSS),.VDD(VDD),.Y(g24468),.A(g10925),.B(g22400));
  OR2 OR2_133(.VSS(VSS),.VDD(VDD),.Y(g32354),.A(g29854),.B(g31285));
  OR2 OR2_134(.VSS(VSS),.VDD(VDD),.Y(g34850),.A(g34841),.B(g18185));
  OR2 OR2_135(.VSS(VSS),.VDD(VDD),.Y(g34412),.A(g34187),.B(g25143));
  OR2 OR2_136(.VSS(VSS),.VDD(VDD),.Y(g28419),.A(g27221),.B(g15884));
  OR2 OR2_137(.VSS(VSS),.VDD(VDD),.Y(g27974),.A(g26544),.B(g25063));
  OR2 OR2_138(.VSS(VSS),.VDD(VDD),.Y(g33946),.A(g32434),.B(g33456));
  OR2 OR2_139(.VSS(VSS),.VDD(VDD),.Y(g25646),.A(g24706),.B(g21739));
  OR2 OR2_140(.VSS(VSS),.VDD(VDD),.Y(g28418),.A(g27220),.B(g15882));
  OR2 OR2_141(.VSS(VSS),.VDD(VDD),.Y(g20187),.A(g16202),.B(g13491));
  OR2 OR2_142(.VSS(VSS),.VDD(VDD),.Y(g26959),.A(g26381),.B(g24299));
  OR2 OR2_143(.VSS(VSS),.VDD(VDD),.Y(g26925),.A(g25939),.B(g18301));
  OR2 OR2_144(.VSS(VSS),.VDD(VDD),.Y(g34011),.A(g33884),.B(g18479));
  OR2 OR2_145(.VSS(VSS),.VDD(VDD),.Y(g26958),.A(g26395),.B(g24297));
  OR2 OR2_146(.VSS(VSS),.VDD(VDD),.Y(g29273),.A(g28269),.B(g18639));
  OR2 OR2_147(.VSS(VSS),.VDD(VDD),.Y(g31291),.A(g29581),.B(g29593));
  OR4 OR4_5(.VSS(VSS),.VDD(VDD),.Y(g17570),.A(g14419),.B(g14397),.C(g11999),.D(I18495));
  OR2 OR2_148(.VSS(VSS),.VDD(VDD),.Y(g33291),.A(g32154),.B(g13477));
  OR2 OR2_149(.VSS(VSS),.VDD(VDD),.Y(g26386),.A(g24719),.B(g23023));
  OR3 OR3_4(.VSS(VSS),.VDD(VDD),.Y(g32426),.A(g26105),.B(g26131),.C(g30613));
  OR2 OR2_150(.VSS(VSS),.VDD(VDD),.Y(g28194),.A(g22540),.B(g27122));
  OR2 OR2_151(.VSS(VSS),.VDD(VDD),.Y(g28589),.A(g27331),.B(g26285));
  OR2 OR2_152(.VSS(VSS),.VDD(VDD),.Y(g26944),.A(g26130),.B(g18658));
  OR2 OR2_153(.VSS(VSS),.VDD(VDD),.Y(g20169),.A(g16184),.B(g13460));
  OR2 OR2_154(.VSS(VSS),.VDD(VDD),.Y(g27579),.A(g26157),.B(g24748));
  OR2 OR2_155(.VSS(VSS),.VDD(VDD),.Y(g29234),.A(g28415),.B(g18239));
  OR2 OR2_156(.VSS(VSS),.VDD(VDD),.Y(g30379),.A(g30089),.B(g18491));
  OR2 OR2_157(.VSS(VSS),.VDD(VDD),.Y(g34627),.A(g34534),.B(g18644));
  OR2 OR2_158(.VSS(VSS),.VDD(VDD),.Y(g27578),.A(g26155),.B(g24747));
  OR4 OR4_6(.VSS(VSS),.VDD(VDD),.Y(g17594),.A(g14450),.B(g14420),.C(g12025),.D(I18543));
  OR2 OR2_159(.VSS(VSS),.VDD(VDD),.Y(g28401),.A(g27212),.B(g15871));
  OR2 OR2_160(.VSS(VSS),.VDD(VDD),.Y(g31760),.A(g30007),.B(g30027));
  OR2 OR2_161(.VSS(VSS),.VDD(VDD),.Y(g34379),.A(g26312),.B(g34143));
  OR2 OR2_162(.VSS(VSS),.VDD(VDD),.Y(g33029),.A(g32332),.B(g21798));
  OR2 OR2_163(.VSS(VSS),.VDD(VDD),.Y(g32211),.A(g31124),.B(g29603));
  OR2 OR2_164(.VSS(VSS),.VDD(VDD),.Y(g30378),.A(g30125),.B(g18487));
  OR2 OR2_165(.VSS(VSS),.VDD(VDD),.Y(g21901),.A(g21251),.B(g15115));
  OR2 OR2_166(.VSS(VSS),.VDD(VDD),.Y(g20217),.A(g16221),.B(g13523));
  OR2 OR2_167(.VSS(VSS),.VDD(VDD),.Y(g33028),.A(g32325),.B(g21797));
  OR2 OR2_168(.VSS(VSS),.VDD(VDD),.Y(g30386),.A(g30139),.B(g18523));
  OR2 OR2_169(.VSS(VSS),.VDD(VDD),.Y(g24363),.A(g7831),.B(g22138));
  OR2 OR2_170(.VSS(VSS),.VDD(VDD),.Y(g26793),.A(g24478),.B(g7520));
  OR2 OR2_171(.VSS(VSS),.VDD(VDD),.Y(g28118),.A(g27821),.B(g26815));
  OR3 OR3_5(.VSS(VSS),.VDD(VDD),.Y(g13526),.A(g209),.B(g10685),.C(g301));
  OR2 OR2_172(.VSS(VSS),.VDD(VDD),.Y(g24478),.A(g11003),.B(g22450));
  OR2 OR2_173(.VSS(VSS),.VDD(VDD),.Y(g34603),.A(g34561),.B(g15075));
  OR2 OR2_174(.VSS(VSS),.VDD(VDD),.Y(g25716),.A(g25088),.B(g21967));
  OR2 OR2_175(.VSS(VSS),.VDD(VDD),.Y(g28749),.A(g27523),.B(g16764));
  OR2 OR2_176(.VSS(VSS),.VDD(VDD),.Y(g26690),.A(g10776),.B(g24433));
  OR2 OR2_177(.VSS(VSS),.VDD(VDD),.Y(g25582),.A(g21662),.B(g24152));
  OR2 OR2_178(.VSS(VSS),.VDD(VDD),.Y(g28748),.A(g27522),.B(g16763));
  OR2 OR2_179(.VSS(VSS),.VDD(VDD),.Y(g28704),.A(g27459),.B(g16671));
  OR2 OR2_180(.VSS(VSS),.VDD(VDD),.Y(g24580),.A(g22340),.B(g13096));
  OR2 OR2_181(.VSS(VSS),.VDD(VDD),.Y(g31927),.A(g31500),.B(g22091));
  OR2 OR2_182(.VSS(VSS),.VDD(VDD),.Y(g30429),.A(g29844),.B(g21813));
  OR2 OR2_183(.VSS(VSS),.VDD(VDD),.Y(g28305),.A(g27103),.B(g15793));
  OR2 OR2_184(.VSS(VSS),.VDD(VDD),.Y(g28053),.A(g27393),.B(g18168));
  OR2 OR2_185(.VSS(VSS),.VDD(VDD),.Y(g32987),.A(g32311),.B(g18323));
  OR2 OR2_186(.VSS(VSS),.VDD(VDD),.Y(g32250),.A(g30598),.B(g29351));
  OR2 OR2_187(.VSS(VSS),.VDD(VDD),.Y(g34802),.A(g34757),.B(g18589));
  OR2 OR2_188(.VSS(VSS),.VDD(VDD),.Y(g25627),.A(g24503),.B(g18247));
  OR2 OR2_189(.VSS(VSS),.VDD(VDD),.Y(g30428),.A(g29807),.B(g21812));
  OR2 OR2_190(.VSS(VSS),.VDD(VDD),.Y(g34730),.A(g34658),.B(g18271));
  OR2 OR2_191(.VSS(VSS),.VDD(VDD),.Y(g34793),.A(g34744),.B(g18570));
  OR4 OR4_7(.VSS(VSS),.VDD(VDD),.Y(I26643),.A(g27073),.B(g27058),.C(g27045),.D(g27040));
  OR2 OR2_192(.VSS(VSS),.VDD(VDD),.Y(g13077),.A(g11330),.B(g943));
  OR3 OR3_6(.VSS(VSS),.VDD(VDD),.Y(I18492),.A(g14538),.B(g14513),.C(g14446));
  OR2 OR2_193(.VSS(VSS),.VDD(VDD),.Y(g28101),.A(g27691),.B(g22062));
  OR2 OR2_194(.VSS(VSS),.VDD(VDD),.Y(g33240),.A(g32052),.B(g32068));
  OR2 OR2_195(.VSS(VSS),.VDD(VDD),.Y(g13597),.A(g9247),.B(g11149));
  OR2 OR2_196(.VSS(VSS),.VDD(VDD),.Y(g28560),.A(g27311),.B(g26249));
  OR2 OR2_197(.VSS(VSS),.VDD(VDD),.Y(g31903),.A(g31374),.B(g21911));
  OR2 OR2_198(.VSS(VSS),.VDD(VDD),.Y(g30549),.A(g30215),.B(g22120));
  OR2 OR2_199(.VSS(VSS),.VDD(VDD),.Y(g25603),.A(g24698),.B(g18114));
  OR2 OR2_200(.VSS(VSS),.VDD(VDD),.Y(g25742),.A(g25093),.B(g22057));
  OR2 OR2_201(.VSS(VSS),.VDD(VDD),.Y(g31755),.A(g29991),.B(g30008));
  OR2 OR2_202(.VSS(VSS),.VDD(VDD),.Y(g33604),.A(g33345),.B(g18520));
  OR2 OR2_203(.VSS(VSS),.VDD(VDD),.Y(g30548),.A(g30204),.B(g22119));
  OR2 OR2_204(.VSS(VSS),.VDD(VDD),.Y(g10589),.A(g7223),.B(g7201));
  OR2 OR2_205(.VSS(VSS),.VDD(VDD),.Y(g29325),.A(g28813),.B(g27820));
  OR2 OR2_206(.VSS(VSS),.VDD(VDD),.Y(g13300),.A(g10656),.B(g10676));
  OR2 OR2_207(.VSS(VSS),.VDD(VDD),.Y(g31770),.A(g30034),.B(g30047));
  OR2 OR2_208(.VSS(VSS),.VDD(VDD),.Y(g30504),.A(g30253),.B(g22025));
  OR2 OR2_209(.VSS(VSS),.VDD(VDD),.Y(g28064),.A(g27298),.B(g21781));
  OR2 OR2_210(.VSS(VSS),.VDD(VDD),.Y(g33563),.A(g33361),.B(g18383));
  OR2 OR2_211(.VSS(VSS),.VDD(VDD),.Y(g33981),.A(g33856),.B(g18371));
  OR2 OR2_212(.VSS(VSS),.VDD(VDD),.Y(g25681),.A(g24710),.B(g18636));
  OR2 OR2_213(.VSS(VSS),.VDD(VDD),.Y(g28733),.A(g27507),.B(g16735));
  OR2 OR2_214(.VSS(VSS),.VDD(VDD),.Y(g26299),.A(g24551),.B(g22665));
  OR3 OR3_7(.VSS(VSS),.VDD(VDD),.Y(g30317),.A(g29208),.B(I28566),.C(I28567));
  OR2 OR2_215(.VSS(VSS),.VDD(VDD),.Y(g25730),.A(g25107),.B(g22013));
  OR2 OR2_216(.VSS(VSS),.VDD(VDD),.Y(g22304),.A(g21347),.B(g17693));
  OR2 OR2_217(.VSS(VSS),.VDD(VDD),.Y(g14119),.A(g10776),.B(g8703));
  OR2 OR2_218(.VSS(VSS),.VDD(VDD),.Y(g31767),.A(g30031),.B(g30043));
  OR2 OR2_219(.VSS(VSS),.VDD(VDD),.Y(g33794),.A(g33126),.B(g32053));
  OR2 OR2_220(.VSS(VSS),.VDD(VDD),.Y(g34002),.A(g33857),.B(g18451));
  OR2 OR2_221(.VSS(VSS),.VDD(VDD),.Y(g33262),.A(g32112),.B(g29528));
  OR2 OR2_222(.VSS(VSS),.VDD(VDD),.Y(g31899),.A(g31470),.B(g21907));
  OR2 OR2_223(.VSS(VSS),.VDD(VDD),.Y(g34057),.A(g33911),.B(g33915));
  OR2 OR2_224(.VSS(VSS),.VDD(VDD),.Y(g28665),.A(g27409),.B(g16614));
  OR2 OR2_225(.VSS(VSS),.VDD(VDD),.Y(g30128),.A(g28495),.B(g11497));
  OR2 OR2_226(.VSS(VSS),.VDD(VDD),.Y(g33990),.A(g33882),.B(g18399));
  OR2 OR2_227(.VSS(VSS),.VDD(VDD),.Y(g24334),.A(g23991),.B(g18676));
  OR2 OR2_228(.VSS(VSS),.VDD(VDD),.Y(g25690),.A(g24864),.B(g21889));
  OR2 OR2_229(.VSS(VSS),.VDD(VDD),.Y(g26737),.A(g24460),.B(g10720));
  OR2 OR2_230(.VSS(VSS),.VDD(VDD),.Y(g29291),.A(g28660),.B(g18767));
  OR2 OR2_231(.VSS(VSS),.VDD(VDD),.Y(g31898),.A(g31707),.B(g21906));
  OR2 OR2_232(.VSS(VSS),.VDD(VDD),.Y(g34626),.A(g34533),.B(g18627));
  OR2 OR2_233(.VSS(VSS),.VDD(VDD),.Y(g30533),.A(g30203),.B(g22079));
  OR2 OR2_234(.VSS(VSS),.VDD(VDD),.Y(g22653),.A(g18993),.B(g15654));
  OR2 OR2_235(.VSS(VSS),.VDD(VDD),.Y(g30298),.A(g28245),.B(g27251));
  OR3 OR3_8(.VSS(VSS),.VDD(VDD),.Y(g23687),.A(g21384),.B(g21363),.C(I22830));
  OR2 OR2_236(.VSS(VSS),.VDD(VDD),.Y(g26880),.A(g26610),.B(g24186));
  OR2 OR2_237(.VSS(VSS),.VDD(VDD),.Y(g24216),.A(g23416),.B(g18197));
  OR2 OR2_238(.VSS(VSS),.VDD(VDD),.Y(g23374),.A(g19767),.B(g13514));
  OR2 OR2_239(.VSS(VSS),.VDD(VDD),.Y(g32202),.A(g31069),.B(g13410));
  OR2 OR2_240(.VSS(VSS),.VDD(VDD),.Y(g22636),.A(g18943),.B(g15611));
  OR2 OR2_241(.VSS(VSS),.VDD(VDD),.Y(g26512),.A(g24786),.B(g23130));
  OR2 OR2_242(.VSS(VSS),.VDD(VDD),.Y(g32257),.A(g31184),.B(g29708));
  OR2 OR2_243(.VSS(VSS),.VDD(VDD),.Y(g13660),.A(g8183),.B(g12527));
  OR2 OR2_244(.VSS(VSS),.VDD(VDD),.Y(g32979),.A(g32181),.B(g18177));
  OR2 OR2_245(.VSS(VSS),.VDD(VDD),.Y(g29506),.A(g28148),.B(g25880));
  OR2 OR2_246(.VSS(VSS),.VDD(VDD),.Y(g34232),.A(g33451),.B(g33944));
  OR2 OR2_247(.VSS(VSS),.VDD(VDD),.Y(g32978),.A(g32197),.B(g18145));
  OR2 OR2_248(.VSS(VSS),.VDD(VDD),.Y(g28074),.A(g27119),.B(g21876));
  OR2 OR2_249(.VSS(VSS),.VDD(VDD),.Y(g33573),.A(g33343),.B(g18415));
  OR2 OR2_250(.VSS(VSS),.VDD(VDD),.Y(g31247),.A(g29513),.B(g13324));
  OR2 OR2_251(.VSS(VSS),.VDD(VDD),.Y(g28594),.A(g27334),.B(g26289));
  OR2 OR2_252(.VSS(VSS),.VDD(VDD),.Y(g31926),.A(g31765),.B(g22090));
  OR2 OR2_253(.VSS(VSS),.VDD(VDD),.Y(g32986),.A(g31996),.B(g18280));
  OR2 OR2_254(.VSS(VSS),.VDD(VDD),.Y(g27253),.A(g24661),.B(g26052));
  OR2 OR2_255(.VSS(VSS),.VDD(VDD),.Y(g33389),.A(g32272),.B(g29964));
  OR2 OR2_256(.VSS(VSS),.VDD(VDD),.Y(g33045),.A(g32206),.B(g24328));
  OR2 OR2_257(.VSS(VSS),.VDD(VDD),.Y(g22664),.A(g19139),.B(g15694));
  OR2 OR2_258(.VSS(VSS),.VDD(VDD),.Y(g34856),.A(g34811),.B(g34743));
  OR2 OR2_259(.VSS(VSS),.VDD(VDD),.Y(g25626),.A(g24499),.B(g18235));
  OR2 OR2_260(.VSS(VSS),.VDD(VDD),.Y(g33612),.A(g33247),.B(g18633));
  OR2 OR2_261(.VSS(VSS),.VDD(VDD),.Y(g34261),.A(g34074),.B(g18688));
  OR2 OR2_262(.VSS(VSS),.VDD(VDD),.Y(g34880),.A(g34867),.B(g18153));
  OR2 OR2_263(.VSS(VSS),.VDD(VDD),.Y(g8921),.A(I12902),.B(I12903));
  OR2 OR2_264(.VSS(VSS),.VDD(VDD),.Y(g30512),.A(g30191),.B(g22033));
  OR2 OR2_265(.VSS(VSS),.VDD(VDD),.Y(g33534),.A(g33186),.B(g21700));
  OR2 OR2_266(.VSS(VSS),.VDD(VDD),.Y(g27236),.A(g24620),.B(g25974));
  OR2 OR2_267(.VSS(VSS),.VDD(VDD),.Y(g32094),.A(g30612),.B(g29363));
  OR2 OR2_268(.VSS(VSS),.VDD(VDD),.Y(g31251),.A(g25973),.B(g29527));
  OR2 OR2_269(.VSS(VSS),.VDD(VDD),.Y(g22585),.A(g20915),.B(g21061));
  OR2 OR2_270(.VSS(VSS),.VDD(VDD),.Y(g33251),.A(g32096),.B(g29509));
  OR2 OR2_271(.VSS(VSS),.VDD(VDD),.Y(g24242),.A(g22834),.B(g18253));
  OR2 OR2_272(.VSS(VSS),.VDD(VDD),.Y(g33272),.A(g32121),.B(g29551));
  OR2 OR2_273(.VSS(VSS),.VDD(VDD),.Y(g28092),.A(g27666),.B(g21924));
  OR4 OR4_8(.VSS(VSS),.VDD(VDD),.Y(I30124),.A(g31070),.B(g31154),.C(g30614),.D(g30673));
  OR2 OR2_274(.VSS(VSS),.VDD(VDD),.Y(g28518),.A(g27281),.B(g26158));
  OR2 OR2_275(.VSS(VSS),.VDD(VDD),.Y(g21893),.A(g20094),.B(g18655));
  OR2 OR2_276(.VSS(VSS),.VDD(VDD),.Y(g29240),.A(g28655),.B(g18328));
  OR2 OR2_277(.VSS(VSS),.VDD(VDD),.Y(g26080),.A(g19393),.B(g24502));
  OR3 OR3_9(.VSS(VSS),.VDD(VDD),.Y(I12583),.A(g1157),.B(g1239),.C(g990));
  OR2 OR2_278(.VSS(VSS),.VDD(VDD),.Y(g25737),.A(g25045),.B(g22052));
  OR2 OR2_279(.VSS(VSS),.VDD(VDD),.Y(g26924),.A(g26153),.B(g18291));
  OR2 OR2_280(.VSS(VSS),.VDD(VDD),.Y(g30445),.A(g29772),.B(g21854));
  OR2 OR2_281(.VSS(VSS),.VDD(VDD),.Y(g33032),.A(g32326),.B(g21842));
  OR2 OR2_282(.VSS(VSS),.VDD(VDD),.Y(g34445),.A(g34382),.B(g18548));
  OR2 OR2_283(.VSS(VSS),.VDD(VDD),.Y(g30499),.A(g30261),.B(g21995));
  OR2 OR2_284(.VSS(VSS),.VDD(VDD),.Y(g33997),.A(g33871),.B(g18427));
  OR2 OR2_285(.VSS(VSS),.VDD(VDD),.Y(g25697),.A(g25086),.B(g21916));
  OR4 OR4_9(.VSS(VSS),.VDD(VDD),.Y(g25856),.A(g25518),.B(g25510),.C(g25488),.D(g25462));
  OR2 OR2_286(.VSS(VSS),.VDD(VDD),.Y(g30498),.A(g30251),.B(g21994));
  OR2 OR2_287(.VSS(VSS),.VDD(VDD),.Y(g25261),.A(g23348),.B(g20193));
  OR2 OR2_288(.VSS(VSS),.VDD(VDD),.Y(g33061),.A(g32334),.B(g22050));
  OR2 OR2_289(.VSS(VSS),.VDD(VDD),.Y(g24265),.A(g22316),.B(g18560));
  OR2 OR2_290(.VSS(VSS),.VDD(VDD),.Y(g26342),.A(g8407),.B(g24591));
  OR2 OR2_291(.VSS(VSS),.VDD(VDD),.Y(g31766),.A(g30029),.B(g30042));
  OR2 OR2_292(.VSS(VSS),.VDD(VDD),.Y(g31871),.A(g30596),.B(g18279));
  OR2 OR2_293(.VSS(VSS),.VDD(VDD),.Y(g30611),.A(g13671),.B(g29743));
  OR2 OR2_294(.VSS(VSS),.VDD(VDD),.Y(g24841),.A(g21420),.B(g23998));
  OR2 OR2_295(.VSS(VSS),.VDD(VDD),.Y(g34611),.A(g34508),.B(g18565));
  OR2 OR2_296(.VSS(VSS),.VDD(VDD),.Y(g23255),.A(g19655),.B(g16122));
  OR2 OR2_297(.VSS(VSS),.VDD(VDD),.Y(g34722),.A(g34707),.B(g18137));
  OR2 OR2_298(.VSS(VSS),.VDD(VDD),.Y(g26887),.A(g26542),.B(g24193));
  OR2 OR2_299(.VSS(VSS),.VDD(VDD),.Y(g28729),.A(g27502),.B(g16732));
  OR2 OR2_300(.VSS(VSS),.VDD(VDD),.Y(g28577),.A(g27326),.B(g26272));
  OR2 OR2_301(.VSS(VSS),.VDD(VDD),.Y(g24510),.A(g22488),.B(g7567));
  OR2 OR2_302(.VSS(VSS),.VDD(VDD),.Y(g30432),.A(g29888),.B(g21816));
  OR2 OR2_303(.VSS(VSS),.VDD(VDD),.Y(g28728),.A(g27501),.B(g16730));
  OR2 OR2_304(.VSS(VSS),.VDD(VDD),.Y(g29262),.A(g28327),.B(g18608));
  OR2 OR2_305(.VSS(VSS),.VDD(VDD),.Y(g27542),.A(g16190),.B(g26094));
  OR2 OR2_306(.VSS(VSS),.VDD(VDD),.Y(g27453),.A(g25976),.B(g24606));
  OR2 OR2_307(.VSS(VSS),.VDD(VDD),.Y(g23383),.A(g19756),.B(g16222));
  OR2 OR2_308(.VSS(VSS),.VDD(VDD),.Y(g24578),.A(g2882),.B(g23825));
  OR2 OR2_309(.VSS(VSS),.VDD(VDD),.Y(g30461),.A(g30219),.B(g21932));
  OR2 OR2_310(.VSS(VSS),.VDD(VDD),.Y(g30342),.A(g29330),.B(g18261));
  OR2 OR2_311(.VSS(VSS),.VDD(VDD),.Y(g34461),.A(g34291),.B(g18681));
  OR2 OR2_312(.VSS(VSS),.VDD(VDD),.Y(g26365),.A(g25504),.B(g25141));
  OR3 OR3_10(.VSS(VSS),.VDD(VDD),.Y(I18452),.A(g14514),.B(g14448),.C(g14418));
  OR2 OR2_313(.VSS(VSS),.VDD(VDD),.Y(g26960),.A(g26258),.B(g24304));
  OR2 OR2_314(.VSS(VSS),.VDD(VDD),.Y(g34031),.A(g33735),.B(g18705));
  OR2 OR2_315(.VSS(VSS),.VDD(VDD),.Y(g31472),.A(g29642),.B(g28352));
  OR2 OR2_316(.VSS(VSS),.VDD(VDD),.Y(g28083),.A(g27249),.B(g18689));
  OR2 OR2_317(.VSS(VSS),.VDD(VDD),.Y(g28348),.A(g27139),.B(g15823));
  OR2 OR2_318(.VSS(VSS),.VDD(VDD),.Y(g34199),.A(g33820),.B(g33828));
  OR2 OR2_319(.VSS(VSS),.VDD(VDD),.Y(g32280),.A(g24790),.B(g31225));
  OR2 OR2_320(.VSS(VSS),.VDD(VDD),.Y(g9984),.A(g4300),.B(g4242));
  OR2 OR2_321(.VSS(VSS),.VDD(VDD),.Y(g34887),.A(g34865),.B(g21670));
  OR2 OR2_322(.VSS(VSS),.VDD(VDD),.Y(g31911),.A(g31784),.B(g21969));
  OR2 OR2_323(.VSS(VSS),.VDD(VDD),.Y(g30529),.A(g30212),.B(g22075));
  OR2 OR2_324(.VSS(VSS),.VDD(VDD),.Y(g33628),.A(g33071),.B(g32450));
  OR2 OR2_325(.VSS(VSS),.VDD(VDD),.Y(g27274),.A(g15779),.B(g25915));
  OR2 OR2_326(.VSS(VSS),.VDD(VDD),.Y(g31246),.A(g25965),.B(g29518));
  OR2 OR2_327(.VSS(VSS),.VDD(VDD),.Y(g25611),.A(g24931),.B(g18128));
  OR2 OR2_328(.VSS(VSS),.VDD(VDD),.Y(g19356),.A(g17784),.B(g14874));
  OR2 OR2_329(.VSS(VSS),.VDD(VDD),.Y(g25722),.A(g25530),.B(g18768));
  OR2 OR2_330(.VSS(VSS),.VDD(VDD),.Y(g28622),.A(g27360),.B(g16519));
  OR2 OR2_331(.VSS(VSS),.VDD(VDD),.Y(g28566),.A(g27316),.B(g26254));
  OR2 OR2_332(.VSS(VSS),.VDD(VDD),.Y(g30528),.A(g30202),.B(g22074));
  OR2 OR2_333(.VSS(VSS),.VDD(VDD),.Y(g9483),.A(g1008),.B(g969));
  OR2 OR2_334(.VSS(VSS),.VDD(VDD),.Y(g30393),.A(g29986),.B(g21748));
  OR2 OR2_335(.VSS(VSS),.VDD(VDD),.Y(g27122),.A(g22537),.B(g25917));
  OR2 OR2_336(.VSS(VSS),.VDD(VDD),.Y(g34843),.A(g33924),.B(g34782));
  OR2 OR2_337(.VSS(VSS),.VDD(VDD),.Y(g34330),.A(g34069),.B(g33717));
  OR2 OR2_338(.VSS(VSS),.VDD(VDD),.Y(g30365),.A(g30158),.B(g18412));
  OR2 OR2_339(.VSS(VSS),.VDD(VDD),.Y(g24275),.A(g23474),.B(g18645));
  OR2 OR2_340(.VSS(VSS),.VDD(VDD),.Y(g29247),.A(g28694),.B(g18410));
  OR2 OR2_341(.VSS(VSS),.VDD(VDD),.Y(g31591),.A(g29358),.B(g29353));
  OR2 OR2_342(.VSS(VSS),.VDD(VDD),.Y(g31785),.A(g30071),.B(g30082));
  OR2 OR2_343(.VSS(VSS),.VDD(VDD),.Y(g33591),.A(g33082),.B(g18474));
  OR2 OR2_344(.VSS(VSS),.VDD(VDD),.Y(g24430),.A(g23151),.B(g8234));
  OR2 OR2_345(.VSS(VSS),.VDD(VDD),.Y(g24746),.A(g22588),.B(g19461));
  OR2 OR2_346(.VSS(VSS),.VDD(VDD),.Y(g32231),.A(g30590),.B(g29346));
  OR2 OR2_347(.VSS(VSS),.VDD(VDD),.Y(g25753),.A(g25165),.B(g22100));
  OR2 OR2_348(.VSS(VSS),.VDD(VDD),.Y(g31754),.A(g29989),.B(g30006));
  OR2 OR2_349(.VSS(VSS),.VDD(VDD),.Y(g28138),.A(g27964),.B(g27968));
  OR2 OR2_350(.VSS(VSS),.VDD(VDD),.Y(g24237),.A(g22515),.B(g18242));
  OR2 OR2_351(.VSS(VSS),.VDD(VDD),.Y(g33950),.A(g32450),.B(g33460));
  OR2 OR2_352(.VSS(VSS),.VDD(VDD),.Y(g29777),.A(g28227),.B(g28234));
  OR2 OR2_353(.VSS(VSS),.VDD(VDD),.Y(g24340),.A(g24016),.B(g18770));
  OR2 OR2_354(.VSS(VSS),.VDD(VDD),.Y(g25650),.A(g24663),.B(g21743));
  OR2 OR2_355(.VSS(VSS),.VDD(VDD),.Y(g25736),.A(g25536),.B(g18785));
  OR2 OR2_356(.VSS(VSS),.VDD(VDD),.Y(g29251),.A(g28679),.B(g18464));
  OR2 OR2_357(.VSS(VSS),.VDD(VDD),.Y(g29272),.A(g28346),.B(g18638));
  OR2 OR2_358(.VSS(VSS),.VDD(VDD),.Y(g28636),.A(g27376),.B(g16538));
  OR2 OR2_359(.VSS(VSS),.VDD(VDD),.Y(g19449),.A(g15567),.B(g12939));
  OR2 OR2_360(.VSS(VSS),.VDD(VDD),.Y(g28852),.A(g27559),.B(g16871));
  OR2 OR2_361(.VSS(VSS),.VDD(VDD),.Y(g34259),.A(g34066),.B(g18679));
  OR2 OR2_362(.VSS(VSS),.VDD(VDD),.Y(g30471),.A(g30175),.B(g21942));
  OR2 OR2_363(.VSS(VSS),.VDD(VDD),.Y(g33996),.A(g33862),.B(g18426));
  OR2 OR2_364(.VSS(VSS),.VDD(VDD),.Y(g34708),.A(g33381),.B(g34572));
  OR4 OR4_10(.VSS(VSS),.VDD(VDD),.Y(g26657),.A(g24908),.B(g24900),.C(g24887),.D(g24861));
  OR2 OR2_365(.VSS(VSS),.VDD(VDD),.Y(g25696),.A(g25012),.B(g21915));
  OR2 OR2_366(.VSS(VSS),.VDD(VDD),.Y(g26955),.A(g26391),.B(g24293));
  OR2 OR2_367(.VSS(VSS),.VDD(VDD),.Y(g34258),.A(g34211),.B(g18675));
  OR2 OR2_368(.VSS(VSS),.VDD(VDD),.Y(g24517),.A(g22158),.B(g18906));
  OR2 OR2_369(.VSS(VSS),.VDD(VDD),.Y(g26879),.A(g25580),.B(g25581));
  OR2 OR2_370(.VSS(VSS),.VDD(VDD),.Y(g26970),.A(g26308),.B(g24332));
  OR2 OR2_371(.VSS(VSS),.VDD(VDD),.Y(g25764),.A(g25551),.B(g18819));
  OR2 OR2_372(.VSS(VSS),.VDD(VDD),.Y(g28664),.A(g27408),.B(g16613));
  OR2 OR2_373(.VSS(VSS),.VDD(VDD),.Y(g26878),.A(g25578),.B(g25579));
  OR2 OR2_374(.VSS(VSS),.VDD(VDD),.Y(g16867),.A(g13493),.B(g11045));
  OR2 OR2_375(.VSS(VSS),.VDD(VDD),.Y(g25960),.A(g24566),.B(g24678));
  OR2 OR2_376(.VSS(VSS),.VDD(VDD),.Y(g34043),.A(g33903),.B(g33905));
  OR2 OR2_377(.VSS(VSS),.VDD(VDD),.Y(g26886),.A(g26651),.B(g24192));
  OR2 OR2_378(.VSS(VSS),.VDD(VDD),.Y(g25868),.A(g25450),.B(g23885));
  OR2 OR2_379(.VSS(VSS),.VDD(VDD),.Y(g28576),.A(g27325),.B(g26271));
  OR2 OR2_380(.VSS(VSS),.VDD(VDD),.Y(g31319),.A(g29612),.B(g28324));
  OR2 OR2_381(.VSS(VSS),.VDD(VDD),.Y(g27575),.A(g26147),.B(g24731));
  OR2 OR2_382(.VSS(VSS),.VDD(VDD),.Y(g26967),.A(g26350),.B(g24319));
  OR2 OR2_383(.VSS(VSS),.VDD(VDD),.Y(g33318),.A(g31969),.B(g32434));
  OR2 OR2_384(.VSS(VSS),.VDD(VDD),.Y(g34602),.A(g34489),.B(g18269));
  OR2 OR2_385(.VSS(VSS),.VDD(VDD),.Y(g25709),.A(g25014),.B(g21960));
  OR2 OR2_386(.VSS(VSS),.VDD(VDD),.Y(g30375),.A(g30149),.B(g18466));
  OR2 OR2_387(.VSS(VSS),.VDD(VDD),.Y(g34657),.A(g33114),.B(g34497));
  OR2 OR2_388(.VSS(VSS),.VDD(VDD),.Y(g28609),.A(g27346),.B(g16483));
  OR2 OR2_389(.VSS(VSS),.VDD(VDD),.Y(g33227),.A(g32029),.B(g32031));
  OR2 OR2_390(.VSS(VSS),.VDD(VDD),.Y(g9536),.A(g1351),.B(g1312));
  OR2 OR2_391(.VSS(VSS),.VDD(VDD),.Y(g33059),.A(g31987),.B(g22021));
  OR2 OR2_392(.VSS(VSS),.VDD(VDD),.Y(g33025),.A(g32162),.B(g21780));
  OR2 OR2_393(.VSS(VSS),.VDD(VDD),.Y(g25708),.A(g25526),.B(g18751));
  OR2 OR2_394(.VSS(VSS),.VDD(VDD),.Y(g34970),.A(g34868),.B(g34961));
  OR4 OR4_11(.VSS(VSS),.VDD(VDD),.Y(I29986),.A(g31070),.B(g31194),.C(g30614),.D(g30673));
  OR2 OR2_395(.VSS(VSS),.VDD(VDD),.Y(g23822),.A(g20218),.B(g16929));
  OR2 OR2_396(.VSS(VSS),.VDD(VDD),.Y(g33540),.A(g33099),.B(g18207));
  OR2 OR2_397(.VSS(VSS),.VDD(VDD),.Y(g27108),.A(g22522),.B(g25911));
  OR2 OR2_398(.VSS(VSS),.VDD(VDD),.Y(g33058),.A(g31976),.B(g22020));
  OR2 OR2_399(.VSS(VSS),.VDD(VDD),.Y(g30337),.A(g29334),.B(g18220));
  OR2 OR2_400(.VSS(VSS),.VDD(VDD),.Y(g32243),.A(g31166),.B(g29683));
  OR2 OR2_401(.VSS(VSS),.VDD(VDD),.Y(g26919),.A(g25951),.B(g18267));
  OR2 OR2_402(.VSS(VSS),.VDD(VDD),.Y(g28052),.A(g27710),.B(g18167));
  OR2 OR2_403(.VSS(VSS),.VDD(VDD),.Y(g27283),.A(g25922),.B(g25924));
  OR2 OR2_404(.VSS(VSS),.VDD(VDD),.Y(g26918),.A(g25931),.B(g18243));
  OR2 OR2_405(.VSS(VSS),.VDD(VDD),.Y(g28745),.A(g27519),.B(g16760));
  OR2 OR2_406(.VSS(VSS),.VDD(VDD),.Y(g15968),.A(g13038),.B(g10677));
  OR4 OR4_12(.VSS(VSS),.VDD(VDD),.Y(I31854),.A(g33492),.B(g33493),.C(g33494),.D(g33495));
  OR2 OR2_407(.VSS(VSS),.VDD(VDD),.Y(g33044),.A(g32199),.B(g24327));
  OR2 OR2_408(.VSS(VSS),.VDD(VDD),.Y(g34792),.A(g34750),.B(g18569));
  OR2 OR2_409(.VSS(VSS),.VDD(VDD),.Y(g32268),.A(g24785),.B(g31219));
  OR2 OR2_410(.VSS(VSS),.VDD(VDD),.Y(g23194),.A(g19564),.B(g19578));
  OR2 OR2_411(.VSS(VSS),.VDD(VDD),.Y(g33281),.A(g32142),.B(g29576));
  OR2 OR2_412(.VSS(VSS),.VDD(VDD),.Y(g31902),.A(g31744),.B(g21910));
  OR2 OR2_413(.VSS(VSS),.VDD(VDD),.Y(g30459),.A(g29314),.B(g21926));
  OR2 OR2_414(.VSS(VSS),.VDD(VDD),.Y(g30425),.A(g29770),.B(g21809));
  OR3 OR3_11(.VSS(VSS),.VDD(VDD),.Y(g33957),.A(g33523),.B(I31868),.C(I31869));
  OR2 OR2_415(.VSS(VSS),.VDD(VDD),.Y(g24347),.A(g23754),.B(g18790));
  OR2 OR2_416(.VSS(VSS),.VDD(VDD),.Y(g34459),.A(g34415),.B(g18673));
  OR2 OR2_417(.VSS(VSS),.VDD(VDD),.Y(g25602),.A(g24673),.B(g18113));
  OR2 OR2_418(.VSS(VSS),.VDD(VDD),.Y(g12982),.A(g12220),.B(g9968));
  OR2 OR2_419(.VSS(VSS),.VDD(VDD),.Y(g25657),.A(g24624),.B(g21782));
  OR2 OR2_420(.VSS(VSS),.VDD(VDD),.Y(g24253),.A(g22525),.B(g18300));
  OR2 OR2_421(.VSS(VSS),.VDD(VDD),.Y(g25774),.A(g25223),.B(g12043));
  OR2 OR2_422(.VSS(VSS),.VDD(VDD),.Y(g29246),.A(g28710),.B(g18406));
  OR2 OR2_423(.VSS(VSS),.VDD(VDD),.Y(g30458),.A(g30005),.B(g24330));
  OR2 OR2_424(.VSS(VSS),.VDD(VDD),.Y(g34458),.A(g34396),.B(g18671));
  OR2 OR2_425(.VSS(VSS),.VDD(VDD),.Y(g33562),.A(g33414),.B(g18379));
  OR2 OR2_426(.VSS(VSS),.VDD(VDD),.Y(g34010),.A(g33872),.B(g18478));
  OR2 OR2_427(.VSS(VSS),.VDD(VDD),.Y(g24236),.A(g22489),.B(g18241));
  OR2 OR2_428(.VSS(VSS),.VDD(VDD),.Y(g25878),.A(g25503),.B(g23920));
  OR2 OR2_429(.VSS(VSS),.VDD(VDD),.Y(g28732),.A(g27505),.B(g16734));
  OR2 OR2_430(.VSS(VSS),.VDD(VDD),.Y(g33699),.A(g32409),.B(g33433));
  OR2 OR2_431(.VSS(VSS),.VDD(VDD),.Y(g32993),.A(g32255),.B(g18352));
  OR2 OR2_432(.VSS(VSS),.VDD(VDD),.Y(g30545),.A(g30268),.B(g22116));
  OR2 OR2_433(.VSS(VSS),.VDD(VDD),.Y(g30444),.A(g29901),.B(g21853));
  OR2 OR2_434(.VSS(VSS),.VDD(VDD),.Y(g29776),.A(g28225),.B(g22846));
  OR3 OR3_12(.VSS(VSS),.VDD(VDD),.Y(g24952),.A(g21326),.B(g21340),.C(I24117));
  OR2 OR2_435(.VSS(VSS),.VDD(VDD),.Y(g24351),.A(g23774),.B(g18807));
  OR2 OR2_436(.VSS(VSS),.VDD(VDD),.Y(g33290),.A(g32149),.B(g29589));
  OR2 OR2_437(.VSS(VSS),.VDD(VDD),.Y(g26901),.A(g26362),.B(g24218));
  OR2 OR2_438(.VSS(VSS),.VDD(VDD),.Y(g34444),.A(g34389),.B(g18546));
  OR2 OR2_439(.VSS(VSS),.VDD(VDD),.Y(g24821),.A(g21404),.B(g23990));
  OR2 OR2_440(.VSS(VSS),.VDD(VDD),.Y(g29754),.A(g28215),.B(g28218));
  OR2 OR2_441(.VSS(VSS),.VDD(VDD),.Y(g34599),.A(g34542),.B(g18149));
  OR2 OR2_442(.VSS(VSS),.VDD(VDD),.Y(g32131),.A(g24495),.B(g30926));
  OR2 OR2_443(.VSS(VSS),.VDD(VDD),.Y(g20063),.A(g15978),.B(g13313));
  OR2 OR2_444(.VSS(VSS),.VDD(VDD),.Y(g34598),.A(g34541),.B(g18136));
  OR2 OR2_445(.VSS(VSS),.VDD(VDD),.Y(g15910),.A(g13025),.B(g10654));
  OR2 OR2_446(.VSS(VSS),.VDD(VDD),.Y(g24264),.A(g22310),.B(g18559));
  OR2 OR2_447(.VSS(VSS),.VDD(VDD),.Y(g23276),.A(g19681),.B(g16161));
  OR2 OR2_448(.VSS(VSS),.VDD(VDD),.Y(g27663),.A(g26323),.B(g24820));
  OR2 OR2_449(.VSS(VSS),.VDD(VDD),.Y(g28400),.A(g27211),.B(g15870));
  OR2 OR2_450(.VSS(VSS),.VDD(VDD),.Y(g32210),.A(g31123),.B(g29600));
  OR2 OR2_451(.VSS(VSS),.VDD(VDD),.Y(g21900),.A(g20977),.B(g15114));
  OR2 OR2_452(.VSS(VSS),.VDD(VDD),.Y(g16866),.A(g13492),.B(g11044));
  OR2 OR2_453(.VSS(VSS),.VDD(VDD),.Y(g28329),.A(g27128),.B(g15813));
  OR2 OR2_454(.VSS(VSS),.VDD(VDD),.Y(g30532),.A(g30193),.B(g22078));
  OR2 OR2_455(.VSS(VSS),.VDD(VDD),.Y(g32279),.A(g31220),.B(g31224));
  OR2 OR2_456(.VSS(VSS),.VDD(VDD),.Y(g34125),.A(g33724),.B(g33124));
  OR2 OR2_457(.VSS(VSS),.VDD(VDD),.Y(g22652),.A(g18992),.B(g15653));
  OR2 OR2_458(.VSS(VSS),.VDD(VDD),.Y(g13762),.A(g499),.B(g12527));
  OR2 OR2_459(.VSS(VSS),.VDD(VDD),.Y(g34977),.A(g34873),.B(g34966));
  OR2 OR2_460(.VSS(VSS),.VDD(VDD),.Y(g25010),.A(g23267),.B(g2932));
  OR2 OR2_461(.VSS(VSS),.VDD(VDD),.Y(g31895),.A(g31505),.B(g24296));
  OR2 OR2_462(.VSS(VSS),.VDD(VDD),.Y(g28328),.A(g27127),.B(g15812));
  OR2 OR2_463(.VSS(VSS),.VDD(VDD),.Y(g33547),.A(g33349),.B(g18331));
  OR2 OR2_464(.VSS(VSS),.VDD(VDD),.Y(g34158),.A(g33784),.B(g19740));
  OR2 OR2_465(.VSS(VSS),.VDD(VDD),.Y(g24209),.A(g23415),.B(g18122));
  OR2 OR2_466(.VSS(VSS),.VDD(VDD),.Y(g34783),.A(g33110),.B(g34667));
  OR2 OR2_467(.VSS(VSS),.VDD(VDD),.Y(g28538),.A(g27294),.B(g26206));
  OR2 OR2_468(.VSS(VSS),.VDD(VDD),.Y(g26966),.A(g26345),.B(g24318));
  OR2 OR2_469(.VSS(VSS),.VDD(VDD),.Y(g25545),.A(g23551),.B(g20658));
  OR2 OR2_470(.VSS(VSS),.VDD(VDD),.Y(g30561),.A(g30284),.B(g22132));
  OR2 OR2_471(.VSS(VSS),.VDD(VDD),.Y(g7673),.A(g4153),.B(g4172));
  OR2 OR2_472(.VSS(VSS),.VDD(VDD),.Y(g30353),.A(g30095),.B(g18355));
  OR2 OR2_473(.VSS(VSS),.VDD(VDD),.Y(g24208),.A(g23404),.B(g18121));
  OR2 OR2_474(.VSS(VSS),.VDD(VDD),.Y(g25599),.A(g24914),.B(g21721));
  OR2 OR2_475(.VSS(VSS),.VDD(VDD),.Y(g34353),.A(g26088),.B(g34114));
  OR2 OR2_476(.VSS(VSS),.VDD(VDD),.Y(g29319),.A(g28812),.B(g14453));
  OR2 OR2_477(.VSS(VSS),.VDD(VDD),.Y(g25598),.A(g24904),.B(g21720));
  OR2 OR2_478(.VSS(VSS),.VDD(VDD),.Y(g33551),.A(g33446),.B(g18342));
  OR2 OR2_479(.VSS(VSS),.VDD(VDD),.Y(g33572),.A(g33339),.B(g18414));
  OR2 OR2_480(.VSS(VSS),.VDD(VDD),.Y(g30336),.A(g29324),.B(g18203));
  OR2 OR2_481(.VSS(VSS),.VDD(VDD),.Y(g29227),.A(g28456),.B(g18169));
  OR2 OR2_482(.VSS(VSS),.VDD(VDD),.Y(g13543),.A(g10543),.B(g10565));
  OR4 OR4_13(.VSS(VSS),.VDD(VDD),.Y(I31839),.A(g33465),.B(g33466),.C(g33467),.D(g33468));
  OR4 OR4_14(.VSS(VSS),.VDD(VDD),.Y(I31838),.A(g33461),.B(g33462),.C(g33463),.D(g33464));
  OR2 OR2_483(.VSS(VSS),.VDD(VDD),.Y(g28100),.A(g27690),.B(g22051));
  OR2 OR2_484(.VSS(VSS),.VDD(VDD),.Y(g20905),.A(g7216),.B(g17264));
  OR2 OR2_485(.VSS(VSS),.VDD(VDD),.Y(g34631),.A(g34562),.B(g15118));
  OR2 OR2_486(.VSS(VSS),.VDD(VDD),.Y(g30364),.A(g30086),.B(g18411));
  OR2 OR2_487(.VSS(VSS),.VDD(VDD),.Y(g34017),.A(g33880),.B(g18504));
  OR2 OR2_488(.VSS(VSS),.VDD(VDD),.Y(g24274),.A(g23187),.B(g18631));
  OR2 OR2_489(.VSS(VSS),.VDD(VDD),.Y(g13242),.A(g11336),.B(g7601));
  OR3 OR3_13(.VSS(VSS),.VDD(VDD),.Y(g33956),.A(g33514),.B(I31863),.C(I31864));
  OR2 OR2_490(.VSS(VSS),.VDD(VDD),.Y(g24346),.A(g23725),.B(g18789));
  OR2 OR2_491(.VSS(VSS),.VDD(VDD),.Y(g33297),.A(g32157),.B(g29621));
  OR2 OR2_492(.VSS(VSS),.VDD(VDD),.Y(g25656),.A(g24945),.B(g18609));
  OR2 OR2_493(.VSS(VSS),.VDD(VDD),.Y(g31889),.A(g31118),.B(g21822));
  OR2 OR2_494(.VSS(VSS),.VDD(VDD),.Y(g33980),.A(g33843),.B(g18370));
  OR2 OR2_495(.VSS(VSS),.VDD(VDD),.Y(g24565),.A(g22309),.B(g19275));
  OR2 OR2_496(.VSS(VSS),.VDD(VDD),.Y(g21892),.A(g19788),.B(g15104));
  OR2 OR2_497(.VSS(VSS),.VDD(VDD),.Y(g25680),.A(g24794),.B(g21839));
  OR3 OR3_14(.VSS(VSS),.VDD(VDD),.Y(g16876),.A(g14028),.B(g11773),.C(g11755));
  OR2 OR2_498(.VSS(VSS),.VDD(VDD),.Y(g29281),.A(g28541),.B(g18743));
  OR2 OR2_499(.VSS(VSS),.VDD(VDD),.Y(g31888),.A(g31067),.B(g21821));
  OR2 OR2_500(.VSS(VSS),.VDD(VDD),.Y(g20034),.A(g15902),.B(g13299));
  OR2 OR2_501(.VSS(VSS),.VDD(VDD),.Y(g29301),.A(g28686),.B(g18797));
  OR2 OR2_502(.VSS(VSS),.VDD(VDD),.Y(g27509),.A(g26023),.B(g24640));
  OR2 OR2_503(.VSS(VSS),.VDD(VDD),.Y(g34289),.A(g26847),.B(g34218));
  OR2 OR2_504(.VSS(VSS),.VDD(VDD),.Y(g24641),.A(g22151),.B(g22159));
  OR2 OR2_505(.VSS(VSS),.VDD(VDD),.Y(g34023),.A(g33796),.B(g24320));
  OR2 OR2_506(.VSS(VSS),.VDD(VDD),.Y(g34288),.A(g26846),.B(g34217));
  OR2 OR2_507(.VSS(VSS),.VDD(VDD),.Y(g32217),.A(g31129),.B(g29616));
  OR2 OR2_508(.VSS(VSS),.VDD(VDD),.Y(g26954),.A(g26380),.B(g24292));
  OR3 OR3_15(.VSS(VSS),.VDD(VDD),.Y(I18449),.A(g14512),.B(g14445),.C(g14415));
  OR2 OR2_509(.VSS(VSS),.VDD(VDD),.Y(g31931),.A(g31494),.B(g22095));
  OR2 OR2_510(.VSS(VSS),.VDD(VDD),.Y(g29290),.A(g28569),.B(g18764));
  OR2 OR2_511(.VSS(VSS),.VDD(VDD),.Y(g25631),.A(g24554),.B(g18275));
  OR2 OR2_512(.VSS(VSS),.VDD(VDD),.Y(g30495),.A(g30222),.B(g21991));
  OR2 OR2_513(.VSS(VSS),.VDD(VDD),.Y(g32223),.A(g31142),.B(g29637));
  OR2 OR2_514(.VSS(VSS),.VDD(VDD),.Y(g29366),.A(g13738),.B(g28439));
  OR2 OR2_515(.VSS(VSS),.VDD(VDD),.Y(g27574),.A(g26145),.B(g24730));
  OR2 OR2_516(.VSS(VSS),.VDD(VDD),.Y(g34976),.A(g34872),.B(g34965));
  OR2 OR2_517(.VSS(VSS),.VDD(VDD),.Y(g26392),.A(g24745),.B(g23050));
  OR2 OR2_518(.VSS(VSS),.VDD(VDD),.Y(g27205),.A(g25833),.B(g24421));
  OR2 OR2_519(.VSS(VSS),.VDD(VDD),.Y(g33546),.A(g33402),.B(g18327));
  OR2 OR2_520(.VSS(VSS),.VDD(VDD),.Y(g30374),.A(g30078),.B(g18465));
  OR2 OR2_521(.VSS(VSS),.VDD(VDD),.Y(g16076),.A(g13081),.B(g10736));
  OR2 OR2_522(.VSS(VSS),.VDD(VDD),.Y(g34374),.A(g26294),.B(g34139));
  OR4 OR4_15(.VSS(VSS),.VDD(VDD),.Y(I30728),.A(g32345),.B(g32350),.C(g32056),.D(g32018));
  OR2 OR2_523(.VSS(VSS),.VDD(VDD),.Y(g33024),.A(g32324),.B(g21752));
  OR2 OR2_524(.VSS(VSS),.VDD(VDD),.Y(g34643),.A(g34554),.B(g18752));
  OR2 OR2_525(.VSS(VSS),.VDD(VDD),.Y(g28435),.A(g27234),.B(g15967));
  OR2 OR2_526(.VSS(VSS),.VDD(VDD),.Y(g28082),.A(g27369),.B(g24315));
  OR2 OR2_527(.VSS(VSS),.VDD(VDD),.Y(g26893),.A(g26753),.B(g24199));
  OR2 OR2_528(.VSS(VSS),.VDD(VDD),.Y(g29226),.A(g28455),.B(g18159));
  OR2 OR2_529(.VSS(VSS),.VDD(VDD),.Y(g28744),.A(g27518),.B(g16759));
  OR2 OR2_530(.VSS(VSS),.VDD(VDD),.Y(g34260),.A(g34113),.B(g18680));
  OR2 OR2_531(.VSS(VSS),.VDD(VDD),.Y(g28345),.A(g27137),.B(g15821));
  OR2 OR2_532(.VSS(VSS),.VDD(VDD),.Y(g29481),.A(g28117),.B(g28125));
  OR2 OR2_533(.VSS(VSS),.VDD(VDD),.Y(g30392),.A(g30091),.B(g18558));
  OR2 OR2_534(.VSS(VSS),.VDD(VDD),.Y(g30489),.A(g30250),.B(g21985));
  OR2 OR2_535(.VSS(VSS),.VDD(VDD),.Y(g33625),.A(g33373),.B(g18809));
  OR2 OR2_536(.VSS(VSS),.VDD(VDD),.Y(g32373),.A(g29894),.B(g31321));
  OR2 OR2_537(.VSS(VSS),.VDD(VDD),.Y(g33987),.A(g33847),.B(g18396));
  OR2 OR2_538(.VSS(VSS),.VDD(VDD),.Y(g31250),.A(g25972),.B(g29526));
  OR2 OR2_539(.VSS(VSS),.VDD(VDD),.Y(g25687),.A(g24729),.B(g21882));
  OR2 OR2_540(.VSS(VSS),.VDD(VDD),.Y(g30559),.A(g30269),.B(g22130));
  OR2 OR2_541(.VSS(VSS),.VDD(VDD),.Y(g30525),.A(g30266),.B(g22071));
  OR2 OR2_542(.VSS(VSS),.VDD(VDD),.Y(g30488),.A(g30197),.B(g21984));
  OR2 OR2_543(.VSS(VSS),.VDD(VDD),.Y(g30424),.A(g29760),.B(g21808));
  OR2 OR2_544(.VSS(VSS),.VDD(VDD),.Y(g25752),.A(g25079),.B(g22099));
  OR2 OR2_545(.VSS(VSS),.VDD(VDD),.Y(g34016),.A(g33867),.B(g18503));
  OR2 OR2_546(.VSS(VSS),.VDD(VDD),.Y(g30558),.A(g30258),.B(g22129));
  OR2 OR2_547(.VSS(VSS),.VDD(VDD),.Y(g27152),.A(g24393),.B(g25817));
  OR2 OR2_548(.VSS(VSS),.VDD(VDD),.Y(g33296),.A(g32156),.B(g29617));
  OR2 OR2_549(.VSS(VSS),.VDD(VDD),.Y(g25643),.A(g24602),.B(g21736));
  OR2 OR2_550(.VSS(VSS),.VDD(VDD),.Y(g29490),.A(g25832),.B(g28136));
  OR2 OR2_551(.VSS(VSS),.VDD(VDD),.Y(g16839),.A(g13473),.B(g11035));
  OR2 OR2_552(.VSS(VSS),.VDD(VDD),.Y(g28332),.A(g27130),.B(g15815));
  OR2 OR2_553(.VSS(VSS),.VDD(VDD),.Y(g30544),.A(g30257),.B(g22115));
  OR2 OR2_554(.VSS(VSS),.VDD(VDD),.Y(g33969),.A(g33864),.B(g18321));
  OR2 OR2_555(.VSS(VSS),.VDD(VDD),.Y(g25669),.A(g24657),.B(g18624));
  OR2 OR2_556(.VSS(VSS),.VDD(VDD),.Y(g28135),.A(g27959),.B(g27963));
  OR2 OR2_557(.VSS(VSS),.VDD(VDD),.Y(g29297),.A(g28683),.B(g18784));
  OR2 OR2_558(.VSS(VSS),.VDD(VDD),.Y(g33060),.A(g31992),.B(g22022));
  OR2 OR2_559(.VSS(VSS),.VDD(VDD),.Y(g33968),.A(g33855),.B(g18320));
  OR2 OR2_560(.VSS(VSS),.VDD(VDD),.Y(g26939),.A(g25907),.B(g21884));
  OR2 OR2_561(.VSS(VSS),.VDD(VDD),.Y(g25668),.A(g24646),.B(g18623));
  OR3 OR3_16(.VSS(VSS),.VDD(VDD),.Y(g33197),.A(g32342),.B(I30745),.C(I30746));
  OR2 OR2_562(.VSS(VSS),.VDD(VDD),.Y(g28361),.A(g27153),.B(g15839));
  OR2 OR2_563(.VSS(VSS),.VDD(VDD),.Y(g32216),.A(g31128),.B(g29615));
  OR2 OR2_564(.VSS(VSS),.VDD(VDD),.Y(g27405),.A(g24572),.B(g25968));
  OR2 OR2_565(.VSS(VSS),.VDD(VDD),.Y(g26938),.A(g26186),.B(g21883));
  OR2 OR2_566(.VSS(VSS),.VDD(VDD),.Y(g31870),.A(g30607),.B(g18262));
  OR3 OR3_17(.VSS(VSS),.VDD(VDD),.Y(I28147),.A(g2946),.B(g24561),.C(g28220));
  OR2 OR2_567(.VSS(VSS),.VDD(VDD),.Y(g24840),.A(g21419),.B(g23996));
  OR2 OR2_568(.VSS(VSS),.VDD(VDD),.Y(g34610),.A(g34507),.B(g18564));
  OR2 OR2_569(.VSS(VSS),.VDD(VDD),.Y(g24390),.A(g23779),.B(g21285));
  OR2 OR2_570(.VSS(VSS),.VDD(VDD),.Y(g30189),.A(g23401),.B(g28543));
  OR2 OR2_571(.VSS(VSS),.VDD(VDD),.Y(g28049),.A(g27684),.B(g18164));
  OR2 OR2_572(.VSS(VSS),.VDD(VDD),.Y(g34255),.A(g34120),.B(g24302));
  OR2 OR2_573(.VSS(VSS),.VDD(VDD),.Y(g34189),.A(g33801),.B(g33808));
  OR2 OR2_574(.VSS(VSS),.VDD(VDD),.Y(g30270),.A(g28624),.B(g27664));
  OR2 OR2_575(.VSS(VSS),.VDD(VDD),.Y(g28048),.A(g27362),.B(g18163));
  OR2 OR2_576(.VSS(VSS),.VDD(VDD),.Y(g20522),.A(g691),.B(g16893));
  OR2 OR2_577(.VSS(VSS),.VDD(VDD),.Y(g26875),.A(g21652),.B(g25575));
  OR2 OR2_578(.VSS(VSS),.VDD(VDD),.Y(g32117),.A(g24482),.B(g30914));
  OR4 OR4_16(.VSS(VSS),.VDD(VDD),.Y(I23163),.A(g20982),.B(g21127),.C(g21193),.D(g21256));
  OR2 OR2_579(.VSS(VSS),.VDD(VDD),.Y(g31894),.A(g30671),.B(g21870));
  OR2 OR2_580(.VSS(VSS),.VDD(VDD),.Y(g31867),.A(g31238),.B(g18175));
  OR2 OR2_581(.VSS(VSS),.VDD(VDD),.Y(g30460),.A(g30207),.B(g21931));
  OR2 OR2_582(.VSS(VSS),.VDD(VDD),.Y(g30383),.A(g30138),.B(g18513));
  OR2 OR2_583(.VSS(VSS),.VDD(VDD),.Y(g34460),.A(g34301),.B(g18677));
  OR2 OR2_584(.VSS(VSS),.VDD(VDD),.Y(g30093),.A(g28467),.B(g11397));
  OR2 OR2_585(.VSS(VSS),.VDD(VDD),.Y(g34030),.A(g33727),.B(g18704));
  OR2 OR2_586(.VSS(VSS),.VDD(VDD),.Y(g25713),.A(g25147),.B(g21964));
  OR2 OR2_587(.VSS(VSS),.VDD(VDD),.Y(g28613),.A(g27350),.B(g26310));
  OR2 OR2_588(.VSS(VSS),.VDD(VDD),.Y(g33581),.A(g33333),.B(g18443));
  OR2 OR2_589(.VSS(VSS),.VDD(VDD),.Y(g33714),.A(g32419),.B(g33450));
  OR4 OR4_17(.VSS(VSS),.VDD(VDD),.Y(g29520),.A(g28291),.B(g28281),.C(g28264),.D(g28254));
  OR2 OR2_590(.VSS(VSS),.VDD(VDD),.Y(g34267),.A(g34079),.B(g18728));
  OR2 OR2_591(.VSS(VSS),.VDD(VDD),.Y(g34294),.A(g26855),.B(g34225));
  OR2 OR2_592(.VSS(VSS),.VDD(VDD),.Y(g31315),.A(g29607),.B(g29623));
  OR2 OR2_593(.VSS(VSS),.VDD(VDD),.Y(g33315),.A(g29665),.B(g32175));
  OR2 OR2_594(.VSS(VSS),.VDD(VDD),.Y(g31910),.A(g31471),.B(g21957));
  OR2 OR2_595(.VSS(VSS),.VDD(VDD),.Y(g13006),.A(g12284),.B(g10034));
  OR2 OR2_596(.VSS(VSS),.VDD(VDD),.Y(g25610),.A(g24923),.B(g18127));
  OR2 OR2_597(.VSS(VSS),.VDD(VDD),.Y(g31257),.A(g29531),.B(g28253));
  OR2 OR2_598(.VSS(VSS),.VDD(VDD),.Y(g25705),.A(g25069),.B(g18744));
  OR2 OR2_599(.VSS(VSS),.VDD(VDD),.Y(g28605),.A(g27341),.B(g26302));
  OR2 OR2_600(.VSS(VSS),.VDD(VDD),.Y(g33257),.A(g32108),.B(g29519));
  OR2 OR2_601(.VSS(VSS),.VDD(VDD),.Y(g32123),.A(g30915),.B(g30919));
  OR2 OR2_602(.VSS(VSS),.VDD(VDD),.Y(g33979),.A(g33942),.B(g18361));
  OR2 OR2_603(.VSS(VSS),.VDD(VDD),.Y(g33055),.A(g31986),.B(g21976));
  OR2 OR2_604(.VSS(VSS),.VDD(VDD),.Y(g16187),.A(g8822),.B(g13486));
  OR2 OR2_605(.VSS(VSS),.VDD(VDD),.Y(g25679),.A(g24728),.B(g21836));
  OR2 OR2_606(.VSS(VSS),.VDD(VDD),.Y(g33070),.A(g32010),.B(g22114));
  OR2 OR2_607(.VSS(VSS),.VDD(VDD),.Y(g33978),.A(g33892),.B(g18356));
  OR2 OR2_608(.VSS(VSS),.VDD(VDD),.Y(g25678),.A(g24709),.B(g21835));
  OR2 OR2_609(.VSS(VSS),.VDD(VDD),.Y(g26915),.A(g25900),.B(g18230));
  OR2 OR2_610(.VSS(VSS),.VDD(VDD),.Y(g33590),.A(g33358),.B(g18470));
  OR2 OR2_611(.VSS(VSS),.VDD(VDD),.Y(g15965),.A(g13035),.B(g10675));
  OR2 OR2_612(.VSS(VSS),.VDD(VDD),.Y(g28371),.A(g27177),.B(g15847));
  OR4 OR4_18(.VSS(VSS),.VDD(VDD),.Y(I30745),.A(g31777),.B(g32321),.C(g32069),.D(g32084));
  OR2 OR2_613(.VSS(VSS),.VDD(VDD),.Y(g32230),.A(g30589),.B(g29345));
  OR2 OR2_614(.VSS(VSS),.VDD(VDD),.Y(g33986),.A(g33639),.B(g18387));
  OR2 OR2_615(.VSS(VSS),.VDD(VDD),.Y(g24252),.A(g22518),.B(g18299));
  OR2 OR2_616(.VSS(VSS),.VDD(VDD),.Y(g25686),.A(g24712),.B(g21881));
  OR2 OR2_617(.VSS(VSS),.VDD(VDD),.Y(g33384),.A(g32248),.B(g29943));
  OR2 OR2_618(.VSS(VSS),.VDD(VDD),.Y(g33067),.A(g31989),.B(g22111));
  OR2 OR2_619(.VSS(VSS),.VDD(VDD),.Y(g12768),.A(g7785),.B(g7202));
  OR2 OR2_620(.VSS(VSS),.VDD(VDD),.Y(g29250),.A(g28695),.B(g18460));
  OR2 OR2_621(.VSS(VSS),.VDD(VDD),.Y(g32992),.A(g32242),.B(g18351));
  OR2 OR2_622(.VSS(VSS),.VDD(VDD),.Y(g32391),.A(g31502),.B(g29982));
  OR2 OR2_623(.VSS(VSS),.VDD(VDD),.Y(g30455),.A(g30041),.B(g21864));
  OR2 OR2_624(.VSS(VSS),.VDD(VDD),.Y(g34455),.A(g34284),.B(g18668));
  OR3 OR3_18(.VSS(VSS),.VDD(VDD),.Y(g11372),.A(g490),.B(g482),.C(g8038));
  OR2 OR2_625(.VSS(VSS),.VDD(VDD),.Y(g31877),.A(g31278),.B(g21732));
  OR2 OR2_626(.VSS(VSS),.VDD(VDD),.Y(g30470),.A(g30165),.B(g21941));
  OR2 OR2_627(.VSS(VSS),.VDD(VDD),.Y(g34617),.A(g34526),.B(g18579));
  OR2 OR2_628(.VSS(VSS),.VDD(VDD),.Y(g22648),.A(g18987),.B(g15652));
  OR3 OR3_19(.VSS(VSS),.VDD(VDD),.Y(I12611),.A(g1500),.B(g1582),.C(g1333));
  OR2 OR2_629(.VSS(VSS),.VDD(VDD),.Y(g29296),.A(g28586),.B(g18781));
  OR2 OR2_630(.VSS(VSS),.VDD(VDD),.Y(g33019),.A(g32339),.B(g18536));
  OR2 OR2_631(.VSS(VSS),.VDD(VDD),.Y(g30201),.A(g23412),.B(g28557));
  OR2 OR2_632(.VSS(VSS),.VDD(VDD),.Y(g33018),.A(g32312),.B(g18525));
  OR4 OR4_19(.VSS(VSS),.VDD(VDD),.Y(I30761),.A(g32071),.B(g32167),.C(g32067),.D(g32082));
  OR2 OR2_633(.VSS(VSS),.VDD(VDD),.Y(g30467),.A(g30185),.B(g21938));
  OR2 OR2_634(.VSS(VSS),.VDD(VDD),.Y(g30494),.A(g30209),.B(g21990));
  OR2 OR2_635(.VSS(VSS),.VDD(VDD),.Y(g34467),.A(g34341),.B(g18717));
  OR2 OR2_636(.VSS(VSS),.VDD(VDD),.Y(g34494),.A(g26849),.B(g34413));
  OR2 OR2_637(.VSS(VSS),.VDD(VDD),.Y(g29197),.A(g27187),.B(g27163));
  OR2 OR2_638(.VSS(VSS),.VDD(VDD),.Y(g34623),.A(g34525),.B(g18585));
  OR2 OR2_639(.VSS(VSS),.VDD(VDD),.Y(g34037),.A(g33803),.B(g18734));
  OR4 OR4_20(.VSS(VSS),.VDD(VDD),.Y(I30400),.A(g31021),.B(g30937),.C(g31327),.D(g30614));
  OR2 OR2_640(.VSS(VSS),.VDD(VDD),.Y(g27248),.A(g24880),.B(g25953));
  OR2 OR2_641(.VSS(VSS),.VDD(VDD),.Y(g30984),.A(g29765),.B(g29755));
  OR2 OR2_642(.VSS(VSS),.VDD(VDD),.Y(g27552),.A(g26092),.B(g24676));
  OR2 OR2_643(.VSS(VSS),.VDD(VDD),.Y(g31917),.A(g31478),.B(g22003));
  OR2 OR2_644(.VSS(VSS),.VDD(VDD),.Y(g30419),.A(g29759),.B(g21803));
  OR2 OR2_645(.VSS(VSS),.VDD(VDD),.Y(g31866),.A(g31252),.B(g18142));
  OR2 OR2_646(.VSS(VSS),.VDD(VDD),.Y(g30352),.A(g30094),.B(g18340));
  OR2 OR2_647(.VSS(VSS),.VDD(VDD),.Y(g27779),.A(g17317),.B(g26694));
  OR2 OR2_648(.VSS(VSS),.VDD(VDD),.Y(g25617),.A(g25466),.B(g18189));
  OR2 OR2_649(.VSS(VSS),.VDD(VDD),.Y(g24213),.A(g23220),.B(g18186));
  OR3 OR3_20(.VSS(VSS),.VDD(VDD),.Y(g23184),.A(g20198),.B(g20185),.C(I22280));
  OR2 OR2_650(.VSS(VSS),.VDD(VDD),.Y(g28724),.A(g27491),.B(g16707));
  OR2 OR2_651(.VSS(VSS),.VDD(VDD),.Y(g34352),.A(g26079),.B(g34109));
  OR2 OR2_652(.VSS(VSS),.VDD(VDD),.Y(g28359),.A(g27151),.B(g15838));
  OR2 OR2_653(.VSS(VSS),.VDD(VDD),.Y(g30418),.A(g29751),.B(g21802));
  OR2 OR2_654(.VSS(VSS),.VDD(VDD),.Y(g32275),.A(g31210),.B(g29732));
  OR2 OR2_655(.VSS(VSS),.VDD(VDD),.Y(g31001),.A(g29360),.B(g28151));
  OR2 OR2_656(.VSS(VSS),.VDD(VDD),.Y(g28358),.A(g27149),.B(g15837));
  OR2 OR2_657(.VSS(VSS),.VDD(VDD),.Y(g34266),.A(g34076),.B(g18719));
  OR2 OR2_658(.VSS(VSS),.VDD(VDD),.Y(g33001),.A(g32282),.B(g18404));
  OR2 OR2_659(.VSS(VSS),.VDD(VDD),.Y(g34170),.A(g33790),.B(g19855));
  OR2 OR2_660(.VSS(VSS),.VDD(VDD),.Y(g24205),.A(g23006),.B(g18109));
  OR2 OR2_661(.VSS(VSS),.VDD(VDD),.Y(g33706),.A(g32412),.B(g33440));
  OR2 OR2_662(.VSS(VSS),.VDD(VDD),.Y(g33597),.A(g33344),.B(g18495));
  OR2 OR2_663(.VSS(VSS),.VDD(VDD),.Y(g32237),.A(g31153),.B(g29667));
  OR2 OR2_664(.VSS(VSS),.VDD(VDD),.Y(g31256),.A(g25983),.B(g29537));
  OR2 OR2_665(.VSS(VSS),.VDD(VDD),.Y(g33256),.A(g32107),.B(g29517));
  OR2 OR2_666(.VSS(VSS),.VDD(VDD),.Y(g25595),.A(g24835),.B(g21717));
  OR2 OR2_667(.VSS(VSS),.VDD(VDD),.Y(g31923),.A(g31763),.B(g22048));
  OR2 OR2_668(.VSS(VSS),.VDD(VDD),.Y(g32983),.A(g31990),.B(g18222));
  OR2 OR2_669(.VSS(VSS),.VDD(VDD),.Y(g19879),.A(g15841),.B(g13265));
  OR2 OR2_670(.VSS(VSS),.VDD(VDD),.Y(g28344),.A(g27136),.B(g15820));
  OR2 OR2_671(.VSS(VSS),.VDD(VDD),.Y(g22832),.A(g19354),.B(g15722));
  OR2 OR2_672(.VSS(VSS),.VDD(VDD),.Y(g33280),.A(g32141),.B(g29574));
  OR2 OR2_673(.VSS(VSS),.VDD(VDD),.Y(g25623),.A(g24552),.B(g18219));
  OR2 OR2_674(.VSS(VSS),.VDD(VDD),.Y(g20051),.A(g15936),.B(g13306));
  OR2 OR2_675(.VSS(VSS),.VDD(VDD),.Y(g25037),.A(g23103),.B(g19911));
  OR2 OR2_676(.VSS(VSS),.VDD(VDD),.Y(g33624),.A(g33371),.B(g18808));
  OR2 OR2_677(.VSS(VSS),.VDD(VDD),.Y(g34167),.A(g33786),.B(g19768));
  OR2 OR2_678(.VSS(VSS),.VDD(VDD),.Y(g34194),.A(g33811),.B(g33815));
  OR4 OR4_21(.VSS(VSS),.VDD(VDD),.Y(g26616),.A(g24881),.B(g24855),.C(g24843),.D(g24822));
  OR2 OR2_679(.VSS(VSS),.VDD(VDD),.Y(g19337),.A(g17770),.B(g17785));
  OR2 OR2_680(.VSS(VSS),.VDD(VDD),.Y(g28682),.A(g27430),.B(g16635));
  OR2 OR2_681(.VSS(VSS),.VDD(VDD),.Y(g29257),.A(g28228),.B(g18600));
  OR4 OR4_22(.VSS(VSS),.VDD(VDD),.Y(I23755),.A(g22904),.B(g22927),.C(g22980),.D(g23444));
  OR2 OR2_682(.VSS(VSS),.VDD(VDD),.Y(g30524),.A(g30255),.B(g22070));
  OR2 OR2_683(.VSS(VSS),.VDD(VDD),.Y(g27233),.A(g25876),.B(g24451));
  OR2 OR2_684(.VSS(VSS),.VDD(VDD),.Y(g16800),.A(g13436),.B(g11027));
  OR2 OR2_685(.VSS(VSS),.VDD(VDD),.Y(g29496),.A(g28567),.B(g27615));
  OR2 OR2_686(.VSS(VSS),.VDD(VDD),.Y(g27182),.A(g25818),.B(g24410));
  OR2 OR2_687(.VSS(VSS),.VDD(VDD),.Y(g30401),.A(g29782),.B(g21760));
  OR2 OR2_688(.VSS(VSS),.VDD(VDD),.Y(g30477),.A(g30239),.B(g21948));
  OR2 OR2_689(.VSS(VSS),.VDD(VDD),.Y(g26305),.A(g24556),.B(g24564));
  OR2 OR2_690(.VSS(VSS),.VDD(VDD),.Y(g24350),.A(g23755),.B(g18806));
  OR2 OR2_691(.VSS(VSS),.VDD(VDD),.Y(g26809),.A(g24930),.B(g24939));
  OR2 OR2_692(.VSS(VSS),.VDD(VDD),.Y(g33066),.A(g32341),.B(g22096));
  OR2 OR2_693(.VSS(VSS),.VDD(VDD),.Y(g26900),.A(g26819),.B(g24217));
  OR2 OR2_694(.VSS(VSS),.VDD(VDD),.Y(g33231),.A(g32032),.B(g32036));
  OR2 OR2_695(.VSS(VSS),.VDD(VDD),.Y(g29741),.A(g28205),.B(g15883));
  OR2 OR2_696(.VSS(VSS),.VDD(VDD),.Y(g32130),.A(g30921),.B(g30925));
  OR2 OR2_697(.VSS(VSS),.VDD(VDD),.Y(g34022),.A(g33873),.B(g18538));
  OR2 OR2_698(.VSS(VSS),.VDD(VDD),.Y(g28134),.A(g27958),.B(g27962));
  OR2 OR2_699(.VSS(VSS),.VDD(VDD),.Y(g31876),.A(g31125),.B(g21731));
  OR2 OR2_700(.VSS(VSS),.VDD(VDD),.Y(g31885),.A(g31017),.B(g21779));
  OR2 OR2_701(.VSS(VSS),.VDD(VDD),.Y(g32362),.A(g29870),.B(g31301));
  OR2 OR2_702(.VSS(VSS),.VDD(VDD),.Y(g34616),.A(g34519),.B(g18577));
  OR2 OR2_703(.VSS(VSS),.VDD(VDD),.Y(g25589),.A(g21690),.B(g24159));
  OR2 OR2_704(.VSS(VSS),.VDD(VDD),.Y(g29801),.A(g25987),.B(g28251));
  OR2 OR2_705(.VSS(VSS),.VDD(VDD),.Y(g29735),.A(g28202),.B(g10898));
  OR2 OR2_706(.VSS(VSS),.VDD(VDD),.Y(g25588),.A(g21686),.B(g24158));
  OR2 OR2_707(.VSS(VSS),.VDD(VDD),.Y(g34305),.A(g25775),.B(g34050));
  OR2 OR2_708(.VSS(VSS),.VDD(VDD),.Y(g25836),.A(g25368),.B(g23856));
  OR2 OR2_709(.VSS(VSS),.VDD(VDD),.Y(g27026),.A(g26828),.B(g17726));
  OR2 OR2_710(.VSS(VSS),.VDD(VDD),.Y(g34254),.A(g34116),.B(g24301));
  OR2 OR2_711(.VSS(VSS),.VDD(VDD),.Y(g30466),.A(g30174),.B(g21937));
  OR2 OR2_712(.VSS(VSS),.VDD(VDD),.Y(g34809),.A(g33677),.B(g34738));
  OR2 OR2_713(.VSS(VSS),.VDD(VDD),.Y(g34900),.A(g34860),.B(g21686));
  OR2 OR2_714(.VSS(VSS),.VDD(VDD),.Y(g26733),.A(g10776),.B(g24447));
  OR2 OR2_715(.VSS(VSS),.VDD(VDD),.Y(g34466),.A(g34337),.B(g18716));
  OR2 OR2_716(.VSS(VSS),.VDD(VDD),.Y(g34808),.A(g34765),.B(g18599));
  OR2 OR2_717(.VSS(VSS),.VDD(VDD),.Y(g32222),.A(g31141),.B(g29636));
  OR3 OR3_21(.VSS(VSS),.VDD(VDD),.Y(g23771),.A(g21432),.B(g21416),.C(I22912));
  OR2 OR2_718(.VSS(VSS),.VDD(VDD),.Y(g26874),.A(I25612),.B(I25613));
  OR2 OR2_719(.VSS(VSS),.VDD(VDD),.Y(g34036),.A(g33722),.B(g18715));
  OR2 OR2_720(.VSS(VSS),.VDD(VDD),.Y(g30560),.A(g30278),.B(g22131));
  OR2 OR2_721(.VSS(VSS),.VDD(VDD),.Y(g34101),.A(g33693),.B(g33700));
  OR2 OR2_722(.VSS(VSS),.VDD(VDD),.Y(g31916),.A(g31756),.B(g22002));
  OR2 OR2_723(.VSS(VSS),.VDD(VDD),.Y(g34642),.A(g34482),.B(g18725));
  OR2 OR2_724(.VSS(VSS),.VDD(VDD),.Y(g25749),.A(g25094),.B(g18800));
  OR2 OR2_725(.VSS(VSS),.VDD(VDD),.Y(g25616),.A(g25096),.B(g18172));
  OR2 OR2_726(.VSS(VSS),.VDD(VDD),.Y(g28649),.A(g27390),.B(g16597));
  OR2 OR2_727(.VSS(VSS),.VDD(VDD),.Y(g33550),.A(g33342),.B(g18338));
  OR2 OR2_728(.VSS(VSS),.VDD(VDD),.Y(g32347),.A(g29839),.B(g31273));
  OR2 OR2_729(.VSS(VSS),.VDD(VDD),.Y(g33314),.A(g29663),.B(g32174));
  OR2 OR2_730(.VSS(VSS),.VDD(VDD),.Y(g31287),.A(g29578),.B(g28292));
  OR2 OR2_731(.VSS(VSS),.VDD(VDD),.Y(g15800),.A(g10821),.B(g13242));
  OR2 OR2_732(.VSS(VSS),.VDD(VDD),.Y(g32253),.A(g24771),.B(g31207));
  OR2 OR2_733(.VSS(VSS),.VDD(VDD),.Y(g25748),.A(g25078),.B(g18799));
  OR2 OR2_734(.VSS(VSS),.VDD(VDD),.Y(g33287),.A(g32146),.B(g29586));
  OR2 OR2_735(.VSS(VSS),.VDD(VDD),.Y(g34064),.A(g33919),.B(g33922));
  OR2 OR2_736(.VSS(VSS),.VDD(VDD),.Y(g30733),.A(g13807),.B(g29773));
  OR2 OR2_737(.VSS(VSS),.VDD(VDD),.Y(g31307),.A(g29596),.B(g28311));
  OR2 OR2_738(.VSS(VSS),.VDD(VDD),.Y(g33076),.A(g32336),.B(g32446));
  OR2 OR2_739(.VSS(VSS),.VDD(VDD),.Y(g34733),.A(g34678),.B(g18651));
  OR2 OR2_740(.VSS(VSS),.VDD(VDD),.Y(g26892),.A(g26719),.B(g24198));
  OR2 OR2_741(.VSS(VSS),.VDD(VDD),.Y(g25704),.A(g25173),.B(g21925));
  OR2 OR2_742(.VSS(VSS),.VDD(VDD),.Y(g22447),.A(g21464),.B(g12761));
  OR2 OR2_743(.VSS(VSS),.VDD(VDD),.Y(g33596),.A(g33341),.B(g18494));
  OR2 OR2_744(.VSS(VSS),.VDD(VDD),.Y(g33054),.A(g31975),.B(g21975));
  OR2 OR2_745(.VSS(VSS),.VDD(VDD),.Y(g32236),.A(g31152),.B(g29664));
  OR2 OR2_746(.VSS(VSS),.VDD(VDD),.Y(g8790),.A(I12782),.B(I12783));
  OR2 OR2_747(.VSS(VSS),.VDD(VDD),.Y(g32351),.A(g29851),.B(g31281));
  OR2 OR2_748(.VSS(VSS),.VDD(VDD),.Y(g32372),.A(g29884),.B(g31314));
  OR2 OR2_749(.VSS(VSS),.VDD(VDD),.Y(g34630),.A(g34560),.B(g15117));
  OR2 OR2_750(.VSS(VSS),.VDD(VDD),.Y(g34693),.A(g34513),.B(g34310));
  OR2 OR2_751(.VSS(VSS),.VDD(VDD),.Y(g24282),.A(g23407),.B(g18657));
  OR2 OR2_752(.VSS(VSS),.VDD(VDD),.Y(g26914),.A(g25949),.B(g18227));
  OR2 OR2_753(.VSS(VSS),.VDD(VDD),.Y(g29706),.A(g28198),.B(g27208));
  OR2 OR2_754(.VSS(VSS),.VDD(VDD),.Y(g8461),.A(g301),.B(g534));
  OR2 OR2_755(.VSS(VSS),.VDD(VDD),.Y(g31269),.A(g26024),.B(g29569));
  OR2 OR2_756(.VSS(VSS),.VDD(VDD),.Y(g34166),.A(g33785),.B(g19752));
  OR2 OR2_757(.VSS(VSS),.VDD(VDD),.Y(g34009),.A(g33863),.B(g18477));
  OR2 OR2_758(.VSS(VSS),.VDD(VDD),.Y(g19336),.A(g17769),.B(g14831));
  OR2 OR2_759(.VSS(VSS),.VDD(VDD),.Y(g26907),.A(g26513),.B(g24224));
  OR2 OR2_760(.VSS(VSS),.VDD(VDD),.Y(g29256),.A(g28597),.B(g18533));
  OR2 OR2_761(.VSS(VSS),.VDD(VDD),.Y(g31773),.A(g30044),.B(g30056));
  OR4 OR4_23(.VSS(VSS),.VDD(VDD),.Y(I30399),.A(g29385),.B(g31376),.C(g30735),.D(g30825));
  OR2 OR2_762(.VSS(VSS),.VDD(VDD),.Y(g31268),.A(g29552),.B(g28266));
  OR2 OR2_763(.VSS(VSS),.VDD(VDD),.Y(g32264),.A(g31187),.B(g29711));
  OR2 OR2_764(.VSS(VSS),.VDD(VDD),.Y(g34008),.A(g33849),.B(g18476));
  OR2 OR2_765(.VSS(VSS),.VDD(VDD),.Y(g29280),.A(g28530),.B(g18742));
  OR2 OR2_766(.VSS(VSS),.VDD(VDD),.Y(g33268),.A(g32116),.B(g29538));
  OR2 OR2_767(.VSS(VSS),.VDD(VDD),.Y(g30476),.A(g30229),.B(g21947));
  OR2 OR2_768(.VSS(VSS),.VDD(VDD),.Y(g30485),.A(g30166),.B(g21981));
  OR2 OR2_769(.VSS(VSS),.VDD(VDD),.Y(g29300),.A(g28666),.B(g18796));
  OR2 OR2_770(.VSS(VSS),.VDD(VDD),.Y(g31670),.A(g29937),.B(g28573));
  OR2 OR2_771(.VSS(VSS),.VDD(VDD),.Y(g8904),.A(g1779),.B(g1798));
  OR4 OR4_24(.VSS(VSS),.VDD(VDD),.Y(I31863),.A(g33506),.B(g33507),.C(g33508),.D(g33509));
  OR2 OR2_772(.VSS(VSS),.VDD(VDD),.Y(g30555),.A(g30227),.B(g22126));
  OR2 OR2_773(.VSS(VSS),.VDD(VDD),.Y(g30454),.A(g29909),.B(g21863));
  OR2 OR2_774(.VSS(VSS),.VDD(VDD),.Y(g34454),.A(g34414),.B(g18667));
  OR2 OR2_775(.VSS(VSS),.VDD(VDD),.Y(g25733),.A(g25108),.B(g18778));
  OR3 OR3_22(.VSS(VSS),.VDD(VDD),.Y(g13091),.A(g329),.B(g319),.C(g10796));
  OR2 OR2_776(.VSS(VSS),.VDD(VDD),.Y(g22591),.A(g18893),.B(g18909));
  OR2 OR2_777(.VSS(VSS),.VDD(VDD),.Y(g27133),.A(g25788),.B(g24392));
  OR2 OR2_778(.VSS(VSS),.VDD(VDD),.Y(g28719),.A(g27485),.B(g16703));
  OR4 OR4_25(.VSS(VSS),.VDD(VDD),.Y(g28191),.A(g27217),.B(g27210),.C(g27186),.D(g27162));
  OR2 OR2_779(.VSS(VSS),.VDD(VDD),.Y(g31930),.A(g31769),.B(g22094));
  OR2 OR2_780(.VSS(VSS),.VDD(VDD),.Y(g32209),.A(g31122),.B(g29599));
  OR2 OR2_781(.VSS(VSS),.VDD(VDD),.Y(g33993),.A(g33646),.B(g18413));
  OR2 OR2_782(.VSS(VSS),.VDD(VDD),.Y(g25630),.A(g24532),.B(g18263));
  OR2 OR2_783(.VSS(VSS),.VDD(VDD),.Y(g28718),.A(g27483),.B(g16702));
  OR2 OR2_784(.VSS(VSS),.VDD(VDD),.Y(g25693),.A(g24627),.B(g18707));
  OR2 OR2_785(.VSS(VSS),.VDD(VDD),.Y(g29231),.A(g28301),.B(g18229));
  OR2 OR2_786(.VSS(VSS),.VDD(VDD),.Y(g33694),.A(g32402),.B(g33429));
  OR2 OR2_787(.VSS(VSS),.VDD(VDD),.Y(g32208),.A(g31120),.B(g29584));
  OR2 OR2_788(.VSS(VSS),.VDD(VDD),.Y(g33965),.A(g33805),.B(g18179));
  OR4 OR4_26(.VSS(VSS),.VDD(VDD),.Y(I12783),.A(g4204),.B(g4207),.C(g4210),.D(g4180));
  OR2 OR2_789(.VSS(VSS),.VDD(VDD),.Y(g25665),.A(g24708),.B(g21790));
  OR2 OR2_790(.VSS(VSS),.VDD(VDD),.Y(g34239),.A(g32845),.B(g33957));
  OR2 OR2_791(.VSS(VSS),.VDD(VDD),.Y(g34238),.A(g32780),.B(g33956));
  OR2 OR2_792(.VSS(VSS),.VDD(VDD),.Y(g23345),.A(g19735),.B(g16203));
  OR2 OR2_793(.VSS(VSS),.VDD(VDD),.Y(g26883),.A(g26670),.B(g24189));
  OR4 OR4_27(.VSS(VSS),.VDD(VDD),.Y(I23162),.A(g19919),.B(g19968),.C(g20014),.D(g20841));
  OR2 OR2_794(.VSS(VSS),.VDD(VDD),.Y(g33619),.A(g33359),.B(g18758));
  OR2 OR2_795(.VSS(VSS),.VDD(VDD),.Y(g33557),.A(g33331),.B(g18363));
  OR2 OR2_796(.VSS(VSS),.VDD(VDD),.Y(g29763),.A(g28217),.B(g22762));
  OR2 OR2_797(.VSS(VSS),.VDD(VDD),.Y(g30382),.A(g30137),.B(g18498));
  OR2 OR2_798(.VSS(VSS),.VDD(VDD),.Y(g30519),.A(g30264),.B(g22040));
  OR2 OR2_799(.VSS(VSS),.VDD(VDD),.Y(g33618),.A(g33353),.B(g18757));
  OR2 OR2_800(.VSS(VSS),.VDD(VDD),.Y(g28389),.A(g27206),.B(g15860));
  OR2 OR2_801(.VSS(VSS),.VDD(VDD),.Y(g30176),.A(g23392),.B(g28531));
  OR2 OR2_802(.VSS(VSS),.VDD(VDD),.Y(g28045),.A(g27378),.B(g18141));
  OR2 OR2_803(.VSS(VSS),.VDD(VDD),.Y(g30092),.A(g28466),.B(g16699));
  OR2 OR2_804(.VSS(VSS),.VDD(VDD),.Y(g31279),.A(g29571),.B(g29579));
  OR2 OR2_805(.VSS(VSS),.VDD(VDD),.Y(g24249),.A(g22624),.B(g18294));
  OR2 OR2_806(.VSS(VSS),.VDD(VDD),.Y(g33279),.A(g32140),.B(g29573));
  OR2 OR2_807(.VSS(VSS),.VDD(VDD),.Y(g25712),.A(g25126),.B(g21963));
  OR2 OR2_808(.VSS(VSS),.VDD(VDD),.Y(g28099),.A(g27992),.B(g22043));
  OR2 OR2_809(.VSS(VSS),.VDD(VDD),.Y(g30518),.A(g30254),.B(g22039));
  OR3 OR3_23(.VSS(VSS),.VDD(VDD),.Y(I22280),.A(g20271),.B(g20150),.C(g20134));
  OR2 OR2_810(.VSS(VSS),.VDD(VDD),.Y(g28388),.A(g27204),.B(g15859));
  OR2 OR2_811(.VSS(VSS),.VDD(VDD),.Y(g16430),.A(g182),.B(g13657));
  OR2 OR2_812(.VSS(VSS),.VDD(VDD),.Y(g28701),.A(g27455),.B(g16669));
  OR2 OR2_813(.VSS(VSS),.VDD(VDD),.Y(g24248),.A(g22710),.B(g18286));
  OR2 OR2_814(.VSS(VSS),.VDD(VDD),.Y(g33278),.A(g32139),.B(g29572));
  OR2 OR2_815(.VSS(VSS),.VDD(VDD),.Y(g12925),.A(g8928),.B(g10511));
  OR2 OR2_816(.VSS(VSS),.VDD(VDD),.Y(g28777),.A(g27539),.B(g16807));
  OR2 OR2_817(.VSS(VSS),.VDD(VDD),.Y(g28534),.A(g27292),.B(g26204));
  OR2 OR2_818(.VSS(VSS),.VDD(VDD),.Y(g28098),.A(g27683),.B(g22016));
  OR2 OR2_819(.VSS(VSS),.VDD(VDD),.Y(g32346),.A(g29838),.B(g31272));
  OR2 OR2_820(.VSS(VSS),.VDD(VDD),.Y(g34637),.A(g34478),.B(g18694));
  OR2 OR2_821(.VSS(VSS),.VDD(VDD),.Y(g24204),.A(g22990),.B(g18108));
  OR2 OR2_822(.VSS(VSS),.VDD(VDD),.Y(g33286),.A(g32145),.B(g29585));
  OR2 OR2_823(.VSS(VSS),.VDD(VDD),.Y(g31468),.A(g29641),.B(g29656));
  OR2 OR2_824(.VSS(VSS),.VDD(VDD),.Y(g31306),.A(g29595),.B(g29610));
  OR4 OR4_28(.VSS(VSS),.VDD(VDD),.Y(I31873),.A(g33524),.B(g33525),.C(g33526),.D(g33527));
  OR2 OR2_825(.VSS(VSS),.VDD(VDD),.Y(g33039),.A(g32187),.B(g24312));
  OR2 OR2_826(.VSS(VSS),.VDD(VDD),.Y(g29480),.A(g28115),.B(g22172));
  OR2 OR2_827(.VSS(VSS),.VDD(VDD),.Y(g27742),.A(g17292),.B(g26673));
  OR2 OR2_828(.VSS(VSS),.VDD(VDD),.Y(g22318),.A(g21394),.B(g17783));
  OR2 OR2_829(.VSS(VSS),.VDD(VDD),.Y(g25594),.A(g24772),.B(g21708));
  OR2 OR2_830(.VSS(VSS),.VDD(VDD),.Y(g33038),.A(g32184),.B(g24311));
  OR2 OR2_831(.VSS(VSS),.VDD(VDD),.Y(g29287),.A(g28555),.B(g18760));
  OR2 OR2_832(.VSS(VSS),.VDD(VDD),.Y(g29307),.A(g28706),.B(g18814));
  OR2 OR2_833(.VSS(VSS),.VDD(VDD),.Y(g28140),.A(I26643),.B(I26644));
  OR2 OR2_834(.VSS(VSS),.VDD(VDD),.Y(g26349),.A(g24630),.B(g13409));
  OR2 OR2_835(.VSS(VSS),.VDD(VDD),.Y(g33601),.A(g33422),.B(g18508));
  OR2 OR2_836(.VSS(VSS),.VDD(VDD),.Y(g25941),.A(g24416),.B(g22219));
  OR3 OR3_24(.VSS(VSS),.VDD(VDD),.Y(g33187),.A(g32014),.B(I30740),.C(I30741));
  OR2 OR2_837(.VSS(VSS),.VDD(VDD),.Y(g33975),.A(g33860),.B(g18346));
  OR2 OR2_838(.VSS(VSS),.VDD(VDD),.Y(g27429),.A(g25969),.B(g24589));
  OR2 OR2_839(.VSS(VSS),.VDD(VDD),.Y(g26906),.A(g26423),.B(g24223));
  OR2 OR2_840(.VSS(VSS),.VDD(VDD),.Y(g25675),.A(g24769),.B(g21832));
  OR2 OR2_841(.VSS(VSS),.VDD(VDD),.Y(g29243),.A(g28657),.B(g18358));
  OR2 OR2_842(.VSS(VSS),.VDD(VDD),.Y(g26348),.A(g8466),.B(g24609));
  OR2 OR2_843(.VSS(VSS),.VDD(VDD),.Y(g30501),.A(g29327),.B(g22018));
  OR2 OR2_844(.VSS(VSS),.VDD(VDD),.Y(g28061),.A(g27287),.B(g21735));
  OR2 OR2_845(.VSS(VSS),.VDD(VDD),.Y(g34729),.A(g34666),.B(g18270));
  OR2 OR2_846(.VSS(VSS),.VDD(VDD),.Y(g32408),.A(g31541),.B(g30073));
  OR2 OR2_847(.VSS(VSS),.VDD(VDD),.Y(g30439),.A(g29761),.B(g21848));
  OR2 OR2_848(.VSS(VSS),.VDD(VDD),.Y(g34728),.A(g34661),.B(g18214));
  OR2 OR2_849(.VSS(VSS),.VDD(VDD),.Y(g34439),.A(g34344),.B(g18181));
  OR2 OR2_850(.VSS(VSS),.VDD(VDD),.Y(g29269),.A(g28249),.B(g18634));
  OR2 OR2_851(.VSS(VSS),.VDD(VDD),.Y(g25637),.A(g24618),.B(g18307));
  OR2 OR2_852(.VSS(VSS),.VDD(VDD),.Y(g24233),.A(g22590),.B(g18236));
  OR2 OR2_853(.VSS(VSS),.VDD(VDD),.Y(g25935),.A(g24402),.B(g22208));
  OR2 OR2_854(.VSS(VSS),.VDD(VDD),.Y(g30438),.A(g29890),.B(g21847));
  OR2 OR2_855(.VSS(VSS),.VDD(VDD),.Y(g19525),.A(g7696),.B(g16811));
  OR2 OR2_856(.VSS(VSS),.VDD(VDD),.Y(g19488),.A(g16965),.B(g14148));
  OR2 OR2_857(.VSS(VSS),.VDD(VDD),.Y(g34438),.A(g34348),.B(g18150));
  OR2 OR2_858(.VSS(VSS),.VDD(VDD),.Y(g29268),.A(g28343),.B(g18625));
  OR4 OR4_29(.VSS(VSS),.VDD(VDD),.Y(I25613),.A(g25571),.B(g25572),.C(g25573),.D(g25574));
  OR2 OR2_859(.VSS(VSS),.VDD(VDD),.Y(g31884),.A(g31290),.B(g21778));
  OR2 OR2_860(.VSS(VSS),.VDD(VDD),.Y(g33791),.A(g33379),.B(g32430));
  OR2 OR2_861(.VSS(VSS),.VDD(VDD),.Y(g30349),.A(g30051),.B(g18333));
  OR2 OR2_862(.VSS(VSS),.VDD(VDD),.Y(g34349),.A(g26019),.B(g34104));
  OR3 OR3_25(.VSS(VSS),.VDD(VDD),.Y(g8417),.A(g1056),.B(g1116),.C(I12583));
  OR2 OR2_863(.VSS(VSS),.VDD(VDD),.Y(g30348),.A(g30083),.B(g18329));
  OR2 OR2_864(.VSS(VSS),.VDD(VDD),.Y(g22645),.A(g18982),.B(g15633));
  OR2 OR2_865(.VSS(VSS),.VDD(VDD),.Y(g34906),.A(g34857),.B(g21694));
  OR2 OR2_866(.VSS(VSS),.VDD(VDD),.Y(g29734),.A(g28201),.B(g15872));
  OR2 OR2_867(.VSS(VSS),.VDD(VDD),.Y(g30304),.A(g28255),.B(g27259));
  OR2 OR2_868(.VSS(VSS),.VDD(VDD),.Y(g33015),.A(g32343),.B(g18507));
  OR2 OR2_869(.VSS(VSS),.VDD(VDD),.Y(g34622),.A(g34520),.B(g18584));
  OR2 OR2_870(.VSS(VSS),.VDD(VDD),.Y(g25729),.A(g25091),.B(g22012));
  OR4 OR4_30(.VSS(VSS),.VDD(VDD),.Y(g26636),.A(g24897),.B(g24884),.C(g24858),.D(g24846));
  OR2 OR2_871(.VSS(VSS),.VDD(VDD),.Y(g28629),.A(g27371),.B(g16532));
  OR2 OR2_872(.VSS(VSS),.VDD(VDD),.Y(g25577),.A(g24143),.B(g24144));
  OR3 OR3_26(.VSS(VSS),.VDD(VDD),.Y(g28220),.A(g23495),.B(I26741),.C(I26742));
  OR2 OR2_873(.VSS(VSS),.VDD(VDD),.Y(g25728),.A(g25076),.B(g22011));
  OR2 OR2_874(.VSS(VSS),.VDD(VDD),.Y(g28628),.A(g27370),.B(g16531));
  OR2 OR2_875(.VSS(VSS),.VDD(VDD),.Y(g33556),.A(g33329),.B(g18362));
  OR2 OR2_876(.VSS(VSS),.VDD(VDD),.Y(g24212),.A(g23280),.B(g18155));
  OR2 OR2_877(.VSS(VSS),.VDD(VDD),.Y(g26963),.A(g26306),.B(g24308));
  OR2 OR2_878(.VSS(VSS),.VDD(VDD),.Y(g33580),.A(g33330),.B(g18442));
  OR2 OR2_879(.VSS(VSS),.VDD(VDD),.Y(g29487),.A(g25815),.B(g28133));
  OR2 OR2_880(.VSS(VSS),.VDD(VDD),.Y(g23795),.A(g20203),.B(g16884));
  OR2 OR2_881(.VSS(VSS),.VDD(VDD),.Y(g28071),.A(g27085),.B(g21873));
  OR2 OR2_882(.VSS(VSS),.VDD(VDD),.Y(g29502),.A(g28139),.B(g25871));
  OR2 OR2_883(.VSS(VSS),.VDD(VDD),.Y(g27533),.A(g26078),.B(g24659));
  OR4 OR4_31(.VSS(VSS),.VDD(VDD),.Y(I29351),.A(g29328),.B(g29323),.C(g29316),.D(g30316));
  OR2 OR2_884(.VSS(VSS),.VDD(VDD),.Y(g28591),.A(g27332),.B(g26286));
  OR2 OR2_885(.VSS(VSS),.VDD(VDD),.Y(g25906),.A(g25559),.B(g24014));
  OR2 OR2_886(.VSS(VSS),.VDD(VDD),.Y(g28776),.A(g27538),.B(g13974));
  OR2 OR2_887(.VSS(VSS),.VDD(VDD),.Y(g30415),.A(g29843),.B(g21799));
  OR2 OR2_888(.VSS(VSS),.VDD(VDD),.Y(g30333),.A(g29834),.B(g21699));
  OR2 OR2_889(.VSS(VSS),.VDD(VDD),.Y(g34636),.A(g34476),.B(g18693));
  OR2 OR2_890(.VSS(VSS),.VDD(VDD),.Y(g22547),.A(g16855),.B(g20215));
  OR2 OR2_891(.VSS(VSS),.VDD(VDD),.Y(g29279),.A(g28442),.B(g18741));
  OR2 OR2_892(.VSS(VSS),.VDD(VDD),.Y(g31922),.A(g31525),.B(g22047));
  OR2 OR2_893(.VSS(VSS),.VDD(VDD),.Y(g32982),.A(g31948),.B(g18208));
  OR2 OR2_894(.VSS(VSS),.VDD(VDD),.Y(g33321),.A(g29712),.B(g32182));
  OR2 OR2_895(.VSS(VSS),.VDD(VDD),.Y(g25622),.A(g24546),.B(g18217));
  OR2 OR2_896(.VSS(VSS),.VDD(VDD),.Y(g29278),.A(g28626),.B(g18740));
  OR2 OR2_897(.VSS(VSS),.VDD(VDD),.Y(g19267),.A(g17752),.B(g17768));
  OR2 OR2_898(.VSS(VSS),.VDD(VDD),.Y(g22226),.A(g21333),.B(g17655));
  OR2 OR2_899(.VSS(VSS),.VDD(VDD),.Y(g24433),.A(g10878),.B(g22400));
  OR2 OR2_900(.VSS(VSS),.VDD(VDD),.Y(g20148),.A(g16128),.B(g13393));
  OR2 OR2_901(.VSS(VSS),.VDD(VDD),.Y(g29286),.A(g28542),.B(g18759));
  OR2 OR2_902(.VSS(VSS),.VDD(VDD),.Y(g27232),.A(g25874),.B(g24450));
  OR2 OR2_903(.VSS(VSS),.VDD(VDD),.Y(g7404),.A(g933),.B(g939));
  OR2 OR2_904(.VSS(VSS),.VDD(VDD),.Y(g29306),.A(g28689),.B(g18813));
  OR4 OR4_32(.VSS(VSS),.VDD(VDD),.Y(g28172),.A(g27469),.B(g27440),.C(g27416),.D(g27395));
  OR2 OR2_905(.VSS(VSS),.VDD(VDD),.Y(g33685),.A(g32396),.B(g33423));
  OR2 OR2_906(.VSS(VSS),.VDD(VDD),.Y(g7764),.A(g2999),.B(g2932));
  OR3 OR3_27(.VSS(VSS),.VDD(VDD),.Y(g33953),.A(g33487),.B(I31848),.C(I31849));
  OR2 OR2_907(.VSS(VSS),.VDD(VDD),.Y(g24343),.A(g23724),.B(g18773));
  OR2 OR2_908(.VSS(VSS),.VDD(VDD),.Y(g26921),.A(g25955),.B(g18285));
  OR2 OR2_909(.VSS(VSS),.VDD(VDD),.Y(g25653),.A(g24664),.B(g18602));
  OR2 OR2_910(.VSS(VSS),.VDD(VDD),.Y(g32390),.A(g31501),.B(g29979));
  OR2 OR2_911(.VSS(VSS),.VDD(VDD),.Y(g27261),.A(g24544),.B(g25996));
  OR2 OR2_912(.VSS(VSS),.VDD(VDD),.Y(g30484),.A(g30154),.B(g21980));
  OR2 OR2_913(.VSS(VSS),.VDD(VDD),.Y(g30554),.A(g30216),.B(g22125));
  OR2 OR2_914(.VSS(VSS),.VDD(VDD),.Y(g22490),.A(g21513),.B(g12795));
  OR3 OR3_28(.VSS(VSS),.VDD(VDD),.Y(g13820),.A(g11184),.B(g9187),.C(g12527));
  OR2 OR2_915(.VSS(VSS),.VDD(VDD),.Y(g26813),.A(g24940),.B(g24949));
  OR4 OR4_33(.VSS(VSS),.VDD(VDD),.Y(g15727),.A(g13383),.B(g13345),.C(g13333),.D(g11010));
  OR2 OR2_916(.VSS(VSS),.VDD(VDD),.Y(g25636),.A(g24507),.B(g18305));
  OR2 OR2_917(.VSS(VSS),.VDD(VDD),.Y(g30609),.A(g13633),.B(g29742));
  OR2 OR2_918(.VSS(VSS),.VDD(VDD),.Y(g34609),.A(g34503),.B(g18563));
  OR2 OR2_919(.VSS(VSS),.VDD(VDD),.Y(g28420),.A(g27222),.B(g13290));
  OR2 OR2_920(.VSS(VSS),.VDD(VDD),.Y(g30608),.A(g13604),.B(g29736));
  OR2 OR2_921(.VSS(VSS),.VDD(VDD),.Y(g28319),.A(g27115),.B(g15807));
  OR2 OR2_922(.VSS(VSS),.VDD(VDD),.Y(g30115),.A(g28489),.B(g11449));
  OR2 OR2_923(.VSS(VSS),.VDD(VDD),.Y(g29143),.A(g27650),.B(g17146));
  OR2 OR2_924(.VSS(VSS),.VDD(VDD),.Y(g34608),.A(g34568),.B(g15082));
  OR4 OR4_34(.VSS(VSS),.VDD(VDD),.Y(g17490),.A(g14364),.B(g14337),.C(g11958),.D(I18421));
  OR2 OR2_925(.VSS(VSS),.VDD(VDD),.Y(g26805),.A(g10776),.B(g24478));
  OR2 OR2_926(.VSS(VSS),.VDD(VDD),.Y(g31762),.A(g30011),.B(g30030));
  OR2 OR2_927(.VSS(VSS),.VDD(VDD),.Y(g23358),.A(g19746),.B(g16212));
  OR4 OR4_35(.VSS(VSS),.VDD(VDD),.Y(I30760),.A(g31778),.B(g32295),.C(g32046),.D(g32050));
  OR2 OR2_928(.VSS(VSS),.VDD(VDD),.Y(g31964),.A(g31654),.B(g14544));
  OR2 OR2_929(.VSS(VSS),.VDD(VDD),.Y(g33964),.A(g33817),.B(g18146));
  OR2 OR2_930(.VSS(VSS),.VDD(VDD),.Y(g25664),.A(g24681),.B(g21789));
  OR2 OR2_931(.VSS(VSS),.VDD(VDD),.Y(g28059),.A(g27042),.B(g18276));
  OR2 OR2_932(.VSS(VSS),.VDD(VDD),.Y(g29791),.A(g28233),.B(g22859));
  OR2 OR2_933(.VSS(VSS),.VDD(VDD),.Y(g16021),.A(g13047),.B(g10706));
  OR2 OR2_934(.VSS(VSS),.VDD(VDD),.Y(g26934),.A(g26845),.B(g18556));
  OR2 OR2_935(.VSS(VSS),.VDD(VDD),.Y(g28058),.A(g27235),.B(g18268));
  OR2 OR2_936(.VSS(VSS),.VDD(VDD),.Y(g29168),.A(g27658),.B(g26613));
  OR2 OR2_937(.VSS(VSS),.VDD(VDD),.Y(g33587),.A(g33363),.B(g18463));
  OR2 OR2_938(.VSS(VSS),.VDD(VDD),.Y(g24896),.A(g22863),.B(g19684));
  OR2 OR2_939(.VSS(VSS),.VDD(VDD),.Y(g34799),.A(g34751),.B(g18578));
  OR2 OR2_940(.VSS(VSS),.VDD(VDD),.Y(g25585),.A(g21674),.B(g24155));
  OR2 OR2_941(.VSS(VSS),.VDD(VDD),.Y(g25576),.A(g24141),.B(g24142));
  OR2 OR2_942(.VSS(VSS),.VDD(VDD),.Y(g29479),.A(g28113),.B(g28116));
  OR2 OR2_943(.VSS(VSS),.VDD(VDD),.Y(g34798),.A(g34754),.B(g18575));
  OR2 OR2_944(.VSS(VSS),.VDD(VDD),.Y(g31909),.A(g31750),.B(g21956));
  OR2 OR2_945(.VSS(VSS),.VDD(VDD),.Y(g28044),.A(g27256),.B(g18130));
  OR2 OR2_946(.VSS(VSS),.VDD(VDD),.Y(g33543),.A(g33106),.B(g18281));
  OR2 OR2_947(.VSS(VSS),.VDD(VDD),.Y(g19595),.A(g17149),.B(g14218));
  OR2 OR2_948(.VSS(VSS),.VDD(VDD),.Y(g29478),.A(g28111),.B(g22160));
  OR2 OR2_949(.VSS(VSS),.VDD(VDD),.Y(g19467),.A(g16896),.B(g14097));
  OR2 OR2_950(.VSS(VSS),.VDD(VDD),.Y(g25609),.A(g24915),.B(g18126));
  OR2 OR2_951(.VSS(VSS),.VDD(VDD),.Y(g34805),.A(g34748),.B(g18594));
  OR2 OR2_952(.VSS(VSS),.VDD(VDD),.Y(g31908),.A(g31519),.B(g21955));
  OR2 OR2_953(.VSS(VSS),.VDD(VDD),.Y(g33000),.A(g32270),.B(g18403));
  OR2 OR2_954(.VSS(VSS),.VDD(VDD),.Y(g29486),.A(g28537),.B(g27595));
  OR2 OR2_955(.VSS(VSS),.VDD(VDD),.Y(g32252),.A(g31183),.B(g31206));
  OR2 OR2_956(.VSS(VSS),.VDD(VDD),.Y(g25608),.A(g24643),.B(g18120));
  OR2 OR2_957(.VSS(VSS),.VDD(VDD),.Y(g33569),.A(g33415),.B(g18402));
  OR2 OR2_958(.VSS(VSS),.VDD(VDD),.Y(g30732),.A(g13778),.B(g29762));
  OR2 OR2_959(.VSS(VSS),.VDD(VDD),.Y(g27271),.A(g24547),.B(g26053));
  OR3 OR3_29(.VSS(VSS),.VDD(VDD),.Y(I18495),.A(g14539),.B(g14515),.C(g14449));
  OR2 OR2_960(.VSS(VSS),.VDD(VDD),.Y(g34732),.A(g34686),.B(g18593));
  OR2 OR2_961(.VSS(VSS),.VDD(VDD),.Y(g26329),.A(g8526),.B(g24609));
  OR2 OR2_962(.VSS(VSS),.VDD(VDD),.Y(g33568),.A(g33409),.B(g18395));
  OR2 OR2_963(.VSS(VSS),.VDD(VDD),.Y(g25745),.A(g25150),.B(g22060));
  OR2 OR2_964(.VSS(VSS),.VDD(VDD),.Y(g29223),.A(g28341),.B(g18131));
  OR2 OR2_965(.VSS(VSS),.VDD(VDD),.Y(g26328),.A(g1183),.B(g24591));
  OR2 OR2_966(.VSS(VSS),.VDD(VDD),.Y(g28562),.A(g27313),.B(g26251));
  OR2 OR2_967(.VSS(VSS),.VDD(VDD),.Y(g14844),.A(g10776),.B(g8703));
  OR2 OR2_968(.VSS(VSS),.VDD(VDD),.Y(g34761),.A(g34679),.B(g34506));
  OR2 OR2_969(.VSS(VSS),.VDD(VDD),.Y(g28699),.A(g27452),.B(g16667));
  OR4 OR4_36(.VSS(VSS),.VDD(VDD),.Y(g27031),.A(g26213),.B(g26190),.C(g26166),.D(g26148));
  OR2 OR2_970(.VSS(VSS),.VDD(VDD),.Y(g33123),.A(g31962),.B(g30577));
  OR4 OR4_37(.VSS(VSS),.VDD(VDD),.Y(I30755),.A(g30564),.B(g32303),.C(g32049),.D(g32055));
  OR2 OR2_971(.VSS(VSS),.VDD(VDD),.Y(g28698),.A(g27451),.B(g16666));
  OR2 OR2_972(.VSS(VSS),.VDD(VDD),.Y(g31751),.A(g29975),.B(g29990));
  OR2 OR2_973(.VSS(VSS),.VDD(VDD),.Y(g31772),.A(g30035),.B(g28654));
  OR2 OR2_974(.VSS(VSS),.VDD(VDD),.Y(g30400),.A(g29766),.B(g21759));
  OR2 OR2_975(.VSS(VSS),.VDD(VDD),.Y(g33974),.A(g33846),.B(g18345));
  OR2 OR2_976(.VSS(VSS),.VDD(VDD),.Y(g30214),.A(g23424),.B(g28572));
  OR2 OR2_977(.VSS(VSS),.VDD(VDD),.Y(g34013),.A(g33901),.B(g18488));
  OR4 OR4_38(.VSS(VSS),.VDD(VDD),.Y(g25805),.A(g25453),.B(g25414),.C(g25374),.D(g25331));
  OR2 OR2_978(.VSS(VSS),.VDD(VDD),.Y(g25674),.A(g24755),.B(g21831));
  OR2 OR2_979(.VSS(VSS),.VDD(VDD),.Y(g31293),.A(g29582),.B(g28299));
  OR2 OR2_980(.VSS(VSS),.VDD(VDD),.Y(g33293),.A(g32151),.B(g29602));
  OR2 OR2_981(.VSS(VSS),.VDD(VDD),.Y(g30539),.A(g30267),.B(g22085));
  OR2 OR2_982(.VSS(VSS),.VDD(VDD),.Y(g34207),.A(g33835),.B(g33304));
  OR2 OR2_983(.VSS(VSS),.VDD(VDD),.Y(g22659),.A(g19062),.B(g15673));
  OR2 OR2_984(.VSS(VSS),.VDD(VDD),.Y(g22625),.A(g18910),.B(g18933));
  OR2 OR2_985(.VSS(VSS),.VDD(VDD),.Y(g25732),.A(g25201),.B(g22017));
  OR2 OR2_986(.VSS(VSS),.VDD(VDD),.Y(g34005),.A(g33883),.B(g18454));
  OR2 OR2_987(.VSS(VSS),.VDD(VDD),.Y(g28632),.A(g27373),.B(g16535));
  OR2 OR2_988(.VSS(VSS),.VDD(VDD),.Y(g33265),.A(g32113),.B(g29530));
  OR2 OR2_989(.VSS(VSS),.VDD(VDD),.Y(g30538),.A(g30256),.B(g22084));
  OR2 OR2_990(.VSS(VSS),.VDD(VDD),.Y(g29373),.A(g13832),.B(g28453));
  OR4 OR4_39(.VSS(VSS),.VDD(VDD),.Y(I30262),.A(g31672),.B(g31710),.C(g31021),.D(g30937));
  OR2 OR2_991(.VSS(VSS),.VDD(VDD),.Y(g33992),.A(g33900),.B(g18408));
  OR2 OR2_992(.VSS(VSS),.VDD(VDD),.Y(g25761),.A(g25152),.B(g18812));
  OR2 OR2_993(.VSS(VSS),.VDD(VDD),.Y(g28661),.A(g27406),.B(g16611));
  OR2 OR2_994(.VSS(VSS),.VDD(VDD),.Y(g28403),.A(g27214),.B(g13282));
  OR2 OR2_995(.VSS(VSS),.VDD(VDD),.Y(g22644),.A(g18981),.B(g15632));
  OR4 OR4_40(.VSS(VSS),.VDD(VDD),.Y(I12782),.A(g4188),.B(g4194),.C(g4197),.D(g4200));
  OR2 OR2_996(.VSS(VSS),.VDD(VDD),.Y(g33579),.A(g33357),.B(g18437));
  OR2 OR2_997(.VSS(VSS),.VDD(VDD),.Y(g14044),.A(g10776),.B(g8703));
  OR2 OR2_998(.VSS(VSS),.VDD(VDD),.Y(g28715),.A(g27480),.B(g16700));
  OR4 OR4_41(.VSS(VSS),.VDD(VDD),.Y(I30718),.A(g32348),.B(g32356),.C(g32097),.D(g32020));
  OR2 OR2_999(.VSS(VSS),.VDD(VDD),.Y(g33578),.A(g33410),.B(g18433));
  OR2 OR2_1000(.VSS(VSS),.VDD(VDD),.Y(g31014),.A(g29367),.B(g28160));
  OR2 OR2_1001(.VSS(VSS),.VDD(VDD),.Y(g27225),.A(g2975),.B(g26364));
  OR2 OR2_1002(.VSS(VSS),.VDD(VDD),.Y(g33014),.A(g32305),.B(g18499));
  OR2 OR2_1003(.VSS(VSS),.VDD(VDD),.Y(g23770),.A(g20188),.B(g16868));
  OR2 OR2_1004(.VSS(VSS),.VDD(VDD),.Y(g26882),.A(g26650),.B(g24188));
  OR2 OR2_1005(.VSS(VSS),.VDD(VDD),.Y(g28551),.A(g27305),.B(g26234));
  OR2 OR2_1006(.VSS(VSS),.VDD(VDD),.Y(g31007),.A(g29364),.B(g28159));
  OR2 OR2_1007(.VSS(VSS),.VDD(VDD),.Y(g27258),.A(g25905),.B(g15749));
  OR2 OR2_1008(.VSS(VSS),.VDD(VDD),.Y(g34100),.A(g33690),.B(g33697));
  OR2 OR2_1009(.VSS(VSS),.VDD(VDD),.Y(g33586),.A(g33416),.B(g18459));
  OR2 OR2_1010(.VSS(VSS),.VDD(VDD),.Y(g33007),.A(g32331),.B(g18455));
  OR2 OR2_1011(.VSS(VSS),.VDD(VDD),.Y(g25539),.A(g23531),.B(g20628));
  OR2 OR2_1012(.VSS(VSS),.VDD(VDD),.Y(g13662),.A(g10896),.B(g10917));
  OR2 OR2_1013(.VSS(VSS),.VDD(VDD),.Y(g34235),.A(g32585),.B(g33953));
  OR2 OR2_1014(.VSS(VSS),.VDD(VDD),.Y(g27244),.A(g24652),.B(g25995));
  OR2 OR2_1015(.VSS(VSS),.VDD(VDD),.Y(g28490),.A(g27262),.B(g16185));
  OR2 OR2_1016(.VSS(VSS),.VDD(VDD),.Y(g33116),.A(g32403),.B(g32411));
  OR2 OR2_1017(.VSS(VSS),.VDD(VDD),.Y(g33615),.A(g33113),.B(g21871));
  OR2 OR2_1018(.VSS(VSS),.VDD(VDD),.Y(g23262),.A(g19661),.B(g16126));
  OR2 OR2_1019(.VSS(VSS),.VDD(VDD),.Y(g21899),.A(g20162),.B(g15113));
  OR2 OR2_1020(.VSS(VSS),.VDD(VDD),.Y(g30515),.A(g30223),.B(g22036));
  OR2 OR2_1021(.VSS(VSS),.VDD(VDD),.Y(g30414),.A(g30002),.B(g21794));
  OR2 OR2_1022(.VSS(VSS),.VDD(VDD),.Y(g28385),.A(g27201),.B(g15857));
  OR2 OR2_1023(.VSS(VSS),.VDD(VDD),.Y(g33041),.A(g32189),.B(g24323));
  OR2 OR2_1024(.VSS(VSS),.VDD(VDD),.Y(g28297),.A(g27096),.B(g15785));
  OR2 OR2_1025(.VSS(VSS),.VDD(VDD),.Y(g21898),.A(g20152),.B(g15112));
  OR2 OR2_1026(.VSS(VSS),.VDD(VDD),.Y(g34882),.A(g34876),.B(g18659));
  OR2 OR2_1027(.VSS(VSS),.VDD(VDD),.Y(g28103),.A(g27696),.B(g22097));
  OR2 OR2_1028(.VSS(VSS),.VDD(VDD),.Y(g24245),.A(g22849),.B(g18256));
  OR2 OR2_1029(.VSS(VSS),.VDD(VDD),.Y(g33275),.A(g32127),.B(g29564));
  OR2 OR2_1030(.VSS(VSS),.VDD(VDD),.Y(g28095),.A(g27674),.B(g21970));
  OR2 OR2_1031(.VSS(VSS),.VDD(VDD),.Y(g30407),.A(g29794),.B(g21766));
  OR2 OR2_1032(.VSS(VSS),.VDD(VDD),.Y(g34407),.A(g34185),.B(g25124));
  OR2 OR2_1033(.VSS(VSS),.VDD(VDD),.Y(g27970),.A(g26514),.B(g25050));
  OR2 OR2_1034(.VSS(VSS),.VDD(VDD),.Y(g31465),.A(g26156),.B(g29647));
  OR2 OR2_1035(.VSS(VSS),.VDD(VDD),.Y(g26759),.A(g24468),.B(g7511));
  OR2 OR2_1036(.VSS(VSS),.VDD(VDD),.Y(g26725),.A(g24457),.B(g10719));
  OR2 OR2_1037(.VSS(VSS),.VDD(VDD),.Y(g28671),.A(g27413),.B(g16619));
  OR2 OR2_1038(.VSS(VSS),.VDD(VDD),.Y(g33983),.A(g33877),.B(g18373));
  OR2 OR2_1039(.VSS(VSS),.VDD(VDD),.Y(g22707),.A(g20559),.B(g17156));
  OR2 OR2_1040(.VSS(VSS),.VDD(VDD),.Y(g33035),.A(g32019),.B(g21872));
  OR2 OR2_1041(.VSS(VSS),.VDD(VDD),.Y(g27886),.A(g14438),.B(g26759));
  OR2 OR2_1042(.VSS(VSS),.VDD(VDD),.Y(g25683),.A(g24669),.B(g18641));
  OR2 OR2_1043(.VSS(VSS),.VDD(VDD),.Y(g29242),.A(g28674),.B(g18354));
  OR2 OR2_1044(.VSS(VSS),.VDD(VDD),.Y(g26082),.A(g2898),.B(g24561));
  OR2 OR2_1045(.VSS(VSS),.VDD(VDD),.Y(g11380),.A(g8583),.B(g8530));
  OR2 OR2_1046(.VSS(VSS),.VDD(VDD),.Y(g30441),.A(g29787),.B(g21850));
  OR2 OR2_1047(.VSS(VSS),.VDD(VDD),.Y(g34441),.A(g34381),.B(g18540));
  OR2 OR2_1048(.VSS(VSS),.VDD(VDD),.Y(g24232),.A(g22686),.B(g18228));
  OR2 OR2_1049(.VSS(VSS),.VDD(VDD),.Y(g34206),.A(g33834),.B(g33836));
  OR2 OR2_1050(.VSS(VSS),.VDD(VDD),.Y(g26940),.A(g25908),.B(g21886));
  OR4 OR4_42(.VSS(VSS),.VDD(VDD),.Y(I25612),.A(g25567),.B(g25568),.C(g25569),.D(g25570));
  OR2 OR2_1051(.VSS(VSS),.VDD(VDD),.Y(g34725),.A(g34700),.B(g18183));
  OR2 OR2_1052(.VSS(VSS),.VDD(VDD),.Y(g24261),.A(g22862),.B(g18314));
  OR2 OR2_1053(.VSS(VSS),.VDD(VDD),.Y(g29230),.A(g28107),.B(g18202));
  OR2 OR2_1054(.VSS(VSS),.VDD(VDD),.Y(g27458),.A(g24590),.B(g25989));
  OR2 OR2_1055(.VSS(VSS),.VDD(VDD),.Y(g29293),.A(g28570),.B(g18777));
  OR2 OR2_1056(.VSS(VSS),.VDD(VDD),.Y(g30114),.A(g28488),.B(g16761));
  OR2 OR2_1057(.VSS(VSS),.VDD(VDD),.Y(g30435),.A(g30025),.B(g21840));
  OR2 OR2_1058(.VSS(VSS),.VDD(VDD),.Y(g29265),.A(g28318),.B(g18620));
  OR2 OR2_1059(.VSS(VSS),.VDD(VDD),.Y(g28546),.A(g27302),.B(g26231));
  OR2 OR2_1060(.VSS(VSS),.VDD(VDD),.Y(g28089),.A(g27269),.B(g18731));
  OR2 OR2_1061(.VSS(VSS),.VDD(VDD),.Y(g23251),.A(g19637),.B(g16098));
  OR2 OR2_1062(.VSS(VSS),.VDD(VDD),.Y(g28211),.A(g27029),.B(g27034));
  OR2 OR2_1063(.VSS(VSS),.VDD(VDD),.Y(g34107),.A(g33710),.B(g33121));
  OR2 OR2_1064(.VSS(VSS),.VDD(VDD),.Y(g19555),.A(g15672),.B(g13030));
  OR2 OR2_1065(.VSS(VSS),.VDD(VDD),.Y(g28088),.A(g27264),.B(g18729));
  OR2 OR2_1066(.VSS(VSS),.VDD(VDD),.Y(g30345),.A(g29644),.B(g18302));
  OR2 OR2_1067(.VSS(VSS),.VDD(VDD),.Y(g30399),.A(g29757),.B(g21758));
  OR2 OR2_1068(.VSS(VSS),.VDD(VDD),.Y(g34849),.A(g34842),.B(g18154));
  OR2 OR2_1069(.VSS(VSS),.VDD(VDD),.Y(g34399),.A(g34178),.B(g25067));
  OR2 OR2_1070(.VSS(VSS),.VDD(VDD),.Y(g25584),.A(g21670),.B(g24154));
  OR2 OR2_1071(.VSS(VSS),.VDD(VDD),.Y(g28497),.A(g27267),.B(g16199));
  OR2 OR2_1072(.VSS(VSS),.VDD(VDD),.Y(g33006),.A(g32291),.B(g18447));
  OR2 OR2_1073(.VSS(VSS),.VDD(VDD),.Y(g30398),.A(g29749),.B(g21757));
  OR2 OR2_1074(.VSS(VSS),.VDD(VDD),.Y(g26962),.A(g26295),.B(g24307));
  OR2 OR2_1075(.VSS(VSS),.VDD(VDD),.Y(g26361),.A(g24674),.B(g22991));
  OR2 OR2_1076(.VSS(VSS),.VDD(VDD),.Y(g23997),.A(g20602),.B(g17191));
  OR2 OR2_1077(.VSS(VSS),.VDD(VDD),.Y(g30141),.A(g28499),.B(g16844));
  OR2 OR2_1078(.VSS(VSS),.VDD(VDD),.Y(g34804),.A(g34740),.B(g18591));
  OR2 OR2_1079(.VSS(VSS),.VDD(VDD),.Y(g28700),.A(g27454),.B(g16668));
  OR2 OR2_1080(.VSS(VSS),.VDD(VDD),.Y(g25759),.A(g25166),.B(g22106));
  OR2 OR2_1081(.VSS(VSS),.VDD(VDD),.Y(g28659),.A(g27404),.B(g16610));
  OR2 OR2_1082(.VSS(VSS),.VDD(VDD),.Y(g25725),.A(g25127),.B(g22008));
  OR2 OR2_1083(.VSS(VSS),.VDD(VDD),.Y(g28625),.A(g27363),.B(g26324));
  OR2 OR2_1084(.VSS(VSS),.VDD(VDD),.Y(g14888),.A(g10776),.B(g8703));
  OR2 OR2_1085(.VSS(VSS),.VDD(VDD),.Y(g32357),.A(g29865),.B(g31296));
  OR2 OR2_1086(.VSS(VSS),.VDD(VDD),.Y(g27159),.A(g25814),.B(g12953));
  OR2 OR2_1087(.VSS(VSS),.VDD(VDD),.Y(g27532),.A(g16176),.B(g26084));
  OR2 OR2_1088(.VSS(VSS),.VDD(VDD),.Y(g25758),.A(g25151),.B(g22105));
  OR2 OR2_1089(.VSS(VSS),.VDD(VDD),.Y(g34263),.A(g34078),.B(g18699));
  OR2 OR2_1090(.VSS(VSS),.VDD(VDD),.Y(g34332),.A(g34071),.B(g33723));
  OR2 OR2_1091(.VSS(VSS),.VDD(VDD),.Y(g33703),.A(g32410),.B(g33434));
  OR2 OR2_1092(.VSS(VSS),.VDD(VDD),.Y(g28296),.A(g27095),.B(g15784));
  OR2 OR2_1093(.VSS(VSS),.VDD(VDD),.Y(g31253),.A(g25980),.B(g29533));
  OR2 OR2_1094(.VSS(VSS),.VDD(VDD),.Y(g27561),.A(g26100),.B(g24702));
  OR2 OR2_1095(.VSS(VSS),.VDD(VDD),.Y(g33253),.A(g32103),.B(g29511));
  OR2 OR2_1096(.VSS(VSS),.VDD(VDD),.Y(g25744),.A(g25129),.B(g22059));
  OR2 OR2_1097(.VSS(VSS),.VDD(VDD),.Y(g28644),.A(g27387),.B(g16593));
  OR2 OR2_1098(.VSS(VSS),.VDD(VDD),.Y(g30406),.A(g29783),.B(g21765));
  OR2 OR2_1099(.VSS(VSS),.VDD(VDD),.Y(g24432),.A(g23900),.B(g21361));
  OR2 OR2_1100(.VSS(VSS),.VDD(VDD),.Y(g30361),.A(g30109),.B(g18391));
  OR2 OR2_1101(.VSS(VSS),.VDD(VDD),.Y(g34406),.A(g34184),.B(g25123));
  OR2 OR2_1102(.VSS(VSS),.VDD(VDD),.Y(g24271),.A(g23451),.B(g18628));
  OR2 OR2_1103(.VSS(VSS),.VDD(VDD),.Y(g33600),.A(g33418),.B(g18501));
  OR2 OR2_1104(.VSS(VSS),.VDD(VDD),.Y(g25940),.A(g24415),.B(g22218));
  OR2 OR2_1105(.VSS(VSS),.VDD(VDD),.Y(g31781),.A(g30058),.B(g30069));
  OR3 OR3_30(.VSS(VSS),.VDD(VDD),.Y(g23162),.A(g20184),.B(g20170),.C(I22267));
  OR2 OR2_1106(.VSS(VSS),.VDD(VDD),.Y(g33236),.A(g32044),.B(g32045));
  OR2 OR2_1107(.VSS(VSS),.VDD(VDD),.Y(g30500),.A(g29326),.B(g21996));
  OR2 OR2_1108(.VSS(VSS),.VDD(VDD),.Y(g29275),.A(g28165),.B(g21868));
  OR2 OR2_1109(.VSS(VSS),.VDD(VDD),.Y(g28060),.A(g27616),.B(g18532));
  OR3 OR3_31(.VSS(VSS),.VDD(VDD),.Y(g33952),.A(g33478),.B(I31843),.C(I31844));
  OR2 OR2_1110(.VSS(VSS),.VDD(VDD),.Y(g24342),.A(g23691),.B(g18772));
  OR2 OR2_1111(.VSS(VSS),.VDD(VDD),.Y(g25652),.A(g24777),.B(g21747));
  OR2 OR2_1112(.VSS(VSS),.VDD(VDD),.Y(g26947),.A(g26394),.B(g24285));
  OR2 OR2_1113(.VSS(VSS),.VDD(VDD),.Y(g8905),.A(g2204),.B(g2223));
  OR2 OR2_1114(.VSS(VSS),.VDD(VDD),.Y(g29237),.A(g28185),.B(g18289));
  OR2 OR2_1115(.VSS(VSS),.VDD(VDD),.Y(g28527),.A(g27286),.B(g26182));
  OR2 OR2_1116(.VSS(VSS),.VDD(VDD),.Y(g33063),.A(g31988),.B(g22066));
  OR2 OR2_1117(.VSS(VSS),.VDD(VDD),.Y(g34004),.A(g33879),.B(g18453));
  OR2 OR2_1118(.VSS(VSS),.VDD(VDD),.Y(g26951),.A(g26390),.B(g24289));
  OR2 OR2_1119(.VSS(VSS),.VDD(VDD),.Y(g26972),.A(g26780),.B(g25229));
  OR2 OR2_1120(.VSS(VSS),.VDD(VDD),.Y(g31873),.A(g31270),.B(g21728));
  OR2 OR2_1121(.VSS(VSS),.VDD(VDD),.Y(g19501),.A(g16986),.B(g14168));
  OR2 OR2_1122(.VSS(VSS),.VDD(VDD),.Y(g34613),.A(g34515),.B(g18567));
  OR2 OR2_1123(.VSS(VSS),.VDD(VDD),.Y(g32249),.A(g31169),.B(g29687));
  OR2 OR2_1124(.VSS(VSS),.VDD(VDD),.Y(g30605),.A(g29529),.B(g29520));
  OR2 OR2_1125(.VSS(VSS),.VDD(VDD),.Y(g27289),.A(g25925),.B(g25927));
  OR2 OR2_1126(.VSS(VSS),.VDD(VDD),.Y(g34273),.A(g27765),.B(g34203));
  OR2 OR2_1127(.VSS(VSS),.VDD(VDD),.Y(g34605),.A(g34566),.B(g15077));
  OR2 OR2_1128(.VSS(VSS),.VDD(VDD),.Y(g18879),.A(g17365),.B(g14423));
  OR2 OR2_1129(.VSS(VSS),.VDD(VDD),.Y(g28581),.A(g27329),.B(g26276));
  OR2 OR2_1130(.VSS(VSS),.VDD(VDD),.Y(g27224),.A(g25870),.B(g15678));
  OR2 OR2_1131(.VSS(VSS),.VDD(VDD),.Y(g30463),.A(g30140),.B(g21934));
  OR2 OR2_1132(.VSS(VSS),.VDD(VDD),.Y(g27571),.A(g26127),.B(g24723));
  OR2 OR2_1133(.VSS(VSS),.VDD(VDD),.Y(g28707),.A(g27461),.B(g16673));
  OR2 OR2_1134(.VSS(VSS),.VDD(VDD),.Y(g34463),.A(g34338),.B(g18686));
  OR2 OR2_1135(.VSS(VSS),.VDD(VDD),.Y(g23825),.A(g20705),.B(g20781));
  OR2 OR2_1136(.VSS(VSS),.VDD(VDD),.Y(g30371),.A(g30099),.B(g18445));
  OR2 OR2_1137(.VSS(VSS),.VDD(VDD),.Y(g28818),.A(g27549),.B(g13998));
  OR2 OR2_1138(.VSS(VSS),.VDD(VDD),.Y(g34033),.A(g33821),.B(g18708));
  OR2 OR2_1139(.VSS(VSS),.VDD(VDD),.Y(g34234),.A(g32520),.B(g33952));
  OR2 OR2_1140(.VSS(VSS),.VDD(VDD),.Y(g28055),.A(g27560),.B(g18190));
  OR2 OR2_1141(.VSS(VSS),.VDD(VDD),.Y(g33542),.A(g33102),.B(g18265));
  OR2 OR2_1142(.VSS(VSS),.VDD(VDD),.Y(g33021),.A(g32302),.B(g21749));
  OR2 OR2_1143(.VSS(VSS),.VDD(VDD),.Y(g24259),.A(g23008),.B(g18312));
  OR2 OR2_1144(.VSS(VSS),.VDD(VDD),.Y(g28070),.A(g27050),.B(g21867));
  OR2 OR2_1145(.VSS(VSS),.VDD(VDD),.Y(g31913),.A(g31485),.B(g21999));
  OR2 OR2_1146(.VSS(VSS),.VDD(VDD),.Y(g18994),.A(g16303),.B(g13632));
  OR2 OR2_1147(.VSS(VSS),.VDD(VDD),.Y(g24471),.A(g10999),.B(g22450));
  OR2 OR2_1148(.VSS(VSS),.VDD(VDD),.Y(g34795),.A(g34753),.B(g18572));
  OR2 OR2_1149(.VSS(VSS),.VDD(VDD),.Y(g25613),.A(g25181),.B(g18140));
  OR2 OR2_1150(.VSS(VSS),.VDD(VDD),.Y(g24258),.A(g22851),.B(g18311));
  OR2 OR2_1151(.VSS(VSS),.VDD(VDD),.Y(g33614),.A(g33249),.B(g18650));
  OR4 OR4_43(.VSS(VSS),.VDD(VDD),.Y(g17511),.A(g14396),.B(g14365),.C(g11976),.D(I18452));
  OR2 OR2_1152(.VSS(VSS),.VDD(VDD),.Y(g32999),.A(g32337),.B(g18401));
  OR2 OR2_1153(.VSS(VSS),.VDD(VDD),.Y(g33607),.A(g33091),.B(g18526));
  OR2 OR2_1154(.VSS(VSS),.VDD(VDD),.Y(g31905),.A(g31746),.B(g21952));
  OR2 OR2_1155(.VSS(VSS),.VDD(VDD),.Y(g31320),.A(g26125),.B(g29632));
  OR2 OR2_1156(.VSS(VSS),.VDD(VDD),.Y(g30514),.A(g30211),.B(g22035));
  OR2 OR2_1157(.VSS(VSS),.VDD(VDD),.Y(g32380),.A(g29907),.B(g31467));
  OR2 OR2_1158(.VSS(VSS),.VDD(VDD),.Y(g31274),.A(g29565),.B(g28280));
  OR2 OR2_1159(.VSS(VSS),.VDD(VDD),.Y(g25605),.A(g24743),.B(g18116));
  OR2 OR2_1160(.VSS(VSS),.VDD(VDD),.Y(g29222),.A(g28252),.B(g18105));
  OR2 OR2_1161(.VSS(VSS),.VDD(VDD),.Y(g24244),.A(g23349),.B(g18255));
  OR2 OR2_1162(.VSS(VSS),.VDD(VDD),.Y(g33274),.A(g32126),.B(g29563));
  OR2 OR2_1163(.VSS(VSS),.VDD(VDD),.Y(g30507),.A(g30190),.B(g22028));
  OR2 OR2_1164(.VSS(VSS),.VDD(VDD),.Y(g32998),.A(g32300),.B(g18393));
  OR2 OR2_1165(.VSS(VSS),.VDD(VDD),.Y(g28094),.A(g27673),.B(g21959));
  OR2 OR2_1166(.VSS(VSS),.VDD(VDD),.Y(g28067),.A(g27309),.B(g21827));
  OR2 OR2_1167(.VSS(VSS),.VDD(VDD),.Y(g33593),.A(g33417),.B(g18482));
  OR2 OR2_1168(.VSS(VSS),.VDD(VDD),.Y(g26789),.A(g10776),.B(g24471));
  OR2 OR2_1169(.VSS(VSS),.VDD(VDD),.Y(g32233),.A(g31150),.B(g29661));
  OR2 OR2_1170(.VSS(VSS),.VDD(VDD),.Y(g12954),.A(g12186),.B(g9906));
  OR2 OR2_1171(.VSS(VSS),.VDD(VDD),.Y(g23319),.A(g19717),.B(g16193));
  OR2 OR2_1172(.VSS(VSS),.VDD(VDD),.Y(g30421),.A(g29784),.B(g21805));
  OR2 OR2_1173(.VSS(VSS),.VDD(VDD),.Y(g33565),.A(g33338),.B(g18389));
  OR2 OR2_1174(.VSS(VSS),.VDD(VDD),.Y(g34421),.A(g27686),.B(g34198));
  OR2 OR2_1175(.VSS(VSS),.VDD(VDD),.Y(g26359),.A(g24651),.B(g22939));
  OR2 OR2_1176(.VSS(VSS),.VDD(VDD),.Y(g28735),.A(g27510),.B(g16737));
  OR2 OR2_1177(.VSS(VSS),.VDD(VDD),.Y(g23318),.A(g19716),.B(g16192));
  OR2 OR2_1178(.VSS(VSS),.VDD(VDD),.Y(g30163),.A(g23381),.B(g28523));
  OR2 OR2_1179(.VSS(VSS),.VDD(VDD),.Y(g33034),.A(g32340),.B(g21844));
  OR2 OR2_1180(.VSS(VSS),.VDD(VDD),.Y(g26920),.A(g25865),.B(g18283));
  OR2 OR2_1181(.VSS(VSS),.VDD(VDD),.Y(g34012),.A(g33886),.B(g18480));
  OR2 OR2_1182(.VSS(VSS),.VDD(VDD),.Y(g29253),.A(g28697),.B(g18490));
  OR2 OR2_1183(.VSS(VSS),.VDD(VDD),.Y(g24879),.A(g21465),.B(g24009));
  OR2 OR2_1184(.VSS(VSS),.VDD(VDD),.Y(g33292),.A(g32150),.B(g29601));
  OR2 OR2_1185(.VSS(VSS),.VDD(VDD),.Y(g26946),.A(g26389),.B(g24284));
  OR2 OR2_1186(.VSS(VSS),.VDD(VDD),.Y(g30541),.A(g30281),.B(g22087));
  OR2 OR2_1187(.VSS(VSS),.VDD(VDD),.Y(g30473),.A(g30196),.B(g21944));
  OR2 OR2_1188(.VSS(VSS),.VDD(VDD),.Y(g24337),.A(g23540),.B(g18754));
  OR2 OR2_1189(.VSS(VSS),.VDD(VDD),.Y(g27489),.A(g24608),.B(g26022));
  OR2 OR2_1190(.VSS(VSS),.VDD(VDD),.Y(g29236),.A(g28313),.B(g18287));
  OR2 OR2_1191(.VSS(VSS),.VDD(VDD),.Y(g28526),.A(g27285),.B(g26178));
  OR2 OR2_1192(.VSS(VSS),.VDD(VDD),.Y(g26344),.A(g2927),.B(g25010));
  OR2 OR2_1193(.VSS(VSS),.VDD(VDD),.Y(g27016),.A(g26821),.B(g14585));
  OR2 OR2_1194(.VSS(VSS),.VDD(VDD),.Y(g30359),.A(g30075),.B(g18385));
  OR2 OR2_1195(.VSS(VSS),.VDD(VDD),.Y(g34724),.A(g34702),.B(g18152));
  OR2 OR2_1196(.VSS(VSS),.VDD(VDD),.Y(g28402),.A(g27213),.B(g15873));
  OR2 OR2_1197(.VSS(VSS),.VDD(VDD),.Y(g30535),.A(g30225),.B(g22081));
  OR2 OR2_1198(.VSS(VSS),.VDD(VDD),.Y(g30434),.A(g30024),.B(g21818));
  OR2 OR2_1199(.VSS(VSS),.VDD(VDD),.Y(g19576),.A(g17138),.B(g14202));
  OR2 OR2_1200(.VSS(VSS),.VDD(VDD),.Y(g30358),.A(g30108),.B(g18381));
  OR2 OR2_1201(.VSS(VSS),.VDD(VDD),.Y(g34535),.A(g34309),.B(g34073));
  OR2 OR2_1202(.VSS(VSS),.VDD(VDD),.Y(g29264),.A(g28248),.B(g18618));
  OR2 OR2_1203(.VSS(VSS),.VDD(VDD),.Y(g29790),.A(g25975),.B(g28242));
  OR2 OR2_1204(.VSS(VSS),.VDD(VDD),.Y(g16928),.A(g13525),.B(g11127));
  OR2 OR2_1205(.VSS(VSS),.VDD(VDD),.Y(g27544),.A(g26087),.B(g24671));
  OR3 OR3_32(.VSS(VSS),.VDD(VDD),.Y(g33164),.A(g32203),.B(I30727),.C(I30728));
  OR2 OR2_1206(.VSS(VSS),.VDD(VDD),.Y(g17268),.A(g9220),.B(g14387));
  OR2 OR2_1207(.VSS(VSS),.VDD(VDD),.Y(g24919),.A(g21606),.B(g22143));
  OR2 OR2_1208(.VSS(VSS),.VDD(VDD),.Y(g30344),.A(g29630),.B(g18298));
  OR2 OR2_1209(.VSS(VSS),.VDD(VDD),.Y(g31891),.A(g31305),.B(g21824));
  OR2 OR2_1210(.VSS(VSS),.VDD(VDD),.Y(g28077),.A(g27120),.B(g21879));
  OR2 OR2_1211(.VSS(VSS),.VDD(VDD),.Y(g33891),.A(g33264),.B(g33269));
  OR2 OR2_1212(.VSS(VSS),.VDD(VDD),.Y(g31474),.A(g29668),.B(g13583));
  OR2 OR2_1213(.VSS(VSS),.VDD(VDD),.Y(g33575),.A(g33086),.B(g18420));
  OR2 OR2_1214(.VSS(VSS),.VDD(VDD),.Y(g24444),.A(g10890),.B(g22400));
  OR2 OR2_1215(.VSS(VSS),.VDD(VDD),.Y(g30291),.A(g28672),.B(g27685));
  OR2 OR2_1216(.VSS(VSS),.VDD(VDD),.Y(g25789),.A(g25285),.B(g14543));
  OR2 OR2_1217(.VSS(VSS),.VDD(VDD),.Y(g32387),.A(g31489),.B(g29952));
  OR2 OR2_1218(.VSS(VSS),.VDD(VDD),.Y(g25724),.A(g25043),.B(g22007));
  OR2 OR2_1219(.VSS(VSS),.VDD(VDD),.Y(g28688),.A(g27435),.B(g16639));
  OR2 OR2_1220(.VSS(VSS),.VDD(VDD),.Y(g33537),.A(g33244),.B(g21716));
  OR2 OR2_1221(.VSS(VSS),.VDD(VDD),.Y(g22487),.A(g21512),.B(g12794));
  OR2 OR2_1222(.VSS(VSS),.VDD(VDD),.Y(g28102),.A(g27995),.B(g22089));
  OR2 OR2_1223(.VSS(VSS),.VDD(VDD),.Y(g33283),.A(g31995),.B(g30318));
  OR2 OR2_1224(.VSS(VSS),.VDD(VDD),.Y(g27383),.A(g24569),.B(g25961));
  OR2 OR2_1225(.VSS(VSS),.VDD(VDD),.Y(g33606),.A(g33369),.B(g18522));
  OR2 OR2_1226(.VSS(VSS),.VDD(VDD),.Y(g31303),.A(g29592),.B(g29606));
  OR2 OR2_1227(.VSS(VSS),.VDD(VDD),.Y(g33303),.A(g32159),.B(g29638));
  OR2 OR2_1228(.VSS(VSS),.VDD(VDD),.Y(g34029),.A(g33798),.B(g18703));
  OR2 OR2_1229(.VSS(VSS),.VDD(VDD),.Y(g26927),.A(g26711),.B(g18539));
  OR2 OR2_1230(.VSS(VSS),.VDD(VDD),.Y(g30506),.A(g30179),.B(g22027));
  OR2 OR2_1231(.VSS(VSS),.VDD(VDD),.Y(g28066),.A(g27553),.B(g21819));
  OR2 OR2_1232(.VSS(VSS),.VDD(VDD),.Y(g21895),.A(g20135),.B(g15108));
  OR2 OR2_1233(.VSS(VSS),.VDD(VDD),.Y(g34028),.A(g33720),.B(g18684));
  OR2 OR2_1234(.VSS(VSS),.VDD(VDD),.Y(g32368),.A(g29881),.B(g31310));
  OR2 OR2_1235(.VSS(VSS),.VDD(VDD),.Y(g33982),.A(g33865),.B(g18372));
  OR2 OR2_1236(.VSS(VSS),.VDD(VDD),.Y(g25682),.A(g24658),.B(g18640));
  OR2 OR2_1237(.VSS(VSS),.VDD(VDD),.Y(g29274),.A(g28360),.B(g18642));
  OR2 OR2_1238(.VSS(VSS),.VDD(VDD),.Y(g24561),.A(I23755),.B(I23756));
  OR2 OR2_1239(.VSS(VSS),.VDD(VDD),.Y(g24353),.A(g23682),.B(g18822));
  OR2 OR2_1240(.VSS(VSS),.VDD(VDD),.Y(g26903),.A(g26388),.B(g24220));
  OR2 OR2_1241(.VSS(VSS),.VDD(VDD),.Y(g35000),.A(g34953),.B(g34999));
  OR2 OR2_1242(.VSS(VSS),.VDD(VDD),.Y(g11737),.A(g8359),.B(g8292));
  OR2 OR2_1243(.VSS(VSS),.VDD(VDD),.Y(g9012),.A(g2047),.B(g2066));
  OR2 OR2_1244(.VSS(VSS),.VDD(VDD),.Y(g26755),.A(g10776),.B(g24457));
  OR2 OR2_1245(.VSS(VSS),.VDD(VDD),.Y(g28511),.A(g27272),.B(g16208));
  OR2 OR2_1246(.VSS(VSS),.VDD(VDD),.Y(g32229),.A(g31148),.B(g29652));
  OR2 OR2_1247(.VSS(VSS),.VDD(VDD),.Y(g26770),.A(g24471),.B(g10732));
  OR2 OR2_1248(.VSS(VSS),.VDD(VDD),.Y(g24336),.A(g24012),.B(g18753));
  OR2 OR2_1249(.VSS(VSS),.VDD(VDD),.Y(g27837),.A(g17401),.B(g26725));
  OR2 OR2_1250(.VSS(VSS),.VDD(VDD),.Y(g33390),.A(g32276),.B(g29968));
  OR2 OR2_1251(.VSS(VSS),.VDD(VDD),.Y(g32228),.A(g31147),.B(g29651));
  OR2 OR2_1252(.VSS(VSS),.VDD(VDD),.Y(g25760),.A(g25238),.B(g22109));
  OR2 OR2_1253(.VSS(VSS),.VDD(VDD),.Y(g29292),.A(g28556),.B(g18776));
  OR2 OR2_1254(.VSS(VSS),.VDD(VDD),.Y(g34649),.A(g33111),.B(g34492));
  OR2 OR2_1255(.VSS(VSS),.VDD(VDD),.Y(g34240),.A(g32910),.B(g33958));
  OR2 OR2_1256(.VSS(VSS),.VDD(VDD),.Y(g30491),.A(g30178),.B(g21987));
  OR2 OR2_1257(.VSS(VSS),.VDD(VDD),.Y(g34903),.A(g34859),.B(g21690));
  OR2 OR2_1258(.VSS(VSS),.VDD(VDD),.Y(g23297),.A(g19692),.B(g16178));
  OR2 OR2_1259(.VSS(VSS),.VDD(VDD),.Y(g34604),.A(g34563),.B(g15076));
  OR2 OR2_1260(.VSS(VSS),.VDD(VDD),.Y(g26899),.A(g26844),.B(g18199));
  OR2 OR2_1261(.VSS(VSS),.VDD(VDD),.Y(g30563),.A(g29347),.B(g22134));
  OR2 OR2_1262(.VSS(VSS),.VDD(VDD),.Y(g26898),.A(g26387),.B(g18194));
  OR2 OR2_1263(.VSS(VSS),.VDD(VDD),.Y(g28085),.A(g27263),.B(g18700));
  OR2 OR2_1264(.VSS(VSS),.VDD(VDD),.Y(g28076),.A(g27098),.B(g21878));
  OR2 OR2_1265(.VSS(VSS),.VDD(VDD),.Y(g28721),.A(g27488),.B(g16705));
  OR2 OR2_1266(.VSS(VSS),.VDD(VDD),.Y(g28596),.A(g27336),.B(g26291));
  OR2 OR2_1267(.VSS(VSS),.VDD(VDD),.Y(g28054),.A(g27723),.B(g18170));
  OR2 OR2_1268(.VSS(VSS),.VDD(VDD),.Y(g33553),.A(g33403),.B(g18350));
  OR2 OR2_1269(.VSS(VSS),.VDD(VDD),.Y(g15803),.A(g12924),.B(g10528));
  OR2 OR2_1270(.VSS(VSS),.VDD(VDD),.Y(g22217),.A(g21302),.B(g17617));
  OR2 OR2_1271(.VSS(VSS),.VDD(VDD),.Y(g33949),.A(g32446),.B(g33459));
  OR2 OR2_1272(.VSS(VSS),.VDD(VDD),.Y(g31326),.A(g29627),.B(g29640));
  OR2 OR2_1273(.VSS(VSS),.VDD(VDD),.Y(g32386),.A(g31488),.B(g29949));
  OR2 OR2_1274(.VSS(VSS),.VDD(VDD),.Y(g30395),.A(g29841),.B(g21754));
  OR2 OR2_1275(.VSS(VSS),.VDD(VDD),.Y(g34794),.A(g34746),.B(g18571));
  OR2 OR2_1276(.VSS(VSS),.VDD(VDD),.Y(g25649),.A(g24654),.B(g21742));
  OR4 OR4_44(.VSS(VSS),.VDD(VDD),.Y(I26644),.A(g27057),.B(g27044),.C(g27039),.D(g27032));
  OR4 OR4_45(.VSS(VSS),.VDD(VDD),.Y(g27037),.A(g26236),.B(g26218),.C(g26195),.D(g26171));
  OR2 OR2_1277(.VSS(VSS),.VDD(VDD),.Y(g34262),.A(g34075),.B(g18697));
  OR2 OR2_1278(.VSS(VSS),.VDD(VDD),.Y(g33536),.A(g33241),.B(g21715));
  OR2 OR2_1279(.VSS(VSS),.VDD(VDD),.Y(g33040),.A(g32164),.B(g24313));
  OR2 OR2_1280(.VSS(VSS),.VDD(VDD),.Y(g33948),.A(g32442),.B(g33458));
  OR2 OR2_1281(.VSS(VSS),.VDD(VDD),.Y(g25648),.A(g24644),.B(g21741));
  OR2 OR2_1282(.VSS(VSS),.VDD(VDD),.Y(g28773),.A(g27535),.B(g16803));
  OR2 OR2_1283(.VSS(VSS),.VDD(VDD),.Y(g31757),.A(g29992),.B(g30010));
  OR2 OR2_1284(.VSS(VSS),.VDD(VDD),.Y(g31904),.A(g31780),.B(g21923));
  OR2 OR2_1285(.VSS(VSS),.VDD(VDD),.Y(g34633),.A(g34481),.B(g18690));
  OR2 OR2_1286(.VSS(VSS),.VDD(VDD),.Y(g25604),.A(g24717),.B(g18115));
  OR2 OR2_1287(.VSS(VSS),.VDD(VDD),.Y(g25755),.A(g25192),.B(g22102));
  OR2 OR2_1288(.VSS(VSS),.VDD(VDD),.Y(g33621),.A(g33365),.B(g18775));
  OR2 OR2_1289(.VSS(VSS),.VDD(VDD),.Y(g34719),.A(g34701),.B(g18133));
  OR2 OR2_1290(.VSS(VSS),.VDD(VDD),.Y(g28180),.A(g20242),.B(g27511));
  OR2 OR2_1291(.VSS(VSS),.VDD(VDD),.Y(g28670),.A(g27412),.B(g16618));
  OR2 OR2_1292(.VSS(VSS),.VDD(VDD),.Y(g26926),.A(g26633),.B(g18531));
  OR2 OR2_1293(.VSS(VSS),.VDD(VDD),.Y(g32429),.A(g30318),.B(g31794));
  OR2 OR2_1294(.VSS(VSS),.VDD(VDD),.Y(g30521),.A(g29331),.B(g22042));
  OR2 OR2_1295(.VSS(VSS),.VDD(VDD),.Y(g14511),.A(g10685),.B(g546));
  OR2 OR2_1296(.VSS(VSS),.VDD(VDD),.Y(g33564),.A(g33332),.B(g18388));
  OR2 OR2_1297(.VSS(VSS),.VDD(VDD),.Y(g26099),.A(g24506),.B(g22538));
  OR2 OR2_1298(.VSS(VSS),.VDD(VDD),.Y(g29283),.A(g28627),.B(g18746));
  OR2 OR2_1299(.VSS(VSS),.VDD(VDD),.Y(g28734),.A(g27508),.B(g16736));
  OR2 OR2_1300(.VSS(VSS),.VDD(VDD),.Y(g28335),.A(g27132),.B(g15818));
  OR2 OR2_1301(.VSS(VSS),.VDD(VDD),.Y(g29303),.A(g28703),.B(g18801));
  OR2 OR2_1302(.VSS(VSS),.VDD(VDD),.Y(g24374),.A(g19345),.B(g24004));
  OR2 OR2_1303(.VSS(VSS),.VDD(VDD),.Y(g30440),.A(g29771),.B(g21849));
  OR2 OR2_1304(.VSS(VSS),.VDD(VDD),.Y(g34440),.A(g34364),.B(g24226));
  OR2 OR2_1305(.VSS(VSS),.VDD(VDD),.Y(g25767),.A(g25207),.B(g12015));
  OR2 OR2_1306(.VSS(VSS),.VDD(VDD),.Y(g28667),.A(g27410),.B(g16616));
  OR2 OR2_1307(.VSS(VSS),.VDD(VDD),.Y(g33062),.A(g31977),.B(g22065));
  OR2 OR2_1308(.VSS(VSS),.VDD(VDD),.Y(g22531),.A(g20773),.B(g20922));
  OR2 OR2_1309(.VSS(VSS),.VDD(VDD),.Y(g27589),.A(g26177),.B(g24763));
  OR2 OR2_1310(.VSS(VSS),.VDD(VDD),.Y(g16448),.A(g13287),.B(g10934));
  OR2 OR2_1311(.VSS(VSS),.VDD(VDD),.Y(g30389),.A(g29969),.B(g18554));
  OR2 OR2_1312(.VSS(VSS),.VDD(VDD),.Y(g24260),.A(g23373),.B(g18313));
  OR2 OR2_1313(.VSS(VSS),.VDD(VDD),.Y(g27524),.A(g26050),.B(g24649));
  OR2 OR2_1314(.VSS(VSS),.VDD(VDD),.Y(g25633),.A(g24420),.B(g18282));
  OR2 OR2_1315(.VSS(VSS),.VDD(VDD),.Y(g31872),.A(g31524),.B(g18535));
  OR2 OR2_1316(.VSS(VSS),.VDD(VDD),.Y(g24842),.A(g7804),.B(g22669));
  OR2 OR2_1317(.VSS(VSS),.VDD(VDD),.Y(g30388),.A(g30023),.B(g18534));
  OR2 OR2_1318(.VSS(VSS),.VDD(VDD),.Y(g34612),.A(g34514),.B(g18566));
  OR2 OR2_1319(.VSS(VSS),.VDD(VDD),.Y(g25719),.A(g25089),.B(g18761));
  OR2 OR2_1320(.VSS(VSS),.VDD(VDD),.Y(g28619),.A(g27358),.B(g16517));
  OR2 OR2_1321(.VSS(VSS),.VDD(VDD),.Y(g34099),.A(g33684),.B(g33689));
  OR2 OR2_1322(.VSS(VSS),.VDD(VDD),.Y(g30534),.A(g30213),.B(g22080));
  OR2 OR2_1323(.VSS(VSS),.VDD(VDD),.Y(g19441),.A(g15507),.B(g12931));
  OR2 OR2_1324(.VSS(VSS),.VDD(VDD),.Y(g25718),.A(g25187),.B(g21971));
  OR2 OR2_1325(.VSS(VSS),.VDD(VDD),.Y(g28618),.A(g27357),.B(g16516));
  OR2 OR2_1326(.VSS(VSS),.VDD(VDD),.Y(g34251),.A(g34157),.B(g18147));
  OR2 OR2_1327(.VSS(VSS),.VDD(VDD),.Y(g28279),.A(g27087),.B(g25909));
  OR2 OR2_1328(.VSS(VSS),.VDD(VDD),.Y(g26766),.A(g10776),.B(g24460));
  OR2 OR2_1329(.VSS(VSS),.VDD(VDD),.Y(g30462),.A(g30228),.B(g21933));
  OR2 OR2_1330(.VSS(VSS),.VDD(VDD),.Y(g23296),.A(g19691),.B(g16177));
  OR2 OR2_1331(.VSS(VSS),.VDD(VDD),.Y(g34462),.A(g34334),.B(g18685));
  OR2 OR2_1332(.VSS(VSS),.VDD(VDD),.Y(g28286),.A(g27090),.B(g15757));
  OR2 OR2_1333(.VSS(VSS),.VDD(VDD),.Y(g32245),.A(g31167),.B(g29684));
  OR2 OR2_1334(.VSS(VSS),.VDD(VDD),.Y(g34032),.A(g33816),.B(g18706));
  OR2 OR2_1335(.VSS(VSS),.VDD(VDD),.Y(g28306),.A(g27104),.B(g15794));
  OR2 OR2_1336(.VSS(VSS),.VDD(VDD),.Y(g33574),.A(g33362),.B(g18416));
  OR2 OR2_1337(.VSS(VSS),.VDD(VDD),.Y(g33047),.A(g31944),.B(g21927));
  OR4 OR4_46(.VSS(VSS),.VDD(VDD),.Y(I26741),.A(g22881),.B(g22905),.C(g22928),.D(g27402));
  OR2 OR2_1338(.VSS(VSS),.VDD(VDD),.Y(g31912),.A(g31752),.B(g21998));
  OR2 OR2_1339(.VSS(VSS),.VDD(VDD),.Y(g31311),.A(g26103),.B(g29618));
  OR2 OR2_1340(.VSS(VSS),.VDD(VDD),.Y(g23197),.A(g19571),.B(g15966));
  OR2 OR2_1341(.VSS(VSS),.VDD(VDD),.Y(g25612),.A(g24941),.B(g18132));
  OR2 OR2_1342(.VSS(VSS),.VDD(VDD),.Y(g28815),.A(g27546),.B(g16842));
  OR2 OR2_1343(.VSS(VSS),.VDD(VDD),.Y(g29483),.A(g25801),.B(g28130));
  OR2 OR2_1344(.VSS(VSS),.VDD(VDD),.Y(g16811),.A(g8690),.B(g13914));
  OR2 OR2_1345(.VSS(VSS),.VDD(VDD),.Y(g25701),.A(g25054),.B(g21920));
  OR4 OR4_47(.VSS(VSS),.VDD(VDD),.Y(I30055),.A(g31070),.B(g31170),.C(g30614),.D(g30673));
  OR2 OR2_1346(.VSS(VSS),.VDD(VDD),.Y(g24705),.A(g2890),.B(g23267));
  OR2 OR2_1347(.VSS(VSS),.VDD(VDD),.Y(g33051),.A(g32316),.B(g21958));
  OR2 OR2_1348(.VSS(VSS),.VDD(VDD),.Y(g24255),.A(g22835),.B(g18308));
  OR2 OR2_1349(.VSS(VSS),.VDD(VDD),.Y(g33592),.A(g33412),.B(g18475));
  OR2 OR2_1350(.VSS(VSS),.VDD(VDD),.Y(g30360),.A(g30145),.B(g18386));
  OR2 OR2_1351(.VSS(VSS),.VDD(VDD),.Y(g24270),.A(g23165),.B(g18614));
  OR2 OR2_1352(.VSS(VSS),.VDD(VDD),.Y(g26911),.A(g26612),.B(g24230));
  OR4 OR4_48(.VSS(VSS),.VDD(VDD),.Y(I30741),.A(g32085),.B(g32030),.C(g32224),.D(g32013));
  OR2 OR2_1353(.VSS(VSS),.VDD(VDD),.Y(g30447),.A(g29798),.B(g21856));
  OR2 OR2_1354(.VSS(VSS),.VDD(VDD),.Y(g21894),.A(g20112),.B(g15107));
  OR2 OR2_1355(.VSS(VSS),.VDD(VDD),.Y(g34447),.A(g34363),.B(g18552));
  OR2 OR2_1356(.VSS(VSS),.VDD(VDD),.Y(g32995),.A(g32330),.B(g18375));
  OR2 OR2_1357(.VSS(VSS),.VDD(VDD),.Y(g24460),.A(g10967),.B(g22450));
  OR2 OR2_1358(.VSS(VSS),.VDD(VDD),.Y(g29904),.A(g28312),.B(g26146));
  OR2 OR2_1359(.VSS(VSS),.VDD(VDD),.Y(g13657),.A(g7251),.B(g10616));
  OR2 OR2_1360(.VSS(VSS),.VDD(VDD),.Y(g29252),.A(g28712),.B(g18486));
  OR2 OR2_1361(.VSS(VSS),.VDD(VDD),.Y(g28884),.A(g27568),.B(g16885));
  OR2 OR2_1362(.VSS(VSS),.VDD(VDD),.Y(g26785),.A(g10776),.B(g24468));
  OR2 OR2_1363(.VSS(VSS),.VDD(VDD),.Y(g24267),.A(g23439),.B(g18611));
  OR2 OR2_1364(.VSS(VSS),.VDD(VDD),.Y(g30451),.A(g29877),.B(g21860));
  OR2 OR2_1365(.VSS(VSS),.VDD(VDD),.Y(g30472),.A(g30186),.B(g21943));
  OR4 OR4_49(.VSS(VSS),.VDD(VDD),.Y(I30735),.A(g32369),.B(g32376),.C(g32089),.D(g32035));
  OR2 OR2_1366(.VSS(VSS),.VDD(VDD),.Y(g34629),.A(g34495),.B(g18654));
  OR4 OR4_50(.VSS(VSS),.VDD(VDD),.Y(g17569),.A(g14416),.B(g14394),.C(g11995),.D(I18492));
  OR2 OR2_1367(.VSS(VSS),.VDD(VDD),.Y(g34451),.A(g34393),.B(g18664));
  OR2 OR2_1368(.VSS(VSS),.VDD(VDD),.Y(g34628),.A(g34493),.B(g18653));
  OR2 OR2_1369(.VSS(VSS),.VDD(VDD),.Y(g34911),.A(g34909),.B(g18188));
  OR2 OR2_1370(.VSS(VSS),.VDD(VDD),.Y(g26950),.A(g26357),.B(g24288));
  OR2 OR2_1371(.VSS(VSS),.VDD(VDD),.Y(g22751),.A(g19333),.B(g15716));
  OR3 OR3_33(.VSS(VSS),.VDD(VDD),.Y(g27008),.A(g26866),.B(g21370),.C(I25736));
  OR2 OR2_1372(.VSS(VSS),.VDD(VDD),.Y(g22639),.A(g18950),.B(g15612));
  OR2 OR2_1373(.VSS(VSS),.VDD(VDD),.Y(g27555),.A(g26095),.B(g24686));
  OR2 OR2_1374(.VSS(VSS),.VDD(VDD),.Y(g28580),.A(g27328),.B(g26275));
  OR2 OR2_1375(.VSS(VSS),.VDD(VDD),.Y(g29508),.A(g28152),.B(g27041));
  OR3 OR3_34(.VSS(VSS),.VDD(VDD),.Y(g8476),.A(g1399),.B(g1459),.C(I12611));
  OR2 OR2_1376(.VSS(VSS),.VDD(VDD),.Y(g20160),.A(g16163),.B(g13415));
  OR2 OR2_1377(.VSS(VSS),.VDD(VDD),.Y(g30355),.A(g30131),.B(g18360));
  OR2 OR2_1378(.VSS(VSS),.VDD(VDD),.Y(g27570),.A(g26126),.B(g24722));
  OR2 OR2_1379(.VSS(VSS),.VDD(VDD),.Y(g31929),.A(g31540),.B(g22093));
  OR2 OR2_1380(.VSS(VSS),.VDD(VDD),.Y(g32989),.A(g32241),.B(g18326));
  OR2 OR2_1381(.VSS(VSS),.VDD(VDD),.Y(g30370),.A(g30135),.B(g18440));
  OR2 OR2_1382(.VSS(VSS),.VDD(VDD),.Y(g25629),.A(g24962),.B(g18258));
  OR2 OR2_1383(.VSS(VSS),.VDD(VDD),.Y(g27907),.A(g17424),.B(g26770));
  OR2 OR2_1384(.VSS(VSS),.VDD(VDD),.Y(g16959),.A(g13542),.B(g11142));
  OR2 OR2_1385(.VSS(VSS),.VDD(VDD),.Y(g31020),.A(g29375),.B(g28164));
  OR2 OR2_1386(.VSS(VSS),.VDD(VDD),.Y(g31928),.A(g31517),.B(g22092));
  OR2 OR2_1387(.VSS(VSS),.VDD(VDD),.Y(g14187),.A(g8871),.B(g11771));
  OR2 OR2_1388(.VSS(VSS),.VDD(VDD),.Y(g32988),.A(g32232),.B(g18325));
  OR2 OR2_1389(.VSS(VSS),.VDD(VDD),.Y(g28084),.A(g27254),.B(g18698));
  OR2 OR2_1390(.VSS(VSS),.VDD(VDD),.Y(g33020),.A(g32160),.B(g21734));
  OR2 OR2_1391(.VSS(VSS),.VDD(VDD),.Y(g33583),.A(g33074),.B(g18448));
  OR2 OR2_1392(.VSS(VSS),.VDD(VDD),.Y(g25628),.A(g24600),.B(g18249));
  OR2 OR2_1393(.VSS(VSS),.VDD(VDD),.Y(g25911),.A(g22514),.B(g24510));
  OR2 OR2_1394(.VSS(VSS),.VDD(VDD),.Y(g27239),.A(g25881),.B(g24465));
  OR2 OR2_1395(.VSS(VSS),.VDD(VDD),.Y(g19605),.A(g15707),.B(g13063));
  OR2 OR2_1396(.VSS(VSS),.VDD(VDD),.Y(g33046),.A(g32308),.B(g21912));
  OR2 OR2_1397(.VSS(VSS),.VDD(VDD),.Y(g32271),.A(g31209),.B(g29731));
  OR2 OR2_1398(.VSS(VSS),.VDD(VDD),.Y(g34172),.A(g33795),.B(g19914));
  OR4 OR4_51(.VSS(VSS),.VDD(VDD),.Y(g28179),.A(g27494),.B(g27474),.C(g27445),.D(g27421));
  OR2 OR2_1399(.VSS(VSS),.VDD(VDD),.Y(g27567),.A(g26121),.B(g24714));
  OR2 OR2_1400(.VSS(VSS),.VDD(VDD),.Y(g27238),.A(g25879),.B(g24464));
  OR4 OR4_52(.VSS(VSS),.VDD(VDD),.Y(g17510),.A(g14393),.B(g14362),.C(g11972),.D(I18449));
  OR2 OR2_1401(.VSS(VSS),.VDD(VDD),.Y(g30394),.A(g29805),.B(g21753));
  OR2 OR2_1402(.VSS(VSS),.VDD(VDD),.Y(g30367),.A(g30133),.B(g18418));
  OR2 OR2_1403(.VSS(VSS),.VDD(VDD),.Y(g24201),.A(g22848),.B(g18104));
  OR2 OR2_1404(.VSS(VSS),.VDD(VDD),.Y(g24277),.A(g23188),.B(g18647));
  OR2 OR2_1405(.VSS(VSS),.VDD(VDD),.Y(g25591),.A(g24642),.B(g21705));
  OR2 OR2_1406(.VSS(VSS),.VDD(VDD),.Y(g33282),.A(g32143),.B(g29577));
  OR4 OR4_53(.VSS(VSS),.VDD(VDD),.Y(g28186),.A(g27209),.B(g27185),.C(g27161),.D(g27146));
  OR2 OR2_1407(.VSS(VSS),.VDD(VDD),.Y(g28685),.A(g27433),.B(g16637));
  OR2 OR2_1408(.VSS(VSS),.VDD(VDD),.Y(g31302),.A(g29590),.B(g28302));
  OR2 OR2_1409(.VSS(VSS),.VDD(VDD),.Y(g28373),.A(g27180),.B(g15849));
  OR2 OR2_1410(.VSS(VSS),.VDD(VDD),.Y(g25754),.A(g25179),.B(g22101));
  OR2 OR2_1411(.VSS(VSS),.VDD(VDD),.Y(g30420),.A(g29769),.B(g21804));
  OR2 OR2_1412(.VSS(VSS),.VDD(VDD),.Y(g28417),.A(g27219),.B(g15881));
  OR2 OR2_1413(.VSS(VSS),.VDD(VDD),.Y(g24782),.A(g23857),.B(g23872));
  OR2 OR2_1414(.VSS(VSS),.VDD(VDD),.Y(g30446),.A(g29788),.B(g21855));
  OR2 OR2_1415(.VSS(VSS),.VDD(VDD),.Y(g34446),.A(g34390),.B(g18550));
  OR2 OR2_1416(.VSS(VSS),.VDD(VDD),.Y(g34318),.A(g25850),.B(g34063));
  OR2 OR2_1417(.VSS(VSS),.VDD(VDD),.Y(g28334),.A(g27131),.B(g15817));
  OR2 OR2_1418(.VSS(VSS),.VDD(VDD),.Y(g29756),.A(g22717),.B(g28223));
  OR2 OR2_1419(.VSS(VSS),.VDD(VDD),.Y(g24352),.A(g22157),.B(g18821));
  OR2 OR2_1420(.VSS(VSS),.VDD(VDD),.Y(g26902),.A(g26378),.B(g24219));
  OR2 OR2_1421(.VSS(VSS),.VDD(VDD),.Y(g26957),.A(g26517),.B(g24295));
  OR2 OR2_1422(.VSS(VSS),.VDD(VDD),.Y(g34025),.A(g33927),.B(g18672));
  OR2 OR2_1423(.VSS(VSS),.VDD(VDD),.Y(g31768),.A(g30033),.B(g30045));
  OR2 OR2_1424(.VSS(VSS),.VDD(VDD),.Y(g26377),.A(g24700),.B(g23007));
  OR2 OR2_1425(.VSS(VSS),.VDD(VDD),.Y(g30540),.A(g30275),.B(g22086));
  OR2 OR2_1426(.VSS(VSS),.VDD(VDD),.Y(g13295),.A(g10625),.B(g10655));
  OR2 OR2_1427(.VSS(VSS),.VDD(VDD),.Y(g15582),.A(g8977),.B(g12925));
  OR2 OR2_1428(.VSS(VSS),.VDD(VDD),.Y(g24266),.A(g22329),.B(g18561));
  OR2 OR2_1429(.VSS(VSS),.VDD(VDD),.Y(g32132),.A(g31487),.B(g31479));
  OR2 OR2_1430(.VSS(VSS),.VDD(VDD),.Y(g9535),.A(g209),.B(g538));
  OR2 OR2_1431(.VSS(VSS),.VDD(VDD),.Y(g31881),.A(g31018),.B(g21775));
  OR2 OR2_1432(.VSS(VSS),.VDD(VDD),.Y(g28216),.A(g27036),.B(g27043));
  OR2 OR2_1433(.VSS(VSS),.VDD(VDD),.Y(g24853),.A(g21452),.B(g24001));
  OR2 OR2_1434(.VSS(VSS),.VDD(VDD),.Y(g22684),.A(g19206),.B(g15703));
  OR2 OR2_1435(.VSS(VSS),.VDD(VDD),.Y(g32259),.A(g31185),.B(g29709));
  OR2 OR2_1436(.VSS(VSS),.VDD(VDD),.Y(g30377),.A(g30124),.B(g18472));
  OR2 OR2_1437(.VSS(VSS),.VDD(VDD),.Y(g32225),.A(g30576),.B(g29336));
  OR2 OR2_1438(.VSS(VSS),.VDD(VDD),.Y(g34957),.A(g34948),.B(g21662));
  OR2 OR2_1439(.VSS(VSS),.VDD(VDD),.Y(g34377),.A(g26304),.B(g34141));
  OR2 OR2_1440(.VSS(VSS),.VDD(VDD),.Y(g33027),.A(g32314),.B(g21796));
  OR3 OR3_35(.VSS(VSS),.VDD(VDD),.Y(I22912),.A(g21555),.B(g21364),.C(g21357));
  OR2 OR2_1441(.VSS(VSS),.VDD(VDD),.Y(g31890),.A(g31143),.B(g21823));
  OR2 OR2_1442(.VSS(VSS),.VDD(VDD),.Y(g24401),.A(g23811),.B(g21298));
  OR2 OR2_1443(.VSS(VSS),.VDD(VDD),.Y(g30562),.A(g30289),.B(g22133));
  OR2 OR2_1444(.VSS(VSS),.VDD(VDD),.Y(g31249),.A(g25971),.B(g29523));
  OR2 OR2_1445(.VSS(VSS),.VDD(VDD),.Y(g19359),.A(g17786),.B(g14875));
  OR2 OR2_1446(.VSS(VSS),.VDD(VDD),.Y(g34645),.A(g34556),.B(g18786));
  OR2 OR2_1447(.VSS(VSS),.VDD(VDD),.Y(g19535),.A(g15651),.B(g13020));
  OR2 OR2_1448(.VSS(VSS),.VDD(VDD),.Y(g31248),.A(g25970),.B(g29522));
  OR2 OR2_1449(.VSS(VSS),.VDD(VDD),.Y(g28747),.A(g27521),.B(g13942));
  OR2 OR2_1450(.VSS(VSS),.VDD(VDD),.Y(g34290),.A(g26848),.B(g34219));
  OR2 OR2_1451(.VSS(VSS),.VDD(VDD),.Y(g33552),.A(g33400),.B(g18343));
  OR2 OR2_1452(.VSS(VSS),.VDD(VDD),.Y(g13289),.A(g10619),.B(g10624));
  OR2 OR2_1453(.VSS(VSS),.VDD(VDD),.Y(g33003),.A(g32323),.B(g18429));
  OR3 OR3_36(.VSS(VSS),.VDD(VDD),.Y(g33204),.A(g32317),.B(I30750),.C(I30751));
  OR2 OR2_1454(.VSS(VSS),.VDD(VDD),.Y(g26895),.A(g26783),.B(g18148));
  OR2 OR2_1455(.VSS(VSS),.VDD(VDD),.Y(g31779),.A(g30050),.B(g28673));
  OR4 OR4_54(.VSS(VSS),.VDD(VDD),.Y(I31843),.A(g33470),.B(g33471),.C(g33472),.D(g33473));
  OR2 OR2_1456(.VSS(VSS),.VDD(VDD),.Y(g10800),.A(g7517),.B(g952));
  OR2 OR2_1457(.VSS(VSS),.VDD(VDD),.Y(g19344),.A(g17771),.B(g14832));
  OR2 OR2_1458(.VSS(VSS),.VDD(VDD),.Y(g27566),.A(g26119),.B(g24713));
  OR2 OR2_1459(.VSS(VSS),.VDD(VDD),.Y(g28814),.A(g27545),.B(g16841));
  OR2 OR2_1460(.VSS(VSS),.VDD(VDD),.Y(g30427),.A(g29796),.B(g21811));
  OR2 OR2_1461(.VSS(VSS),.VDD(VDD),.Y(g20276),.A(g16243),.B(g13566));
  OR2 OR2_1462(.VSS(VSS),.VDD(VDD),.Y(g29583),.A(g28182),.B(g27099));
  OR2 OR2_1463(.VSS(VSS),.VDD(VDD),.Y(g32375),.A(g29896),.B(g31324));
  OR2 OR2_1464(.VSS(VSS),.VDD(VDD),.Y(g14936),.A(g10776),.B(g8703));
  OR2 OR2_1465(.VSS(VSS),.VDD(VDD),.Y(g30366),.A(g30122),.B(g18417));
  OR4 OR4_55(.VSS(VSS),.VDD(VDD),.Y(I30054),.A(g29385),.B(g31376),.C(g30735),.D(g30825));
  OR2 OR2_1466(.VSS(VSS),.VDD(VDD),.Y(g24276),.A(g23083),.B(g18646));
  OR2 OR2_1467(.VSS(VSS),.VDD(VDD),.Y(g28751),.A(g27526),.B(g16766));
  OR2 OR2_1468(.VSS(VSS),.VDD(VDD),.Y(g28772),.A(g27534),.B(g16802));
  OR2 OR2_1469(.VSS(VSS),.VDD(VDD),.Y(g34366),.A(g26257),.B(g34133));
  OR4 OR4_56(.VSS(VSS),.VDD(VDD),.Y(I31869),.A(g33519),.B(g33520),.C(g33521),.D(g33522));
  OR2 OR2_1470(.VSS(VSS),.VDD(VDD),.Y(g34632),.A(g34565),.B(g15119));
  OR2 OR2_1471(.VSS(VSS),.VDD(VDD),.Y(g25739),.A(g25149),.B(g22054));
  OR2 OR2_1472(.VSS(VSS),.VDD(VDD),.Y(g24254),.A(g23265),.B(g18306));
  OR4 OR4_57(.VSS(VSS),.VDD(VDD),.Y(I31868),.A(g33515),.B(g33516),.C(g33517),.D(g33518));
  OR2 OR2_1473(.VSS(VSS),.VDD(VDD),.Y(g28230),.A(g27669),.B(g14261));
  OR2 OR2_1474(.VSS(VSS),.VDD(VDD),.Y(g33945),.A(g32430),.B(g33455));
  OR2 OR2_1475(.VSS(VSS),.VDD(VDD),.Y(g25738),.A(g25059),.B(g22053));
  OR2 OR2_1476(.VSS(VSS),.VDD(VDD),.Y(g25645),.A(g24679),.B(g21738));
  OR2 OR2_1477(.VSS(VSS),.VDD(VDD),.Y(g30547),.A(g30194),.B(g22118));
  OR2 OR2_1478(.VSS(VSS),.VDD(VDD),.Y(g30403),.A(g29750),.B(g21762));
  OR2 OR2_1479(.VSS(VSS),.VDD(VDD),.Y(g33999),.A(g33893),.B(g18436));
  OR2 OR2_1480(.VSS(VSS),.VDD(VDD),.Y(g33380),.A(g32234),.B(g29926));
  OR2 OR2_1481(.VSS(VSS),.VDD(VDD),.Y(g25699),.A(g25125),.B(g21918));
  OR2 OR2_1482(.VSS(VSS),.VDD(VDD),.Y(g34403),.A(g34180),.B(g25085));
  OR2 OR2_1483(.VSS(VSS),.VDD(VDD),.Y(g29282),.A(g28617),.B(g18745));
  OR2 OR2_1484(.VSS(VSS),.VDD(VDD),.Y(g28416),.A(g27218),.B(g15880));
  OR2 OR2_1485(.VSS(VSS),.VDD(VDD),.Y(g16261),.A(g7898),.B(g13469));
  OR2 OR2_1486(.VSS(VSS),.VDD(VDD),.Y(g32994),.A(g32290),.B(g18367));
  OR2 OR2_1487(.VSS(VSS),.VDD(VDD),.Y(g33998),.A(g33878),.B(g18428));
  OR2 OR2_1488(.VSS(VSS),.VDD(VDD),.Y(g29302),.A(g28601),.B(g18798));
  OR2 OR2_1489(.VSS(VSS),.VDD(VDD),.Y(g25698),.A(g25104),.B(g21917));
  OR2 OR2_1490(.VSS(VSS),.VDD(VDD),.Y(g29105),.A(g27645),.B(g17134));
  OR2 OR2_1491(.VSS(VSS),.VDD(VDD),.Y(g30481),.A(g30221),.B(g21977));
  OR2 OR2_1492(.VSS(VSS),.VDD(VDD),.Y(g7932),.A(g4072),.B(g4153));
  OR2 OR2_1493(.VSS(VSS),.VDD(VDD),.Y(g26956),.A(g26487),.B(g24294));
  OR2 OR2_1494(.VSS(VSS),.VDD(VDD),.Y(g30551),.A(g30235),.B(g22122));
  OR4 OR4_58(.VSS(VSS),.VDD(VDD),.Y(I30734),.A(g31790),.B(g32191),.C(g32086),.D(g32095));
  OR2 OR2_1495(.VSS(VSS),.VDD(VDD),.Y(g26889),.A(g26689),.B(g24195));
  OR2 OR2_1496(.VSS(VSS),.VDD(VDD),.Y(g31932),.A(g31792),.B(g22107));
  OR2 OR2_1497(.VSS(VSS),.VDD(VDD),.Y(g26888),.A(g26671),.B(g24194));
  OR3 OR3_37(.VSS(VSS),.VDD(VDD),.Y(g23721),.A(g21401),.B(g21385),.C(I22852));
  OR2 OR2_1498(.VSS(VSS),.VDD(VDD),.Y(g25632),.A(g24558),.B(g18277));
  OR2 OR2_1499(.VSS(VSS),.VDD(VDD),.Y(g28578),.A(g27327),.B(g26273));
  OR2 OR2_1500(.VSS(VSS),.VDD(VDD),.Y(g30127),.A(g28494),.B(g16805));
  OR2 OR2_1501(.VSS(VSS),.VDD(VDD),.Y(g29768),.A(g22760),.B(g28229));
  OR2 OR2_1502(.VSS(VSS),.VDD(VDD),.Y(g34127),.A(g33657),.B(g32438));
  OR2 OR2_1503(.VSS(VSS),.VDD(VDD),.Y(g31897),.A(g31237),.B(g24322));
  OR2 OR2_1504(.VSS(VSS),.VDD(VDD),.Y(g30490),.A(g30167),.B(g21986));
  OR2 OR2_1505(.VSS(VSS),.VDD(VDD),.Y(g33961),.A(g33789),.B(g21712));
  OR2 OR2_1506(.VSS(VSS),.VDD(VDD),.Y(g25661),.A(g24754),.B(g21786));
  OR2 OR2_1507(.VSS(VSS),.VDD(VDD),.Y(g27484),.A(g25988),.B(g24628));
  OR2 OR2_1508(.VSS(VSS),.VDD(VDD),.Y(g30376),.A(g30112),.B(g18471));
  OR2 OR2_1509(.VSS(VSS),.VDD(VDD),.Y(g30385),.A(g30172),.B(g18518));
  OR2 OR2_1510(.VSS(VSS),.VDD(VDD),.Y(g26931),.A(g26778),.B(g18547));
  OR2 OR2_1511(.VSS(VSS),.VDD(VDD),.Y(g30103),.A(g28477),.B(g16731));
  OR2 OR2_1512(.VSS(VSS),.VDD(VDD),.Y(g34376),.A(g26301),.B(g34140));
  OR2 OR2_1513(.VSS(VSS),.VDD(VDD),.Y(g34297),.A(g26858),.B(g34228));
  OR2 OR2_1514(.VSS(VSS),.VDD(VDD),.Y(g34103),.A(g33701),.B(g33707));
  OR2 OR2_1515(.VSS(VSS),.VDD(VDD),.Y(g33026),.A(g32307),.B(g21795));
  OR2 OR2_1516(.VSS(VSS),.VDD(VDD),.Y(g30354),.A(g30064),.B(g18359));
  OR2 OR2_1517(.VSS(VSS),.VDD(VDD),.Y(g22516),.A(g21559),.B(g12817));
  OR2 OR2_1518(.VSS(VSS),.VDD(VDD),.Y(g34980),.A(g34969),.B(g18587));
  OR3 OR3_38(.VSS(VSS),.VDD(VDD),.Y(g33212),.A(g32328),.B(I30755),.C(I30756));
  OR2 OR2_1519(.VSS(VSS),.VDD(VDD),.Y(g25715),.A(g25071),.B(g21966));
  OR2 OR2_1520(.VSS(VSS),.VDD(VDD),.Y(g8679),.A(g222),.B(g199));
  OR2 OR2_1521(.VSS(VSS),.VDD(VDD),.Y(g34095),.A(g33681),.B(g33687));
  OR2 OR2_1522(.VSS(VSS),.VDD(VDD),.Y(g30824),.A(g13833),.B(g29789));
  OR2 OR2_1523(.VSS(VSS),.VDD(VDD),.Y(g28720),.A(g27486),.B(g16704));
  OR2 OR2_1524(.VSS(VSS),.VDD(VDD),.Y(g28041),.A(g24145),.B(g26878));
  OR2 OR2_1525(.VSS(VSS),.VDD(VDD),.Y(g17264),.A(g7118),.B(g14309));
  OR2 OR2_1526(.VSS(VSS),.VDD(VDD),.Y(g28430),.A(g27229),.B(g15914));
  OR2 OR2_1527(.VSS(VSS),.VDD(VDD),.Y(g32125),.A(g30918),.B(g29376));
  OR2 OR2_1528(.VSS(VSS),.VDD(VDD),.Y(g28746),.A(g27520),.B(g16762));
  OR2 OR2_1529(.VSS(VSS),.VDD(VDD),.Y(g32977),.A(g32169),.B(g21710));
  OR2 OR2_1530(.VSS(VSS),.VDD(VDD),.Y(g19604),.A(g15704),.B(g13059));
  OR4 OR4_59(.VSS(VSS),.VDD(VDD),.Y(I30469),.A(g31672),.B(g31710),.C(g31021),.D(g30937));
  OR2 OR2_1531(.VSS(VSS),.VDD(VDD),.Y(g29249),.A(g28658),.B(g18438));
  OR2 OR2_1532(.VSS(VSS),.VDD(VDD),.Y(g26089),.A(g24501),.B(g22534));
  OR2 OR2_1533(.VSS(VSS),.VDD(VDD),.Y(g24907),.A(g21558),.B(g24015));
  OR4 OR4_60(.VSS(VSS),.VDD(VDD),.Y(I30468),.A(g29385),.B(g31376),.C(g30735),.D(g30825));
  OR2 OR2_1534(.VSS(VSS),.VDD(VDD),.Y(g29482),.A(g28524),.B(g27588));
  OR2 OR2_1535(.VSS(VSS),.VDD(VDD),.Y(g34931),.A(g2984),.B(g34912));
  OR2 OR2_1536(.VSS(VSS),.VDD(VDD),.Y(g29248),.A(g28677),.B(g18434));
  OR3 OR3_39(.VSS(VSS),.VDD(VDD),.Y(g33149),.A(g32204),.B(I30717),.C(I30718));
  OR2 OR2_1537(.VSS(VSS),.VDD(VDD),.Y(g30426),.A(g29785),.B(g21810));
  OR2 OR2_1538(.VSS(VSS),.VDD(VDD),.Y(g32353),.A(g29853),.B(g31283));
  OR2 OR2_1539(.VSS(VSS),.VDD(VDD),.Y(g33387),.A(g32263),.B(g29954));
  OR2 OR2_1540(.VSS(VSS),.VDD(VDD),.Y(g24239),.A(g22752),.B(g18250));
  OR2 OR2_1541(.VSS(VSS),.VDD(VDD),.Y(g9055),.A(g2606),.B(g2625));
  OR2 OR2_1542(.VSS(VSS),.VDD(VDD),.Y(g28684),.A(g27432),.B(g16636));
  OR2 OR2_1543(.VSS(VSS),.VDD(VDD),.Y(g32144),.A(g30927),.B(g30930));
  OR2 OR2_1544(.VSS(VSS),.VDD(VDD),.Y(g33620),.A(g33360),.B(g18774));
  OR2 OR2_1545(.VSS(VSS),.VDD(VDD),.Y(g34190),.A(g33802),.B(g33810));
  OR2 OR2_1546(.VSS(VSS),.VDD(VDD),.Y(g24238),.A(g23254),.B(g18248));
  OR2 OR2_1547(.VSS(VSS),.VDD(VDD),.Y(g30520),.A(g30272),.B(g22041));
  OR2 OR2_1548(.VSS(VSS),.VDD(VDD),.Y(g28517),.A(g27280),.B(g26154));
  OR2 OR2_1549(.VSS(VSS),.VDD(VDD),.Y(g30546),.A(g30277),.B(g22117));
  OR2 OR2_1550(.VSS(VSS),.VDD(VDD),.Y(g33971),.A(g33890),.B(g18330));
  OR2 OR2_1551(.VSS(VSS),.VDD(VDD),.Y(g29786),.A(g22843),.B(g28240));
  OR2 OR2_1552(.VSS(VSS),.VDD(VDD),.Y(g25671),.A(g24637),.B(g21828));
  OR2 OR2_1553(.VSS(VSS),.VDD(VDD),.Y(g34024),.A(g33807),.B(g24331));
  OR2 OR2_1554(.VSS(VSS),.VDD(VDD),.Y(g13938),.A(g11213),.B(g11191));
  OR2 OR2_1555(.VSS(VSS),.VDD(VDD),.Y(g24518),.A(g22517),.B(g7601));
  OR2 OR2_1556(.VSS(VSS),.VDD(VDD),.Y(g22530),.A(g16751),.B(g20171));
  OR2 OR2_1557(.VSS(VSS),.VDD(VDD),.Y(g28362),.A(g27154),.B(g15840));
  OR2 OR2_1558(.VSS(VSS),.VDD(VDD),.Y(g30497),.A(g30242),.B(g21993));
  OR2 OR2_1559(.VSS(VSS),.VDD(VDD),.Y(g24935),.A(g22937),.B(g19749));
  OR4 OR4_61(.VSS(VSS),.VDD(VDD),.Y(I12903),.A(g4222),.B(g4219),.C(g4216),.D(g4213));
  OR2 OR2_1560(.VSS(VSS),.VDD(VDD),.Y(g29233),.A(g28171),.B(g18234));
  OR2 OR2_1561(.VSS(VSS),.VDD(VDD),.Y(g26969),.A(g26313),.B(g24329));
  OR3 OR3_40(.VSS(VSS),.VDD(VDD),.Y(I18421),.A(g14447),.B(g14417),.C(g14395));
  OR2 OR2_1562(.VSS(VSS),.VDD(VDD),.Y(g32289),.A(g24796),.B(g31230));
  OR2 OR2_1563(.VSS(VSS),.VDD(VDD),.Y(g22641),.A(g18974),.B(g15631));
  OR2 OR2_1564(.VSS(VSS),.VDD(VDD),.Y(g34625),.A(g34532),.B(g18610));
  OR2 OR2_1565(.VSS(VSS),.VDD(VDD),.Y(g26968),.A(g26307),.B(g24321));
  OR4 OR4_62(.VSS(VSS),.VDD(VDD),.Y(g17464),.A(g14334),.B(g14313),.C(g11935),.D(I18385));
  OR2 OR2_1566(.VSS(VSS),.VDD(VDD),.Y(g31896),.A(g31242),.B(g24305));
  OR2 OR2_1567(.VSS(VSS),.VDD(VDD),.Y(g34250),.A(g34111),.B(g21713));
  OR2 OR2_1568(.VSS(VSS),.VDD(VDD),.Y(g32288),.A(g31226),.B(g31229));
  OR2 OR2_1569(.VSS(VSS),.VDD(VDD),.Y(g28727),.A(g27500),.B(g16729));
  OR2 OR2_1570(.VSS(VSS),.VDD(VDD),.Y(g16258),.A(g13247),.B(g10856));
  OR2 OR2_1571(.VSS(VSS),.VDD(VDD),.Y(g33011),.A(g32338),.B(g18481));
  OR2 OR2_1572(.VSS(VSS),.VDD(VDD),.Y(g30339),.A(g29629),.B(g18244));
  OR2 OR2_1573(.VSS(VSS),.VDD(VDD),.Y(g24215),.A(g23484),.B(g18196));
  OR2 OR2_1574(.VSS(VSS),.VDD(VDD),.Y(g24577),.A(g2856),.B(g22531));
  OR2 OR2_1575(.VSS(VSS),.VDD(VDD),.Y(g30338),.A(g29613),.B(g18240));
  OR2 OR2_1576(.VSS(VSS),.VDD(VDD),.Y(g34644),.A(g34555),.B(g18769));
  OR2 OR2_1577(.VSS(VSS),.VDD(VDD),.Y(g33582),.A(g33351),.B(g18444));
  OR2 OR2_1578(.VSS(VSS),.VDD(VDD),.Y(g19534),.A(g15650),.B(g13019));
  OR2 OR2_1579(.VSS(VSS),.VDD(VDD),.Y(g27241),.A(g24584),.B(g25984));
  OR2 OR2_1580(.VSS(VSS),.VDD(VDD),.Y(g28347),.A(g27138),.B(g15822));
  OR2 OR2_1581(.VSS(VSS),.VDD(VDD),.Y(g29717),.A(g28200),.B(g10883));
  OR2 OR2_1582(.VSS(VSS),.VDD(VDD),.Y(g33310),.A(g29631),.B(g32165));
  OR2 OR2_1583(.VSS(VSS),.VDD(VDD),.Y(g26894),.A(g25979),.B(g18129));
  OR2 OR2_1584(.VSS(VSS),.VDD(VDD),.Y(g33627),.A(g33376),.B(g18826));
  OR2 OR2_1585(.VSS(VSS),.VDD(VDD),.Y(g31925),.A(g31789),.B(g22061));
  OR2 OR2_1586(.VSS(VSS),.VDD(VDD),.Y(g32976),.A(g32207),.B(g21704));
  OR2 OR2_1587(.VSS(VSS),.VDD(VDD),.Y(g32985),.A(g31963),.B(g18266));
  OR2 OR2_1588(.VSS(VSS),.VDD(VDD),.Y(g24349),.A(g23646),.B(g18805));
  OR2 OR2_1589(.VSS(VSS),.VDD(VDD),.Y(g16810),.A(g13461),.B(g11032));
  OR2 OR2_1590(.VSS(VSS),.VDD(VDD),.Y(g25700),.A(g25040),.B(g21919));
  OR2 OR2_1591(.VSS(VSS),.VDD(VDD),.Y(g28600),.A(g27339),.B(g16427));
  OR2 OR2_1592(.VSS(VSS),.VDD(VDD),.Y(g25659),.A(g24707),.B(g21784));
  OR2 OR2_1593(.VSS(VSS),.VDD(VDD),.Y(g25625),.A(g24553),.B(g18226));
  OR2 OR2_1594(.VSS(VSS),.VDD(VDD),.Y(g20083),.A(g2902),.B(g17058));
  OR2 OR2_1595(.VSS(VSS),.VDD(VDD),.Y(g30527),.A(g30192),.B(g22073));
  OR2 OR2_1596(.VSS(VSS),.VDD(VDD),.Y(g30411),.A(g29872),.B(g21770));
  OR2 OR2_1597(.VSS(VSS),.VDD(VDD),.Y(g33050),.A(g31974),.B(g21930));
  OR2 OR2_1598(.VSS(VSS),.VDD(VDD),.Y(g32374),.A(g29895),.B(g31323));
  OR3 OR3_41(.VSS(VSS),.VDD(VDD),.Y(g33958),.A(g33532),.B(I31873),.C(I31874));
  OR2 OR2_1599(.VSS(VSS),.VDD(VDD),.Y(g24348),.A(g22149),.B(g18804));
  OR2 OR2_1600(.VSS(VSS),.VDD(VDD),.Y(g34411),.A(g34186),.B(g25142));
  OR2 OR2_1601(.VSS(VSS),.VDD(VDD),.Y(g16970),.A(g13567),.B(g11163));
  OR2 OR2_1602(.VSS(VSS),.VDD(VDD),.Y(g25658),.A(g24635),.B(g21783));
  OR2 OR2_1603(.VSS(VSS),.VDD(VDD),.Y(g28372),.A(g27178),.B(g15848));
  OR2 OR2_1604(.VSS(VSS),.VDD(VDD),.Y(g23217),.A(g19588),.B(g16023));
  OR2 OR2_1605(.VSS(VSS),.VDD(VDD),.Y(g33386),.A(g32258),.B(g29951));
  OR2 OR2_1606(.VSS(VSS),.VDD(VDD),.Y(g26910),.A(g26571),.B(g24228));
  OR2 OR2_1607(.VSS(VSS),.VDD(VDD),.Y(g33603),.A(g33372),.B(g18515));
  OR2 OR2_1608(.VSS(VSS),.VDD(VDD),.Y(g25943),.A(g24423),.B(g22299));
  OR4 OR4_63(.VSS(VSS),.VDD(VDD),.Y(I30740),.A(g31776),.B(g32188),.C(g32083),.D(g32087));
  OR2 OR2_1609(.VSS(VSS),.VDD(VDD),.Y(g13623),.A(g482),.B(g12527));
  OR2 OR2_1610(.VSS(VSS),.VDD(VDD),.Y(g25644),.A(g24622),.B(g21737));
  OR2 OR2_1611(.VSS(VSS),.VDD(VDD),.Y(g30503),.A(g30243),.B(g22024));
  OR2 OR2_1612(.VSS(VSS),.VDD(VDD),.Y(g28063),.A(g27541),.B(g21773));
  OR2 OR2_1613(.VSS(VSS),.VDD(VDD),.Y(g34894),.A(g34862),.B(g21678));
  OR2 OR2_1614(.VSS(VSS),.VDD(VDD),.Y(g29148),.A(g27651),.B(g26606));
  OR2 OR2_1615(.VSS(VSS),.VDD(VDD),.Y(g32392),.A(g31513),.B(g30000));
  OR2 OR2_1616(.VSS(VSS),.VDD(VDD),.Y(g27515),.A(g26051),.B(g13431));
  OR2 OR2_1617(.VSS(VSS),.VDD(VDD),.Y(g30450),.A(g29861),.B(g21859));
  OR2 OR2_1618(.VSS(VSS),.VDD(VDD),.Y(g24653),.A(g2848),.B(g22585));
  OR2 OR2_1619(.VSS(VSS),.VDD(VDD),.Y(g34450),.A(g34281),.B(g18663));
  OR2 OR2_1620(.VSS(VSS),.VDD(VDD),.Y(g13155),.A(g11496),.B(g11546));
  OR2 OR2_1621(.VSS(VSS),.VDD(VDD),.Y(g31793),.A(g28031),.B(g30317));
  OR2 OR2_1622(.VSS(VSS),.VDD(VDD),.Y(g34819),.A(g34741),.B(g34684));
  OR2 OR2_1623(.VSS(VSS),.VDD(VDD),.Y(g34257),.A(g34226),.B(g18674));
  OR2 OR2_1624(.VSS(VSS),.VDD(VDD),.Y(g28209),.A(g27223),.B(g27141));
  OR2 OR2_1625(.VSS(VSS),.VDD(VDD),.Y(g30496),.A(g30231),.B(g21992));
  OR2 OR2_1626(.VSS(VSS),.VDD(VDD),.Y(g8956),.A(g1913),.B(g1932));
  OR2 OR2_1627(.VSS(VSS),.VDD(VDD),.Y(g34979),.A(g34875),.B(g34968));
  OR2 OR2_1628(.VSS(VSS),.VDD(VDD),.Y(g34055),.A(g33909),.B(g33910));
  OR2 OR2_1629(.VSS(VSS),.VDD(VDD),.Y(g33549),.A(g33328),.B(g18337));
  OR2 OR2_1630(.VSS(VSS),.VDD(VDD),.Y(g28208),.A(g27025),.B(g27028));
  OR2 OR2_1631(.VSS(VSS),.VDD(VDD),.Y(g26877),.A(g21658),.B(g25577));
  OR2 OR2_1632(.VSS(VSS),.VDD(VDD),.Y(g34978),.A(g34874),.B(g34967));
  OR2 OR2_1633(.VSS(VSS),.VDD(VDD),.Y(g33548),.A(g33327),.B(g18336));
  OR2 OR2_1634(.VSS(VSS),.VDD(VDD),.Y(g27584),.A(g26165),.B(g24758));
  OR2 OR2_1635(.VSS(VSS),.VDD(VDD),.Y(g25867),.A(g25449),.B(g23884));
  OR2 OR2_1636(.VSS(VSS),.VDD(VDD),.Y(g25894),.A(g24817),.B(g23229));
  OR2 OR2_1637(.VSS(VSS),.VDD(VDD),.Y(g30384),.A(g30101),.B(g18517));
  OR2 OR2_1638(.VSS(VSS),.VDD(VDD),.Y(g31317),.A(g29611),.B(g29626));
  OR2 OR2_1639(.VSS(VSS),.VDD(VDD),.Y(g33317),.A(g29688),.B(g32179));
  OR2 OR2_1640(.VSS(VSS),.VDD(VDD),.Y(g29229),.A(g28532),.B(g18191));
  OR2 OR2_1641(.VSS(VSS),.VDD(VDD),.Y(g25714),.A(g25056),.B(g21965));
  OR2 OR2_1642(.VSS(VSS),.VDD(VDD),.Y(g28614),.A(g27351),.B(g26311));
  OR2 OR2_1643(.VSS(VSS),.VDD(VDD),.Y(g25707),.A(g25041),.B(g18749));
  OR2 OR2_1644(.VSS(VSS),.VDD(VDD),.Y(g25819),.A(g25323),.B(g23836));
  OR2 OR2_1645(.VSS(VSS),.VDD(VDD),.Y(g28607),.A(g27342),.B(g26303));
  OR2 OR2_1646(.VSS(VSS),.VDD(VDD),.Y(g29228),.A(g28426),.B(g18173));
  OR2 OR2_1647(.VSS(VSS),.VDD(VDD),.Y(g25910),.A(g25565),.B(g22142));
  OR2 OR2_1648(.VSS(VSS),.VDD(VDD),.Y(g28320),.A(g27116),.B(g15808));
  OR2 OR2_1649(.VSS(VSS),.VDD(VDD),.Y(g31002),.A(g29362),.B(g28154));
  OR2 OR2_1650(.VSS(VSS),.VDD(VDD),.Y(g28073),.A(g27097),.B(g21875));
  OR2 OR2_1651(.VSS(VSS),.VDD(VDD),.Y(g33002),.A(g32304),.B(g18419));
  OR2 OR2_1652(.VSS(VSS),.VDD(VDD),.Y(g33057),.A(g31968),.B(g22019));
  OR2 OR2_1653(.VSS(VSS),.VDD(VDD),.Y(g34801),.A(g34756),.B(g18588));
  OR2 OR2_1654(.VSS(VSS),.VDD(VDD),.Y(g34735),.A(g34709),.B(g15116));
  OR2 OR2_1655(.VSS(VSS),.VDD(VDD),.Y(g32124),.A(g24488),.B(g30920));
  OR2 OR2_1656(.VSS(VSS),.VDD(VDD),.Y(g29716),.A(g28199),.B(g15856));
  OR2 OR2_1657(.VSS(VSS),.VDD(VDD),.Y(g24200),.A(g22831),.B(g18103));
  OR2 OR2_1658(.VSS(VSS),.VDD(VDD),.Y(g31245),.A(g25964),.B(g29516));
  OR2 OR2_1659(.VSS(VSS),.VDD(VDD),.Y(g34019),.A(g33889),.B(g18506));
  OR2 OR2_1660(.VSS(VSS),.VDD(VDD),.Y(g26917),.A(g26122),.B(g18233));
  OR2 OR2_1661(.VSS(VSS),.VDD(VDD),.Y(g15792),.A(g12920),.B(g10501));
  OR3 OR3_42(.VSS(VSS),.VDD(VDD),.Y(g26866),.A(g20204),.B(g20242),.C(g24363));
  OR2 OR2_1662(.VSS(VSS),.VDD(VDD),.Y(g28565),.A(g27315),.B(g26253));
  OR2 OR2_1663(.VSS(VSS),.VDD(VDD),.Y(g33626),.A(g33374),.B(g18825));
  OR2 OR2_1664(.VSS(VSS),.VDD(VDD),.Y(g33323),.A(g31936),.B(g32442));
  OR2 OR2_1665(.VSS(VSS),.VDD(VDD),.Y(g34695),.A(g34523),.B(g34322));
  OR2 OR2_1666(.VSS(VSS),.VDD(VDD),.Y(g25590),.A(g21694),.B(g24160));
  OR2 OR2_1667(.VSS(VSS),.VDD(VDD),.Y(g34018),.A(g33887),.B(g18505));
  OR2 OR2_1668(.VSS(VSS),.VDD(VDD),.Y(g30526),.A(g30181),.B(g22072));
  OR2 OR2_1669(.VSS(VSS),.VDD(VDD),.Y(g32267),.A(g31208),.B(g31218));
  OR2 OR2_1670(.VSS(VSS),.VDD(VDD),.Y(g32294),.A(g31231),.B(g31232));
  OR2 OR2_1671(.VSS(VSS),.VDD(VDD),.Y(g33298),.A(g32158),.B(g29622));
  OR2 OR2_1672(.VSS(VSS),.VDD(VDD),.Y(g25741),.A(g25178),.B(g22056));
  OR2 OR2_1673(.VSS(VSS),.VDD(VDD),.Y(g28641),.A(g27385),.B(g16591));
  OR2 OR2_1674(.VSS(VSS),.VDD(VDD),.Y(g31775),.A(g30048),.B(g30059));
  OR4 OR4_64(.VSS(VSS),.VDD(VDD),.Y(I30123),.A(g29385),.B(g31376),.C(g30735),.D(g30825));
  OR2 OR2_1675(.VSS(VSS),.VDD(VDD),.Y(g8957),.A(g2338),.B(g2357));
  OR2 OR2_1676(.VSS(VSS),.VDD(VDD),.Y(g24799),.A(g23901),.B(g23921));
  OR2 OR2_1677(.VSS(VSS),.VDD(VDD),.Y(g30402),.A(g29871),.B(g21761));
  OR2 OR2_1678(.VSS(VSS),.VDD(VDD),.Y(g24813),.A(g22685),.B(g19594));
  OR4 OR4_65(.VSS(VSS),.VDD(VDD),.Y(I30751),.A(g32042),.B(g32161),.C(g31943),.D(g31959));
  OR2 OR2_1679(.VSS(VSS),.VDD(VDD),.Y(g30457),.A(g29369),.B(g21885));
  OR2 OR2_1680(.VSS(VSS),.VDD(VDD),.Y(g34402),.A(g34179),.B(g25084));
  OR2 OR2_1681(.VSS(VSS),.VDD(VDD),.Y(g34457),.A(g34394),.B(g18670));
  OR2 OR2_1682(.VSS(VSS),.VDD(VDD),.Y(g26923),.A(g25923),.B(g18290));
  OR2 OR2_1683(.VSS(VSS),.VDD(VDD),.Y(g32219),.A(g31131),.B(g29620));
  OR2 OR2_1684(.VSS(VSS),.VDD(VDD),.Y(g33232),.A(g32034),.B(g30936));
  OR2 OR2_1685(.VSS(VSS),.VDD(VDD),.Y(g25735),.A(g25077),.B(g18783));
  OR2 OR2_1686(.VSS(VSS),.VDD(VDD),.Y(g25877),.A(g25502),.B(g23919));
  OR2 OR2_1687(.VSS(VSS),.VDD(VDD),.Y(g28635),.A(g27375),.B(g16537));
  OR2 OR2_1688(.VSS(VSS),.VDD(VDD),.Y(g32218),.A(g31130),.B(g29619));
  OR2 OR2_1689(.VSS(VSS),.VDD(VDD),.Y(g27135),.A(g24387),.B(g25803));
  OR2 OR2_1690(.VSS(VSS),.VDD(VDD),.Y(g33995),.A(g33848),.B(g18425));
  OR2 OR2_1691(.VSS(VSS),.VDD(VDD),.Y(g34001),.A(g33844),.B(g18450));
  OR2 OR2_1692(.VSS(VSS),.VDD(VDD),.Y(g33261),.A(g32111),.B(g29525));
  OR2 OR2_1693(.VSS(VSS),.VDD(VDD),.Y(g25695),.A(g24998),.B(g21914));
  OR2 OR2_1694(.VSS(VSS),.VDD(VDD),.Y(g31880),.A(g31280),.B(g21774));
  OR2 OR2_1695(.VSS(VSS),.VDD(VDD),.Y(g30597),.A(g13564),.B(g29693));
  OR2 OR2_1696(.VSS(VSS),.VDD(VDD),.Y(g34256),.A(g34173),.B(g24303));
  OR2 OR2_1697(.VSS(VSS),.VDD(VDD),.Y(g29802),.A(g28243),.B(g22871));
  OR2 OR2_1698(.VSS(VSS),.VDD(VDD),.Y(g34280),.A(g26833),.B(g34213));
  OR2 OR2_1699(.VSS(VSS),.VDD(VDD),.Y(g29730),.A(g28150),.B(g28141));
  OR2 OR2_1700(.VSS(VSS),.VDD(VDD),.Y(g30300),.A(g28246),.B(g27252));
  OR2 OR2_1701(.VSS(VSS),.VDD(VDD),.Y(g29793),.A(g28237),.B(g27247));
  OR2 OR2_1702(.VSS(VSS),.VDD(VDD),.Y(g34624),.A(g34509),.B(g18592));
  OR2 OR2_1703(.VSS(VSS),.VDD(VDD),.Y(g34300),.A(g26864),.B(g34230));
  OR2 OR2_1704(.VSS(VSS),.VDD(VDD),.Y(g15125),.A(g10363),.B(g13605));
  OR2 OR2_1705(.VSS(VSS),.VDD(VDD),.Y(g26876),.A(g21655),.B(g25576));
  OR2 OR2_1706(.VSS(VSS),.VDD(VDD),.Y(g26885),.A(g26541),.B(g24191));
  OR3 OR3_43(.VSS(VSS),.VDD(VDD),.Y(g23751),.A(g21415),.B(g21402),.C(I22880));
  OR2 OR2_1707(.VSS(VSS),.VDD(VDD),.Y(g25917),.A(g22524),.B(g24518));
  OR2 OR2_1708(.VSS(VSS),.VDD(VDD),.Y(g32277),.A(g31211),.B(g29733));
  OR2 OR2_1709(.VSS(VSS),.VDD(VDD),.Y(g24214),.A(g23471),.B(g18195));
  OR2 OR2_1710(.VSS(VSS),.VDD(VDD),.Y(g31316),.A(g29609),.B(g29624));
  OR2 OR2_1711(.VSS(VSS),.VDD(VDD),.Y(g33316),.A(g29685),.B(g32178));
  OR2 OR2_1712(.VSS(VSS),.VDD(VDD),.Y(g22634),.A(g18934),.B(g15590));
  OR2 OR2_1713(.VSS(VSS),.VDD(VDD),.Y(g24207),.A(g23396),.B(g18119));
  OR2 OR2_1714(.VSS(VSS),.VDD(VDD),.Y(g22872),.A(g19372),.B(g19383));
  OR4 OR4_66(.VSS(VSS),.VDD(VDD),.Y(I29985),.A(g29385),.B(g31376),.C(g30735),.D(g30825));
  OR3 OR3_44(.VSS(VSS),.VDD(VDD),.Y(I22958),.A(g21603),.B(g21386),.C(g21365));
  OR2 OR2_1715(.VSS(VSS),.VDD(VDD),.Y(g34231),.A(g33898),.B(g33902));
  OR2 OR2_1716(.VSS(VSS),.VDD(VDD),.Y(g29504),.A(g28143),.B(g25875));
  OR2 OR2_1717(.VSS(VSS),.VDD(VDD),.Y(g25706),.A(g25030),.B(g18748));
  OR2 OR2_1718(.VSS(VSS),.VDD(VDD),.Y(g25597),.A(g24892),.B(g21719));
  OR2 OR2_1719(.VSS(VSS),.VDD(VDD),.Y(g32037),.A(g30566),.B(g29329));
  OR2 OR2_1720(.VSS(VSS),.VDD(VDD),.Y(g33989),.A(g33870),.B(g18398));
  OR2 OR2_1721(.VSS(VSS),.VDD(VDD),.Y(g33056),.A(g32327),.B(g22004));
  OR2 OR2_1722(.VSS(VSS),.VDD(VDD),.Y(g13570),.A(g9223),.B(g11130));
  OR2 OR2_1723(.VSS(VSS),.VDD(VDD),.Y(g25689),.A(g24849),.B(g21888));
  OR2 OR2_1724(.VSS(VSS),.VDD(VDD),.Y(g13914),.A(g8643),.B(g11380));
  OR2 OR2_1725(.VSS(VSS),.VDD(VDD),.Y(g33611),.A(g33243),.B(g18632));
  OR2 OR2_1726(.VSS(VSS),.VDD(VDD),.Y(g31924),.A(g31486),.B(g22049));
  OR2 OR2_1727(.VSS(VSS),.VDD(VDD),.Y(g32984),.A(g31934),.B(g18264));
  OR2 OR2_1728(.VSS(VSS),.VDD(VDD),.Y(g33988),.A(g33861),.B(g18397));
  OR2 OR2_1729(.VSS(VSS),.VDD(VDD),.Y(g25688),.A(g24812),.B(g21887));
  OR2 OR2_1730(.VSS(VSS),.VDD(VDD),.Y(g28750),.A(g27525),.B(g16765));
  OR2 OR2_1731(.VSS(VSS),.VDD(VDD),.Y(g25624),.A(g24408),.B(g18224));
  OR2 OR2_1732(.VSS(VSS),.VDD(VDD),.Y(g26916),.A(g25916),.B(g18232));
  OR2 OR2_1733(.VSS(VSS),.VDD(VDD),.Y(g30511),.A(g30180),.B(g22032));
  OR2 OR2_1734(.VSS(VSS),.VDD(VDD),.Y(g20241),.A(g16233),.B(g13541));
  OR2 OR2_1735(.VSS(VSS),.VDD(VDD),.Y(g32352),.A(g29852),.B(g31282));
  OR4 OR4_67(.VSS(VSS),.VDD(VDD),.Y(I30746),.A(g32047),.B(g31985),.C(g31991),.D(g32309));
  OR2 OR2_1736(.VSS(VSS),.VDD(VDD),.Y(g24241),.A(g22920),.B(g18252));
  OR2 OR2_1737(.VSS(VSS),.VDD(VDD),.Y(g33271),.A(g32120),.B(g29549));
  OR2 OR2_1738(.VSS(VSS),.VDD(VDD),.Y(g27972),.A(g26131),.B(g26105));
  OR2 OR2_1739(.VSS(VSS),.VDD(VDD),.Y(g32155),.A(g30935),.B(g29475));
  OR2 OR2_1740(.VSS(VSS),.VDD(VDD),.Y(g15017),.A(g10776),.B(g8703));
  OR2 OR2_1741(.VSS(VSS),.VDD(VDD),.Y(g28091),.A(g27665),.B(g21913));
  OR2 OR2_1742(.VSS(VSS),.VDD(VDD),.Y(g32266),.A(g30604),.B(g29354));
  OR2 OR2_1743(.VSS(VSS),.VDD(VDD),.Y(g29245),.A(g28676),.B(g18384));
  OR2 OR2_1744(.VSS(VSS),.VDD(VDD),.Y(g26721),.A(g10776),.B(g24444));
  OR2 OR2_1745(.VSS(VSS),.VDD(VDD),.Y(g29299),.A(g28587),.B(g18794));
  OR2 OR2_1746(.VSS(VSS),.VDD(VDD),.Y(g33031),.A(g32315),.B(g21841));
  OR2 OR2_1747(.VSS(VSS),.VDD(VDD),.Y(g30456),.A(g29378),.B(g21869));
  OR2 OR2_1748(.VSS(VSS),.VDD(VDD),.Y(g34456),.A(g34395),.B(g18669));
  OR2 OR2_1749(.VSS(VSS),.VDD(VDD),.Y(g29298),.A(g28571),.B(g18793));
  OR2 OR2_1750(.VSS(VSS),.VDD(VDD),.Y(g24235),.A(g22632),.B(g18238));
  OR2 OR2_1751(.VSS(VSS),.VDD(VDD),.Y(g13941),.A(g11019),.B(g11023));
  OR2 OR2_1752(.VSS(VSS),.VDD(VDD),.Y(g31887),.A(g31292),.B(g21820));
  OR2 OR2_1753(.VSS(VSS),.VDD(VDD),.Y(g28390),.A(g27207),.B(g15861));
  OR2 OR2_1754(.VSS(VSS),.VDD(VDD),.Y(g30480),.A(g29321),.B(g21972));
  OR2 OR2_1755(.VSS(VSS),.VDD(VDD),.Y(g30916),.A(g13853),.B(g29799));
  OR2 OR2_1756(.VSS(VSS),.VDD(VDD),.Y(g29775),.A(g25966),.B(g28232));
  OR4 OR4_68(.VSS(VSS),.VDD(VDD),.Y(I26523),.A(g20720),.B(g20857),.C(g20998),.D(g21143));
  OR2 OR2_1757(.VSS(VSS),.VDD(VDD),.Y(g25885),.A(g25522),.B(g23957));
  OR2 OR2_1758(.VSS(VSS),.VDD(VDD),.Y(g30550),.A(g30226),.B(g22121));
  OR2 OR2_1759(.VSS(VSS),.VDD(VDD),.Y(g30314),.A(g28268),.B(g27266));
  OR2 OR2_1760(.VSS(VSS),.VDD(VDD),.Y(g23615),.A(g20109),.B(g20131));
  OR2 OR2_1761(.VSS(VSS),.VDD(VDD),.Y(g30287),.A(g28653),.B(g27677));
  OR2 OR2_1762(.VSS(VSS),.VDD(VDD),.Y(g34314),.A(g25831),.B(g34061));
  OR2 OR2_1763(.VSS(VSS),.VDD(VDD),.Y(g30307),.A(g28256),.B(g27260));
  OR2 OR2_1764(.VSS(VSS),.VDD(VDD),.Y(g33393),.A(g32286),.B(g29984));
  OR2 OR2_1765(.VSS(VSS),.VDD(VDD),.Y(g23720),.A(g20165),.B(g16801));
  OR4 OR4_69(.VSS(VSS),.VDD(VDD),.Y(I12902),.A(g4235),.B(g4232),.C(g4229),.D(g4226));
  OR2 OR2_1766(.VSS(VSS),.VDD(VDD),.Y(g25763),.A(g25113),.B(g18817));
  OR2 OR2_1767(.VSS(VSS),.VDD(VDD),.Y(g29232),.A(g28183),.B(g18231));
  OR2 OR2_1768(.VSS(VSS),.VDD(VDD),.Y(g31764),.A(g30015),.B(g30032));
  OR2 OR2_1769(.VSS(VSS),.VDD(VDD),.Y(g23275),.A(g19680),.B(g16160));
  OR2 OR2_1770(.VSS(VSS),.VDD(VDD),.Y(g34721),.A(g34696),.B(g18135));
  OR2 OR2_1771(.VSS(VSS),.VDD(VDD),.Y(g31869),.A(g30592),.B(g18221));
  OR4 OR4_70(.VSS(VSS),.VDD(VDD),.Y(I30193),.A(g31070),.B(g30614),.C(g30673),.D(g31528));
  OR2 OR2_1772(.VSS(VSS),.VDD(VDD),.Y(g30431),.A(g29875),.B(g21815));
  OR2 OR2_1773(.VSS(VSS),.VDD(VDD),.Y(g33960),.A(g33759),.B(g21701));
  OR2 OR2_1774(.VSS(VSS),.VDD(VDD),.Y(g25660),.A(g24726),.B(g21785));
  OR2 OR2_1775(.VSS(VSS),.VDD(VDD),.Y(g29261),.A(g28247),.B(g18605));
  OR2 OR2_1776(.VSS(VSS),.VDD(VDD),.Y(g31868),.A(g30600),.B(g18204));
  OR2 OR2_1777(.VSS(VSS),.VDD(VDD),.Y(g26335),.A(g1526),.B(g24609));
  OR2 OR2_1778(.VSS(VSS),.VDD(VDD),.Y(g19572),.A(g17133),.B(g14193));
  OR2 OR2_1779(.VSS(VSS),.VDD(VDD),.Y(g22152),.A(g21188),.B(g17469));
  OR2 OR2_1780(.VSS(VSS),.VDD(VDD),.Y(g26930),.A(g26799),.B(g18544));
  OR2 OR2_1781(.VSS(VSS),.VDD(VDD),.Y(g34269),.A(g34083),.B(g18732));
  OR2 OR2_1782(.VSS(VSS),.VDD(VDD),.Y(g30341),.A(g29380),.B(g18246));
  OR2 OR2_1783(.VSS(VSS),.VDD(VDD),.Y(g26694),.A(g24444),.B(g10704));
  OR2 OR2_1784(.VSS(VSS),.VDD(VDD),.Y(g26965),.A(g26336),.B(g24317));
  OR2 OR2_1785(.VSS(VSS),.VDD(VDD),.Y(g33709),.A(g32414),.B(g33441));
  OR2 OR2_1786(.VSS(VSS),.VDD(VDD),.Y(g34268),.A(g34082),.B(g18730));
  OR2 OR2_1787(.VSS(VSS),.VDD(VDD),.Y(g31259),.A(g25992),.B(g29554));
  OR2 OR2_1788(.VSS(VSS),.VDD(VDD),.Y(g32285),.A(g31222),.B(g29740));
  OR2 OR2_1789(.VSS(VSS),.VDD(VDD),.Y(g33259),.A(g32109),.B(g29521));
  OR2 OR2_1790(.VSS(VSS),.VDD(VDD),.Y(g28536),.A(g27293),.B(g26205));
  OR4 OR4_71(.VSS(VSS),.VDD(VDD),.Y(I30727),.A(g31759),.B(g32196),.C(g31933),.D(g31941));
  OR2 OR2_1791(.VSS(VSS),.VDD(VDD),.Y(g31258),.A(g25991),.B(g29550));
  OR2 OR2_1792(.VSS(VSS),.VDD(VDD),.Y(g24206),.A(g23386),.B(g18110));
  OR2 OR2_1793(.VSS(VSS),.VDD(VDD),.Y(g13728),.A(g6804),.B(g12527));
  OR2 OR2_1794(.VSS(VSS),.VDD(VDD),.Y(g28702),.A(g27457),.B(g16670));
  OR2 OR2_1795(.VSS(VSS),.VDD(VDD),.Y(g30734),.A(g13808),.B(g29774));
  OR3 OR3_45(.VSS(VSS),.VDD(VDD),.Y(I22298),.A(g20371),.B(g20161),.C(g20151));
  OR2 OR2_1796(.VSS(VSS),.VDD(VDD),.Y(g30335),.A(g29746),.B(g18174));
  OR2 OR2_1797(.VSS(VSS),.VDD(VDD),.Y(g34734),.A(g34681),.B(g18652));
  OR2 OR2_1798(.VSS(VSS),.VDD(VDD),.Y(g25721),.A(g25057),.B(g18766));
  OR2 OR2_1799(.VSS(VSS),.VDD(VDD),.Y(g28621),.A(g27359),.B(g16518));
  OR2 OR2_1800(.VSS(VSS),.VDD(VDD),.Y(g25596),.A(g24865),.B(g21718));
  OR4 OR4_72(.VSS(VSS),.VDD(VDD),.Y(I31853),.A(g33488),.B(g33489),.C(g33490),.D(g33491));
  OR2 OR2_1801(.VSS(VSS),.VDD(VDD),.Y(g33043),.A(g32195),.B(g24325));
  OR2 OR2_1802(.VSS(VSS),.VDD(VDD),.Y(g31244),.A(g25963),.B(g29515));
  OR2 OR2_1803(.VSS(VSS),.VDD(VDD),.Y(g20082),.A(g16026),.B(g13321));
  OR2 OR2_1804(.VSS(VSS),.VDD(VDD),.Y(g28564),.A(g27314),.B(g26252));
  OR2 OR2_1805(.VSS(VSS),.VDD(VDD),.Y(g23193),.A(g19556),.B(g15937));
  OR4 OR4_73(.VSS(VSS),.VDD(VDD),.Y(I23756),.A(g23457),.B(g23480),.C(g23494),.D(g23511));
  OR2 OR2_1806(.VSS(VSS),.VDD(VDD),.Y(g26278),.A(g24545),.B(g24549));
  OR2 OR2_1807(.VSS(VSS),.VDD(VDD),.Y(g33069),.A(g32009),.B(g22113));
  OR2 OR2_1808(.VSS(VSS),.VDD(VDD),.Y(g33602),.A(g33425),.B(g18511));
  OR2 OR2_1809(.VSS(VSS),.VDD(VDD),.Y(g25942),.A(g24422),.B(g22298));
  OR2 OR2_1810(.VSS(VSS),.VDD(VDD),.Y(g31774),.A(g30046),.B(g30057));
  OR2 OR2_1811(.VSS(VSS),.VDD(VDD),.Y(g7834),.A(g2886),.B(g2946));
  OR2 OR2_1812(.VSS(VSS),.VDD(VDD),.Y(g30487),.A(g30187),.B(g21983));
  OR2 OR2_1813(.VSS(VSS),.VDD(VDD),.Y(g31375),.A(g29628),.B(g28339));
  OR2 OR2_1814(.VSS(VSS),.VDD(VDD),.Y(g33068),.A(g31994),.B(g22112));
  OR3 OR3_46(.VSS(VSS),.VDD(VDD),.Y(g33955),.A(g33505),.B(I31858),.C(I31859));
  OR2 OR2_1815(.VSS(VSS),.VDD(VDD),.Y(g24345),.A(g23606),.B(g18788));
  OR2 OR2_1816(.VSS(VSS),.VDD(VDD),.Y(g25655),.A(g24645),.B(g18607));
  OR2 OR2_1817(.VSS(VSS),.VDD(VDD),.Y(g31879),.A(g31475),.B(g21745));
  OR2 OR2_1818(.VSS(VSS),.VDD(VDD),.Y(g30502),.A(g30232),.B(g22023));
  OR2 OR2_1819(.VSS(VSS),.VDD(VDD),.Y(g28062),.A(g27288),.B(g21746));
  OR2 OR2_1820(.VSS(VSS),.VDD(VDD),.Y(g30557),.A(g30247),.B(g22128));
  OR2 OR2_1821(.VSS(VSS),.VDD(VDD),.Y(g33970),.A(g33868),.B(g18322));
  OR2 OR2_1822(.VSS(VSS),.VDD(VDD),.Y(g34619),.A(g34528),.B(g18581));
  OR3 OR3_47(.VSS(VSS),.VDD(VDD),.Y(I22880),.A(g21509),.B(g21356),.C(g21351));
  OR2 OR2_1823(.VSS(VSS),.VDD(VDD),.Y(g25670),.A(g24967),.B(g18626));
  OR2 OR2_1824(.VSS(VSS),.VDD(VDD),.Y(g29271),.A(g28333),.B(g18637));
  OR2 OR2_1825(.VSS(VSS),.VDD(VDD),.Y(g31878),.A(g31015),.B(g21733));
  OR4 OR4_74(.VSS(VSS),.VDD(VDD),.Y(I31864),.A(g33510),.B(g33511),.C(g33512),.D(g33513));
  OR2 OR2_1826(.VSS(VSS),.VDD(VDD),.Y(g30443),.A(g29808),.B(g21852));
  OR2 OR2_1827(.VSS(VSS),.VDD(VDD),.Y(g34618),.A(g34527),.B(g18580));
  OR2 OR2_1828(.VSS(VSS),.VDD(VDD),.Y(g24398),.A(g23801),.B(g21296));
  OR2 OR2_1829(.VSS(VSS),.VDD(VDD),.Y(g30279),.A(g28637),.B(g27668));
  OR2 OR2_1830(.VSS(VSS),.VDD(VDD),.Y(g34443),.A(g34385),.B(g18545));
  OR2 OR2_1831(.VSS(VSS),.VDD(VDD),.Y(g25734),.A(g25058),.B(g18782));
  OR2 OR2_1832(.VSS(VSS),.VDD(VDD),.Y(g28634),.A(g27374),.B(g16536));
  OR2 OR2_1833(.VSS(VSS),.VDD(VDD),.Y(g28851),.A(g27558),.B(g16870));
  OR2 OR2_1834(.VSS(VSS),.VDD(VDD),.Y(g31886),.A(g31481),.B(g21791));
  OR2 OR2_1835(.VSS(VSS),.VDD(VDD),.Y(g29753),.A(g28213),.B(g22720));
  OR4 OR4_75(.VSS(VSS),.VDD(VDD),.Y(g25839),.A(g25507),.B(g25485),.C(g25459),.D(g25420));
  OR2 OR2_1836(.VSS(VSS),.VDD(VDD),.Y(g34278),.A(g26829),.B(g34212));
  OR2 OR2_1837(.VSS(VSS),.VDD(VDD),.Y(g30469),.A(g30153),.B(g21940));
  OR2 OR2_1838(.VSS(VSS),.VDD(VDD),.Y(g33967),.A(g33842),.B(g18319));
  OR2 OR2_1839(.VSS(VSS),.VDD(VDD),.Y(g33994),.A(g33841),.B(g18424));
  OR2 OR2_1840(.VSS(VSS),.VDD(VDD),.Y(g27506),.A(g26021),.B(g24639));
  OR2 OR2_1841(.VSS(VSS),.VDD(VDD),.Y(g30286),.A(g28191),.B(g28186));
  OR2 OR2_1842(.VSS(VSS),.VDD(VDD),.Y(g25694),.A(g24638),.B(g18738));
  OR2 OR2_1843(.VSS(VSS),.VDD(VDD),.Y(g25667),.A(g24682),.B(g18619));
  OR2 OR2_1844(.VSS(VSS),.VDD(VDD),.Y(g24263),.A(g23497),.B(g18529));
  OR2 OR2_1845(.VSS(VSS),.VDD(VDD),.Y(g34286),.A(g26842),.B(g34216));
  OR2 OR2_1846(.VSS(VSS),.VDD(VDD),.Y(g30468),.A(g30238),.B(g21939));
  OR2 OR2_1847(.VSS(VSS),.VDD(VDD),.Y(g34468),.A(g34342),.B(g18718));
  OR2 OR2_1848(.VSS(VSS),.VDD(VDD),.Y(g34039),.A(g33743),.B(g18736));
  OR2 OR2_1849(.VSS(VSS),.VDD(VDD),.Y(g34306),.A(g25782),.B(g34054));
  OR4 OR4_76(.VSS(VSS),.VDD(VDD),.Y(g29529),.A(g28303),.B(g28293),.C(g28283),.D(g28267));
  OR2 OR2_1850(.VSS(VSS),.VDD(VDD),.Y(g22640),.A(g18951),.B(g15613));
  OR2 OR2_1851(.VSS(VSS),.VDD(VDD),.Y(g34038),.A(g33731),.B(g18735));
  OR2 OR2_1852(.VSS(VSS),.VDD(VDD),.Y(g31919),.A(g31758),.B(g22044));
  OR2 OR2_1853(.VSS(VSS),.VDD(VDD),.Y(g32454),.A(g30322),.B(g31795));
  OR2 OR2_1854(.VSS(VSS),.VDD(VDD),.Y(g25619),.A(g24961),.B(g18193));
  OR2 OR2_1855(.VSS(VSS),.VDD(VDD),.Y(g15124),.A(g13605),.B(g4581));
  OR2 OR2_1856(.VSS(VSS),.VDD(VDD),.Y(g26884),.A(g26511),.B(g24190));
  OR2 OR2_1857(.VSS(VSS),.VDD(VDD),.Y(g28574),.A(g27324),.B(g26270));
  OR2 OR2_1858(.VSS(VSS),.VDD(VDD),.Y(g31918),.A(g31786),.B(g22015));
  OR2 OR2_1859(.VSS(VSS),.VDD(VDD),.Y(g28047),.A(g27676),.B(g18160));
  OR2 OR2_1860(.VSS(VSS),.VDD(VDD),.Y(g33010),.A(g32301),.B(g18473));
  OR2 OR2_1861(.VSS(VSS),.VDD(VDD),.Y(g34601),.A(g34488),.B(g18211));
  OR2 OR2_1862(.VSS(VSS),.VDD(VDD),.Y(g29764),.A(g28219),.B(g28226));
  OR2 OR2_1863(.VSS(VSS),.VDD(VDD),.Y(g25618),.A(g25491),.B(g18192));
  OR2 OR2_1864(.VSS(VSS),.VDD(VDD),.Y(g34975),.A(g34871),.B(g34964));
  OR2 OR2_1865(.VSS(VSS),.VDD(VDD),.Y(g24500),.A(g24011),.B(g21605));
  OR2 OR2_1866(.VSS(VSS),.VDD(VDD),.Y(g33545),.A(g33399),.B(g18324));
  OR2 OR2_1867(.VSS(VSS),.VDD(VDD),.Y(g9013),.A(g2472),.B(g2491));
  OR2 OR2_1868(.VSS(VSS),.VDD(VDD),.Y(g26363),.A(g2965),.B(g24965));
  OR2 OR2_1869(.VSS(VSS),.VDD(VDD),.Y(g33599),.A(g33087),.B(g18500));
  OR2 OR2_1870(.VSS(VSS),.VDD(VDD),.Y(g32239),.A(g30595),.B(g29350));
  OR2 OR2_1871(.VSS(VSS),.VDD(VDD),.Y(g28051),.A(g27699),.B(g18166));
  OR2 OR2_1872(.VSS(VSS),.VDD(VDD),.Y(g27240),.A(g25883),.B(g24467));
  OR2 OR2_1873(.VSS(VSS),.VDD(VDD),.Y(g28072),.A(g27086),.B(g21874));
  OR2 OR2_1874(.VSS(VSS),.VDD(VDD),.Y(g33598),.A(g33364),.B(g18496));
  OR2 OR2_1875(.VSS(VSS),.VDD(VDD),.Y(g32238),.A(g30594),.B(g29349));
  OR4 OR4_77(.VSS(VSS),.VDD(VDD),.Y(I29352),.A(g29322),.B(g29315),.C(g30315),.D(g30308));
  OR2 OR2_1876(.VSS(VSS),.VDD(VDD),.Y(g28592),.A(g27333),.B(g26288));
  OR4 OR4_78(.VSS(VSS),.VDD(VDD),.Y(I31874),.A(g33528),.B(g33529),.C(g33530),.D(g33531));
  OR2 OR2_1877(.VSS(VSS),.VDD(VDD),.Y(g34791),.A(g34771),.B(g18184));
  OR2 OR2_1878(.VSS(VSS),.VDD(VDD),.Y(g22662),.A(g19069),.B(g15679));
  OR2 OR2_1879(.VSS(VSS),.VDD(VDD),.Y(g34884),.A(g34858),.B(g21666));
  OR2 OR2_1880(.VSS(VSS),.VDD(VDD),.Y(g29259),.A(g28304),.B(g18603));
  OR2 OR2_1881(.VSS(VSS),.VDD(VDD),.Y(g29225),.A(g28451),.B(g18158));
  OR2 OR2_1882(.VSS(VSS),.VDD(VDD),.Y(g30410),.A(g29857),.B(g21769));
  OR2 OR2_1883(.VSS(VSS),.VDD(VDD),.Y(g31322),.A(g26128),.B(g29635));
  OR2 OR2_1884(.VSS(VSS),.VDD(VDD),.Y(g14062),.A(g11047),.B(g11116));
  OR2 OR2_1885(.VSS(VSS),.VDD(VDD),.Y(g34168),.A(g33787),.B(g19784));
  OR2 OR2_1886(.VSS(VSS),.VDD(VDD),.Y(g27563),.A(g26104),.B(g24704));
  OR2 OR2_1887(.VSS(VSS),.VDD(VDD),.Y(g29258),.A(g28238),.B(g18601));
  OR2 OR2_1888(.VSS(VSS),.VDD(VDD),.Y(g31901),.A(g31516),.B(g21909));
  OR2 OR2_1889(.VSS(VSS),.VDD(VDD),.Y(g33159),.A(g32016),.B(g30730));
  OR2 OR2_1890(.VSS(VSS),.VDD(VDD),.Y(g30479),.A(g29320),.B(g21950));
  OR2 OR2_1891(.VSS(VSS),.VDD(VDD),.Y(g33977),.A(g33876),.B(g18348));
  OR2 OR2_1892(.VSS(VSS),.VDD(VDD),.Y(g30363),.A(g30121),.B(g18407));
  OR2 OR2_1893(.VSS(VSS),.VDD(VDD),.Y(g25601),.A(g24660),.B(g18112));
  OR2 OR2_1894(.VSS(VSS),.VDD(VDD),.Y(g12981),.A(g12219),.B(g9967));
  OR2 OR2_1895(.VSS(VSS),.VDD(VDD),.Y(g24273),.A(g23166),.B(g18630));
  OR2 OR2_1896(.VSS(VSS),.VDD(VDD),.Y(g25677),.A(g24684),.B(g21834));
  OR2 OR2_1897(.VSS(VSS),.VDD(VDD),.Y(g31783),.A(I29351),.B(I29352));
  OR2 OR2_1898(.VSS(VSS),.VDD(VDD),.Y(g23209),.A(g19585),.B(g19601));
  OR2 OR2_1899(.VSS(VSS),.VDD(VDD),.Y(g30478),.A(g30248),.B(g21949));
  OR2 OR2_1900(.VSS(VSS),.VDD(VDD),.Y(g34015),.A(g33858),.B(g18502));
  OR2 OR2_1901(.VSS(VSS),.VDD(VDD),.Y(g29244),.A(g28692),.B(g18380));
  OR2 OR2_1902(.VSS(VSS),.VDD(VDD),.Y(g33561),.A(g33408),.B(g18376));
  OR2 OR2_1903(.VSS(VSS),.VDD(VDD),.Y(g30486),.A(g30177),.B(g21982));
  OR2 OR2_1904(.VSS(VSS),.VDD(VDD),.Y(g31295),.A(g26090),.B(g29598));
  OR2 OR2_1905(.VSS(VSS),.VDD(VDD),.Y(g26922),.A(g25902),.B(g18288));
  OR2 OR2_1906(.VSS(VSS),.VDD(VDD),.Y(g28731),.A(g27504),.B(g16733));
  OR2 OR2_1907(.VSS(VSS),.VDD(VDD),.Y(g33295),.A(g32153),.B(g29605));
  OR2 OR2_1908(.VSS(VSS),.VDD(VDD),.Y(g31144),.A(g29477),.B(g28193));
  OR2 OR2_1909(.VSS(VSS),.VDD(VDD),.Y(g25937),.A(g24406),.B(g22216));
  OR2 OR2_1910(.VSS(VSS),.VDD(VDD),.Y(g30556),.A(g30236),.B(g22127));
  OR2 OR2_1911(.VSS(VSS),.VDD(VDD),.Y(g24234),.A(g22622),.B(g18237));
  OR2 OR2_1912(.VSS(VSS),.VDD(VDD),.Y(g13973),.A(g11024),.B(g11028));
  OR2 OR2_1913(.VSS(VSS),.VDD(VDD),.Y(g29068),.A(g27628),.B(g17119));
  OR4 OR4_79(.VSS(VSS),.VDD(VDD),.Y(g25791),.A(g25411),.B(g25371),.C(g25328),.D(g25290));
  OR2 OR2_1914(.VSS(VSS),.VDD(VDD),.Y(g28691),.A(g27437),.B(g16642));
  OR2 OR2_1915(.VSS(VSS),.VDD(VDD),.Y(g29879),.A(g28289),.B(g26096));
  OR2 OR2_1916(.VSS(VSS),.VDD(VDD),.Y(g26953),.A(g26486),.B(g24291));
  OR2 OR2_1917(.VSS(VSS),.VDD(VDD),.Y(g28405),.A(g27216),.B(g15875));
  OR2 OR2_1918(.VSS(VSS),.VDD(VDD),.Y(g33966),.A(g33837),.B(g18318));
  OR2 OR2_1919(.VSS(VSS),.VDD(VDD),.Y(g25666),.A(g24788),.B(g21793));
  OR2 OR2_1920(.VSS(VSS),.VDD(VDD),.Y(g33017),.A(g32292),.B(g18510));
  OR2 OR2_1921(.VSS(VSS),.VDD(VDD),.Y(g26800),.A(g24922),.B(g24929));
  OR2 OR2_1922(.VSS(VSS),.VDD(VDD),.Y(g34321),.A(g25866),.B(g34065));
  OR2 OR2_1923(.VSS(VSS),.VDD(VDD),.Y(g30531),.A(g30274),.B(g22077));
  OR2 OR2_1924(.VSS(VSS),.VDD(VDD),.Y(g23346),.A(g19736),.B(g16204));
  OR2 OR2_1925(.VSS(VSS),.VDD(VDD),.Y(g29792),.A(g28235),.B(g28244));
  OR2 OR2_1926(.VSS(VSS),.VDD(VDD),.Y(g12832),.A(g10347),.B(g10348));
  OR2 OR2_1927(.VSS(VSS),.VDD(VDD),.Y(g13761),.A(g490),.B(g12527));
  OR2 OR2_1928(.VSS(VSS),.VDD(VDD),.Y(g16022),.A(g13048),.B(g10707));
  OR2 OR2_1929(.VSS(VSS),.VDD(VDD),.Y(g26334),.A(g1171),.B(g24591));
  OR2 OR2_1930(.VSS(VSS),.VDD(VDD),.Y(g28046),.A(g27667),.B(g18157));
  OR2 OR2_1931(.VSS(VSS),.VDD(VDD),.Y(g32349),.A(g29840),.B(g31275));
  OR2 OR2_1932(.VSS(VSS),.VDD(VDD),.Y(g31289),.A(g29580),.B(g29591));
  OR2 OR2_1933(.VSS(VSS),.VDD(VDD),.Y(g30373),.A(g30111),.B(g18461));
  OR2 OR2_1934(.VSS(VSS),.VDD(VDD),.Y(g33289),.A(g32148),.B(g29588));
  OR2 OR2_1935(.VSS(VSS),.VDD(VDD),.Y(g22331),.A(g21405),.B(g17809));
  OR2 OR2_1936(.VSS(VSS),.VDD(VDD),.Y(g26964),.A(g26259),.B(g24316));
  OR2 OR2_1937(.VSS(VSS),.VDD(VDD),.Y(g34373),.A(g26292),.B(g34138));
  OR2 OR2_1938(.VSS(VSS),.VDD(VDD),.Y(g33023),.A(g32313),.B(g21751));
  OR2 OR2_1939(.VSS(VSS),.VDD(VDD),.Y(g31288),.A(g2955),.B(g29914));
  OR2 OR2_1940(.VSS(VSS),.VDD(VDD),.Y(g23153),.A(g19521),.B(g15876));
  OR2 OR2_1941(.VSS(VSS),.VDD(VDD),.Y(g33288),.A(g32147),.B(g29587));
  OR2 OR2_1942(.VSS(VSS),.VDD(VDD),.Y(g31308),.A(g26101),.B(g29614));
  OR2 OR2_1943(.VSS(VSS),.VDD(VDD),.Y(g33571),.A(g33367),.B(g18409));
  OR2 OR2_1944(.VSS(VSS),.VDD(VDD),.Y(g30417),.A(g29874),.B(g21801));
  OR2 OR2_1945(.VSS(VSS),.VDD(VDD),.Y(g34800),.A(g34752),.B(g18586));
  OR2 OR2_1946(.VSS(VSS),.VDD(VDD),.Y(g34417),.A(g27678),.B(g34196));
  OR2 OR2_1947(.VSS(VSS),.VDD(VDD),.Y(g28357),.A(g27148),.B(g15836));
  OR2 OR2_1948(.VSS(VSS),.VDD(VDD),.Y(g30334),.A(g29837),.B(g18143));
  OR2 OR2_1949(.VSS(VSS),.VDD(VDD),.Y(g28105),.A(g27997),.B(g22135));
  OR2 OR2_1950(.VSS(VSS),.VDD(VDD),.Y(g28743),.A(g27517),.B(g16758));
  OR2 OR2_1951(.VSS(VSS),.VDD(VDD),.Y(g29078),.A(g27633),.B(g26572));
  OR2 OR2_1952(.VSS(VSS),.VDD(VDD),.Y(g26909),.A(g26543),.B(g24227));
  OR3 OR3_48(.VSS(VSS),.VDD(VDD),.Y(I18385),.A(g14413),.B(g14391),.C(g14360));
  OR2 OR2_1953(.VSS(VSS),.VDD(VDD),.Y(g34762),.A(g34687),.B(g34524));
  OR2 OR2_1954(.VSS(VSS),.VDD(VDD),.Y(g25740),.A(g25164),.B(g22055));
  OR2 OR2_1955(.VSS(VSS),.VDD(VDD),.Y(g26908),.A(g26358),.B(g24225));
  OR2 OR2_1956(.VSS(VSS),.VDD(VDD),.Y(g28640),.A(g27384),.B(g16590));
  OR2 OR2_1957(.VSS(VSS),.VDD(VDD),.Y(g30423),.A(g29887),.B(g21807));
  OR2 OR2_1958(.VSS(VSS),.VDD(VDD),.Y(g33976),.A(g33869),.B(g18347));
  OR2 OR2_1959(.VSS(VSS),.VDD(VDD),.Y(g33985),.A(g33896),.B(g18382));
  OR3 OR3_49(.VSS(VSS),.VDD(VDD),.Y(g24946),.A(g22360),.B(g22409),.C(g8130));
  OR2 OR2_1960(.VSS(VSS),.VDD(VDD),.Y(g25676),.A(g24668),.B(g21833));
  OR2 OR2_1961(.VSS(VSS),.VDD(VDD),.Y(g25685),.A(g24476),.B(g21866));
  OR4 OR4_80(.VSS(VSS),.VDD(VDD),.Y(I30750),.A(g31788),.B(g32310),.C(g32054),.D(g32070));
  OR3 OR3_50(.VSS(VSS),.VDD(VDD),.Y(g33954),.A(g33496),.B(I31853),.C(I31854));
  OR2 OR2_1962(.VSS(VSS),.VDD(VDD),.Y(g21891),.A(g19948),.B(g15103));
  OR2 OR2_1963(.VSS(VSS),.VDD(VDD),.Y(g24344),.A(g22145),.B(g18787));
  OR2 OR2_1964(.VSS(VSS),.VDD(VDD),.Y(g25654),.A(g24634),.B(g18606));
  OR2 OR2_1965(.VSS(VSS),.VDD(VDD),.Y(g25936),.A(g24403),.B(g22209));
  OR2 OR2_1966(.VSS(VSS),.VDD(VDD),.Y(g30543),.A(g29338),.B(g22110));
  OR4 OR4_81(.VSS(VSS),.VDD(VDD),.Y(I26522),.A(g19890),.B(g19935),.C(g19984),.D(g26365));
  OR2 OR2_1967(.VSS(VSS),.VDD(VDD),.Y(g31260),.A(g25993),.B(g29555));
  OR2 OR2_1968(.VSS(VSS),.VDD(VDD),.Y(g34000),.A(g33943),.B(g18441));
  OR2 OR2_1969(.VSS(VSS),.VDD(VDD),.Y(g26751),.A(g24903),.B(g24912));
  OR2 OR2_1970(.VSS(VSS),.VDD(VDD),.Y(g33260),.A(g32110),.B(g29524));
  OR2 OR2_1971(.VSS(VSS),.VDD(VDD),.Y(g29295),.A(g28663),.B(g18780));
  OR2 OR2_1972(.VSS(VSS),.VDD(VDD),.Y(g31668),.A(g29924),.B(g28558));
  OR2 OR2_1973(.VSS(VSS),.VDD(VDD),.Y(g14583),.A(g10685),.B(g542));
  OR2 OR2_1974(.VSS(VSS),.VDD(VDD),.Y(g25762),.A(g25095),.B(g18816));
  OR2 OR2_1975(.VSS(VSS),.VDD(VDD),.Y(g28662),.A(g27407),.B(g16612));
  OR2 OR2_1976(.VSS(VSS),.VDD(VDD),.Y(g26293),.A(g24550),.B(g24555));
  OR2 OR2_1977(.VSS(VSS),.VDD(VDD),.Y(g33559),.A(g33073),.B(g18368));
  OR4 OR4_82(.VSS(VSS),.VDD(VDD),.Y(I30192),.A(g29385),.B(g31376),.C(g30735),.D(g30825));
  OR2 OR2_1978(.VSS(VSS),.VDD(VDD),.Y(g33016),.A(g32284),.B(g18509));
  OR2 OR2_1979(.VSS(VSS),.VDD(VDD),.Y(g25587),.A(g21682),.B(g24157));
  OR2 OR2_1980(.VSS(VSS),.VDD(VDD),.Y(g33558),.A(g33350),.B(g18364));
  OR2 OR2_1981(.VSS(VSS),.VDD(VDD),.Y(g23750),.A(g20174),.B(g16840));
  OR2 OR2_1982(.VSS(VSS),.VDD(VDD),.Y(g31893),.A(g31490),.B(g21837));
  OR2 OR2_1983(.VSS(VSS),.VDD(VDD),.Y(g34807),.A(g34764),.B(g18596));
  OR2 OR2_1984(.VSS(VSS),.VDD(VDD),.Y(g34974),.A(g34870),.B(g34963));
  OR2 OR2_1985(.VSS(VSS),.VDD(VDD),.Y(g31865),.A(g31149),.B(g21709));
  OR2 OR2_1986(.VSS(VSS),.VDD(VDD),.Y(g33544),.A(g33392),.B(g18317));
  OR2 OR2_1987(.VSS(VSS),.VDD(VDD),.Y(g34639),.A(g34486),.B(g18722));
  OR2 OR2_1988(.VSS(VSS),.VDD(VDD),.Y(g12911),.A(g10278),.B(g12768));
  OR2 OR2_1989(.VSS(VSS),.VDD(VDD),.Y(g30293),.A(g28236),.B(g27246));
  OR3 OR3_51(.VSS(VSS),.VDD(VDD),.Y(g23796),.A(g21462),.B(g21433),.C(I22958));
  OR2 OR2_1990(.VSS(VSS),.VDD(VDD),.Y(g28778),.A(g27540),.B(g16808));
  OR2 OR2_1991(.VSS(VSS),.VDD(VDD),.Y(g16239),.A(g7892),.B(g13432));
  OR2 OR2_1992(.VSS(VSS),.VDD(VDD),.Y(g34293),.A(g26854),.B(g34224));
  OR2 OR2_1993(.VSS(VSS),.VDD(VDD),.Y(g34638),.A(g34484),.B(g18721));
  OR2 OR2_1994(.VSS(VSS),.VDD(VDD),.Y(g34265),.A(g34117),.B(g18711));
  OR2 OR2_1995(.VSS(VSS),.VDD(VDD),.Y(g30416),.A(g29858),.B(g21800));
  OR2 OR2_1996(.VSS(VSS),.VDD(VDD),.Y(g27591),.A(g26181),.B(g24765));
  OR2 OR2_1997(.VSS(VSS),.VDD(VDD),.Y(g34416),.A(g34191),.B(g25159));
  OR2 OR2_1998(.VSS(VSS),.VDD(VDD),.Y(g29289),.A(g28642),.B(g18763));
  OR2 OR2_1999(.VSS(VSS),.VDD(VDD),.Y(g25747),.A(g25130),.B(g18795));
  OR2 OR2_2000(.VSS(VSS),.VDD(VDD),.Y(g28647),.A(g27389),.B(g16596));
  OR2 OR2_2001(.VSS(VSS),.VDD(VDD),.Y(g33610),.A(g33242),.B(g18616));
  OR2 OR2_2002(.VSS(VSS),.VDD(VDD),.Y(g29309),.A(g28722),.B(g18818));
  OR2 OR2_2003(.VSS(VSS),.VDD(VDD),.Y(g30391),.A(g30080),.B(g18557));
  OR2 OR2_2004(.VSS(VSS),.VDD(VDD),.Y(g33042),.A(g32193),.B(g24324));
  OR2 OR2_2005(.VSS(VSS),.VDD(VDD),.Y(g27147),.A(g25802),.B(g24399));
  OR2 OR2_2006(.VSS(VSS),.VDD(VDD),.Y(g31255),.A(g25982),.B(g29536));
  OR2 OR2_2007(.VSS(VSS),.VDD(VDD),.Y(g29288),.A(g28630),.B(g18762));
  OR2 OR2_2008(.VSS(VSS),.VDD(VDD),.Y(g33255),.A(g32106),.B(g29514));
  OR2 OR2_2009(.VSS(VSS),.VDD(VDD),.Y(g29224),.A(g28919),.B(g18156));
  OR2 OR2_2010(.VSS(VSS),.VDD(VDD),.Y(g30510),.A(g30263),.B(g22031));
  OR2 OR2_2011(.VSS(VSS),.VDD(VDD),.Y(g29308),.A(g28612),.B(g18815));
  OR2 OR2_2012(.VSS(VSS),.VDD(VDD),.Y(g24240),.A(g22861),.B(g18251));
  OR2 OR2_2013(.VSS(VSS),.VDD(VDD),.Y(g33270),.A(g32119),.B(g29547));
  OR2 OR2_2014(.VSS(VSS),.VDD(VDD),.Y(g28090),.A(g27275),.B(g18733));
  OR2 OR2_2015(.VSS(VSS),.VDD(VDD),.Y(g30579),.A(g30173),.B(g14571));
  OR2 OR2_2016(.VSS(VSS),.VDD(VDD),.Y(g27858),.A(g17405),.B(g26737));
  OR2 OR2_2017(.VSS(VSS),.VDD(VDD),.Y(g25751),.A(g25061),.B(g22098));
  OR2 OR2_2018(.VSS(VSS),.VDD(VDD),.Y(g28651),.A(g27392),.B(g16599));
  OR2 OR2_2019(.VSS(VSS),.VDD(VDD),.Y(g29495),.A(g28563),.B(g27614));
  OR2 OR2_2020(.VSS(VSS),.VDD(VDD),.Y(g33383),.A(g32244),.B(g29940));
  OR2 OR2_2021(.VSS(VSS),.VDD(VDD),.Y(g25639),.A(g25122),.B(g18530));
  OR2 OR2_2022(.VSS(VSS),.VDD(VDD),.Y(g34014),.A(g33647),.B(g18493));
  OR2 OR2_2023(.VSS(VSS),.VDD(VDD),.Y(g33030),.A(g32166),.B(g21826));
  OR2 OR2_2024(.VSS(VSS),.VDD(VDD),.Y(g31267),.A(g29548),.B(g28263));
  OR2 OR2_2025(.VSS(VSS),.VDD(VDD),.Y(g25638),.A(g24977),.B(g18316));
  OR2 OR2_2026(.VSS(VSS),.VDD(VDD),.Y(g34007),.A(g33640),.B(g18467));
  OR2 OR2_2027(.VSS(VSS),.VDD(VDD),.Y(g16883),.A(g13509),.B(g11115));
  OR2 OR2_2028(.VSS(VSS),.VDD(VDD),.Y(g33267),.A(g32115),.B(g29535));
  OR2 OR2_2029(.VSS(VSS),.VDD(VDD),.Y(g33294),.A(g32152),.B(g29604));
  OR2 OR2_2030(.VSS(VSS),.VDD(VDD),.Y(g27394),.A(g25957),.B(g24573));
  OR2 OR2_2031(.VSS(VSS),.VDD(VDD),.Y(g28331),.A(g27129),.B(g15814));
  OR2 OR2_2032(.VSS(VSS),.VDD(VDD),.Y(g30442),.A(g29797),.B(g21851));
  OR2 OR2_2033(.VSS(VSS),.VDD(VDD),.Y(g33065),.A(g32008),.B(g22068));
  OR2 OR2_2034(.VSS(VSS),.VDD(VDD),.Y(g34442),.A(g34380),.B(g18542));
  OR2 OR2_2035(.VSS(VSS),.VDD(VDD),.Y(g28513),.A(g27276),.B(g26123));
  OR2 OR2_2036(.VSS(VSS),.VDD(VDD),.Y(g31875),.A(g31066),.B(g21730));
  OR2 OR2_2037(.VSS(VSS),.VDD(VDD),.Y(g29643),.A(g28192),.B(g27145));
  OR2 OR2_2038(.VSS(VSS),.VDD(VDD),.Y(g34615),.A(g34516),.B(g18576));
  OR3 OR3_52(.VSS(VSS),.VDD(VDD),.Y(g33219),.A(g32335),.B(I30760),.C(I30761));
  OR2 OR2_2039(.VSS(VSS),.VDD(VDD),.Y(g24262),.A(g23387),.B(g18315));
  OR2 OR2_2040(.VSS(VSS),.VDD(VDD),.Y(g28404),.A(g27215),.B(g15874));
  OR2 OR2_2041(.VSS(VSS),.VDD(VDD),.Y(g34720),.A(g34694),.B(g18134));
  OR2 OR2_2042(.VSS(VSS),.VDD(VDD),.Y(g34041),.A(g33829),.B(g18739));
  OR2 OR2_2043(.VSS(VSS),.VDD(VDD),.Y(g28717),.A(g27482),.B(g16701));
  OR2 OR2_2044(.VSS(VSS),.VDD(VDD),.Y(g30430),.A(g29859),.B(g21814));
  OR2 OR2_2045(.VSS(VSS),.VDD(VDD),.Y(g30493),.A(g30198),.B(g21989));
  OR2 OR2_2046(.VSS(VSS),.VDD(VDD),.Y(g28212),.A(g27030),.B(g27035));
  OR2 OR2_2047(.VSS(VSS),.VDD(VDD),.Y(g29260),.A(g28315),.B(g18604));
  OR2 OR2_2048(.VSS(VSS),.VDD(VDD),.Y(g25835),.A(g25367),.B(g23855));
  OR2 OR2_2049(.VSS(VSS),.VDD(VDD),.Y(g30465),.A(g30164),.B(g21936));
  OR2 OR2_2050(.VSS(VSS),.VDD(VDD),.Y(g34465),.A(g34295),.B(g18712));
  OR2 OR2_2051(.VSS(VSS),.VDD(VDD),.Y(g25586),.A(g21678),.B(g24156));
  OR2 OR2_2052(.VSS(VSS),.VDD(VDD),.Y(g34237),.A(g32715),.B(g33955));
  OR2 OR2_2053(.VSS(VSS),.VDD(VDD),.Y(g30340),.A(g29377),.B(g18245));
  OR2 OR2_2054(.VSS(VSS),.VDD(VDD),.Y(g29489),.A(g28550),.B(g27601));
  OR2 OR2_2055(.VSS(VSS),.VDD(VDD),.Y(g34035),.A(g33721),.B(g18714));
  OR2 OR2_2056(.VSS(VSS),.VDD(VDD),.Y(g29488),.A(g28547),.B(g27600));
  OR2 OR2_2057(.VSS(VSS),.VDD(VDD),.Y(g34806),.A(g34763),.B(g18595));
  OR2 OR2_2058(.VSS(VSS),.VDD(VDD),.Y(g23183),.A(g19545),.B(g15911));
  OR2 OR2_2059(.VSS(VSS),.VDD(VDD),.Y(g28723),.A(g27490),.B(g16706));
  OR2 OR2_2060(.VSS(VSS),.VDD(VDD),.Y(g33617),.A(g33263),.B(g24326));
  OR2 OR2_2061(.VSS(VSS),.VDD(VDD),.Y(g31915),.A(g31520),.B(g22001));
  OR2 OR2_2062(.VSS(VSS),.VDD(VDD),.Y(g25615),.A(g24803),.B(g18162));
  OR2 OR2_2063(.VSS(VSS),.VDD(VDD),.Y(g30517),.A(g30244),.B(g22038));
  OR2 OR2_2064(.VSS(VSS),.VDD(VDD),.Y(g28387),.A(g27203),.B(g15858));
  OR2 OR2_2065(.VSS(VSS),.VDD(VDD),.Y(g31277),.A(g29570),.B(g28285));
  OR2 OR2_2066(.VSS(VSS),.VDD(VDD),.Y(g25720),.A(g25042),.B(g18765));
  OR2 OR2_2067(.VSS(VSS),.VDD(VDD),.Y(g24247),.A(g22623),.B(g18259));
  OR2 OR2_2068(.VSS(VSS),.VDD(VDD),.Y(g33277),.A(g32129),.B(g29568));
  OR3 OR3_53(.VSS(VSS),.VDD(VDD),.Y(g14182),.A(g11741),.B(g11721),.C(g753));
  OR2 OR2_2069(.VSS(VSS),.VDD(VDD),.Y(g15935),.A(g13029),.B(g10665));
  OR2 OR2_2070(.VSS(VSS),.VDD(VDD),.Y(g28097),.A(g27682),.B(g22005));
  OR2 OR2_2071(.VSS(VSS),.VDD(VDD),.Y(g28104),.A(g27697),.B(g22108));
  OR2 OR2_2072(.VSS(VSS),.VDD(VDD),.Y(g25746),.A(g25217),.B(g22063));
  OR2 OR2_2073(.VSS(VSS),.VDD(VDD),.Y(g28646),.A(g27388),.B(g16595));
  OR2 OR2_2074(.VSS(VSS),.VDD(VDD),.Y(g33595),.A(g33368),.B(g18489));
  OR2 OR2_2075(.VSS(VSS),.VDD(VDD),.Y(g32235),.A(g31151),.B(g29662));
  OR2 OR2_2076(.VSS(VSS),.VDD(VDD),.Y(g27562),.A(g26102),.B(g24703));
  OR2 OR2_2077(.VSS(VSS),.VDD(VDD),.Y(g33623),.A(g33370),.B(g18792));
  OR4 OR4_83(.VSS(VSS),.VDD(VDD),.Y(I30756),.A(g32088),.B(g32163),.C(g32098),.D(g32105));
  OR2 OR2_2078(.VSS(VSS),.VDD(VDD),.Y(g33037),.A(g32177),.B(g24310));
  OR2 OR2_2079(.VSS(VSS),.VDD(VDD),.Y(g30362),.A(g30120),.B(g18392));
  OR2 OR2_2080(.VSS(VSS),.VDD(VDD),.Y(g34193),.A(g33809),.B(g33814));
  OR2 OR2_2081(.VSS(VSS),.VDD(VDD),.Y(g24251),.A(g22637),.B(g18296));
  OR2 OR2_2082(.VSS(VSS),.VDD(VDD),.Y(g24272),.A(g23056),.B(g18629));
  OR2 OR2_2083(.VSS(VSS),.VDD(VDD),.Y(g31782),.A(g30060),.B(g30070));
  OR2 OR2_2084(.VSS(VSS),.VDD(VDD),.Y(g27290),.A(g25926),.B(g25928));
  OR2 OR2_2085(.VSS(VSS),.VDD(VDD),.Y(g28369),.A(g27160),.B(g25938));
  OR2 OR2_2086(.VSS(VSS),.VDD(VDD),.Y(g30523),.A(g30245),.B(g22069));
  OR2 OR2_2087(.VSS(VSS),.VDD(VDD),.Y(g33984),.A(g33881),.B(g18374));
  OR2 OR2_2088(.VSS(VSS),.VDD(VDD),.Y(g25684),.A(g24983),.B(g18643));
  OR2 OR2_2089(.VSS(VSS),.VDD(VDD),.Y(g29255),.A(g28714),.B(g18516));
  OR2 OR2_2090(.VSS(VSS),.VDD(VDD),.Y(g28368),.A(g27158),.B(g27184));
  OR2 OR2_2091(.VSS(VSS),.VDD(VDD),.Y(g26703),.A(g24447),.B(g10705));
  OR2 OR2_2092(.VSS(VSS),.VDD(VDD),.Y(g29270),.A(g28258),.B(g18635));
  OR2 OR2_2093(.VSS(VSS),.VDD(VDD),.Y(g32991),.A(g32322),.B(g18349));
  OR2 OR2_2094(.VSS(VSS),.VDD(VDD),.Y(g30475),.A(g30220),.B(g21946));
  OR2 OR2_2095(.VSS(VSS),.VDD(VDD),.Y(g34006),.A(g33897),.B(g18462));
  OR2 OR2_2096(.VSS(VSS),.VDD(VDD),.Y(g28850),.A(g27557),.B(g16869));
  OR2 OR2_2097(.VSS(VSS),.VDD(VDD),.Y(g33266),.A(g32114),.B(g29532));
  OR2 OR2_2098(.VSS(VSS),.VDD(VDD),.Y(g23574),.A(g20093),.B(g20108));
  OR2 OR2_2099(.VSS(VSS),.VDD(VDD),.Y(g13972),.A(g11232),.B(g11203));
  OR2 OR2_2100(.VSS(VSS),.VDD(VDD),.Y(g34727),.A(g34655),.B(g18213));
  OR2 OR2_2101(.VSS(VSS),.VDD(VDD),.Y(g26781),.A(g24913),.B(g24921));
  OR2 OR2_2102(.VSS(VSS),.VDD(VDD),.Y(g30437),.A(g29876),.B(g21846));
  OR2 OR2_2103(.VSS(VSS),.VDD(VDD),.Y(g26952),.A(g26360),.B(g24290));
  OR2 OR2_2104(.VSS(VSS),.VDD(VDD),.Y(g29294),.A(g28645),.B(g18779));
  OR2 OR2_2105(.VSS(VSS),.VDD(VDD),.Y(g29267),.A(g28257),.B(g18622));
  OR2 OR2_2106(.VSS(VSS),.VDD(VDD),.Y(g19619),.A(g15712),.B(g13080));
  OR2 OR2_2107(.VSS(VSS),.VDD(VDD),.Y(g8863),.A(g1644),.B(g1664));
  OR2 OR2_2108(.VSS(VSS),.VDD(VDD),.Y(g19557),.A(g17123),.B(g14190));
  OR3 OR3_54(.VSS(VSS),.VDD(VDD),.Y(I22830),.A(g21429),.B(g21338),.C(g21307));
  OR2 OR2_2109(.VSS(VSS),.VDD(VDD),.Y(g27403),.A(g25962),.B(g24581));
  OR2 OR2_2110(.VSS(VSS),.VDD(VDD),.Y(g33589),.A(g33340),.B(g18469));
  OR2 OR2_2111(.VSS(VSS),.VDD(VDD),.Y(g30347),.A(g29383),.B(g18304));
  OR2 OR2_2112(.VSS(VSS),.VDD(VDD),.Y(g28716),.A(g27481),.B(g13887));
  OR2 OR2_2113(.VSS(VSS),.VDD(VDD),.Y(g34347),.A(g25986),.B(g34102));
  OR2 OR2_2114(.VSS(VSS),.VDD(VDD),.Y(g33588),.A(g33334),.B(g18468));
  OR2 OR2_2115(.VSS(VSS),.VDD(VDD),.Y(g34253),.A(g34171),.B(g24300));
  OR2 OR2_2116(.VSS(VSS),.VDD(VDD),.Y(g27226),.A(g25872),.B(g24436));
  OR2 OR2_2117(.VSS(VSS),.VDD(VDD),.Y(g28582),.A(g27330),.B(g26277));
  OR2 OR2_2118(.VSS(VSS),.VDD(VDD),.Y(g34600),.A(g34538),.B(g18182));
  OR2 OR2_2119(.VSS(VSS),.VDD(VDD),.Y(g24447),.A(g10948),.B(g22450));
  OR2 OR2_2120(.VSS(VSS),.VDD(VDD),.Y(g14387),.A(g9086),.B(g11048));
  OR2 OR2_2121(.VSS(VSS),.VDD(VDD),.Y(g34781),.A(g33431),.B(g34715));
  OR2 OR2_2122(.VSS(VSS),.VDD(VDD),.Y(g27551),.A(g26091),.B(g24675));
  OR2 OR2_2123(.VSS(VSS),.VDD(VDD),.Y(g27572),.A(g26129),.B(g24724));
  OR2 OR2_2124(.VSS(VSS),.VDD(VDD),.Y(g33119),.A(g32420),.B(g32428));
  OR2 OR2_2125(.VSS(VSS),.VDD(VDD),.Y(g28310),.A(g27107),.B(g15797));
  OR2 OR2_2126(.VSS(VSS),.VDD(VDD),.Y(g34236),.A(g32650),.B(g33954));
  OR2 OR2_2127(.VSS(VSS),.VDD(VDD),.Y(g30351),.A(g30084),.B(g18339));
  OR2 OR2_2128(.VSS(VSS),.VDD(VDD),.Y(g30372),.A(g30110),.B(g18446));
  OR2 OR2_2129(.VSS(VSS),.VDD(VDD),.Y(g25727),.A(g25163),.B(g22010));
  OR2 OR2_2130(.VSS(VSS),.VDD(VDD),.Y(g33118),.A(g32413),.B(g32418));
  OR2 OR2_2131(.VSS(VSS),.VDD(VDD),.Y(g34372),.A(g26287),.B(g34137));
  OR2 OR2_2132(.VSS(VSS),.VDD(VDD),.Y(g31864),.A(g31271),.B(g21703));
  OR2 OR2_2133(.VSS(VSS),.VDD(VDD),.Y(g33022),.A(g32306),.B(g21750));
  OR2 OR2_2134(.VSS(VSS),.VDD(VDD),.Y(g26422),.A(g24774),.B(g23104));
  OR2 OR2_2135(.VSS(VSS),.VDD(VDD),.Y(g31749),.A(g29974),.B(g29988));
  OR2 OR2_2136(.VSS(VSS),.VDD(VDD),.Y(g16052),.A(g13060),.B(g10724));
  OR2 OR2_2137(.VSS(VSS),.VDD(VDD),.Y(g7450),.A(g1277),.B(g1283));
  OR2 OR2_2138(.VSS(VSS),.VDD(VDD),.Y(g28050),.A(g27692),.B(g18165));
  OR2 OR2_2139(.VSS(VSS),.VDD(VDD),.Y(g33616),.A(g33237),.B(g24314));
  OR2 OR2_2140(.VSS(VSS),.VDD(VDD),.Y(g33313),.A(g29649),.B(g32171));
  OR2 OR2_2141(.VSS(VSS),.VDD(VDD),.Y(g30516),.A(g30233),.B(g22037));
  OR2 OR2_2142(.VSS(VSS),.VDD(VDD),.Y(g34264),.A(g34081),.B(g18701));
  OR2 OR2_2143(.VSS(VSS),.VDD(VDD),.Y(g28386),.A(g27202),.B(g13277));
  OR2 OR2_2144(.VSS(VSS),.VDD(VDD),.Y(g34790),.A(g34774),.B(g18151));
  OR2 OR2_2145(.VSS(VSS),.VDD(VDD),.Y(g31276),.A(g29567),.B(g28282));
  OR2 OR2_2146(.VSS(VSS),.VDD(VDD),.Y(g25703),.A(g25087),.B(g21922));
  OR2 OR2_2147(.VSS(VSS),.VDD(VDD),.Y(g28603),.A(g27340),.B(g26300));
  OR2 OR2_2148(.VSS(VSS),.VDD(VDD),.Y(g24246),.A(g23372),.B(g18257));
  OR2 OR2_2149(.VSS(VSS),.VDD(VDD),.Y(g33276),.A(g32128),.B(g29566));
  OR2 OR2_2150(.VSS(VSS),.VDD(VDD),.Y(g28096),.A(g27988),.B(g21997));
  OR2 OR2_2151(.VSS(VSS),.VDD(VDD),.Y(g32399),.A(g31527),.B(g30062));
  OR2 OR2_2152(.VSS(VSS),.VDD(VDD),.Y(g33053),.A(g31967),.B(g21974));
  OR2 OR2_2153(.VSS(VSS),.VDD(VDD),.Y(g31254),.A(g25981),.B(g29534));
  OR2 OR2_2154(.VSS(VSS),.VDD(VDD),.Y(g27980),.A(g26105),.B(g26131));
  OR2 OR2_2155(.VSS(VSS),.VDD(VDD),.Y(g33254),.A(g32104),.B(g29512));
  OR2 OR2_2156(.VSS(VSS),.VDD(VDD),.Y(g31900),.A(g31484),.B(g21908));
  OR2 OR2_2157(.VSS(VSS),.VDD(VDD),.Y(g31466),.A(g26160),.B(g29650));
  OR2 OR2_2158(.VSS(VSS),.VDD(VDD),.Y(g32398),.A(g31526),.B(g30061));
  OR3 OR3_55(.VSS(VSS),.VDD(VDD),.Y(I22267),.A(g20236),.B(g20133),.C(g20111));
  OR2 OR2_2159(.VSS(VSS),.VDD(VDD),.Y(g25600),.A(g24650),.B(g18111));
  OR2 OR2_2160(.VSS(VSS),.VDD(VDD),.Y(g26913),.A(g25848),.B(g18225));
  OR2 OR2_2161(.VSS(VSS),.VDD(VDD),.Y(g28681),.A(g27428),.B(g16634));
  OR2 OR2_2162(.VSS(VSS),.VDD(VDD),.Y(g23405),.A(g19791),.B(g16245));
  OR2 OR2_2163(.VSS(VSS),.VDD(VDD),.Y(g29277),.A(g28440),.B(g18710));
  OR2 OR2_2164(.VSS(VSS),.VDD(VDD),.Y(g30422),.A(g29795),.B(g21806));
  OR2 OR2_2165(.VSS(VSS),.VDD(VDD),.Y(g33036),.A(g32168),.B(g24309));
  OR2 OR2_2166(.VSS(VSS),.VDD(VDD),.Y(g28429),.A(g27228),.B(g15913));
  OR2 OR2_2167(.VSS(VSS),.VDD(VDD),.Y(g33560),.A(g33404),.B(g18369));
  OR2 OR2_2168(.VSS(VSS),.VDD(VDD),.Y(g24355),.A(g23799),.B(g18824));
  OR2 OR2_2169(.VSS(VSS),.VDD(VDD),.Y(g28730),.A(g27503),.B(g13912));
  OR2 OR2_2170(.VSS(VSS),.VDD(VDD),.Y(g26905),.A(g26397),.B(g24222));
  OR4 OR4_84(.VSS(VSS),.VDD(VDD),.Y(g25821),.A(g25482),.B(g25456),.C(g25417),.D(g25377));
  OR2 OR2_2171(.VSS(VSS),.VDD(VDD),.Y(g28428),.A(g27227),.B(g15912));
  OR2 OR2_2172(.VSS(VSS),.VDD(VDD),.Y(g30542),.A(g29337),.B(g22088));
  OR2 OR2_2173(.VSS(VSS),.VDD(VDD),.Y(g30453),.A(g29902),.B(g21862));
  OR2 OR2_2174(.VSS(VSS),.VDD(VDD),.Y(g33064),.A(g31993),.B(g22067));
  OR2 OR2_2175(.VSS(VSS),.VDD(VDD),.Y(g19363),.A(g17810),.B(g14913));
  OR2 OR2_2176(.VSS(VSS),.VDD(VDD),.Y(g28690),.A(g27436),.B(g16641));
  OR2 OR2_2177(.VSS(VSS),.VDD(VDD),.Y(g34021),.A(g33652),.B(g18519));
  OR2 OR2_2178(.VSS(VSS),.VDD(VDD),.Y(g34453),.A(g34410),.B(g18666));
  OR2 OR2_2179(.VSS(VSS),.VDD(VDD),.Y(g27426),.A(g25967),.B(g24588));
  OR2 OR2_2180(.VSS(VSS),.VDD(VDD),.Y(g28549),.A(g27304),.B(g26233));
  OR2 OR2_2181(.VSS(VSS),.VDD(VDD),.Y(g24151),.A(g18088),.B(g21661));
  OR2 OR2_2182(.VSS(VSS),.VDD(VDD),.Y(g33733),.A(g33105),.B(g32012));
  OR2 OR2_2183(.VSS(VSS),.VDD(VDD),.Y(g32361),.A(g29869),.B(g31300));
  OR2 OR2_2184(.VSS(VSS),.VDD(VDD),.Y(g34726),.A(g34665),.B(g18212));
  OR2 OR2_2185(.VSS(VSS),.VDD(VDD),.Y(g28548),.A(g27303),.B(g26232));
  OR2 OR2_2186(.VSS(VSS),.VDD(VDD),.Y(g31874),.A(g31016),.B(g21729));
  OR2 OR2_2187(.VSS(VSS),.VDD(VDD),.Y(g30436),.A(g29860),.B(g21845));
  OR2 OR2_2188(.VSS(VSS),.VDD(VDD),.Y(g19486),.A(g15589),.B(g12979));
  OR2 OR2_2189(.VSS(VSS),.VDD(VDD),.Y(g34614),.A(g34518),.B(g18568));
  OR2 OR2_2190(.VSS(VSS),.VDD(VDD),.Y(g29266),.A(g28330),.B(g18621));
  OR2 OR2_2191(.VSS(VSS),.VDD(VDD),.Y(g34607),.A(g34567),.B(g15081));
  OR2 OR2_2192(.VSS(VSS),.VDD(VDD),.Y(g30530),.A(g30224),.B(g22076));
  OR2 OR2_2193(.VSS(VSS),.VDD(VDD),.Y(g28317),.A(g27114),.B(g15805));
  OR2 OR2_2194(.VSS(VSS),.VDD(VDD),.Y(g33009),.A(g32273),.B(g18458));
  OR2 OR2_2195(.VSS(VSS),.VDD(VDD),.Y(g34274),.A(g27822),.B(g34205));
  OR2 OR2_2196(.VSS(VSS),.VDD(VDD),.Y(g30346),.A(g29381),.B(g18303));
  OR2 OR2_2197(.VSS(VSS),.VDD(VDD),.Y(g25834),.A(g25366),.B(g23854));
  OR2 OR2_2198(.VSS(VSS),.VDD(VDD),.Y(g27024),.A(g26826),.B(g17692));
  OR4 OR4_85(.VSS(VSS),.VDD(VDD),.Y(I31849),.A(g33483),.B(g33484),.C(g33485),.D(g33486));
  OR2 OR2_2199(.VSS(VSS),.VDD(VDD),.Y(g33008),.A(g32261),.B(g18457));
  OR2 OR2_2200(.VSS(VSS),.VDD(VDD),.Y(g30464),.A(g30152),.B(g21935));
  OR2 OR2_2201(.VSS(VSS),.VDD(VDD),.Y(g32221),.A(g31140),.B(g29634));
  OR2 OR2_2202(.VSS(VSS),.VDD(VDD),.Y(g34464),.A(g34340),.B(g18687));
  OR2 OR2_2203(.VSS(VSS),.VDD(VDD),.Y(g31892),.A(g31019),.B(g21825));
  OR4 OR4_86(.VSS(VSS),.VDD(VDD),.Y(I31848),.A(g33479),.B(g33480),.C(g33481),.D(g33482));
  OR2 OR2_2204(.VSS(VSS),.VDD(VDD),.Y(g28057),.A(g27033),.B(g18218));
  OR2 OR2_2205(.VSS(VSS),.VDD(VDD),.Y(g34034),.A(g33719),.B(g18713));
  OR2 OR2_2206(.VSS(VSS),.VDD(VDD),.Y(g33555),.A(g33355),.B(g18357));
  OR2 OR2_2207(.VSS(VSS),.VDD(VDD),.Y(g34641),.A(g34479),.B(g18724));
  OR2 OR2_2208(.VSS(VSS),.VDD(VDD),.Y(g34797),.A(g34747),.B(g18574));
  OR2 OR2_2209(.VSS(VSS),.VDD(VDD),.Y(g25726),.A(g25148),.B(g22009));
  OR2 OR2_2210(.VSS(VSS),.VDD(VDD),.Y(g33570),.A(g33420),.B(g18405));
  OR2 OR2_2211(.VSS(VSS),.VDD(VDD),.Y(g31914),.A(g31499),.B(g22000));
  OR2 OR2_2212(.VSS(VSS),.VDD(VDD),.Y(g34292),.A(g26853),.B(g34223));
  OR2 OR2_2213(.VSS(VSS),.VDD(VDD),.Y(g28323),.A(g27118),.B(g15810));
  OR2 OR2_2214(.VSS(VSS),.VDD(VDD),.Y(g33914),.A(g33305),.B(g33311));
  OR2 OR2_2215(.VSS(VSS),.VDD(VDD),.Y(g34153),.A(g33899),.B(g33451));
  OR2 OR2_2216(.VSS(VSS),.VDD(VDD),.Y(g27126),.A(g24378),.B(g25787));
  OR2 OR2_2217(.VSS(VSS),.VDD(VDD),.Y(g25614),.A(g24797),.B(g18161));
  OR2 OR2_2218(.VSS(VSS),.VDD(VDD),.Y(g28533),.A(g27291),.B(g26203));
  OR2 OR2_2219(.VSS(VSS),.VDD(VDD),.Y(g31907),.A(g31492),.B(g21954));
  OR2 OR2_2220(.VSS(VSS),.VDD(VDD),.Y(g30409),.A(g29842),.B(g21768));
  OR2 OR2_2221(.VSS(VSS),.VDD(VDD),.Y(g27250),.A(g25901),.B(g15738));
  OR2 OR2_2222(.VSS(VSS),.VDD(VDD),.Y(g26891),.A(g26652),.B(g24197));
  OR2 OR2_2223(.VSS(VSS),.VDD(VDD),.Y(g24203),.A(g22982),.B(g18107));
  OR2 OR2_2224(.VSS(VSS),.VDD(VDD),.Y(g25607),.A(g24773),.B(g18118));
  OR2 OR2_2225(.VSS(VSS),.VDD(VDD),.Y(g10802),.A(g7533),.B(g1296));
  OR4 OR4_87(.VSS(VSS),.VDD(VDD),.Y(g15732),.A(g13411),.B(g13384),.C(g13349),.D(g11016));
  OR2 OR2_2226(.VSS(VSS),.VDD(VDD),.Y(g28775),.A(g27537),.B(g16806));
  OR2 OR2_2227(.VSS(VSS),.VDD(VDD),.Y(g30408),.A(g29806),.B(g21767));
  OR2 OR2_2228(.VSS(VSS),.VDD(VDD),.Y(g29864),.A(g28272),.B(g26086));
  OR2 OR2_2229(.VSS(VSS),.VDD(VDD),.Y(g34635),.A(g34485),.B(g18692));
  OR2 OR2_2230(.VSS(VSS),.VDD(VDD),.Y(g25593),.A(g24716),.B(g21707));
  OR2 OR2_2231(.VSS(VSS),.VDD(VDD),.Y(g33567),.A(g33081),.B(g18394));
  OR2 OR2_2232(.VSS(VSS),.VDD(VDD),.Y(g33594),.A(g33421),.B(g18485));
  OR2 OR2_2233(.VSS(VSS),.VDD(VDD),.Y(g32371),.A(g29883),.B(g31313));
  OR2 OR2_2234(.VSS(VSS),.VDD(VDD),.Y(g29313),.A(g28284),.B(g27270));
  OR2 OR2_2235(.VSS(VSS),.VDD(VDD),.Y(g24281),.A(g23397),.B(g18656));
  OR2 OR2_2236(.VSS(VSS),.VDD(VDD),.Y(g33238),.A(g32048),.B(g32051));
  OR2 OR2_2237(.VSS(VSS),.VDD(VDD),.Y(g26327),.A(g8462),.B(g24591));
  OR2 OR2_2238(.VSS(VSS),.VDD(VDD),.Y(g22225),.A(g21332),.B(g17654));
  OR2 OR2_2239(.VSS(VSS),.VDD(VDD),.Y(g29748),.A(g28210),.B(g28214));
  OR2 OR2_2240(.VSS(VSS),.VDD(VDD),.Y(g22708),.A(g19266),.B(g15711));
  OR2 OR2_2241(.VSS(VSS),.VDD(VDD),.Y(g29276),.A(g28616),.B(g18709));
  OR2 OR2_2242(.VSS(VSS),.VDD(VDD),.Y(g29285),.A(g28639),.B(g18750));
  OR2 OR2_2243(.VSS(VSS),.VDD(VDD),.Y(g29305),.A(g28602),.B(g18811));
  OR2 OR2_2244(.VSS(VSS),.VDD(VDD),.Y(g29254),.A(g28725),.B(g18512));
  OR3 OR3_56(.VSS(VSS),.VDD(VDD),.Y(g33176),.A(g32198),.B(I30734),.C(I30735));
  OR2 OR2_2245(.VSS(VSS),.VDD(VDD),.Y(g16882),.A(g13508),.B(g11114));
  OR2 OR2_2246(.VSS(VSS),.VDD(VDD),.Y(g30474),.A(g30208),.B(g21945));
  OR2 OR2_2247(.VSS(VSS),.VDD(VDD),.Y(g25635),.A(g24504),.B(g18293));
  OR2 OR2_2248(.VSS(VSS),.VDD(VDD),.Y(g31883),.A(g31132),.B(g21777));
  OR2 OR2_2249(.VSS(VSS),.VDD(VDD),.Y(g30537),.A(g30246),.B(g22083));
  OR2 OR2_2250(.VSS(VSS),.VDD(VDD),.Y(g19587),.A(g15700),.B(g13046));
  OR4 OR4_88(.VSS(VSS),.VDD(VDD),.Y(I30331),.A(g31672),.B(g31710),.C(g31021),.D(g30937));
  OR2 OR2_2251(.VSS(VSS),.VDD(VDD),.Y(g34537),.A(g34324),.B(g34084));
  OR2 OR2_2252(.VSS(VSS),.VDD(VDD),.Y(g13794),.A(g7396),.B(g10684));
  OR2 OR2_2253(.VSS(VSS),.VDD(VDD),.Y(g34283),.A(g26839),.B(g34215));
  OR2 OR2_2254(.VSS(VSS),.VDD(VDD),.Y(g30492),.A(g30188),.B(g21988));
  OR2 OR2_2255(.VSS(VSS),.VDD(VDD),.Y(g34606),.A(g34564),.B(g15080));
  OR2 OR2_2256(.VSS(VSS),.VDD(VDD),.Y(g34303),.A(g25768),.B(g34045));
  OR2 OR2_2257(.VSS(VSS),.VDD(VDD),.Y(g28316),.A(g27113),.B(g15804));
  OR2 OR2_2258(.VSS(VSS),.VDD(VDD),.Y(g27581),.A(g26161),.B(g24750));
  OR2 OR2_2259(.VSS(VSS),.VDD(VDD),.Y(g27450),.A(g2917),.B(g26483));
  OR4 OR4_89(.VSS(VSS),.VDD(VDD),.Y(I30717),.A(g31787),.B(g32200),.C(g31940),.D(g31949));
  OR2 OR2_2260(.VSS(VSS),.VDD(VDD),.Y(g33577),.A(g33405),.B(g18430));
  OR2 OR2_2261(.VSS(VSS),.VDD(VDD),.Y(g30381),.A(g30126),.B(g18497));
  OR2 OR2_2262(.VSS(VSS),.VDD(VDD),.Y(g25575),.A(g24139),.B(g24140));
  OR2 OR2_2263(.VSS(VSS),.VDD(VDD),.Y(g28056),.A(g27230),.B(g18210));
  OR2 OR2_2264(.VSS(VSS),.VDD(VDD),.Y(g32359),.A(g29867),.B(g31298));
  OR2 OR2_2265(.VSS(VSS),.VDD(VDD),.Y(g27257),.A(g25904),.B(g24498));
  OR2 OR2_2266(.VSS(VSS),.VDD(VDD),.Y(g29166),.A(g27653),.B(g17153));
  OR2 OR2_2267(.VSS(VSS),.VDD(VDD),.Y(g25711),.A(g25105),.B(g21962));
  OR2 OR2_2268(.VSS(VSS),.VDD(VDD),.Y(g28611),.A(g27348),.B(g16485));
  OR2 OR2_2269(.VSS(VSS),.VDD(VDD),.Y(g24715),.A(g22189),.B(g22207));
  OR2 OR2_2270(.VSS(VSS),.VDD(VDD),.Y(g32358),.A(g29866),.B(g31297));
  OR2 OR2_2271(.VSS(VSS),.VDD(VDD),.Y(g34796),.A(g34745),.B(g18573));
  OR2 OR2_2272(.VSS(VSS),.VDD(VDD),.Y(g29892),.A(g28300),.B(g26120));
  OR2 OR2_2273(.VSS(VSS),.VDD(VDD),.Y(g27590),.A(g26179),.B(g24764));
  OR2 OR2_2274(.VSS(VSS),.VDD(VDD),.Y(g29476),.A(g28108),.B(g28112));
  OR2 OR2_2275(.VSS(VSS),.VDD(VDD),.Y(g29485),.A(g28535),.B(g27594));
  OR2 OR2_2276(.VSS(VSS),.VDD(VDD),.Y(g31906),.A(g31477),.B(g21953));
  OR2 OR2_2277(.VSS(VSS),.VDD(VDD),.Y(g30390),.A(g29985),.B(g18555));
  OR2 OR2_2278(.VSS(VSS),.VDD(VDD),.Y(g32344),.A(g29804),.B(g31266));
  OR2 OR2_2279(.VSS(VSS),.VDD(VDD),.Y(g31284),.A(g29575),.B(g28290));
  OR2 OR2_2280(.VSS(VSS),.VDD(VDD),.Y(g25606),.A(g24761),.B(g18117));
  OR2 OR2_2281(.VSS(VSS),.VDD(VDD),.Y(g28342),.A(g27134),.B(g15819));
  OR2 OR2_2282(.VSS(VSS),.VDD(VDD),.Y(g31304),.A(g29594),.B(g29608));
  OR3 OR3_57(.VSS(VSS),.VDD(VDD),.Y(g29914),.A(g22531),.B(g22585),.C(I28147));
  OR2 OR2_2283(.VSS(VSS),.VDD(VDD),.Y(g21897),.A(g20095),.B(g15111));
  OR2 OR2_2284(.VSS(VSS),.VDD(VDD),.Y(g33622),.A(g33366),.B(g18791));
  OR2 OR2_2285(.VSS(VSS),.VDD(VDD),.Y(g33566),.A(g33356),.B(g18390));
  OR2 OR2_2286(.VSS(VSS),.VDD(VDD),.Y(g25750),.A(g25543),.B(g18802));
  OR2 OR2_2287(.VSS(VSS),.VDD(VDD),.Y(g26949),.A(g26356),.B(g24287));
  OR2 OR2_2288(.VSS(VSS),.VDD(VDD),.Y(g28650),.A(g27391),.B(g16598));
  OR2 OR2_2289(.VSS(VSS),.VDD(VDD),.Y(g30522),.A(g29332),.B(g22064));
  OR2 OR2_2290(.VSS(VSS),.VDD(VDD),.Y(g27150),.A(g25804),.B(g24400));
  OR2 OR2_2291(.VSS(VSS),.VDD(VDD),.Y(g34663),.A(g32028),.B(g34500));
  OR2 OR2_2292(.VSS(VSS),.VDD(VDD),.Y(g29239),.A(g28427),.B(g18297));
  OR2 OR2_2293(.VSS(VSS),.VDD(VDD),.Y(g26948),.A(g26399),.B(g24286));
  OR2 OR2_2294(.VSS(VSS),.VDD(VDD),.Y(g24354),.A(g23775),.B(g18823));
  OR2 OR2_2295(.VSS(VSS),.VDD(VDD),.Y(g27019),.A(g26822),.B(g14610));
  OR2 OR2_2296(.VSS(VSS),.VDD(VDD),.Y(g26904),.A(g26393),.B(g24221));
  OR2 OR2_2297(.VSS(VSS),.VDD(VDD),.Y(g29238),.A(g28178),.B(g18292));
  OR2 OR2_2298(.VSS(VSS),.VDD(VDD),.Y(g30483),.A(g30241),.B(g21979));
  OR2 OR2_2299(.VSS(VSS),.VDD(VDD),.Y(g30553),.A(g30205),.B(g22124));
  OR2 OR2_2300(.VSS(VSS),.VDD(VDD),.Y(g22901),.A(g19384),.B(g15745));
  OR2 OR2_2301(.VSS(VSS),.VDD(VDD),.Y(g28132),.A(g27932),.B(g27957));
  OR2 OR2_2302(.VSS(VSS),.VDD(VDD),.Y(g13997),.A(g11029),.B(g11036));
  OR2 OR2_2303(.VSS(VSS),.VDD(VDD),.Y(g29176),.A(g27661),.B(g17177));
  OR2 OR2_2304(.VSS(VSS),.VDD(VDD),.Y(g30536),.A(g30234),.B(g22082));
  OR2 OR2_2305(.VSS(VSS),.VDD(VDD),.Y(g26673),.A(g24433),.B(g10674));
  OR2 OR2_2306(.VSS(VSS),.VDD(VDD),.Y(g34040),.A(g33818),.B(g18737));
  OR2 OR2_2307(.VSS(VSS),.VDD(VDD),.Y(g33963),.A(g33830),.B(g18124));
  OR2 OR2_2308(.VSS(VSS),.VDD(VDD),.Y(g25663),.A(g24666),.B(g21788));
  OR2 OR2_2309(.VSS(VSS),.VDD(VDD),.Y(g34252),.A(g34146),.B(g18180));
  OR2 OR2_2310(.VSS(VSS),.VDD(VDD),.Y(g34621),.A(g34517),.B(g18583));
  OR2 OR2_2311(.VSS(VSS),.VDD(VDD),.Y(g28708),.A(g27462),.B(g16674));
  OR2 OR2_2312(.VSS(VSS),.VDD(VDD),.Y(g26933),.A(g26808),.B(g18551));
  OR2 OR2_2313(.VSS(VSS),.VDD(VDD),.Y(g28087),.A(g27255),.B(g18720));
  OR2 OR2_2314(.VSS(VSS),.VDD(VDD),.Y(g33576),.A(g33401),.B(g18423));
  OR2 OR2_2315(.VSS(VSS),.VDD(VDD),.Y(g33585),.A(g33411),.B(g18456));
  OR2 OR2_2316(.VSS(VSS),.VDD(VDD),.Y(g24211),.A(g23572),.B(g18138));
  OR2 OR2_2317(.VSS(VSS),.VDD(VDD),.Y(g28043),.A(g27323),.B(g21714));
  OR2 OR2_2318(.VSS(VSS),.VDD(VDD),.Y(g33554),.A(g33407),.B(g18353));
  OR2 OR2_2319(.VSS(VSS),.VDD(VDD),.Y(g32240),.A(g24757),.B(g31182));
  OR2 OR2_2320(.VSS(VSS),.VDD(VDD),.Y(g30397),.A(g29747),.B(g21756));
  OR4 OR4_90(.VSS(VSS),.VDD(VDD),.Y(I26742),.A(g23430),.B(g23445),.C(g23458),.D(g23481));
  OR2 OR2_2321(.VSS(VSS),.VDD(VDD),.Y(g33609),.A(g33239),.B(g18615));
  OR2 OR2_2322(.VSS(VSS),.VDD(VDD),.Y(g29501),.A(g28583),.B(g27634));
  OR2 OR2_2323(.VSS(VSS),.VDD(VDD),.Y(g33312),.A(g29646),.B(g32170));
  OR2 OR2_2324(.VSS(VSS),.VDD(VDD),.Y(g30509),.A(g30210),.B(g22030));
  OR2 OR2_2325(.VSS(VSS),.VDD(VDD),.Y(g33608),.A(g33322),.B(g18537));
  OR2 OR2_2326(.VSS(VSS),.VDD(VDD),.Y(g28069),.A(g27564),.B(g21865));
  OR2 OR2_2327(.VSS(VSS),.VDD(VDD),.Y(g33115),.A(g32397),.B(g32401));
  OR2 OR2_2328(.VSS(VSS),.VDD(VDD),.Y(g25702),.A(g25068),.B(g21921));
  OR2 OR2_2329(.VSS(VSS),.VDD(VDD),.Y(g25757),.A(g25132),.B(g22104));
  OR2 OR2_2330(.VSS(VSS),.VDD(VDD),.Y(g28774),.A(g27536),.B(g16804));
  OR2 OR2_2331(.VSS(VSS),.VDD(VDD),.Y(g30508),.A(g30199),.B(g22029));
  OR2 OR2_2332(.VSS(VSS),.VDD(VDD),.Y(g31921),.A(g31508),.B(g22046));
  OR2 OR2_2333(.VSS(VSS),.VDD(VDD),.Y(g28068),.A(g27310),.B(g21838));
  OR2 OR2_2334(.VSS(VSS),.VDD(VDD),.Y(g32981),.A(g32425),.B(g18206));
  OR2 OR2_2335(.VSS(VSS),.VDD(VDD),.Y(g28375),.A(g27183),.B(g15851));
  OR2 OR2_2336(.VSS(VSS),.VDD(VDD),.Y(g33052),.A(g31961),.B(g21973));
  OR2 OR2_2337(.VSS(VSS),.VDD(VDD),.Y(g34634),.A(g34483),.B(g18691));
  OR2 OR2_2338(.VSS(VSS),.VDD(VDD),.Y(g25621),.A(g24523),.B(g18205));
  OR2 OR2_2339(.VSS(VSS),.VDD(VDD),.Y(g31745),.A(g29959),.B(g29973));
  OR2 OR2_2340(.VSS(VSS),.VDD(VDD),.Y(g21896),.A(g20084),.B(g15110));
  OR2 OR2_2341(.VSS(VSS),.VDD(VDD),.Y(g24250),.A(g22633),.B(g18295));
  OR2 OR2_2342(.VSS(VSS),.VDD(VDD),.Y(g26912),.A(g25946),.B(g18209));
  OR2 OR2_2343(.VSS(VSS),.VDD(VDD),.Y(g27231),.A(g25873),.B(g15699));
  OR2 OR2_2344(.VSS(VSS),.VDD(VDD),.Y(g29284),.A(g28554),.B(g18747));
  OR2 OR2_2345(.VSS(VSS),.VDD(VDD),.Y(g32395),.A(g31523),.B(g30049));
  OR2 OR2_2346(.VSS(VSS),.VDD(VDD),.Y(g24339),.A(g23690),.B(g18756));
  OR2 OR2_2347(.VSS(VSS),.VDD(VDD),.Y(g33973),.A(g33840),.B(g18344));
  OR2 OR2_2348(.VSS(VSS),.VDD(VDD),.Y(g29304),.A(g28588),.B(g18810));
  OR2 OR2_2349(.VSS(VSS),.VDD(VDD),.Y(g32262),.A(g31186),.B(g29710));
  OR2 OR2_2350(.VSS(VSS),.VDD(VDD),.Y(g23716),.A(g9194),.B(g20905));
  OR2 OR2_2351(.VSS(VSS),.VDD(VDD),.Y(g25673),.A(g24727),.B(g21830));
  OR2 OR2_2352(.VSS(VSS),.VDD(VDD),.Y(g32990),.A(g32281),.B(g18341));
  OR3 OR3_58(.VSS(VSS),.VDD(VDD),.Y(I18417),.A(g14444),.B(g14414),.C(g14392));
  OR2 OR2_2353(.VSS(VSS),.VDD(VDD),.Y(g24338),.A(g23658),.B(g18755));
  OR2 OR2_2354(.VSS(VSS),.VDD(VDD),.Y(g11370),.A(g8807),.B(g550));
  OR2 OR2_2355(.VSS(VSS),.VDD(VDD),.Y(g30452),.A(g29891),.B(g21861));
  OR2 OR2_2356(.VSS(VSS),.VDD(VDD),.Y(g34452),.A(g34401),.B(g18665));
  OR2 OR2_2357(.VSS(VSS),.VDD(VDD),.Y(g13858),.A(g209),.B(g10685));
  OR2 OR2_2358(.VSS(VSS),.VDD(VDD),.Y(g33732),.A(g33104),.B(g32011));
  OR2 OR2_2359(.VSS(VSS),.VDD(VDD),.Y(g30311),.A(g28265),.B(g27265));
  OR3 OR3_59(.VSS(VSS),.VDD(VDD),.Y(g24968),.A(g22360),.B(g22409),.C(g23389));
  OR2 OR2_2360(.VSS(VSS),.VDD(VDD),.Y(g25634),.A(g24559),.B(g18284));
  OR2 OR2_2361(.VSS(VSS),.VDD(VDD),.Y(g31761),.A(g30009),.B(g30028));
  OR2 OR2_2362(.VSS(VSS),.VDD(VDD),.Y(g33692),.A(g32400),.B(g33428));
  OR2 OR2_2363(.VSS(VSS),.VDD(VDD),.Y(g19475),.A(g16930),.B(g14126));
  OR2 OR2_2364(.VSS(VSS),.VDD(VDD),.Y(g27456),.A(g25978),.B(g24607));
  OR2 OR2_2365(.VSS(VSS),.VDD(VDD),.Y(g26396),.A(g24762),.B(g23062));
  OR2 OR2_2366(.VSS(VSS),.VDD(VDD),.Y(g28545),.A(g27301),.B(g26230));
  OR2 OR2_2367(.VSS(VSS),.VDD(VDD),.Y(g28078),.A(g27140),.B(g21880));
  OR2 OR2_2368(.VSS(VSS),.VDD(VDD),.Y(g33013),.A(g32283),.B(g18484));
  OR2 OR2_2369(.VSS(VSS),.VDD(VDD),.Y(g22669),.A(g7763),.B(g19525));
  OR2 OR2_2370(.VSS(VSS),.VDD(VDD),.Y(g32247),.A(g31168),.B(g29686));
  OR3 OR3_60(.VSS(VSS),.VDD(VDD),.Y(I18543),.A(g14568),.B(g14540),.C(g14516));
  OR2 OR2_2371(.VSS(VSS),.VDD(VDD),.Y(g28086),.A(g27268),.B(g18702));
  OR2 OR2_2372(.VSS(VSS),.VDD(VDD),.Y(g32389),.A(g31496),.B(g29966));
  OR2 OR2_2373(.VSS(VSS),.VDD(VDD),.Y(g30350),.A(g30118),.B(g18334));
  OR2 OR2_2374(.VSS(VSS),.VDD(VDD),.Y(g34350),.A(g26048),.B(g34106));
  OR2 OR2_2375(.VSS(VSS),.VDD(VDD),.Y(g33539),.A(g33245),.B(g18178));
  OR2 OR2_2376(.VSS(VSS),.VDD(VDD),.Y(g32388),.A(g31495),.B(g29962));
  OR2 OR2_2377(.VSS(VSS),.VDD(VDD),.Y(g33005),.A(g32260),.B(g18432));
  OR2 OR2_2378(.VSS(VSS),.VDD(VDD),.Y(g27596),.A(g26207),.B(g24775));
  OR2 OR2_2379(.VSS(VSS),.VDD(VDD),.Y(g11025),.A(g2980),.B(g7831));
  OR2 OR2_2380(.VSS(VSS),.VDD(VDD),.Y(g28817),.A(g27548),.B(g16845));
  OR2 OR2_2381(.VSS(VSS),.VDD(VDD),.Y(g33538),.A(g33252),.B(g18144));
  OR2 OR2_2382(.VSS(VSS),.VDD(VDD),.Y(g28322),.A(g27117),.B(g15809));
  OR2 OR2_2383(.VSS(VSS),.VDD(VDD),.Y(g27243),.A(g25884),.B(g24475));
  OR2 OR2_2384(.VSS(VSS),.VDD(VDD),.Y(g30396),.A(g29856),.B(g21755));
  OR2 OR2_2385(.VSS(VSS),.VDD(VDD),.Y(g32251),.A(g30599),.B(g29352));
  OR2 OR2_2386(.VSS(VSS),.VDD(VDD),.Y(g13540),.A(g10822),.B(g10827));
  OR2 OR2_2387(.VSS(VSS),.VDD(VDD),.Y(g27431),.A(g24582),.B(g25977));
  OR2 OR2_2388(.VSS(VSS),.VDD(VDD),.Y(g20202),.A(g16211),.B(g13507));
  OR2 OR2_2389(.VSS(VSS),.VDD(VDD),.Y(g34731),.A(g34662),.B(g18272));
  OR2 OR2_2390(.VSS(VSS),.VDD(VDD),.Y(g29484),.A(g28124),.B(g22191));
  OR2 OR2_2391(.VSS(VSS),.VDD(VDD),.Y(g24202),.A(g22899),.B(g18106));
  OR2 OR2_2392(.VSS(VSS),.VDD(VDD),.Y(g26929),.A(g26635),.B(g18543));
  OR2 OR2_2393(.VSS(VSS),.VDD(VDD),.Y(g24257),.A(g22938),.B(g18310));
  OR2 OR2_2394(.VSS(VSS),.VDD(VDD),.Y(g30413),.A(g30001),.B(g21772));
  OR2 OR2_2395(.VSS(VSS),.VDD(VDD),.Y(g24496),.A(g24008),.B(g21557));
  OR2 OR2_2396(.VSS(VSS),.VDD(VDD),.Y(g31241),.A(g25959),.B(g29510));
  OR2 OR2_2397(.VSS(VSS),.VDD(VDD),.Y(g26928),.A(g26713),.B(g18541));
  OR4 OR4_91(.VSS(VSS),.VDD(VDD),.Y(g17488),.A(g14361),.B(g14335),.C(g11954),.D(I18417));
  OR2 OR2_2398(.VSS(VSS),.VDD(VDD),.Y(g25592),.A(g24672),.B(g21706));
  OR2 OR2_2399(.VSS(VSS),.VDD(VDD),.Y(g25756),.A(g25112),.B(g22103));
  OR2 OR2_2400(.VSS(VSS),.VDD(VDD),.Y(g28561),.A(g27312),.B(g26250));
  OR2 OR2_2401(.VSS(VSS),.VDD(VDD),.Y(g28295),.A(g27094),.B(g15783));
  OR2 OR2_2402(.VSS(VSS),.VDD(VDD),.Y(g28680),.A(g27427),.B(g16633));
  OR2 OR2_2403(.VSS(VSS),.VDD(VDD),.Y(g32997),.A(g32269),.B(g18378));
  OR2 OR2_2404(.VSS(VSS),.VDD(VDD),.Y(g30405),.A(g29767),.B(g21764));
  OR2 OR2_2405(.VSS(VSS),.VDD(VDD),.Y(g16173),.A(g8796),.B(g13464));
  OR2 OR2_2406(.VSS(VSS),.VDD(VDD),.Y(g34405),.A(g34183),.B(g25103));
  OR2 OR2_2407(.VSS(VSS),.VDD(VDD),.Y(g33235),.A(g32040),.B(g30982));
  OR2 OR2_2408(.VSS(VSS),.VDD(VDD),.Y(g23317),.A(g19715),.B(g16191));
  OR3 OR3_61(.VSS(VSS),.VDD(VDD),.Y(I22852),.A(g21459),.B(g21350),.C(g21339));
  OR2 OR2_2409(.VSS(VSS),.VDD(VDD),.Y(g29813),.A(g26020),.B(g28261));
  OR2 OR2_2410(.VSS(VSS),.VDD(VDD),.Y(g22679),.A(g19145),.B(g15701));
  OR2 OR2_2411(.VSS(VSS),.VDD(VDD),.Y(g23129),.A(g19500),.B(g15863));
  OR2 OR2_2412(.VSS(VSS),.VDD(VDD),.Y(g13699),.A(g10921),.B(g10947));
  OR2 OR2_2413(.VSS(VSS),.VDD(VDD),.Y(g34020),.A(g33904),.B(g18514));
  OR2 OR2_2414(.VSS(VSS),.VDD(VDD),.Y(g25731),.A(g25128),.B(g22014));
  OR2 OR2_2415(.VSS(VSS),.VDD(VDD),.Y(g28631),.A(g27372),.B(g16534));
  OR4 OR4_92(.VSS(VSS),.VDD(VDD),.Y(I28567),.A(g29204),.B(g29205),.C(g29206),.D(g29207));
  OR3 OR3_62(.VSS(VSS),.VDD(VDD),.Y(I24117),.A(g23088),.B(g23154),.C(g23172));
  OR2 OR2_2416(.VSS(VSS),.VDD(VDD),.Y(g32360),.A(g29868),.B(g31299));
  OR2 OR2_2417(.VSS(VSS),.VDD(VDD),.Y(g16506),.A(g13294),.B(g10966));
  OR2 OR2_2418(.VSS(VSS),.VDD(VDD),.Y(g15789),.A(g10819),.B(g13211));
  OR4 OR4_93(.VSS(VSS),.VDD(VDD),.Y(I30261),.A(g29385),.B(g31376),.C(g30735),.D(g30825));
  OR2 OR2_2419(.VSS(VSS),.VDD(VDD),.Y(g34046),.A(g33906),.B(g33908));
  OR2 OR2_2420(.VSS(VSS),.VDD(VDD),.Y(g31882),.A(g31115),.B(g21776));
  OR2 OR2_2421(.VSS(VSS),.VDD(VDD),.Y(g33991),.A(g33885),.B(g18400));
  OR2 OR2_2422(.VSS(VSS),.VDD(VDD),.Y(g14078),.A(g10776),.B(g8703));
  OR2 OR2_2423(.VSS(VSS),.VDD(VDD),.Y(g20196),.A(g16207),.B(g13497));
  OR2 OR2_2424(.VSS(VSS),.VDD(VDD),.Y(g25691),.A(g24536),.B(g21890));
  OR2 OR2_2425(.VSS(VSS),.VDD(VDD),.Y(g27487),.A(g25990),.B(g24629));
  OR2 OR2_2426(.VSS(VSS),.VDD(VDD),.Y(g34282),.A(g26838),.B(g34214));
  OR2 OR2_2427(.VSS(VSS),.VDD(VDD),.Y(g23298),.A(g19693),.B(g16179));
  OR2 OR2_2428(.VSS(VSS),.VDD(VDD),.Y(g30357),.A(g30107),.B(g18366));
  OR2 OR2_2429(.VSS(VSS),.VDD(VDD),.Y(g28309),.A(g27106),.B(g15796));
  OR2 OR2_2430(.VSS(VSS),.VDD(VDD),.Y(g32220),.A(g31139),.B(g29633));
  OR2 OR2_2431(.VSS(VSS),.VDD(VDD),.Y(g26881),.A(g26629),.B(g24187));
  OR2 OR2_2432(.VSS(VSS),.VDD(VDD),.Y(g16927),.A(g13524),.B(g11126));
  OR2 OR2_2433(.VSS(VSS),.VDD(VDD),.Y(g25929),.A(g24395),.B(g22193));
  OR2 OR2_2434(.VSS(VSS),.VDD(VDD),.Y(g28308),.A(g27105),.B(g15795));
  OR2 OR2_2435(.VSS(VSS),.VDD(VDD),.Y(g27278),.A(g15786),.B(g25921));
  OR2 OR2_2436(.VSS(VSS),.VDD(VDD),.Y(g29692),.A(g28197),.B(g10873));
  OR2 OR2_2437(.VSS(VSS),.VDD(VDD),.Y(g24457),.A(g10902),.B(g22400));
  OR2 OR2_2438(.VSS(VSS),.VDD(VDD),.Y(g14977),.A(g10776),.B(g8703));
  OR2 OR2_2439(.VSS(VSS),.VDD(VDD),.Y(g25583),.A(g21666),.B(g24153));
  OR2 OR2_2440(.VSS(VSS),.VDD(VDD),.Y(g33584),.A(g33406),.B(g18449));
  OR2 OR2_2441(.VSS(VSS),.VDD(VDD),.Y(g34640),.A(g34487),.B(g18723));
  OR2 OR2_2442(.VSS(VSS),.VDD(VDD),.Y(g19274),.A(g17753),.B(g14791));
  OR2 OR2_2443(.VSS(VSS),.VDD(VDD),.Y(g19593),.A(g17145),.B(g14210));
  OR2 OR2_2444(.VSS(VSS),.VDD(VDD),.Y(g34803),.A(g34758),.B(g18590));
  OR2 OR2_2445(.VSS(VSS),.VDD(VDD),.Y(g28816),.A(g27547),.B(g16843));
  OR2 OR2_2446(.VSS(VSS),.VDD(VDD),.Y(g20077),.A(g16025),.B(g13320));
  OR2 OR2_2447(.VSS(VSS),.VDD(VDD),.Y(g23261),.A(g19660),.B(g16125));
  OR2 OR2_2448(.VSS(VSS),.VDD(VDD),.Y(g26890),.A(g26630),.B(g24196));
  OR2 OR2_2449(.VSS(VSS),.VDD(VDD),.Y(g28687),.A(g27434),.B(g16638));
  OR2 OR2_2450(.VSS(VSS),.VDD(VDD),.Y(g29539),.A(g2864),.B(g28220));
  OR2 OR2_2451(.VSS(VSS),.VDD(VDD),.Y(g32355),.A(g29855),.B(g31286));
  OR2 OR2_2452(.VSS(VSS),.VDD(VDD),.Y(g34881),.A(g34866),.B(g18187));
  OR2 OR2_2453(.VSS(VSS),.VDD(VDD),.Y(g24256),.A(g22873),.B(g18309));
  OR2 OR2_2454(.VSS(VSS),.VDD(VDD),.Y(g32370),.A(g29882),.B(g31312));
  OR2 OR2_2455(.VSS(VSS),.VDD(VDD),.Y(g28374),.A(g27181),.B(g15850));
  OR2 OR2_2456(.VSS(VSS),.VDD(VDD),.Y(g24280),.A(g23292),.B(g15109));
  OR2 OR2_2457(.VSS(VSS),.VDD(VDD),.Y(g25743),.A(g25110),.B(g22058));
  OR2 OR2_2458(.VSS(VSS),.VDD(VDD),.Y(g28643),.A(g27386),.B(g16592));
  OR2 OR2_2459(.VSS(VSS),.VDD(VDD),.Y(g27937),.A(g14506),.B(g26793));
  OR2 OR2_2460(.VSS(VSS),.VDD(VDD),.Y(g32996),.A(g32256),.B(g18377));
  OR2 OR2_2461(.VSS(VSS),.VDD(VDD),.Y(g34027),.A(g33718),.B(g18683));
  OR2 OR2_2462(.VSS(VSS),.VDD(VDD),.Y(g29241),.A(g28638),.B(g18332));
  OR2 OR2_2463(.VSS(VSS),.VDD(VDD),.Y(g13385),.A(g11967),.B(g9479));
//
  NAND2 NAND2_0(.VSS(VSS),.VDD(VDD),.Y(g11980),.A(I14817),.B(I14818));
  NAND2 NAND2_1(.VSS(VSS),.VDD(VDD),.Y(g13889),.A(g11566),.B(g11435));
  NAND2 NAND2_2(.VSS(VSS),.VDD(VDD),.Y(g13980),.A(g10295),.B(g11435));
  NAND2 NAND2_3(.VSS(VSS),.VDD(VDD),.Y(g12169),.A(g9804),.B(g5448));
  NAND2 NAND2_4(.VSS(VSS),.VDD(VDD),.Y(I22761),.A(g11939),.B(I22760));
  NAND2 NAND2_5(.VSS(VSS),.VDD(VDD),.Y(I13443),.A(g262),.B(I13442));
  NAND2 NAND2_6(.VSS(VSS),.VDD(VDD),.Y(I14185),.A(g8442),.B(g3470));
  NAND4 NAND4_0(.VSS(VSS),.VDD(VDD),.Y(g16719),.A(g3243),.B(g13700),.C(g3310),.D(g11350));
  NAND2 NAND2_7(.VSS(VSS),.VDD(VDD),.Y(I14518),.A(g661),.B(I14516));
  NAND4 NAND4_1(.VSS(VSS),.VDD(VDD),.Y(g10224),.A(g6661),.B(g6704),.C(g6675),.D(g6697));
  NAND2 NAND2_8(.VSS(VSS),.VDD(VDD),.Y(g17595),.A(g8616),.B(g14367));
  NAND2 NAND2_9(.VSS(VSS),.VDD(VDD),.Y(g22984),.A(g20114),.B(g2868));
  NAND2 NAND2_10(.VSS(VSS),.VDD(VDD),.Y(I12346),.A(g3111),.B(I12344));
  NAND2 NAND2_11(.VSS(VSS),.VDD(VDD),.Y(g12478),.A(I15299),.B(I15300));
  NAND4 NAND4_2(.VSS(VSS),.VDD(VDD),.Y(g21432),.A(g17790),.B(g14820),.C(g17761),.D(g14780));
  NAND3 NAND3_0(.VSS(VSS),.VDD(VDD),.Y(g28830),.A(g27886),.B(g7451),.C(g7369));
  NAND2 NAND2_12(.VSS(VSS),.VDD(VDD),.Y(I14883),.A(g9500),.B(g5489));
  NAND2 NAND2_13(.VSS(VSS),.VDD(VDD),.Y(g19474),.A(g11609),.B(g17794));
  NAND2 NAND2_14(.VSS(VSS),.VDD(VDD),.Y(g11426),.A(g8742),.B(g4878));
  NAND2 NAND2_15(.VSS(VSS),.VDD(VDD),.Y(g11190),.A(g8539),.B(g3447));
  NAND2 NAND2_16(.VSS(VSS),.VDD(VDD),.Y(g9852),.A(g3684),.B(g4871));
  NAND2 NAND2_17(.VSS(VSS),.VDD(VDD),.Y(g23342),.A(g6928),.B(g21163));
  NAND2 NAND2_18(.VSS(VSS),.VDD(VDD),.Y(g27223),.A(I25908),.B(I25909));
  NAND2 NAND2_19(.VSS(VSS),.VDD(VDD),.Y(I15089),.A(g2393),.B(I15087));
  NAND2 NAND2_20(.VSS(VSS),.VDD(VDD),.Y(g22853),.A(g20219),.B(g2922));
  NAND2 NAND2_21(.VSS(VSS),.VDD(VDD),.Y(g25003),.A(g21353),.B(g23462));
  NAND2 NAND2_22(.VSS(VSS),.VDD(VDD),.Y(I15088),.A(g9832),.B(I15087));
  NAND2 NAND2_23(.VSS(VSS),.VDD(VDD),.Y(g24916),.A(g19450),.B(g23154));
  NAND2 NAND2_24(.VSS(VSS),.VDD(VDD),.Y(g25779),.A(g19694),.B(g24362));
  NAND2 NAND2_25(.VSS(VSS),.VDD(VDD),.Y(g12084),.A(g2342),.B(g8211));
  NAND3 NAND3_1(.VSS(VSS),.VDD(VDD),.Y(g28270),.A(g10504),.B(g26105),.C(g26987));
  NAND2 NAND2_26(.VSS(VSS),.VDD(VDD),.Y(g22836),.A(g18918),.B(g2852));
  NAND2 NAND2_27(.VSS(VSS),.VDD(VDD),.Y(g21330),.A(g11401),.B(g17157));
  NAND2 NAND2_28(.VSS(VSS),.VDD(VDD),.Y(g20076),.A(g13795),.B(g16521));
  NAND4 NAND4_3(.VSS(VSS),.VDD(VDD),.Y(g21365),.A(g15744),.B(g13119),.C(g15730),.D(g13100));
  NAND2 NAND2_29(.VSS(VSS),.VDD(VDD),.Y(g23132),.A(g8155),.B(g19932));
  NAND2 NAND2_30(.VSS(VSS),.VDD(VDD),.Y(I22683),.A(g11893),.B(g21434));
  NAND2 NAND2_31(.VSS(VSS),.VDD(VDD),.Y(g28938),.A(g27796),.B(g8205));
  NAND2 NAND2_32(.VSS(VSS),.VDD(VDD),.Y(g9825),.A(I13391),.B(I13392));
  NAND2 NAND2_33(.VSS(VSS),.VDD(VDD),.Y(g7201),.A(I11865),.B(I11866));
  NAND4 NAND4_4(.VSS(VSS),.VDD(VDD),.Y(g15719),.A(g5256),.B(g14490),.C(g5335),.D(g9780));
  NAND3 NAND3_2(.VSS(VSS),.VDD(VDD),.Y(g27654),.A(g164),.B(g26598),.C(g23042));
  NAND2 NAND2_34(.VSS(VSS),.VDD(VDD),.Y(g22864),.A(g7780),.B(g21156));
  NAND2 NAND2_35(.VSS(VSS),.VDD(VDD),.Y(I20165),.A(g16246),.B(g990));
  NAND2 NAND2_36(.VSS(VSS),.VDD(VDD),.Y(g14489),.A(g12126),.B(g5084));
  NAND2 NAND2_37(.VSS(VSS),.VDD(VDD),.Y(g29082),.A(g27837),.B(g9694));
  NAND2 NAND2_38(.VSS(VSS),.VDD(VDD),.Y(g25233),.A(g20838),.B(g23623));
  NAND2 NAND2_39(.VSS(VSS),.VDD(VDD),.Y(g24942),.A(g20039),.B(g23172));
  NAND2 NAND2_40(.VSS(VSS),.VDD(VDD),.Y(I26459),.A(g26576),.B(g14306));
  NAND3 NAND3_3(.VSS(VSS),.VDD(VDD),.Y(g15832),.A(g7903),.B(g7479),.C(g13256));
  NAND4 NAND4_5(.VSS(VSS),.VDD(VDD),.Y(g14830),.A(g6605),.B(g12211),.C(g6723),.D(g12721));
  NAND2 NAND2_41(.VSS(VSS),.VDD(VDD),.Y(I32431),.A(g34056),.B(g34051));
  NAND2 NAND2_42(.VSS(VSS),.VDD(VDD),.Y(g9972),.A(I13510),.B(I13511));
  NAND2 NAND2_43(.VSS(VSS),.VDD(VDD),.Y(I20222),.A(g16272),.B(I20221));
  NAND3 NAND3_4(.VSS(VSS),.VDD(VDD),.Y(g17748),.A(g562),.B(g14708),.C(g12323));
  NAND2 NAND2_44(.VSS(VSS),.VDD(VDD),.Y(g11969),.A(g7252),.B(g1636));
  NAND2 NAND2_45(.VSS(VSS),.VDD(VDD),.Y(g20734),.A(g14408),.B(g17312));
  NAND3 NAND3_5(.VSS(VSS),.VDD(VDD),.Y(g28837),.A(g27800),.B(g7374),.C(g2197));
  NAND2 NAND2_46(.VSS(VSS),.VDD(VDD),.Y(I25244),.A(g24744),.B(I25242));
  NAND3 NAND3_6(.VSS(VSS),.VDD(VDD),.Y(g11968),.A(g837),.B(g9334),.C(g9086));
  NAND4 NAND4_6(.VSS(VSS),.VDD(VDD),.Y(g13968),.A(g3913),.B(g11255),.C(g4031),.D(g11631));
  NAND2 NAND2_47(.VSS(VSS),.VDD(VDD),.Y(g15045),.A(g12716),.B(g7142));
  NAND2 NAND2_48(.VSS(VSS),.VDD(VDD),.Y(g12423),.A(I15242),.B(I15243));
  NAND4 NAND4_7(.VSS(VSS),.VDD(VDD),.Y(g27587),.A(g24917),.B(g25018),.C(g24918),.D(g26857));
  NAND2 NAND2_49(.VSS(VSS),.VDD(VDD),.Y(g20838),.A(g5041),.B(g17284));
  NAND2 NAND2_50(.VSS(VSS),.VDD(VDD),.Y(g13855),.A(g4944),.B(g11804));
  NAND3 NAND3_7(.VSS(VSS),.VDD(VDD),.Y(g19483),.A(g15969),.B(g10841),.C(g10922));
  NAND2 NAND2_51(.VSS(VSS),.VDD(VDD),.Y(g10610),.A(g7462),.B(g7490));
  NAND2 NAND2_52(.VSS(VSS),.VDD(VDD),.Y(g11411),.A(g9713),.B(g3625));
  NAND2 NAND2_53(.VSS(VSS),.VDD(VDD),.Y(I13110),.A(g5808),.B(I13109));
  NAND2 NAND2_54(.VSS(VSS),.VDD(VDD),.Y(g22642),.A(g7870),.B(g19560));
  NAND2 NAND2_55(.VSS(VSS),.VDD(VDD),.Y(g12587),.A(g7497),.B(g6315));
  NAND2 NAND2_56(.VSS(VSS),.VDD(VDD),.Y(g13870),.A(g11773),.B(g4732));
  NAND4 NAND4_8(.VSS(VSS),.VDD(VDD),.Y(g13527),.A(g182),.B(g168),.C(g203),.D(g12812));
  NAND2 NAND2_57(.VSS(VSS),.VDD(VDD),.Y(g23810),.A(I22973),.B(I22974));
  NAND2 NAND2_58(.VSS(VSS),.VDD(VDD),.Y(g20619),.A(g14317),.B(g17217));
  NAND4 NAND4_9(.VSS(VSS),.VDD(VDD),.Y(g16628),.A(g3602),.B(g11207),.C(g3618),.D(g13902));
  NAND2 NAND2_59(.VSS(VSS),.VDD(VDD),.Y(I23119),.A(g20076),.B(I23118));
  NAND4 NAND4_10(.VSS(VSS),.VDD(VDD),.Y(g10124),.A(g5276),.B(g5320),.C(g5290),.D(g5313));
  NAND2 NAND2_60(.VSS(VSS),.VDD(VDD),.Y(g12000),.A(g8418),.B(g2610));
  NAND2 NAND2_61(.VSS(VSS),.VDD(VDD),.Y(I23118),.A(g20076),.B(g417));
  NAND2 NAND2_62(.VSS(VSS),.VDD(VDD),.Y(g22874),.A(g18918),.B(g2844));
  NAND2 NAND2_63(.VSS(VSS),.VDD(VDD),.Y(g10939),.A(g7352),.B(g1459));
  NAND2 NAND2_64(.VSS(VSS),.VDD(VDD),.Y(g13867),.A(g11312),.B(g8449));
  NAND4 NAND4_11(.VSS(VSS),.VDD(VDD),.Y(g14686),.A(g5268),.B(g12059),.C(g5276),.D(g12239));
  NAND2 NAND2_65(.VSS(VSS),.VDD(VDD),.Y(I12840),.A(g4222),.B(g4235));
  NAND2 NAND2_66(.VSS(VSS),.VDD(VDD),.Y(g29049),.A(g9640),.B(g27779));
  NAND4 NAND4_12(.VSS(VSS),.VDD(VDD),.Y(g16776),.A(g3945),.B(g13772),.C(g4012),.D(g11419));
  NAND2 NAND2_67(.VSS(VSS),.VDD(VDD),.Y(g13315),.A(g1459),.B(g10715));
  NAND2 NAND2_68(.VSS(VSS),.VDD(VDD),.Y(g11707),.A(g8718),.B(g4864));
  NAND2 NAND2_69(.VSS(VSS),.VDD(VDD),.Y(I18530),.A(g1811),.B(I18529));
  NAND2 NAND2_70(.VSS(VSS),.VDD(VDD),.Y(g20039),.A(g11250),.B(g17794));
  NAND2 NAND2_71(.VSS(VSS),.VDD(VDD),.Y(I14609),.A(g8993),.B(g8678));
  NAND2 NAND2_72(.VSS(VSS),.VDD(VDD),.Y(I13334),.A(g1687),.B(g1691));
  NAND2 NAND2_73(.VSS(VSS),.VDD(VDD),.Y(g13257),.A(g1389),.B(g10544));
  NAND2 NAND2_74(.VSS(VSS),.VDD(VDD),.Y(g29004),.A(g27933),.B(g8330));
  NAND4 NAND4_13(.VSS(VSS),.VDD(VDD),.Y(g21459),.A(g17814),.B(g14854),.C(g17605),.D(g17581));
  NAND2 NAND2_75(.VSS(VSS),.VDD(VDD),.Y(g11979),.A(g9861),.B(g5452));
  NAND3 NAND3_8(.VSS(VSS),.VDD(VDD),.Y(g13496),.A(g1351),.B(g11336),.C(g11815));
  NAND3 NAND3_9(.VSS(VSS),.VDD(VDD),.Y(g11590),.A(g6928),.B(g3990),.C(g4049));
  NAND3 NAND3_10(.VSS(VSS),.VDD(VDD),.Y(g12639),.A(g10194),.B(g6682),.C(g6732));
  NAND2 NAND2_76(.VSS(VSS),.VDD(VDD),.Y(g22712),.A(g18957),.B(g2864));
  NAND2 NAND2_77(.VSS(VSS),.VDD(VDD),.Y(g23010),.A(g20516),.B(g2984));
  NAND2 NAND2_78(.VSS(VSS),.VDD(VDD),.Y(g7897),.A(I12288),.B(I12289));
  NAND2 NAND2_79(.VSS(VSS),.VDD(VDD),.Y(g24601),.A(g22957),.B(g2965));
  NAND2 NAND2_80(.VSS(VSS),.VDD(VDD),.Y(g13986),.A(g10323),.B(g11747));
  NAND2 NAND2_81(.VSS(VSS),.VDD(VDD),.Y(g12293),.A(g7436),.B(g5283));
  NAND2 NAND2_82(.VSS(VSS),.VDD(VDD),.Y(g24677),.A(g22957),.B(g2975));
  NAND2 NAND2_83(.VSS(VSS),.VDD(VDD),.Y(g12638),.A(g7514),.B(g6661));
  NAND2 NAND2_84(.VSS(VSS),.VDD(VDD),.Y(g24975),.A(g21388),.B(g23363));
  NAND4 NAND4_14(.VSS(VSS),.VDD(VDD),.Y(g10160),.A(g5623),.B(g5666),.C(g5637),.D(g5659));
  NAND4 NAND4_15(.VSS(VSS),.VDD(VDD),.Y(g17712),.A(g5599),.B(g14425),.C(g5666),.D(g12301));
  NAND3 NAND3_11(.VSS(VSS),.VDD(VDD),.Y(g12416),.A(g10133),.B(g7064),.C(g10166));
  NAND2 NAND2_85(.VSS(VSS),.VDD(VDD),.Y(g14160),.A(g11626),.B(g8958));
  NAND3 NAND3_12(.VSS(VSS),.VDD(VDD),.Y(g28853),.A(g27742),.B(g1636),.C(g7252));
  NAND4 NAND4_16(.VSS(VSS),.VDD(VDD),.Y(g13067),.A(g5240),.B(g12059),.C(g5331),.D(g9780));
  NAND2 NAND2_86(.VSS(VSS),.VDD(VDD),.Y(g28167),.A(g925),.B(g27046));
  NAND2 NAND2_87(.VSS(VSS),.VDD(VDD),.Y(I18635),.A(g14713),.B(I18633));
  NAND2 NAND2_88(.VSS(VSS),.VDD(VDD),.Y(g10617),.A(g10151),.B(g9909));
  NAND3 NAND3_13(.VSS(VSS),.VDD(VDD),.Y(g16319),.A(g8224),.B(g8170),.C(g13736));
  NAND2 NAND2_89(.VSS(VSS),.VDD(VDD),.Y(I32187),.A(g33661),.B(I32185));
  NAND2 NAND2_90(.VSS(VSS),.VDD(VDD),.Y(I12252),.A(g1124),.B(I12251));
  NAND2 NAND2_91(.VSS(VSS),.VDD(VDD),.Y(g14915),.A(g12553),.B(g10266));
  NAND2 NAND2_92(.VSS(VSS),.VDD(VDD),.Y(g22941),.A(g20219),.B(g2970));
  NAND2 NAND2_93(.VSS(VSS),.VDD(VDD),.Y(I17406),.A(g1472),.B(I17404));
  NAND2 NAND2_94(.VSS(VSS),.VDD(VDD),.Y(g12578),.A(g7791),.B(g10341));
  NAND4 NAND4_17(.VSS(VSS),.VDD(VDD),.Y(g27586),.A(g24924),.B(g24916),.C(g24905),.D(g26863));
  NAND2 NAND2_95(.VSS(VSS),.VDD(VDD),.Y(g12014),.A(g7197),.B(g703));
  NAND2 NAND2_96(.VSS(VSS),.VDD(VDD),.Y(g14075),.A(g11658),.B(g11527));
  NAND3 NAND3_14(.VSS(VSS),.VDD(VDD),.Y(g15591),.A(g4332),.B(g4322),.C(g13202));
  NAND3 NAND3_15(.VSS(VSS),.VDD(VDD),.Y(g28864),.A(g27886),.B(g7411),.C(g1996));
  NAND2 NAND2_97(.VSS(VSS),.VDD(VDD),.Y(g10623),.A(g10181),.B(g9976));
  NAND4 NAND4_18(.VSS(VSS),.VDD(VDD),.Y(g17675),.A(g5252),.B(g14399),.C(g5320),.D(g12239));
  NAND2 NAND2_98(.VSS(VSS),.VDD(VDD),.Y(g23656),.A(I22800),.B(I22801));
  NAND2 NAND2_99(.VSS(VSS),.VDD(VDD),.Y(g21353),.A(g11467),.B(g17157));
  NAND2 NAND2_100(.VSS(VSS),.VDD(VDD),.Y(I13751),.A(g4584),.B(I13749));
  NAND2 NAND2_101(.VSS(VSS),.VDD(VDD),.Y(g14782),.A(g12755),.B(g10491));
  NAND2 NAND2_102(.VSS(VSS),.VDD(VDD),.Y(I14400),.A(g3654),.B(I14398));
  NAND2 NAND2_103(.VSS(VSS),.VDD(VDD),.Y(g12116),.A(g2051),.B(g8255));
  NAND2 NAND2_104(.VSS(VSS),.VDD(VDD),.Y(g14984),.A(g7812),.B(g12680));
  NAND4 NAND4_19(.VSS(VSS),.VDD(VDD),.Y(g13866),.A(g3239),.B(g11194),.C(g3321),.D(g11519));
  NAND2 NAND2_105(.VSS(VSS),.VDD(VDD),.Y(I18537),.A(g2236),.B(I18536));
  NAND3 NAND3_16(.VSS(VSS),.VDD(VDD),.Y(g16281),.A(g4754),.B(g13937),.C(g12054));
  NAND3 NAND3_17(.VSS(VSS),.VDD(VDD),.Y(g28900),.A(g27886),.B(g7451),.C(g2040));
  NAND2 NAND2_106(.VSS(VSS),.VDD(VDD),.Y(g14822),.A(g12755),.B(g12632));
  NAND2 NAND2_107(.VSS(VSS),.VDD(VDD),.Y(g14170),.A(g11715),.B(g11537));
  NAND3 NAND3_18(.VSS(VSS),.VDD(VDD),.Y(g15844),.A(g14714),.B(g9340),.C(g12378));
  NAND2 NAND2_108(.VSS(VSS),.VDD(VDD),.Y(I22972),.A(g9657),.B(g19638));
  NAND4 NAND4_20(.VSS(VSS),.VDD(VDD),.Y(g21364),.A(g15787),.B(g15781),.C(g15753),.D(g13131));
  NAND2 NAND2_109(.VSS(VSS),.VDD(VDD),.Y(I13391),.A(g1821),.B(I13390));
  NAND3 NAND3_19(.VSS(VSS),.VDD(VDD),.Y(g13256),.A(g11846),.B(g11294),.C(g11812));
  NAND2 NAND2_110(.VSS(VSS),.VDD(VDD),.Y(I13510),.A(g2089),.B(I13509));
  NAND2 NAND2_111(.VSS(VSS),.VDD(VDD),.Y(g11923),.A(I14734),.B(I14735));
  NAND2 NAND2_112(.VSS(VSS),.VDD(VDD),.Y(g12340),.A(g4888),.B(g8984));
  NAND2 NAND2_113(.VSS(VSS),.VDD(VDD),.Y(g12035),.A(g10000),.B(g6144));
  NAND2 NAND2_114(.VSS(VSS),.VDD(VDD),.Y(g13923),.A(g11692),.B(g11527));
  NAND2 NAND2_115(.VSS(VSS),.VDD(VDD),.Y(I15300),.A(g1982),.B(I15298));
  NAND2 NAND2_116(.VSS(VSS),.VDD(VDD),.Y(g9830),.A(I13402),.B(I13403));
  NAND2 NAND2_117(.VSS(VSS),.VDD(VDD),.Y(g20186),.A(g16926),.B(g8177));
  NAND2 NAND2_118(.VSS(VSS),.VDD(VDD),.Y(g20676),.A(g14379),.B(g17287));
  NAND2 NAND2_119(.VSS(VSS),.VDD(VDD),.Y(g21289),.A(g14616),.B(g17493));
  NAND2 NAND2_120(.VSS(VSS),.VDD(VDD),.Y(I12205),.A(g1135),.B(I12203));
  NAND2 NAND2_121(.VSS(VSS),.VDD(VDD),.Y(g13102),.A(g7523),.B(g10759));
  NAND3 NAND3_20(.VSS(VSS),.VDD(VDD),.Y(g25429),.A(g22417),.B(g1917),.C(g8302));
  NAND2 NAND2_122(.VSS(VSS),.VDD(VDD),.Y(g23309),.A(g6905),.B(g21024));
  NAND3 NAND3_21(.VSS(VSS),.VDD(VDD),.Y(g28874),.A(g27907),.B(g7424),.C(g2421));
  NAND2 NAND2_123(.VSS(VSS),.VDD(VDD),.Y(g29121),.A(g9755),.B(g27886));
  NAND2 NAND2_124(.VSS(VSS),.VDD(VDD),.Y(g21288),.A(g14616),.B(g17492));
  NAND2 NAND2_125(.VSS(VSS),.VDD(VDD),.Y(g7582),.A(g1361),.B(g1373));
  NAND2 NAND2_126(.VSS(VSS),.VDD(VDD),.Y(I13442),.A(g262),.B(g239));
  NAND3 NAND3_22(.VSS(VSS),.VDD(VDD),.Y(g13066),.A(g4430),.B(g7178),.C(g10590));
  NAND4 NAND4_21(.VSS(VSS),.VDD(VDD),.Y(g24936),.A(g20186),.B(g20173),.C(g23379),.D(g14029));
  NAND3 NAND3_23(.VSS(VSS),.VDD(VDD),.Y(g31262),.A(g767),.B(g29916),.C(g11679));
  NAND2 NAND2_127(.VSS(VSS),.VDD(VDD),.Y(g10022),.A(g6474),.B(g6466));
  NAND2 NAND2_128(.VSS(VSS),.VDD(VDD),.Y(g14864),.A(g7791),.B(g10421));
  NAND2 NAND2_129(.VSS(VSS),.VDD(VDD),.Y(g8769),.A(g691),.B(g714));
  NAND2 NAND2_130(.VSS(VSS),.VDD(VDD),.Y(g7227),.A(g4584),.B(g4593));
  NAND2 NAND2_131(.VSS(VSS),.VDD(VDD),.Y(I32186),.A(g33665),.B(I32185));
  NAND2 NAND2_132(.VSS(VSS),.VDD(VDD),.Y(g12523),.A(g7563),.B(g6346));
  NAND3 NAND3_24(.VSS(VSS),.VDD(VDD),.Y(g28892),.A(g27779),.B(g1772),.C(g7275));
  NAND2 NAND2_133(.VSS(VSS),.VDD(VDD),.Y(g13854),.A(g4765),.B(g11797));
  NAND2 NAND2_134(.VSS(VSS),.VDD(VDD),.Y(g11511),.A(I14481),.B(I14482));
  NAND2 NAND2_135(.VSS(VSS),.VDD(VDD),.Y(I14991),.A(g9685),.B(g6527));
  NAND2 NAND2_136(.VSS(VSS),.VDD(VDD),.Y(g8967),.A(g4264),.B(g4258));
  NAND4 NAND4_22(.VSS(VSS),.VDD(VDD),.Y(g13511),.A(g182),.B(g174),.C(g203),.D(g12812));
  NAND2 NAND2_137(.VSS(VSS),.VDD(VDD),.Y(g20216),.A(I20487),.B(I20488));
  NAND3 NAND3_25(.VSS(VSS),.VDD(VDD),.Y(g14254),.A(g11968),.B(g11933),.C(g11951));
  NAND3 NAND3_26(.VSS(VSS),.VDD(VDD),.Y(g28914),.A(g27937),.B(g7462),.C(g2555));
  NAND2 NAND2_138(.VSS(VSS),.VDD(VDD),.Y(g29134),.A(g9762),.B(g27907));
  NAND3 NAND3_27(.VSS(VSS),.VDD(VDD),.Y(g28907),.A(g27858),.B(g2361),.C(g2287));
  NAND2 NAND2_139(.VSS(VSS),.VDD(VDD),.Y(g12222),.A(g8310),.B(g2028));
  NAND2 NAND2_140(.VSS(VSS),.VDD(VDD),.Y(g29028),.A(g27933),.B(g8381));
  NAND2 NAND2_141(.VSS(VSS),.VDD(VDD),.Y(g22852),.A(g18957),.B(g2856));
  NAND2 NAND2_142(.VSS(VSS),.VDD(VDD),.Y(g14101),.A(g11653),.B(g11729));
  NAND2 NAND2_143(.VSS(VSS),.VDD(VDD),.Y(g25002),.A(g19474),.B(g23154));
  NAND2 NAND2_144(.VSS(VSS),.VDD(VDD),.Y(I29297),.A(g12117),.B(I29295));
  NAND3 NAND3_28(.VSS(VSS),.VDD(VDD),.Y(g14177),.A(g11741),.B(g11721),.C(g753));
  NAND2 NAND2_145(.VSS(VSS),.VDD(VDD),.Y(g11480),.A(g10323),.B(g8906));
  NAND2 NAND2_146(.VSS(VSS),.VDD(VDD),.Y(I26460),.A(g26576),.B(I26459));
  NAND2 NAND2_147(.VSS(VSS),.VDD(VDD),.Y(I22946),.A(g19620),.B(I22944));
  NAND2 NAND2_148(.VSS(VSS),.VDD(VDD),.Y(I18536),.A(g2236),.B(g14642));
  NAND2 NAND2_149(.VSS(VSS),.VDD(VDD),.Y(I15287),.A(g10061),.B(g6697));
  NAND2 NAND2_150(.VSS(VSS),.VDD(VDD),.Y(I14206),.A(g3821),.B(I14204));
  NAND4 NAND4_23(.VSS(VSS),.VDD(VDD),.Y(g16956),.A(g3925),.B(g13824),.C(g4019),.D(g11631));
  NAND2 NAND2_151(.VSS(VSS),.VDD(VDD),.Y(I26093),.A(g26055),.B(g13539));
  NAND2 NAND2_152(.VSS(VSS),.VDD(VDD),.Y(I15307),.A(g10116),.B(I15306));
  NAND2 NAND2_153(.VSS(VSS),.VDD(VDD),.Y(g23195),.A(g20136),.B(g37));
  NAND2 NAND2_154(.VSS(VSS),.VDD(VDD),.Y(g13307),.A(g1116),.B(g10695));
  NAND2 NAND2_155(.VSS(VSS),.VDD(VDD),.Y(I15243),.A(g6351),.B(I15241));
  NAND4 NAND4_24(.VSS(VSS),.VDD(VDD),.Y(g16181),.A(g13475),.B(g13495),.C(g13057),.D(g13459));
  NAND2 NAND2_156(.VSS(VSS),.VDD(VDD),.Y(g12351),.A(I15194),.B(I15195));
  NAND2 NAND2_157(.VSS(VSS),.VDD(VDD),.Y(g24814),.A(g20011),.B(g23167));
  NAND2 NAND2_158(.VSS(VSS),.VDD(VDD),.Y(g22312),.A(g907),.B(g19063));
  NAND3 NAND3_29(.VSS(VSS),.VDD(VDD),.Y(g28935),.A(g27800),.B(g2227),.C(g7328));
  NAND2 NAND2_159(.VSS(VSS),.VDD(VDD),.Y(g24807),.A(I23979),.B(I23980));
  NAND2 NAND2_160(.VSS(VSS),.VDD(VDD),.Y(I15341),.A(g10154),.B(I15340));
  NAND2 NAND2_161(.VSS(VSS),.VDD(VDD),.Y(g14665),.A(g12604),.B(g12798));
  NAND2 NAND2_162(.VSS(VSS),.VDD(VDD),.Y(g24974),.A(g21301),.B(g23363));
  NAND2 NAND2_163(.VSS(VSS),.VDD(VDD),.Y(g31997),.A(g22306),.B(g30580));
  NAND2 NAND2_164(.VSS(VSS),.VDD(VDD),.Y(g14008),.A(g11610),.B(g11435));
  NAND2 NAND2_165(.VSS(VSS),.VDD(VDD),.Y(I14399),.A(g8542),.B(I14398));
  NAND2 NAND2_166(.VSS(VSS),.VDD(VDD),.Y(I22760),.A(g11939),.B(g21434));
  NAND2 NAND2_167(.VSS(VSS),.VDD(VDD),.Y(g9258),.A(I13044),.B(I13045));
  NAND2 NAND2_168(.VSS(VSS),.VDD(VDD),.Y(g22921),.A(g20219),.B(g2950));
  NAND3 NAND3_30(.VSS(VSS),.VDD(VDD),.Y(g15715),.A(g336),.B(g305),.C(g13385));
  NAND2 NAND2_169(.VSS(VSS),.VDD(VDD),.Y(g17312),.A(g7297),.B(g14248));
  NAND2 NAND2_170(.VSS(VSS),.VDD(VDD),.Y(g25995),.A(g24621),.B(g22853));
  NAND2 NAND2_171(.VSS(VSS),.VDD(VDD),.Y(g14892),.A(g12700),.B(g12515));
  NAND4 NAND4_25(.VSS(VSS),.VDD(VDD),.Y(g17608),.A(g5953),.B(g12067),.C(g5969),.D(g14701));
  NAND2 NAND2_172(.VSS(VSS),.VDD(VDD),.Y(I14398),.A(g8542),.B(g3654));
  NAND2 NAND2_173(.VSS(VSS),.VDD(VDD),.Y(g15572),.A(g12969),.B(g7219));
  NAND2 NAND2_174(.VSS(VSS),.VDD(VDD),.Y(I18634),.A(g2504),.B(I18633));
  NAND2 NAND2_175(.VSS(VSS),.VDD(VDD),.Y(I15335),.A(g2116),.B(I15333));
  NAND2 NAND2_176(.VSS(VSS),.VDD(VDD),.Y(g34056),.A(I31984),.B(I31985));
  NAND4 NAND4_26(.VSS(VSS),.VDD(VDD),.Y(g14570),.A(g3933),.B(g11255),.C(g4023),.D(g8595));
  NAND2 NAND2_177(.VSS(VSS),.VDD(VDD),.Y(g11993),.A(g1894),.B(g8302));
  NAND4 NAND4_27(.VSS(VSS),.VDD(VDD),.Y(g13993),.A(g3961),.B(g11255),.C(g3969),.D(g11419));
  NAND2 NAND2_178(.VSS(VSS),.VDD(VDD),.Y(I23963),.A(g13631),.B(I23961));
  NAND2 NAND2_179(.VSS(VSS),.VDD(VDD),.Y(g9975),.A(I13519),.B(I13520));
  NAND2 NAND2_180(.VSS(VSS),.VDD(VDD),.Y(g21124),.A(g5731),.B(g17393));
  NAND2 NAND2_181(.VSS(VSS),.VDD(VDD),.Y(I14332),.A(g9966),.B(I14330));
  NAND2 NAND2_182(.VSS(VSS),.VDD(VDD),.Y(g13667),.A(g3723),.B(g11119));
  NAND4 NAND4_28(.VSS(VSS),.VDD(VDD),.Y(g13131),.A(g6243),.B(g12101),.C(g6377),.D(g10003));
  NAND2 NAND2_183(.VSS(VSS),.VDD(VDD),.Y(g10567),.A(g1862),.B(g7405));
  NAND2 NAND2_184(.VSS(VSS),.VDD(VDD),.Y(g20007),.A(g11512),.B(g17794));
  NAND2 NAND2_185(.VSS(VSS),.VDD(VDD),.Y(I23585),.A(g22409),.B(g4332));
  NAND4 NAND4_29(.VSS(VSS),.VDD(VDD),.Y(g28349),.A(g27074),.B(g24770),.C(g27187),.D(g19644));
  NAND2 NAND2_186(.VSS(VSS),.VDD(VDD),.Y(g29719),.A(g28406),.B(g13739));
  NAND2 NAND2_187(.VSS(VSS),.VDD(VDD),.Y(g21294),.A(g11324),.B(g17157));
  NAND3 NAND3_31(.VSS(VSS),.VDD(VDD),.Y(g25498),.A(g22498),.B(g2610),.C(g8418));
  NAND2 NAND2_188(.VSS(VSS),.VDD(VDD),.Y(g28906),.A(g27796),.B(g8150));
  NAND2 NAND2_189(.VSS(VSS),.VDD(VDD),.Y(g13210),.A(g7479),.B(g10521));
  NAND2 NAND2_190(.VSS(VSS),.VDD(VDD),.Y(g34650),.A(I32757),.B(I32758));
  NAND4 NAND4_30(.VSS(VSS),.VDD(VDD),.Y(g16625),.A(g3203),.B(g13700),.C(g3274),.D(g11519));
  NAND4 NAND4_31(.VSS(VSS),.VDD(VDD),.Y(g17732),.A(g3937),.B(g13824),.C(g4012),.D(g13933));
  NAND4 NAND4_32(.VSS(VSS),.VDD(VDD),.Y(g10185),.A(g5969),.B(g6012),.C(g5983),.D(g6005));
  NAND2 NAND2_191(.VSS(VSS),.VDD(VDD),.Y(g11443),.A(g9916),.B(g3649));
  NAND2 NAND2_192(.VSS(VSS),.VDD(VDD),.Y(g12436),.A(I15263),.B(I15264));
  NAND2 NAND2_193(.VSS(VSS),.VDD(VDD),.Y(g11279),.A(g8504),.B(g3443));
  NAND4 NAND4_33(.VSS(VSS),.VDD(VDD),.Y(g14519),.A(g3889),.B(g11225),.C(g4000),.D(g8595));
  NAND2 NAND2_194(.VSS(VSS),.VDD(VDD),.Y(I29296),.A(g29495),.B(I29295));
  NAND2 NAND2_195(.VSS(VSS),.VDD(VDD),.Y(g14675),.A(g12317),.B(g9898));
  NAND2 NAND2_196(.VSS(VSS),.VDD(VDD),.Y(I25219),.A(g482),.B(g24718));
  NAND4 NAND4_34(.VSS(VSS),.VDD(VDD),.Y(g27593),.A(g24972),.B(g24950),.C(g24906),.D(g26861));
  NAND2 NAND2_197(.VSS(VSS),.VDD(VDD),.Y(I26419),.A(g14247),.B(I26417));
  NAND2 NAND2_198(.VSS(VSS),.VDD(VDD),.Y(I22755),.A(g21434),.B(I22753));
  NAND2 NAND2_199(.VSS(VSS),.VDD(VDD),.Y(g12073),.A(g10058),.B(g6490));
  NAND2 NAND2_200(.VSS(VSS),.VDD(VDD),.Y(g14154),.A(g11669),.B(g8958));
  NAND4 NAND4_35(.VSS(VSS),.VDD(VDD),.Y(g17761),.A(g6291),.B(g14529),.C(g6358),.D(g12423));
  NAND2 NAND2_201(.VSS(VSS),.VDD(VDD),.Y(I26418),.A(g26519),.B(I26417));
  NAND2 NAND2_202(.VSS(VSS),.VDD(VDD),.Y(g13469),.A(g4983),.B(g10862));
  NAND2 NAND2_203(.VSS(VSS),.VDD(VDD),.Y(g25432),.A(g12374),.B(g22384));
  NAND2 NAND2_204(.VSS(VSS),.VDD(VDD),.Y(g10935),.A(g1459),.B(g7352));
  NAND2 NAND2_205(.VSS(VSS),.VDD(VDD),.Y(g14637),.A(g12255),.B(g9815));
  NAND2 NAND2_206(.VSS(VSS),.VDD(VDD),.Y(I15306),.A(g10116),.B(g2407));
  NAND2 NAND2_207(.VSS(VSS),.VDD(VDD),.Y(g16296),.A(g9360),.B(g13501));
  NAND2 NAND2_208(.VSS(VSS),.VDD(VDD),.Y(g25271),.A(I24462),.B(I24463));
  NAND2 NAND2_209(.VSS(VSS),.VDD(VDD),.Y(g7133),.A(I11825),.B(I11826));
  NAND3 NAND3_32(.VSS(VSS),.VDD(VDD),.Y(g12464),.A(g10169),.B(g7087),.C(g10191));
  NAND2 NAND2_210(.VSS(VSS),.VDD(VDD),.Y(g7846),.A(g4843),.B(g4878));
  NAND4 NAND4_36(.VSS(VSS),.VDD(VDD),.Y(g12797),.A(g10275),.B(g7655),.C(g7643),.D(g7627));
  NAND2 NAND2_211(.VSS(VSS),.VDD(VDD),.Y(I22794),.A(g21434),.B(I22792));
  NAND2 NAND2_212(.VSS(VSS),.VDD(VDD),.Y(I22845),.A(g12113),.B(I22844));
  NAND2 NAND2_213(.VSS(VSS),.VDD(VDD),.Y(g7803),.A(I12204),.B(I12205));
  NAND2 NAND2_214(.VSS(VSS),.VDD(VDD),.Y(g31950),.A(g7285),.B(g30573));
  NAND2 NAND2_215(.VSS(VSS),.VDD(VDD),.Y(g12292),.A(g4698),.B(g8933));
  NAND2 NAND2_216(.VSS(VSS),.VDD(VDD),.Y(g9461),.A(I13140),.B(I13141));
  NAND2 NAND2_217(.VSS(VSS),.VDD(VDD),.Y(g12153),.A(g2610),.B(g8330));
  NAND2 NAND2_218(.VSS(VSS),.VDD(VDD),.Y(g25199),.A(I24364),.B(I24365));
  NAND2 NAND2_219(.VSS(VSS),.VDD(VDD),.Y(I22899),.A(g12193),.B(g21228));
  NAND2 NAND2_220(.VSS(VSS),.VDD(VDD),.Y(g8829),.A(g5011),.B(g4836));
  NAND2 NAND2_221(.VSS(VSS),.VDD(VDD),.Y(g11975),.A(g8267),.B(g8316));
  NAND2 NAND2_222(.VSS(VSS),.VDD(VDD),.Y(I12204),.A(g1094),.B(I12203));
  NAND3 NAND3_33(.VSS(VSS),.VDD(VDD),.Y(g19513),.A(g15969),.B(g10841),.C(g10922));
  NAND2 NAND2_223(.VSS(VSS),.VDD(VDD),.Y(g23617),.A(I22761),.B(I22762));
  NAND2 NAND2_224(.VSS(VSS),.VDD(VDD),.Y(g15024),.A(g12780),.B(g10421));
  NAND2 NAND2_225(.VSS(VSS),.VDD(VDD),.Y(I20205),.A(g11147),.B(I20203));
  NAND2 NAND2_226(.VSS(VSS),.VDD(VDD),.Y(g12136),.A(I14992),.B(I14993));
  NAND2 NAND2_227(.VSS(VSS),.VDD(VDD),.Y(I22719),.A(g21434),.B(I22717));
  NAND2 NAND2_228(.VSS(VSS),.VDD(VDD),.Y(g9904),.A(I13443),.B(I13444));
  NAND4 NAND4_37(.VSS(VSS),.VDD(VDD),.Y(g13143),.A(g10695),.B(g7661),.C(g979),.D(g1061));
  NAND2 NAND2_229(.VSS(VSS),.VDD(VDD),.Y(I13453),.A(g1955),.B(I13452));
  NAND2 NAND2_230(.VSS(VSS),.VDD(VDD),.Y(I22718),.A(g11916),.B(I22717));
  NAND3 NAND3_34(.VSS(VSS),.VDD(VDD),.Y(g33394),.A(g10159),.B(g4474),.C(g32426));
  NAND2 NAND2_231(.VSS(VSS),.VDD(VDD),.Y(g11169),.A(I14229),.B(I14230));
  NAND2 NAND2_232(.VSS(VSS),.VDD(VDD),.Y(I29315),.A(g12154),.B(I29313));
  NAND2 NAND2_233(.VSS(VSS),.VDD(VDD),.Y(I15168),.A(g9823),.B(I15166));
  NAND2 NAND2_234(.VSS(VSS),.VDD(VDD),.Y(g13884),.A(g11797),.B(g4727));
  NAND3 NAND3_35(.VSS(VSS),.VDD(VDD),.Y(g11410),.A(g6875),.B(g6895),.C(g8696));
  NAND2 NAND2_235(.VSS(VSS),.VDD(VDD),.Y(g23623),.A(g9364),.B(g20717));
  NAND2 NAND2_236(.VSS(VSS),.VDD(VDD),.Y(g9391),.A(I13110),.B(I13111));
  NAND2 NAND2_237(.VSS(VSS),.VDD(VDD),.Y(I15363),.A(g10182),.B(g2675));
  NAND2 NAND2_238(.VSS(VSS),.VDD(VDD),.Y(g8124),.A(I12402),.B(I12403));
  NAND2 NAND2_239(.VSS(VSS),.VDD(VDD),.Y(g24362),.A(g21370),.B(g22136));
  NAND3 NAND3_36(.VSS(VSS),.VDD(VDD),.Y(g11479),.A(g6875),.B(g3288),.C(g3347));
  NAND2 NAND2_240(.VSS(VSS),.VDD(VDD),.Y(g23782),.A(g2741),.B(g21062));
  NAND2 NAND2_241(.VSS(VSS),.VDD(VDD),.Y(g13666),.A(g11190),.B(g8441));
  NAND4 NAND4_38(.VSS(VSS),.VDD(VDD),.Y(g13479),.A(g12686),.B(g12639),.C(g12590),.D(g12526));
  NAND2 NAND2_242(.VSS(VSS),.VDD(VDD),.Y(g8069),.A(I12373),.B(I12374));
  NAND2 NAND2_243(.VSS(VSS),.VDD(VDD),.Y(I32517),.A(g34424),.B(I32516));
  NAND2 NAND2_244(.VSS(VSS),.VDD(VDD),.Y(g13217),.A(g4082),.B(g10808));
  NAND2 NAND2_245(.VSS(VSS),.VDD(VDD),.Y(g10622),.A(g10178),.B(g9973));
  NAND2 NAND2_246(.VSS(VSS),.VDD(VDD),.Y(g10566),.A(g7315),.B(g7356));
  NAND4 NAND4_39(.VSS(VSS),.VDD(VDD),.Y(g13478),.A(g12511),.B(g12460),.C(g12414),.D(g12344));
  NAND2 NAND2_247(.VSS(VSS),.VDD(VDD),.Y(I13565),.A(g2648),.B(I13564));
  NAND2 NAND2_248(.VSS(VSS),.VDD(VDD),.Y(I13464),.A(g2384),.B(I13462));
  NAND3 NAND3_37(.VSS(VSS),.VDD(VDD),.Y(g13486),.A(g10862),.B(g4983),.C(g4966));
  NAND2 NAND2_249(.VSS(VSS),.VDD(VDD),.Y(g25258),.A(I24439),.B(I24440));
  NAND2 NAND2_250(.VSS(VSS),.VDD(VDD),.Y(g23266),.A(g18918),.B(g2894));
  NAND4 NAND4_40(.VSS(VSS),.VDD(VDD),.Y(g13580),.A(g11849),.B(g7503),.C(g7922),.D(g10544));
  NAND2 NAND2_251(.VSS(VSS),.VDD(VDD),.Y(g10653),.A(g10204),.B(g10042));
  NAND2 NAND2_252(.VSS(VSS),.VDD(VDD),.Y(g14139),.A(g11626),.B(g11584));
  NAND4 NAND4_41(.VSS(VSS),.VDD(VDD),.Y(g16741),.A(g3207),.B(g13765),.C(g3303),.D(g11519));
  NAND2 NAND2_253(.VSS(VSS),.VDD(VDD),.Y(I14789),.A(g9891),.B(I14788));
  NAND2 NAND2_254(.VSS(VSS),.VDD(VDD),.Y(g23167),.A(g8219),.B(g19981));
  NAND4 NAND4_42(.VSS(VSS),.VDD(VDD),.Y(g13084),.A(g5587),.B(g12093),.C(g5677),.D(g9864));
  NAND3 NAND3_38(.VSS(VSS),.VDD(VDD),.Y(g28973),.A(g27907),.B(g2465),.C(g7387));
  NAND4 NAND4_43(.VSS(VSS),.VDD(VDD),.Y(g14636),.A(g5595),.B(g12029),.C(g5677),.D(g12563));
  NAND2 NAND2_255(.VSS(VSS),.VDD(VDD),.Y(I14788),.A(g9891),.B(g6167));
  NAND4 NAND4_44(.VSS(VSS),.VDD(VDD),.Y(g14333),.A(g12042),.B(g12014),.C(g11990),.D(g11892));
  NAND2 NAND2_256(.VSS(VSS),.VDD(VDD),.Y(I17462),.A(g1300),.B(I17460));
  NAND4 NAND4_45(.VSS(VSS),.VDD(VDD),.Y(g21401),.A(g17755),.B(g14730),.C(g17712),.D(g14695));
  NAND4 NAND4_46(.VSS(VSS),.VDD(VDD),.Y(g27796),.A(g21228),.B(g25263),.C(g26424),.D(g26171));
  NAND4 NAND4_47(.VSS(VSS),.VDD(VDD),.Y(g20236),.A(g16875),.B(g14014),.C(g16625),.D(g16604));
  NAND2 NAND2_257(.VSS(VSS),.VDD(VDD),.Y(g12796),.A(g4467),.B(g6961));
  NAND2 NAND2_258(.VSS(VSS),.VDD(VDD),.Y(g9654),.A(g2485),.B(g2453));
  NAND3 NAND3_39(.VSS(VSS),.VDD(VDD),.Y(g15867),.A(g14714),.B(g9417),.C(g9340));
  NAND3 NAND3_40(.VSS(VSS),.VDD(VDD),.Y(g25337),.A(g22342),.B(g1648),.C(g8187));
  NAND2 NAND2_259(.VSS(VSS),.VDD(VDD),.Y(g28934),.A(g27882),.B(g14641));
  NAND4 NAND4_48(.VSS(VSS),.VDD(VDD),.Y(g14664),.A(g5220),.B(g12059),.C(g5339),.D(g12497));
  NAND4 NAND4_49(.VSS(VSS),.VDD(VDD),.Y(g16196),.A(g13496),.B(g13513),.C(g13079),.D(g13476));
  NAND4 NAND4_50(.VSS(VSS),.VDD(VDD),.Y(g11676),.A(g358),.B(g8944),.C(g376),.D(g385));
  NAND3 NAND3_41(.VSS(VSS),.VDD(VDD),.Y(g34545),.A(g11679),.B(g794),.C(g34354));
  NAND2 NAND2_260(.VSS(VSS),.VDD(VDD),.Y(I22871),.A(g12150),.B(g21228));
  NAND2 NAND2_261(.VSS(VSS),.VDD(VDD),.Y(g11953),.A(g8195),.B(g8241));
  NAND2 NAND2_262(.VSS(VSS),.VDD(VDD),.Y(g13676),.A(g11834),.B(g11283));
  NAND2 NAND2_263(.VSS(VSS),.VDD(VDD),.Y(g23616),.A(I22754),.B(I22755));
  NAND2 NAND2_264(.VSS(VSS),.VDD(VDD),.Y(g29355),.A(g24383),.B(g28109));
  NAND2 NAND2_265(.VSS(VSS),.VDD(VDD),.Y(g15581),.A(g7232),.B(g12999));
  NAND2 NAND2_266(.VSS(VSS),.VDD(VDD),.Y(g10585),.A(g1996),.B(g7451));
  NAND2 NAND2_267(.VSS(VSS),.VDD(VDD),.Y(g9595),.A(g2351),.B(g2319));
  NAND2 NAND2_268(.VSS(VSS),.VDD(VDD),.Y(g23748),.A(I22872),.B(I22873));
  NAND2 NAND2_269(.VSS(VSS),.VDD(VDD),.Y(I14291),.A(g3835),.B(I14289));
  NAND2 NAND2_270(.VSS(VSS),.VDD(VDD),.Y(g11936),.A(g8241),.B(g1783));
  NAND2 NAND2_271(.VSS(VSS),.VDD(VDD),.Y(I15334),.A(g10152),.B(I15333));
  NAND2 NAND2_272(.VSS(VSS),.VDD(VDD),.Y(g12192),.A(g8267),.B(g2319));
  NAND2 NAND2_273(.VSS(VSS),.VDD(VDD),.Y(g10609),.A(g10111),.B(g9826));
  NAND2 NAND2_274(.VSS(VSS),.VDD(VDD),.Y(I13109),.A(g5808),.B(g5813));
  NAND2 NAND2_275(.VSS(VSS),.VDD(VDD),.Y(g22940),.A(g18918),.B(g2860));
  NAND2 NAND2_276(.VSS(VSS),.VDD(VDD),.Y(I12097),.A(g1339),.B(I12096));
  NAND2 NAND2_277(.VSS(VSS),.VDD(VDD),.Y(g25425),.A(g20081),.B(g23172));
  NAND3 NAND3_42(.VSS(VSS),.VDD(VDD),.Y(g12522),.A(g10133),.B(g5990),.C(g6040));
  NAND2 NAND2_278(.VSS(VSS),.VDD(VDD),.Y(g23809),.A(I22966),.B(I22967));
  NAND4 NAND4_51(.VSS(VSS),.VDD(VDD),.Y(g17744),.A(g6303),.B(g14529),.C(g6373),.D(g12672));
  NAND2 NAND2_279(.VSS(VSS),.VDD(VDD),.Y(I17447),.A(g13336),.B(I17446));
  NAND3 NAND3_43(.VSS(VSS),.VDD(VDD),.Y(g28207),.A(g12546),.B(g26131),.C(g27977));
  NAND3 NAND3_44(.VSS(VSS),.VDD(VDD),.Y(g17399),.A(g9626),.B(g9574),.C(g14535));
  NAND2 NAND2_280(.VSS(VSS),.VDD(VDD),.Y(g14921),.A(g12492),.B(g10266));
  NAND4 NAND4_52(.VSS(VSS),.VDD(VDD),.Y(g15741),.A(g5244),.B(g14490),.C(g5320),.D(g14631));
  NAND2 NAND2_281(.VSS(VSS),.VDD(VDD),.Y(I32516),.A(g34424),.B(g34422));
  NAND2 NAND2_282(.VSS(VSS),.VDD(VDD),.Y(g9629),.A(g6462),.B(g6466));
  NAND2 NAND2_283(.VSS(VSS),.VDD(VDD),.Y(I13750),.A(g4608),.B(I13749));
  NAND2 NAND2_284(.VSS(VSS),.VDD(VDD),.Y(g14813),.A(g7766),.B(g12824));
  NAND2 NAND2_285(.VSS(VSS),.VDD(VDD),.Y(g11543),.A(g9714),.B(g3969));
  NAND2 NAND2_286(.VSS(VSS),.VDD(VDD),.Y(I12850),.A(g4277),.B(I12848));
  NAND4 NAND4_53(.VSS(VSS),.VDD(VDD),.Y(g13909),.A(g11396),.B(g8847),.C(g11674),.D(g8803));
  NAND2 NAND2_287(.VSS(VSS),.VDD(VDD),.Y(g23733),.A(g20751),.B(g11178));
  NAND4 NAND4_54(.VSS(VSS),.VDD(VDD),.Y(g15735),.A(g5547),.B(g14425),.C(g5659),.D(g9864));
  NAND3 NAND3_45(.VSS(VSS),.VDD(VDD),.Y(g15877),.A(g14833),.B(g9340),.C(g12543));
  NAND2 NAND2_288(.VSS(VSS),.VDD(VDD),.Y(g9800),.A(g5436),.B(g5428));
  NAND4 NAND4_55(.VSS(VSS),.VDD(VDD),.Y(g14674),.A(g5941),.B(g12067),.C(g6023),.D(g12614));
  NAND3 NAND3_46(.VSS(VSS),.VDD(VDD),.Y(g11117),.A(g8087),.B(g8186),.C(g8239));
  NAND3 NAND3_47(.VSS(VSS),.VDD(VDD),.Y(g29025),.A(g27937),.B(g2629),.C(g7462));
  NAND2 NAND2_289(.VSS(VSS),.VDD(VDD),.Y(g13000),.A(g7228),.B(g10598));
  NAND2 NAND2_290(.VSS(VSS),.VDD(VDD),.Y(I22754),.A(g11937),.B(I22753));
  NAND2 NAND2_291(.VSS(VSS),.VDD(VDD),.Y(g29540),.A(g28336),.B(g13464));
  NAND2 NAND2_292(.VSS(VSS),.VDD(VDD),.Y(g23630),.A(g20739),.B(g11123));
  NAND3 NAND3_48(.VSS(VSS),.VDD(VDD),.Y(g22833),.A(g1193),.B(g19560),.C(g10666));
  NAND2 NAND2_293(.VSS(VSS),.VDD(VDD),.Y(g15695),.A(g1266),.B(g13125));
  NAND2 NAND2_294(.VSS(VSS),.VDD(VDD),.Y(g25532),.A(g21360),.B(g23363));
  NAND2 NAND2_295(.VSS(VSS),.VDD(VDD),.Y(g15018),.A(g12739),.B(g12515));
  NAND2 NAND2_296(.VSS(VSS),.VDD(VDD),.Y(I13390),.A(g1821),.B(g1825));
  NAND2 NAND2_297(.VSS(VSS),.VDD(VDD),.Y(g14732),.A(g12662),.B(g12515));
  NAND2 NAND2_298(.VSS(VSS),.VDD(VDD),.Y(g24905),.A(g534),.B(g23088));
  NAND2 NAND2_299(.VSS(VSS),.VDD(VDD),.Y(I15242),.A(g10003),.B(I15241));
  NAND2 NAND2_300(.VSS(VSS),.VDD(VDD),.Y(g19857),.A(g13628),.B(g16296));
  NAND2 NAND2_301(.VSS(VSS),.VDD(VDD),.Y(g17500),.A(g14573),.B(g14548));
  NAND2 NAND2_302(.VSS(VSS),.VDD(VDD),.Y(I15123),.A(g2102),.B(I15121));
  NAND2 NAND2_303(.VSS(VSS),.VDD(VDD),.Y(g14761),.A(g12651),.B(g10281));
  NAND2 NAND2_304(.VSS(VSS),.VDD(VDD),.Y(I22844),.A(g12113),.B(g21228));
  NAND4 NAND4_56(.VSS(VSS),.VDD(VDD),.Y(g21555),.A(g17846),.B(g14946),.C(g17686),.D(g17650));
  NAND4 NAND4_57(.VSS(VSS),.VDD(VDD),.Y(g16854),.A(g3965),.B(g13824),.C(g3976),.D(g8595));
  NAND2 NAND2_305(.VSS(VSS),.VDD(VDD),.Y(g11974),.A(g2185),.B(g8259));
  NAND2 NAND2_306(.VSS(VSS),.VDD(VDD),.Y(g31671),.A(I29262),.B(I29263));
  NAND4 NAND4_58(.VSS(VSS),.VDD(VDD),.Y(g27933),.A(g21228),.B(g25356),.C(g26424),.D(g26236));
  NAND3 NAND3_49(.VSS(VSS),.VDD(VDD),.Y(g19549),.A(g15969),.B(g10841),.C(g10899));
  NAND4 NAND4_59(.VSS(VSS),.VDD(VDD),.Y(g8806),.A(g358),.B(g370),.C(g376),.D(g385));
  NAND2 NAND2_307(.VSS(VSS),.VDD(VDD),.Y(g11639),.A(g8933),.B(g4722));
  NAND2 NAND2_308(.VSS(VSS),.VDD(VDD),.Y(g9823),.A(I13383),.B(I13384));
  NAND2 NAND2_309(.VSS(VSS),.VDD(VDD),.Y(g12933),.A(g7150),.B(g10515));
  NAND2 NAND2_310(.VSS(VSS),.VDD(VDD),.Y(I25907),.A(g26256),.B(g24782));
  NAND4 NAND4_60(.VSS(VSS),.VDD(VDD),.Y(g10207),.A(g6315),.B(g6358),.C(g6329),.D(g6351));
  NAND2 NAND2_311(.VSS(VSS),.VDD(VDD),.Y(I20204),.A(g16246),.B(I20203));
  NAND2 NAND2_312(.VSS(VSS),.VDD(VDD),.Y(g26752),.A(g9397),.B(g25189));
  NAND2 NAND2_313(.VSS(VSS),.VDD(VDD),.Y(g14005),.A(g11514),.B(g11729));
  NAND4 NAND4_61(.VSS(VSS),.VDD(VDD),.Y(g16660),.A(g3953),.B(g11225),.C(g3969),.D(g13933));
  NAND2 NAND2_314(.VSS(VSS),.VDD(VDD),.Y(I26439),.A(g26549),.B(I26438));
  NAND4 NAND4_62(.VSS(VSS),.VDD(VDD),.Y(g17605),.A(g5559),.B(g14425),.C(g5630),.D(g12563));
  NAND2 NAND2_315(.VSS(VSS),.VDD(VDD),.Y(g11992),.A(g7275),.B(g1772));
  NAND2 NAND2_316(.VSS(VSS),.VDD(VDD),.Y(I29314),.A(g29501),.B(I29313));
  NAND2 NAND2_317(.VSS(VSS),.VDD(VDD),.Y(I26438),.A(g26549),.B(g14271));
  NAND2 NAND2_318(.VSS(VSS),.VDD(VDD),.Y(I12096),.A(g1339),.B(g1322));
  NAND2 NAND2_319(.VSS(VSS),.VDD(VDD),.Y(I23962),.A(g23184),.B(I23961));
  NAND2 NAND2_320(.VSS(VSS),.VDD(VDD),.Y(I17446),.A(g13336),.B(g956));
  NAND3 NAND3_50(.VSS(VSS),.VDD(VDD),.Y(g28206),.A(g12546),.B(g26105),.C(g27985));
  NAND2 NAND2_321(.VSS(VSS),.VDD(VDD),.Y(g25309),.A(g22384),.B(g12021));
  NAND2 NAND2_322(.VSS(VSS),.VDD(VDD),.Y(I13564),.A(g2648),.B(g2652));
  NAND2 NAND2_323(.VSS(VSS),.VDD(VDD),.Y(I12730),.A(g4287),.B(I12728));
  NAND2 NAND2_324(.VSS(VSS),.VDD(VDD),.Y(g7857),.A(I12241),.B(I12242));
  NAND3 NAND3_51(.VSS(VSS),.VDD(VDD),.Y(g28758),.A(g27779),.B(g7356),.C(g7275));
  NAND2 NAND2_325(.VSS(VSS),.VDD(VDD),.Y(I29269),.A(g29486),.B(g12050));
  NAND4 NAND4_63(.VSS(VSS),.VDD(VDD),.Y(g14771),.A(g5961),.B(g12129),.C(g5969),.D(g12351));
  NAND2 NAND2_326(.VSS(VSS),.VDD(VDD),.Y(g8913),.A(I12877),.B(I12878));
  NAND3 NAND3_52(.VSS(VSS),.VDD(VDD),.Y(g11442),.A(g8644),.B(g3288),.C(g3343));
  NAND2 NAND2_327(.VSS(VSS),.VDD(VDD),.Y(I13183),.A(g6500),.B(I13182));
  NAND2 NAND2_328(.VSS(VSS),.VDD(VDD),.Y(g14683),.A(g12553),.B(g12443));
  NAND4 NAND4_64(.VSS(VSS),.VDD(VDD),.Y(g17514),.A(g3917),.B(g13772),.C(g4019),.D(g8595));
  NAND2 NAND2_329(.VSS(VSS),.VDD(VDD),.Y(g25495),.A(g12483),.B(g22472));
  NAND2 NAND2_330(.VSS(VSS),.VDD(VDD),.Y(g12592),.A(I15364),.B(I15365));
  NAND2 NAND2_331(.VSS(VSS),.VDD(VDD),.Y(I13509),.A(g2089),.B(g2093));
  NAND2 NAND2_332(.VSS(VSS),.VDD(VDD),.Y(I14247),.A(g1322),.B(g8091));
  NAND2 NAND2_333(.VSS(VSS),.VDD(VDD),.Y(I15041),.A(g9752),.B(g1834));
  NAND2 NAND2_334(.VSS(VSS),.VDD(VDD),.Y(g10515),.A(g10337),.B(g5022));
  NAND2 NAND2_335(.VSS(VSS),.VDD(VDD),.Y(I13851),.A(g862),.B(I13850));
  NAND2 NAND2_336(.VSS(VSS),.VDD(VDD),.Y(g25985),.A(g24631),.B(g23956));
  NAND2 NAND2_337(.VSS(VSS),.VDD(VDD),.Y(g14882),.A(g12558),.B(g12453));
  NAND2 NAND2_338(.VSS(VSS),.VDD(VDD),.Y(g34424),.A(I32440),.B(I32441));
  NAND2 NAND2_339(.VSS(VSS),.VDD(VDD),.Y(g14407),.A(g12008),.B(g9807));
  NAND3 NAND3_53(.VSS(VSS),.VDD(VDD),.Y(g19856),.A(g13626),.B(g16278),.C(g8105));
  NAND2 NAND2_340(.VSS(VSS),.VDD(VDD),.Y(I23951),.A(g13603),.B(I23949));
  NAND2 NAND2_341(.VSS(VSS),.VDD(VDD),.Y(I15340),.A(g10154),.B(g2541));
  NAND2 NAND2_342(.VSS(VSS),.VDD(VDD),.Y(g26255),.A(g8075),.B(g24779));
  NAND2 NAND2_343(.VSS(VSS),.VDD(VDD),.Y(g12152),.A(g2485),.B(g8324));
  NAND2 NAND2_344(.VSS(VSS),.VDD(VDD),.Y(g22325),.A(g1252),.B(g19140));
  NAND2 NAND2_345(.VSS(VSS),.VDD(VDD),.Y(g13983),.A(g11658),.B(g8906));
  NAND4 NAND4_65(.VSS(VSS),.VDD(VDD),.Y(g16694),.A(g3905),.B(g13772),.C(g3976),.D(g11631));
  NAND4 NAND4_66(.VSS(VSS),.VDD(VDD),.Y(g17788),.A(g5232),.B(g14490),.C(g5327),.D(g12497));
  NAND2 NAND2_346(.VSS(VSS),.VDD(VDD),.Y(g12413),.A(g7521),.B(g5654));
  NAND2 NAND2_347(.VSS(VSS),.VDD(VDD),.Y(g10584),.A(g7362),.B(g7405));
  NAND2 NAND2_348(.VSS(VSS),.VDD(VDD),.Y(g28406),.A(g27064),.B(g13675));
  NAND2 NAND2_349(.VSS(VSS),.VDD(VDD),.Y(I13452),.A(g1955),.B(g1959));
  NAND3 NAND3_54(.VSS(VSS),.VDD(VDD),.Y(g28962),.A(g27886),.B(g2040),.C(g7369));
  NAND2 NAND2_350(.VSS(VSS),.VDD(VDD),.Y(I29279),.A(g12081),.B(I29277));
  NAND3 NAND3_55(.VSS(VSS),.VDD(VDD),.Y(g28500),.A(g590),.B(g27629),.C(g12323));
  NAND2 NAND2_351(.VSS(VSS),.VDD(VDD),.Y(g10759),.A(g7537),.B(g324));
  NAND3 NAND3_56(.VSS(VSS),.VDD(VDD),.Y(g15721),.A(g7564),.B(g311),.C(g13385));
  NAND2 NAND2_352(.VSS(VSS),.VDD(VDD),.Y(I29278),.A(g29488),.B(I29277));
  NAND2 NAND2_353(.VSS(VSS),.VDD(VDD),.Y(I14766),.A(g5821),.B(I14764));
  NAND2 NAND2_354(.VSS(VSS),.VDD(VDD),.Y(I15130),.A(g2527),.B(I15128));
  NAND2 NAND2_355(.VSS(VSS),.VDD(VDD),.Y(I15193),.A(g9935),.B(g6005));
  NAND2 NAND2_356(.VSS(VSS),.VDD(VDD),.Y(I29286),.A(g12085),.B(I29284));
  NAND2 NAND2_357(.VSS(VSS),.VDD(VDD),.Y(g14758),.A(g7704),.B(g12405));
  NAND2 NAND2_358(.VSS(VSS),.VDD(VDD),.Y(g11130),.A(g1221),.B(g7918));
  NAND2 NAND2_359(.VSS(VSS),.VDD(VDD),.Y(g14082),.A(g11697),.B(g11537));
  NAND2 NAND2_360(.VSS(VSS),.VDD(VDD),.Y(g11193),.A(I14258),.B(I14259));
  NAND3 NAND3_57(.VSS(VSS),.VDD(VDD),.Y(g13130),.A(g1351),.B(g11815),.C(g11336));
  NAND2 NAND2_361(.VSS(VSS),.VDD(VDD),.Y(g14107),.A(g11571),.B(g11527));
  NAND3 NAND3_58(.VSS(VSS),.VDD(VDD),.Y(g16278),.A(g8102),.B(g8057),.C(g13664));
  NAND2 NAND2_362(.VSS(VSS),.VDD(VDD),.Y(g12020),.A(g2028),.B(g8365));
  NAND3 NAND3_59(.VSS(VSS),.VDD(VDD),.Y(g19611),.A(g1070),.B(g1199),.C(g15995));
  NAND2 NAND2_363(.VSS(VSS),.VDD(VDD),.Y(g23139),.A(g21163),.B(g10756));
  NAND3 NAND3_60(.VSS(VSS),.VDD(VDD),.Y(g16306),.A(g4944),.B(g13971),.C(g12088));
  NAND2 NAND2_364(.VSS(VSS),.VDD(VDD),.Y(I12261),.A(g1454),.B(g1448));
  NAND2 NAND2_365(.VSS(VSS),.VDD(VDD),.Y(g14940),.A(g12744),.B(g12581));
  NAND2 NAND2_366(.VSS(VSS),.VDD(VDD),.Y(I18627),.A(g14712),.B(I18625));
  NAND3 NAND3_61(.VSS(VSS),.VDD(VDD),.Y(g13475),.A(g1008),.B(g11294),.C(g11786));
  NAND2 NAND2_367(.VSS(VSS),.VDD(VDD),.Y(g14848),.A(g12651),.B(g12453));
  NAND4 NAND4_67(.VSS(VSS),.VDD(VDD),.Y(g27282),.A(g11192),.B(g26269),.C(g26248),.D(g479));
  NAND4 NAND4_68(.VSS(VSS),.VDD(VDD),.Y(g21415),.A(g17773),.B(g14771),.C(g17740),.D(g14739));
  NAND4 NAND4_69(.VSS(VSS),.VDD(VDD),.Y(g16815),.A(g3909),.B(g13824),.C(g4005),.D(g11631));
  NAND4 NAND4_70(.VSS(VSS),.VDD(VDD),.Y(g13727),.A(g174),.B(g203),.C(g168),.D(g12812));
  NAND4 NAND4_71(.VSS(VSS),.VDD(VDD),.Y(g15734),.A(g5228),.B(g12059),.C(g5290),.D(g14631));
  NAND2 NAND2_368(.VSS(VSS),.VDD(VDD),.Y(g14804),.A(g12651),.B(g12798));
  NAND2 NAND2_369(.VSS(VSS),.VDD(VDD),.Y(g25255),.A(g20979),.B(g23659));
  NAND2 NAND2_370(.VSS(VSS),.VDD(VDD),.Y(I13731),.A(g4537),.B(I13729));
  NAND2 NAND2_371(.VSS(VSS),.VDD(VDD),.Y(g12357),.A(g7439),.B(g6329));
  NAND2 NAND2_372(.VSS(VSS),.VDD(VDD),.Y(g31978),.A(g30580),.B(g15591));
  NAND2 NAND2_373(.VSS(VSS),.VDD(VDD),.Y(I22824),.A(g21434),.B(I22822));
  NAND2 NAND2_374(.VSS(VSS),.VDD(VDD),.Y(I15253),.A(g10078),.B(g1848));
  NAND2 NAND2_375(.VSS(VSS),.VDD(VDD),.Y(g24621),.A(g22957),.B(g2927));
  NAND2 NAND2_376(.VSS(VSS),.VDD(VDD),.Y(I18681),.A(g2638),.B(I18680));
  NAND2 NAND2_377(.VSS(VSS),.VDD(VDD),.Y(g14962),.A(g12558),.B(g10281));
  NAND2 NAND2_378(.VSS(VSS),.VDD(VDD),.Y(g13600),.A(g3021),.B(g11039));
  NAND2 NAND2_379(.VSS(VSS),.VDD(VDD),.Y(I22931),.A(g21228),.B(I22929));
  NAND2 NAND2_380(.VSS(VSS),.VDD(VDD),.Y(g9645),.A(g2060),.B(g2028));
  NAND2 NAND2_381(.VSS(VSS),.VDD(VDD),.Y(g23576),.A(I22718),.B(I22719));
  NAND2 NAND2_382(.VSS(VSS),.VDD(VDD),.Y(g19764),.A(I20166),.B(I20167));
  NAND2 NAND2_383(.VSS(VSS),.VDD(VDD),.Y(g11952),.A(g1624),.B(g8187));
  NAND2 NAND2_384(.VSS(VSS),.VDD(VDD),.Y(I15175),.A(g9977),.B(I15174));
  NAND2 NAND2_385(.VSS(VSS),.VDD(VDD),.Y(I32757),.A(g34469),.B(I32756));
  NAND2 NAND2_386(.VSS(VSS),.VDD(VDD),.Y(I14370),.A(g3303),.B(I14368));
  NAND2 NAND2_387(.VSS(VSS),.VDD(VDD),.Y(g26782),.A(g9467),.B(g25203));
  NAND2 NAND2_388(.VSS(VSS),.VDD(VDD),.Y(g13821),.A(g11251),.B(g8340));
  NAND2 NAND2_389(.VSS(VSS),.VDD(VDD),.Y(g14048),.A(g11658),.B(g11483));
  NAND2 NAND2_390(.VSS(VSS),.VDD(VDD),.Y(I15264),.A(g2273),.B(I15262));
  NAND2 NAND2_391(.VSS(VSS),.VDD(VDD),.Y(g22755),.A(g20136),.B(g18984));
  NAND2 NAND2_392(.VSS(VSS),.VDD(VDD),.Y(g28421),.A(g27074),.B(g13715));
  NAND3 NAND3_62(.VSS(VSS),.VDD(VDD),.Y(g26352),.A(g744),.B(g24875),.C(g11679));
  NAND2 NAND2_393(.VSS(VSS),.VDD(VDD),.Y(I12271),.A(g956),.B(I12269));
  NAND3 NAND3_63(.VSS(VSS),.VDD(VDD),.Y(g13264),.A(g11869),.B(g11336),.C(g11849));
  NAND2 NAND2_394(.VSS(VSS),.VDD(VDD),.Y(g24933),.A(g19466),.B(g23154));
  NAND4 NAND4_72(.VSS(VSS),.VDD(VDD),.Y(g13137),.A(g10699),.B(g7675),.C(g1322),.D(g1404));
  NAND4 NAND4_73(.VSS(VSS),.VDD(VDD),.Y(g13516),.A(g11533),.B(g11490),.C(g11444),.D(g11412));
  NAND2 NAND2_395(.VSS(VSS),.VDD(VDD),.Y(g15039),.A(g12755),.B(g7142));
  NAND2 NAND2_396(.VSS(VSS),.VDD(VDD),.Y(g29060),.A(g9649),.B(g27800));
  NAND4 NAND4_74(.VSS(VSS),.VDD(VDD),.Y(g17755),.A(g5619),.B(g14522),.C(g5630),.D(g9864));
  NAND2 NAND2_397(.VSS(VSS),.VDD(VDD),.Y(g13873),.A(g11566),.B(g11729));
  NAND2 NAND2_398(.VSS(VSS),.VDD(VDD),.Y(I31974),.A(g33631),.B(I31972));
  NAND2 NAND2_399(.VSS(VSS),.VDD(VDD),.Y(g14947),.A(g12785),.B(g10491));
  NAND2 NAND2_400(.VSS(VSS),.VDD(VDD),.Y(g10605),.A(g2555),.B(g7490));
  NAND2 NAND2_401(.VSS(VSS),.VDD(VDD),.Y(g12482),.A(I15307),.B(I15308));
  NAND3 NAND3_64(.VSS(VSS),.VDD(VDD),.Y(g25470),.A(g22457),.B(g2051),.C(g8365));
  NAND2 NAND2_402(.VSS(VSS),.VDD(VDD),.Y(g13834),.A(g4754),.B(g11773));
  NAND3 NAND3_65(.VSS(VSS),.VDD(VDD),.Y(g16321),.A(g4955),.B(g13996),.C(g12088));
  NAND2 NAND2_403(.VSS(VSS),.VDD(VDD),.Y(g10951),.A(g7845),.B(g7868));
  NAND3 NAND3_66(.VSS(VSS),.VDD(VDD),.Y(g28920),.A(g27779),.B(g1802),.C(g7315));
  NAND2 NAND2_404(.VSS(VSS),.VDD(VDD),.Y(g24574),.A(g22709),.B(g22687));
  NAND2 NAND2_405(.VSS(VSS),.VDD(VDD),.Y(g14234),.A(g9177),.B(g11881));
  NAND2 NAND2_406(.VSS(VSS),.VDD(VDD),.Y(g31706),.A(I29270),.B(I29271));
  NAND2 NAND2_407(.VSS(VSS),.VDD(VDD),.Y(I18626),.A(g2079),.B(I18625));
  NAND3 NAND3_67(.VSS(VSS),.VDD(VDD),.Y(g28946),.A(g27907),.B(g2495),.C(g2421));
  NAND2 NAND2_408(.VSS(VSS),.VDD(VDD),.Y(g25467),.A(g12432),.B(g22417));
  NAND2 NAND2_409(.VSS(VSS),.VDD(VDD),.Y(g23761),.A(I22893),.B(I22894));
  NAND2 NAND2_410(.VSS(VSS),.VDD(VDD),.Y(g23692),.A(g9501),.B(g20995));
  NAND2 NAND2_411(.VSS(VSS),.VDD(VDD),.Y(g27380),.A(I26071),.B(I26072));
  NAND2 NAND2_412(.VSS(VSS),.VDD(VDD),.Y(g12356),.A(g7438),.B(g6012));
  NAND2 NAND2_413(.VSS(VSS),.VDD(VDD),.Y(g9591),.A(g1926),.B(g1894));
  NAND3 NAND3_68(.VSS(VSS),.VDD(VDD),.Y(g12999),.A(g4392),.B(g10476),.C(g4401));
  NAND3 NAND3_69(.VSS(VSS),.VDD(VDD),.Y(g11320),.A(g4633),.B(g4621),.C(g7202));
  NAND2 NAND2_414(.VSS(VSS),.VDD(VDD),.Y(g25984),.A(g24567),.B(g22668));
  NAND2 NAND2_415(.VSS(VSS),.VDD(VDD),.Y(g19886),.A(g11403),.B(g17794));
  NAND2 NAND2_416(.VSS(VSS),.VDD(VDD),.Y(I15122),.A(g9910),.B(I15121));
  NAND2 NAND2_417(.VSS(VSS),.VDD(VDD),.Y(g13346),.A(g4854),.B(g11012));
  NAND2 NAND2_418(.VSS(VSS),.VDD(VDD),.Y(g19792),.A(I20204),.B(I20205));
  NAND2 NAND2_419(.VSS(VSS),.VDD(VDD),.Y(I14957),.A(g6181),.B(I14955));
  NAND3 NAND3_70(.VSS(VSS),.VDD(VDD),.Y(g26053),.A(g22875),.B(g24677),.C(g22941));
  NAND3 NAND3_71(.VSS(VSS),.VDD(VDD),.Y(g13464),.A(g10831),.B(g4793),.C(g4776));
  NAND2 NAND2_420(.VSS(VSS),.VDD(VDD),.Y(g13797),.A(g8102),.B(g11273));
  NAND2 NAND2_421(.VSS(VSS),.VDD(VDD),.Y(g11292),.A(I14331),.B(I14332));
  NAND2 NAND2_422(.VSS(VSS),.VDD(VDD),.Y(I32756),.A(g34469),.B(g25779));
  NAND2 NAND2_423(.VSS(VSS),.VDD(VDD),.Y(g11153),.A(I14205),.B(I14206));
  NAND2 NAND2_424(.VSS(VSS),.VDD(VDD),.Y(g29094),.A(g27858),.B(g9700));
  NAND3 NAND3_72(.VSS(VSS),.VDD(VDD),.Y(g12449),.A(g7004),.B(g5297),.C(g5352));
  NAND2 NAND2_425(.VSS(VSS),.VDD(VDD),.Y(I14290),.A(g8282),.B(I14289));
  NAND2 NAND2_426(.VSS(VSS),.VDD(VDD),.Y(g11409),.A(g9842),.B(g3298));
  NAND2 NAND2_427(.VSS(VSS),.VDD(VDD),.Y(I22894),.A(g21228),.B(I22892));
  NAND2 NAND2_428(.VSS(VSS),.VDD(VDD),.Y(I14427),.A(g8595),.B(g4005));
  NAND4 NAND4_75(.VSS(VSS),.VDD(VDD),.Y(g14829),.A(g6621),.B(g12137),.C(g6675),.D(g12471));
  NAND2 NAND2_429(.VSS(VSS),.VDD(VDD),.Y(I31983),.A(g33653),.B(g33648));
  NAND2 NAND2_430(.VSS(VSS),.VDD(VDD),.Y(g14434),.A(g6415),.B(g11945));
  NAND2 NAND2_431(.VSS(VSS),.VDD(VDD),.Y(g29018),.A(g9586),.B(g27742));
  NAND2 NAND2_432(.VSS(VSS),.VDD(VDD),.Y(I12878),.A(g4180),.B(I12876));
  NAND2 NAND2_433(.VSS(VSS),.VDD(VDD),.Y(g10946),.A(g1489),.B(g7876));
  NAND3 NAND3_73(.VSS(VSS),.VDD(VDD),.Y(g28927),.A(g27837),.B(g1906),.C(g7322));
  NAND4 NAND4_76(.VSS(VSS),.VDD(VDD),.Y(g14946),.A(g6247),.B(g12173),.C(g6346),.D(g12672));
  NAND2 NAND2_434(.VSS(VSS),.VDD(VDD),.Y(g9750),.A(I13335),.B(I13336));
  NAND2 NAND2_435(.VSS(VSS),.VDD(VDD),.Y(I11826),.A(g4601),.B(I11824));
  NAND2 NAND2_436(.VSS(VSS),.VDD(VDD),.Y(g14344),.A(g5377),.B(g11885));
  NAND2 NAND2_437(.VSS(VSS),.VDD(VDD),.Y(g24583),.A(g22753),.B(g22711));
  NAND2 NAND2_438(.VSS(VSS),.VDD(VDD),.Y(I13182),.A(g6500),.B(g6505));
  NAND2 NAND2_439(.VSS(VSS),.VDD(VDD),.Y(I17496),.A(g1448),.B(I17494));
  NAND3 NAND3_74(.VSS(VSS),.VDD(VDD),.Y(g28903),.A(g27800),.B(g2197),.C(g7280));
  NAND2 NAND2_440(.VSS(VSS),.VDD(VDD),.Y(g14682),.A(g4933),.B(g11780));
  NAND2 NAND2_441(.VSS(VSS),.VDD(VDD),.Y(g12149),.A(g8205),.B(g2185));
  NAND2 NAND2_442(.VSS(VSS),.VDD(VDD),.Y(I14481),.A(g10074),.B(I14480));
  NAND3 NAND3_75(.VSS(VSS),.VDD(VDD),.Y(g28755),.A(g27742),.B(g7268),.C(g1592));
  NAND2 NAND2_443(.VSS(VSS),.VDD(VDD),.Y(g12148),.A(g2060),.B(g8310));
  NAND4 NAND4_77(.VSS(VSS),.VDD(VDD),.Y(g13109),.A(g6279),.B(g12173),.C(g6369),.D(g10003));
  NAND4 NAND4_78(.VSS(VSS),.VDD(VDD),.Y(g16772),.A(g3558),.B(g13799),.C(g3654),.D(g11576));
  NAND2 NAND2_444(.VSS(VSS),.VDD(VDD),.Y(g24787),.A(g3391),.B(g23079));
  NAND3 NAND3_76(.VSS(VSS),.VDD(VDD),.Y(g29001),.A(g27937),.B(g2599),.C(g7431));
  NAND4 NAND4_79(.VSS(VSS),.VDD(VDD),.Y(g13108),.A(g5551),.B(g12029),.C(g5685),.D(g9864));
  NAND2 NAND2_445(.VSS(VSS),.VDD(VDD),.Y(g12343),.A(g7470),.B(g5630));
  NAND3 NAND3_77(.VSS(VSS),.VDD(VDD),.Y(g13283),.A(g12440),.B(g12399),.C(g9843));
  NAND2 NAND2_446(.VSS(VSS),.VDD(VDD),.Y(I22801),.A(g21434),.B(I22799));
  NAND3 NAND3_78(.VSS(VSS),.VDD(VDD),.Y(g11492),.A(g6928),.B(g6941),.C(g8756));
  NAND3 NAND3_79(.VSS(VSS),.VDD(VDD),.Y(g12971),.A(g9024),.B(g8977),.C(g10664));
  NAND2 NAND2_447(.VSS(VSS),.VDD(VDD),.Y(I12545),.A(g191),.B(I12544));
  NAND2 NAND2_448(.VSS(VSS),.VDD(VDD),.Y(g9528),.A(I13183),.B(I13184));
  NAND2 NAND2_449(.VSS(VSS),.VDD(VDD),.Y(g12369),.A(g9049),.B(g637));
  NAND2 NAND2_450(.VSS(VSS),.VDD(VDD),.Y(g28395),.A(g27074),.B(g13655));
  NAND2 NAND2_451(.VSS(VSS),.VDD(VDD),.Y(I14956),.A(g9620),.B(I14955));
  NAND2 NAND2_452(.VSS(VSS),.VDD(VDD),.Y(g11381),.A(g9660),.B(g3274));
  NAND2 NAND2_453(.VSS(VSS),.VDD(VDD),.Y(g28899),.A(g27833),.B(g14612));
  NAND2 NAND2_454(.VSS(VSS),.VDD(VDD),.Y(I18529),.A(g1811),.B(g14640));
  NAND2 NAND2_455(.VSS(VSS),.VDD(VDD),.Y(g28990),.A(g27882),.B(g8310));
  NAND3 NAND3_80(.VSS(VSS),.VDD(VDD),.Y(g17220),.A(g9369),.B(g9298),.C(g14376));
  NAND2 NAND2_456(.VSS(VSS),.VDD(VDD),.Y(I15174),.A(g9977),.B(g2661));
  NAND2 NAND2_457(.VSS(VSS),.VDD(VDD),.Y(g29157),.A(g9835),.B(g27937));
  NAND3 NAND3_81(.VSS(VSS),.VDD(VDD),.Y(g17246),.A(g9439),.B(g9379),.C(g14405));
  NAND3 NAND3_82(.VSS(VSS),.VDD(VDD),.Y(g12412),.A(g10044),.B(g5297),.C(g5348));
  NAND2 NAND2_458(.VSS(VSS),.VDD(VDD),.Y(I26049),.A(g25997),.B(g13500));
  NAND3 NAND3_83(.VSS(VSS),.VDD(VDD),.Y(g26382),.A(g577),.B(g24953),.C(g12323));
  NAND3 NAND3_84(.VSS(VSS),.VDD(VDD),.Y(g33930),.A(g33394),.B(g12767),.C(g9848));
  NAND2 NAND2_459(.VSS(VSS),.VDD(VDD),.Y(g22754),.A(g20114),.B(g19376));
  NAND2 NAND2_460(.VSS(VSS),.VDD(VDD),.Y(g33838),.A(g33083),.B(g4369));
  NAND2 NAND2_461(.VSS(VSS),.VDD(VDD),.Y(g14927),.A(g12695),.B(g10281));
  NAND2 NAND2_462(.VSS(VSS),.VDD(VDD),.Y(g16586),.A(g13851),.B(g13823));
  NAND2 NAND2_463(.VSS(VSS),.VDD(VDD),.Y(I22866),.A(g21228),.B(I22864));
  NAND2 NAND2_464(.VSS(VSS),.VDD(VDD),.Y(g21345),.A(g11429),.B(g17157));
  NAND3 NAND3_85(.VSS(VSS),.VDD(VDD),.Y(g27582),.A(g10857),.B(g26131),.C(g26105));
  NAND2 NAND2_465(.VSS(VSS),.VDD(VDD),.Y(g9372),.A(g5080),.B(g5084));
  NAND3 NAND3_86(.VSS(VSS),.VDD(VDD),.Y(g28861),.A(g27837),.B(g7405),.C(g1906));
  NAND2 NAND2_466(.VSS(VSS),.VDD(VDD),.Y(I20461),.A(g17515),.B(I20460));
  NAND3 NAND3_87(.VSS(VSS),.VDD(VDD),.Y(g25476),.A(g22472),.B(g2476),.C(g8373));
  NAND2 NAND2_467(.VSS(VSS),.VDD(VDD),.Y(g8359),.A(I12545),.B(I12546));
  NAND2 NAND2_468(.VSS(VSS),.VDD(VDD),.Y(g24662),.A(g22957),.B(g2955));
  NAND2 NAND2_469(.VSS(VSS),.VDD(VDD),.Y(I24461),.A(g23796),.B(g14437));
  NAND2 NAND2_470(.VSS(VSS),.VDD(VDD),.Y(g10604),.A(g7424),.B(g7456));
  NAND4 NAND4_80(.VSS(VSS),.VDD(VDD),.Y(g15751),.A(g5591),.B(g14522),.C(g5666),.D(g14669));
  NAND4 NAND4_81(.VSS(VSS),.VDD(VDD),.Y(g10755),.A(g7352),.B(g7675),.C(g1322),.D(g1404));
  NAND2 NAND2_471(.VSS(VSS),.VDD(VDD),.Y(g24890),.A(g13852),.B(g22929));
  NAND2 NAND2_472(.VSS(VSS),.VDD(VDD),.Y(g14755),.A(g12593),.B(g12772));
  NAND3 NAND3_88(.VSS(VSS),.VDD(VDD),.Y(g19495),.A(g15969),.B(g10841),.C(g7781));
  NAND2 NAND2_473(.VSS(VSS),.VDD(VDD),.Y(g27925),.A(I26439),.B(I26440));
  NAND2 NAND2_474(.VSS(VSS),.VDD(VDD),.Y(I22923),.A(g21284),.B(I22921));
  NAND2 NAND2_475(.VSS(VSS),.VDD(VDD),.Y(g29660),.A(g28448),.B(g9582));
  NAND3 NAND3_89(.VSS(VSS),.VDD(VDD),.Y(g20248),.A(g17056),.B(g14146),.C(g14123));
  NAND2 NAND2_476(.VSS(VSS),.VDD(VDD),.Y(g16275),.A(g9291),.B(g13480));
  NAND2 NAND2_477(.VSS(VSS),.VDD(VDD),.Y(g14981),.A(g12785),.B(g12632));
  NAND2 NAND2_478(.VSS(VSS),.VDD(VDD),.Y(I14211),.A(g9252),.B(g9295));
  NAND2 NAND2_479(.VSS(VSS),.VDD(VDD),.Y(g9334),.A(g827),.B(g832));
  NAND2 NAND2_480(.VSS(VSS),.VDD(VDD),.Y(g12112),.A(g8139),.B(g1624));
  NAND2 NAND2_481(.VSS(VSS),.VDD(VDD),.Y(I17923),.A(g13378),.B(g1478));
  NAND3 NAND3_90(.VSS(VSS),.VDD(VDD),.Y(g33306),.A(g776),.B(g32212),.C(g11679));
  NAND4 NAND4_82(.VSS(VSS),.VDD(VDD),.Y(g11326),.A(g8993),.B(g376),.C(g365),.D(g370));
  NAND2 NAND2_482(.VSS(VSS),.VDD(VDD),.Y(g20081),.A(g11325),.B(g17794));
  NAND2 NAND2_483(.VSS(VSS),.VDD(VDD),.Y(g14794),.A(g12492),.B(g12772));
  NAND2 NAND2_484(.VSS(VSS),.VDD(VDD),.Y(g14845),.A(g12558),.B(g12798));
  NAND2 NAND2_485(.VSS(VSS),.VDD(VDD),.Y(I14497),.A(g9020),.B(g8737));
  NAND2 NAND2_486(.VSS(VSS),.VDD(VDD),.Y(I24365),.A(g14320),.B(I24363));
  NAND2 NAND2_487(.VSS(VSS),.VDD(VDD),.Y(I13850),.A(g862),.B(g7397));
  NAND4 NAND4_83(.VSS(VSS),.VDD(VDD),.Y(g13040),.A(g5196),.B(g12002),.C(g5308),.D(g9780));
  NAND2 NAND2_488(.VSS(VSS),.VDD(VDD),.Y(g13948),.A(g11610),.B(g8864));
  NAND2 NAND2_489(.VSS(VSS),.VDD(VDD),.Y(g14899),.A(g12744),.B(g10421));
  NAND2 NAND2_490(.VSS(VSS),.VDD(VDD),.Y(g29085),.A(g9694),.B(g27837));
  NAND2 NAND2_491(.VSS(VSS),.VDD(VDD),.Y(g28997),.A(g27903),.B(g8324));
  NAND2 NAND2_492(.VSS(VSS),.VDD(VDD),.Y(g25382),.A(g12333),.B(g22342));
  NAND2 NAND2_493(.VSS(VSS),.VDD(VDD),.Y(I12289),.A(g1300),.B(I12287));
  NAND4 NAND4_84(.VSS(VSS),.VDD(VDD),.Y(g14898),.A(g5901),.B(g12129),.C(g6000),.D(g12614));
  NAND2 NAND2_494(.VSS(VSS),.VDD(VDD),.Y(I32204),.A(g33670),.B(I32202));
  NAND2 NAND2_495(.VSS(VSS),.VDD(VDD),.Y(I23950),.A(g23162),.B(I23949));
  NAND2 NAND2_496(.VSS(VSS),.VDD(VDD),.Y(g15014),.A(g12785),.B(g12680));
  NAND2 NAND2_497(.VSS(VSS),.VDD(VDD),.Y(I12288),.A(g1484),.B(I12287));
  NAND2 NAND2_498(.VSS(VSS),.VDD(VDD),.Y(g24380),.A(I23601),.B(I23602));
  NAND2 NAND2_499(.VSS(VSS),.VDD(VDD),.Y(g12429),.A(g7473),.B(g6675));
  NAND2 NAND2_500(.VSS(VSS),.VDD(VDD),.Y(g14521),.A(g12170),.B(g5428));
  NAND2 NAND2_501(.VSS(VSS),.VDD(VDD),.Y(I25221),.A(g24718),.B(I25219));
  NAND2 NAND2_502(.VSS(VSS),.VDD(VDD),.Y(g12428),.A(g7472),.B(g6358));
  NAND3 NAND3_91(.VSS(VSS),.VDD(VDD),.Y(g28871),.A(g27858),.B(g7418),.C(g2331));
  NAND2 NAND2_503(.VSS(VSS),.VDD(VDD),.Y(I17885),.A(g1135),.B(I17883));
  NAND2 NAND2_504(.VSS(VSS),.VDD(VDD),.Y(g9908),.A(I13453),.B(I13454));
  NAND2 NAND2_505(.VSS(VSS),.VDD(VDD),.Y(g22902),.A(g18957),.B(g2848));
  NAND2 NAND2_506(.VSS(VSS),.VDD(VDD),.Y(I16780),.A(g12332),.B(I16778));
  NAND2 NAND2_507(.VSS(VSS),.VDD(VDD),.Y(g10573),.A(g7992),.B(g8179));
  NAND2 NAND2_508(.VSS(VSS),.VDD(VDD),.Y(g9567),.A(g6116),.B(g6120));
  NAND2 NAND2_509(.VSS(VSS),.VDD(VDD),.Y(g14861),.A(g12744),.B(g10341));
  NAND2 NAND2_510(.VSS(VSS),.VDD(VDD),.Y(g14573),.A(g9506),.B(g12249));
  NAND2 NAND2_511(.VSS(VSS),.VDD(VDD),.Y(g24932),.A(g19886),.B(g23172));
  NAND4 NAND4_85(.VSS(VSS),.VDD(VDD),.Y(g15720),.A(g5917),.B(g14497),.C(g6019),.D(g9935));
  NAND3 NAND3_92(.VSS(VSS),.VDD(VDD),.Y(g11933),.A(g837),.B(g9334),.C(g7197));
  NAND2 NAND2_512(.VSS(VSS),.VDD(VDD),.Y(I14855),.A(g5142),.B(I14853));
  NAND2 NAND2_513(.VSS(VSS),.VDD(VDD),.Y(g14045),.A(g11571),.B(g11747));
  NAND2 NAND2_514(.VSS(VSS),.VDD(VDD),.Y(g29335),.A(g25540),.B(g28131));
  NAND2 NAND2_515(.VSS(VSS),.VDD(VDD),.Y(g13634),.A(g11797),.B(g11261));
  NAND2 NAND2_516(.VSS(VSS),.VDD(VDD),.Y(g13851),.A(g8224),.B(g11360));
  NAND2 NAND2_517(.VSS(VSS),.VDD(VDD),.Y(g27317),.A(g24793),.B(g26255));
  NAND2 NAND2_518(.VSS(VSS),.VDD(VDD),.Y(I12374),.A(g3462),.B(I12372));
  NAND2 NAND2_519(.VSS(VSS),.VDD(VDD),.Y(g25215),.A(I24384),.B(I24385));
  NAND2 NAND2_520(.VSS(VSS),.VDD(VDD),.Y(g7850),.A(g554),.B(g807));
  NAND2 NAND2_521(.VSS(VSS),.VDD(VDD),.Y(g12317),.A(g10026),.B(g6486));
  NAND2 NAND2_522(.VSS(VSS),.VDD(VDD),.Y(g29694),.A(g28391),.B(g13709));
  NAND2 NAND2_523(.VSS(VSS),.VDD(VDD),.Y(g14098),.A(g11566),.B(g8864));
  NAND2 NAND2_524(.VSS(VSS),.VDD(VDD),.Y(g17699),.A(I18681),.B(I18682));
  NAND2 NAND2_525(.VSS(VSS),.VDD(VDD),.Y(g25439),.A(g22498),.B(g12122));
  NAND3 NAND3_93(.VSS(VSS),.VDD(VDD),.Y(g28911),.A(g27907),.B(g7456),.C(g2465));
  NAND2 NAND2_526(.VSS(VSS),.VDD(VDD),.Y(g23972),.A(g7097),.B(g20751));
  NAND3 NAND3_94(.VSS(VSS),.VDD(VDD),.Y(g17290),.A(g9506),.B(g9449),.C(g14431));
  NAND2 NAND2_527(.VSS(VSS),.VDD(VDD),.Y(I29253),.A(g29482),.B(g12017));
  NAND2 NAND2_528(.VSS(VSS),.VDD(VDD),.Y(g29131),.A(g27907),.B(g9762));
  NAND2 NAND2_529(.VSS(VSS),.VDD(VDD),.Y(I15213),.A(g10035),.B(I15212));
  NAND2 NAND2_530(.VSS(VSS),.VDD(VDD),.Y(I12842),.A(g4235),.B(I12840));
  NAND2 NAND2_531(.VSS(VSS),.VDD(VDD),.Y(g25349),.A(g22432),.B(g12051));
  NAND2 NAND2_532(.VSS(VSS),.VDD(VDD),.Y(g12245),.A(g7344),.B(g5637));
  NAND2 NAND2_533(.VSS(VSS),.VDD(VDD),.Y(g12323),.A(g9480),.B(g640));
  NAND2 NAND2_534(.VSS(VSS),.VDD(VDD),.Y(I14714),.A(g5128),.B(I14712));
  NAND2 NAND2_535(.VSS(VSS),.VDD(VDD),.Y(g22661),.A(g20136),.B(g94));
  NAND2 NAND2_536(.VSS(VSS),.VDD(VDD),.Y(I13730),.A(g4534),.B(I13729));
  NAND4 NAND4_86(.VSS(VSS),.VDD(VDD),.Y(g27775),.A(g21228),.B(g25262),.C(g26424),.D(g26166));
  NAND3 NAND3_95(.VSS(VSS),.VDD(VDD),.Y(g16236),.A(g13573),.B(g13554),.C(g13058));
  NAND2 NAND2_537(.VSS(VSS),.VDD(VDD),.Y(I14257),.A(g8154),.B(g3133));
  NAND3 NAND3_96(.VSS(VSS),.VDD(VDD),.Y(g28950),.A(g27937),.B(g7490),.C(g2599));
  NAND2 NAND2_538(.VSS(VSS),.VDD(VDD),.Y(I15051),.A(g9759),.B(g2259));
  NAND2 NAND2_539(.VSS(VSS),.VDD(VDD),.Y(I14818),.A(g6513),.B(I14816));
  NAND2 NAND2_540(.VSS(VSS),.VDD(VDD),.Y(g9724),.A(g5092),.B(g5084));
  NAND2 NAND2_541(.VSS(VSS),.VDD(VDD),.Y(g22715),.A(g20114),.B(g2999));
  NAND2 NAND2_542(.VSS(VSS),.VDD(VDD),.Y(I23120),.A(g417),.B(I23118));
  NAND2 NAND2_543(.VSS(VSS),.VDD(VDD),.Y(g24620),.A(g22902),.B(g22874));
  NAND4 NAND4_87(.VSS(VSS),.VDD(VDD),.Y(g14871),.A(g6653),.B(g12211),.C(g6661),.D(g12471));
  NAND2 NAND2_544(.VSS(VSS),.VDD(VDD),.Y(I12544),.A(g191),.B(g194));
  NAND2 NAND2_545(.VSS(VSS),.VDD(VDD),.Y(g13756),.A(g203),.B(g12812));
  NAND2 NAND2_546(.VSS(VSS),.VDD(VDD),.Y(I18680),.A(g2638),.B(g14752));
  NAND2 NAND2_547(.VSS(VSS),.VDD(VDD),.Y(g12232),.A(g8804),.B(g4878));
  NAND3 NAND3_97(.VSS(VSS),.VDD(VDD),.Y(g16264),.A(g518),.B(g9158),.C(g13223));
  NAND2 NAND2_548(.VSS(VSS),.VDD(VDD),.Y(g19875),.A(g13667),.B(g16316));
  NAND2 NAND2_549(.VSS(VSS),.VDD(VDD),.Y(I22930),.A(g12223),.B(I22929));
  NAND3 NAND3_98(.VSS(VSS),.VDD(VDD),.Y(g26052),.A(g22714),.B(g24662),.C(g22921));
  NAND2 NAND2_550(.VSS(VSS),.VDD(VDD),.Y(g26745),.A(g6856),.B(g25317));
  NAND4 NAND4_88(.VSS(VSS),.VDD(VDD),.Y(g17572),.A(g3598),.B(g13799),.C(g3676),.D(g8542));
  NAND2 NAND2_551(.VSS(VSS),.VDD(VDD),.Y(g11350),.A(I14369),.B(I14370));
  NAND2 NAND2_552(.VSS(VSS),.VDD(VDD),.Y(I22965),.A(g12288),.B(g21228));
  NAND2 NAND2_553(.VSS(VSS),.VDD(VDD),.Y(I32433),.A(g34051),.B(I32431));
  NAND2 NAND2_554(.VSS(VSS),.VDD(VDD),.Y(g24369),.A(I23586),.B(I23587));
  NAND2 NAND2_555(.VSS(VSS),.VDD(VDD),.Y(g12512),.A(g7766),.B(g10312));
  NAND2 NAND2_556(.VSS(VSS),.VDD(VDD),.Y(g21359),.A(g11509),.B(g17157));
  NAND2 NAND2_557(.VSS(VSS),.VDD(VDD),.Y(g13846),.A(g1116),.B(g10649));
  NAND2 NAND2_558(.VSS(VSS),.VDD(VDD),.Y(g10472),.A(I13851),.B(I13852));
  NAND2 NAND2_559(.VSS(VSS),.VDD(VDD),.Y(g11396),.A(g8713),.B(g4688));
  NAND2 NAND2_560(.VSS(VSS),.VDD(VDD),.Y(I12270),.A(g1141),.B(I12269));
  NAND2 NAND2_561(.VSS(VSS),.VDD(VDD),.Y(I14735),.A(g5475),.B(I14733));
  NAND3 NAND3_99(.VSS(VSS),.VDD(VDD),.Y(g19455),.A(g15969),.B(g10841),.C(g7781));
  NAND4 NAND4_89(.VSS(VSS),.VDD(VDD),.Y(g20133),.A(g17668),.B(g17634),.C(g17597),.D(g14569));
  NAND2 NAND2_562(.VSS(VSS),.VDD(VDD),.Y(g17297),.A(g2729),.B(g14291));
  NAND2 NAND2_563(.VSS(VSS),.VDD(VDD),.Y(g21344),.A(g11428),.B(g17157));
  NAND4 NAND4_90(.VSS(VSS),.VDD(VDD),.Y(g11405),.A(g2741),.B(g2735),.C(g6856),.D(g2748));
  NAND4 NAND4_91(.VSS(VSS),.VDD(VDD),.Y(g15781),.A(g6267),.B(g12173),.C(g6329),.D(g14745));
  NAND2 NAND2_564(.VSS(VSS),.VDD(VDD),.Y(g20011),.A(g3731),.B(g16476));
  NAND2 NAND2_565(.VSS(VSS),.VDD(VDD),.Y(g14776),.A(g12780),.B(g12622));
  NAND3 NAND3_100(.VSS(VSS),.VDD(VDD),.Y(g28203),.A(g12546),.B(g27985),.C(g27977));
  NAND3 NAND3_101(.VSS(VSS),.VDD(VDD),.Y(g10754),.A(g7936),.B(g7913),.C(g8411));
  NAND2 NAND2_566(.VSS(VSS),.VDD(VDD),.Y(g29015),.A(g27742),.B(g9586));
  NAND2 NAND2_567(.VSS(VSS),.VDD(VDD),.Y(g13929),.A(g11669),.B(g11763));
  NAND2 NAND2_568(.VSS(VSS),.VDD(VDD),.Y(I12219),.A(g1478),.B(I12217));
  NAND2 NAND2_569(.VSS(VSS),.VDD(VDD),.Y(g25200),.A(g5742),.B(g23642));
  NAND2 NAND2_570(.VSS(VSS),.VDD(VDD),.Y(g14825),.A(g12806),.B(g12680));
  NAND2 NAND2_571(.VSS(VSS),.VDD(VDD),.Y(g14950),.A(g7812),.B(g12632));
  NAND2 NAND2_572(.VSS(VSS),.VDD(VDD),.Y(g11020),.A(g9187),.B(g9040));
  NAND2 NAND2_573(.VSS(VSS),.VDD(VDD),.Y(g12080),.A(g1917),.B(g8201));
  NAND4 NAND4_92(.VSS(VSS),.VDD(VDD),.Y(g13928),.A(g3562),.B(g11238),.C(g3680),.D(g11576));
  NAND2 NAND2_574(.VSS(VSS),.VDD(VDD),.Y(I12218),.A(g1437),.B(I12217));
  NAND2 NAND2_575(.VSS(VSS),.VDD(VDD),.Y(g14858),.A(g7766),.B(g12515));
  NAND2 NAND2_576(.VSS(VSS),.VDD(VDD),.Y(g19782),.A(I20188),.B(I20189));
  NAND2 NAND2_577(.VSS(VSS),.VDD(VDD),.Y(g29556),.A(g28349),.B(g13486));
  NAND2 NAND2_578(.VSS(VSS),.VDD(VDD),.Y(g31747),.A(I29296),.B(I29297));
  NAND2 NAND2_579(.VSS(VSS),.VDD(VDD),.Y(g14151),.A(g11692),.B(g11483));
  NAND2 NAND2_580(.VSS(VSS),.VDD(VDD),.Y(g14996),.A(g12662),.B(g10312));
  NAND2 NAND2_581(.VSS(VSS),.VDD(VDD),.Y(g24925),.A(g20092),.B(g23154));
  NAND2 NAND2_582(.VSS(VSS),.VDD(VDD),.Y(g24958),.A(g21330),.B(g23462));
  NAND4 NAND4_93(.VSS(VSS),.VDD(VDD),.Y(g17520),.A(g5260),.B(g12002),.C(g5276),.D(g14631));
  NAND2 NAND2_583(.VSS(VSS),.VDD(VDD),.Y(g12461),.A(g7536),.B(g6000));
  NAND2 NAND2_584(.VSS(VSS),.VDD(VDD),.Y(I24364),.A(g23687),.B(I24363));
  NAND3 NAND3_102(.VSS(VSS),.VDD(VDD),.Y(g12342),.A(g7004),.B(g7018),.C(g10129));
  NAND2 NAND2_585(.VSS(VSS),.VDD(VDD),.Y(I22937),.A(g12226),.B(I22936));
  NAND2 NAND2_586(.VSS(VSS),.VDD(VDD),.Y(I26395),.A(g14227),.B(I26393));
  NAND2 NAND2_587(.VSS(VSS),.VDD(VDD),.Y(I14923),.A(g9558),.B(g5835));
  NAND2 NAND2_588(.VSS(VSS),.VDD(VDD),.Y(g12145),.A(g8195),.B(g1760));
  NAND2 NAND2_589(.VSS(VSS),.VDD(VDD),.Y(g11302),.A(g9496),.B(g3281));
  NAND2 NAND2_590(.VSS(VSS),.VDD(VDD),.Y(I15105),.A(g9780),.B(g5313));
  NAND2 NAND2_591(.VSS(VSS),.VDD(VDD),.Y(I23980),.A(g13670),.B(I23978));
  NAND2 NAND2_592(.VSS(VSS),.VDD(VDD),.Y(g24944),.A(g21354),.B(g23363));
  NAND4 NAND4_94(.VSS(VSS),.VDD(VDD),.Y(g13105),.A(g10671),.B(g7675),.C(g1322),.D(g1404));
  NAND2 NAND2_593(.VSS(VSS),.VDD(VDD),.Y(I16779),.A(g11292),.B(I16778));
  NAND2 NAND2_594(.VSS(VSS),.VDD(VDD),.Y(I12470),.A(g392),.B(I12468));
  NAND2 NAND2_595(.VSS(VSS),.VDD(VDD),.Y(g9092),.A(g3004),.B(g3050));
  NAND2 NAND2_596(.VSS(VSS),.VDD(VDD),.Y(I16778),.A(g11292),.B(g12332));
  NAND3 NAND3_103(.VSS(VSS),.VDD(VDD),.Y(g19589),.A(g15969),.B(g10841),.C(g10884));
  NAND2 NAND2_597(.VSS(VSS),.VDD(VDD),.Y(I12277),.A(g1467),.B(g1472));
  NAND2 NAND2_598(.VSS(VSS),.VDD(VDD),.Y(I13499),.A(g232),.B(I13497));
  NAND2 NAND2_599(.VSS(VSS),.VDD(VDD),.Y(I17884),.A(g13336),.B(I17883));
  NAND2 NAND2_600(.VSS(VSS),.VDD(VDD),.Y(g15021),.A(g12711),.B(g10341));
  NAND2 NAND2_601(.VSS(VSS),.VDD(VDD),.Y(I12075),.A(g996),.B(I12074));
  NAND2 NAND2_602(.VSS(VSS),.VDD(VDD),.Y(g27365),.A(I26050),.B(I26051));
  NAND2 NAND2_603(.VSS(VSS),.VDD(VDD),.Y(g24802),.A(I23970),.B(I23971));
  NAND2 NAND2_604(.VSS(VSS),.VDD(VDD),.Y(g29186),.A(g27051),.B(g4507));
  NAND2 NAND2_605(.VSS(VSS),.VDD(VDD),.Y(g29676),.A(g28381),.B(g13676));
  NAND3 NAND3_104(.VSS(VSS),.VDD(VDD),.Y(g7690),.A(g4669),.B(g4659),.C(g4653));
  NAND4 NAND4_95(.VSS(VSS),.VDD(VDD),.Y(g15726),.A(g6263),.B(g14529),.C(g6365),.D(g10003));
  NAND2 NAND2_606(.VSS(VSS),.VDD(VDD),.Y(I13498),.A(g255),.B(I13497));
  NAND2 NAND2_607(.VSS(VSS),.VDD(VDD),.Y(g24793),.A(g3742),.B(g23124));
  NAND2 NAND2_608(.VSS(VSS),.VDD(VDD),.Y(g26235),.A(g8016),.B(g24766));
  NAND2 NAND2_609(.VSS(VSS),.VDD(VDD),.Y(g14058),.A(g7121),.B(g11537));
  NAND2 NAND2_610(.VSS(VSS),.VDD(VDD),.Y(I26440),.A(g14271),.B(I26438));
  NAND2 NAND2_611(.VSS(VSS),.VDD(VDD),.Y(g28895),.A(g27775),.B(g8146));
  NAND2 NAND2_612(.VSS(VSS),.VDD(VDD),.Y(I14885),.A(g5489),.B(I14883));
  NAND2 NAND2_613(.VSS(VSS),.VDD(VDD),.Y(g11881),.A(g9060),.B(g3361));
  NAND2 NAND2_614(.VSS(VSS),.VDD(VDD),.Y(I14854),.A(g9433),.B(I14853));
  NAND2 NAND2_615(.VSS(VSS),.VDD(VDD),.Y(g25400),.A(g22472),.B(g12086));
  NAND2 NAND2_616(.VSS(VSS),.VDD(VDD),.Y(g12225),.A(g8324),.B(g2453));
  NAND2 NAND2_617(.VSS(VSS),.VDD(VDD),.Y(g14902),.A(g7791),.B(g12581));
  NAND2 NAND2_618(.VSS(VSS),.VDD(VDD),.Y(g12471),.A(I15288),.B(I15289));
  NAND2 NAND2_619(.VSS(VSS),.VDD(VDD),.Y(I29303),.A(g29496),.B(I29302));
  NAND2 NAND2_620(.VSS(VSS),.VDD(VDD),.Y(g12087),.A(g7431),.B(g2599));
  NAND2 NAND2_621(.VSS(VSS),.VDD(VDD),.Y(g14120),.A(g11780),.B(g4907));
  NAND4 NAND4_96(.VSS(VSS),.VDD(VDD),.Y(g14739),.A(g5929),.B(g12067),.C(g5983),.D(g12351));
  NAND2 NAND2_622(.VSS(VSS),.VDD(VDD),.Y(g10738),.A(g6961),.B(g10308));
  NAND2 NAND2_623(.VSS(VSS),.VDD(VDD),.Y(I22922),.A(g14677),.B(I22921));
  NAND2 NAND2_624(.VSS(VSS),.VDD(VDD),.Y(I25845),.A(g26212),.B(g24799));
  NAND2 NAND2_625(.VSS(VSS),.VDD(VDD),.Y(g14146),.A(g11020),.B(g691));
  NAND2 NAND2_626(.VSS(VSS),.VDD(VDD),.Y(g32072),.A(g31009),.B(g13301));
  NAND2 NAND2_627(.VSS(VSS),.VDD(VDD),.Y(g19466),.A(g11562),.B(g17794));
  NAND2 NAND2_628(.VSS(VSS),.VDD(VDD),.Y(I15003),.A(g9691),.B(I15002));
  NAND2 NAND2_629(.VSS(VSS),.VDD(VDD),.Y(g12244),.A(g7343),.B(g5320));
  NAND3 NAND3_105(.VSS(VSS),.VDD(VDD),.Y(g13248),.A(g9985),.B(g12399),.C(g9843));
  NAND2 NAND2_630(.VSS(VSS),.VDD(VDD),.Y(I14480),.A(g10074),.B(g655));
  NAND2 NAND2_631(.VSS(VSS),.VDD(VDD),.Y(g28376),.A(g27064),.B(g13620));
  NAND2 NAND2_632(.VSS(VSS),.VDD(VDD),.Y(g13779),.A(g11804),.B(g11283));
  NAND2 NAND2_633(.VSS(VSS),.VDD(VDD),.Y(I22685),.A(g21434),.B(I22683));
  NAND2 NAND2_634(.VSS(VSS),.VDD(VDD),.Y(g27955),.A(I26460),.B(I26461));
  NAND2 NAND2_635(.VSS(VSS),.VDD(VDD),.Y(g28980),.A(g27933),.B(g14680));
  NAND2 NAND2_636(.VSS(VSS),.VDD(VDD),.Y(I23987),.A(g482),.B(I23985));
  NAND2 NAND2_637(.VSS(VSS),.VDD(VDD),.Y(g23719),.A(I22845),.B(I22846));
  NAND2 NAND2_638(.VSS(VSS),.VDD(VDD),.Y(I12401),.A(g3808),.B(g3813));
  NAND2 NAND2_639(.VSS(VSS),.VDD(VDD),.Y(g28888),.A(g27738),.B(g8139));
  NAND3 NAND3_106(.VSS(VSS),.VDD(VDD),.Y(g28824),.A(g27779),.B(g7356),.C(g1772));
  NAND2 NAND2_640(.VSS(VSS),.VDD(VDD),.Y(I20488),.A(g16757),.B(I20486));
  NAND2 NAND2_641(.VSS(VSS),.VDD(VDD),.Y(I22800),.A(g11960),.B(I22799));
  NAND2 NAND2_642(.VSS(VSS),.VDD(VDD),.Y(I22936),.A(g12226),.B(g21228));
  NAND2 NAND2_643(.VSS(VSS),.VDD(VDD),.Y(g11356),.A(g9552),.B(g3632));
  NAND4 NAND4_97(.VSS(VSS),.VDD(VDD),.Y(g8691),.A(g3267),.B(g3310),.C(g3281),.D(g3303));
  NAND2 NAND2_644(.VSS(VSS),.VDD(VDD),.Y(g13945),.A(g691),.B(g11740));
  NAND3 NAND3_107(.VSS(VSS),.VDD(VDD),.Y(g19874),.A(g13665),.B(g16299),.C(g8163));
  NAND4 NAND4_98(.VSS(VSS),.VDD(VDD),.Y(g17581),.A(g5607),.B(g12029),.C(g5623),.D(g14669));
  NAND3 NAND3_108(.VSS(VSS),.VDD(VDD),.Y(g17315),.A(g9564),.B(g9516),.C(g14503));
  NAND3 NAND3_109(.VSS(VSS),.VDD(VDD),.Y(g28931),.A(g27886),.B(g2070),.C(g1996));
  NAND2 NAND2_645(.VSS(VSS),.VDD(VDD),.Y(I23969),.A(g22202),.B(g490));
  NAND2 NAND2_646(.VSS(VSS),.VDD(VDD),.Y(g14547),.A(g9439),.B(g12201));
  NAND2 NAND2_647(.VSS(VSS),.VDD(VDD),.Y(g14895),.A(g7766),.B(g12571));
  NAND2 NAND2_648(.VSS(VSS),.VDD(VDD),.Y(g11998),.A(g8324),.B(g8373));
  NAND2 NAND2_649(.VSS(VSS),.VDD(VDD),.Y(I22762),.A(g21434),.B(I22760));
  NAND2 NAND2_650(.VSS(VSS),.VDD(VDD),.Y(g13672),.A(g8933),.B(g11261));
  NAND2 NAND2_651(.VSS(VSS),.VDD(VDD),.Y(g12459),.A(g7437),.B(g5623));
  NAND4 NAND4_99(.VSS(VSS),.VDD(VDD),.Y(g16663),.A(g13854),.B(g13834),.C(g14655),.D(g12292));
  NAND2 NAND2_652(.VSS(VSS),.VDD(VDD),.Y(g10551),.A(g1728),.B(g7356));
  NAND2 NAND2_653(.VSS(VSS),.VDD(VDD),.Y(g21388),.A(g11608),.B(g17157));
  NAND3 NAND3_110(.VSS(VSS),.VDD(VDD),.Y(g24880),.A(g23281),.B(g23266),.C(g22839));
  NAND2 NAND2_654(.VSS(VSS),.VDD(VDD),.Y(g23324),.A(g703),.B(g20181));
  NAND2 NAND2_655(.VSS(VSS),.VDD(VDD),.Y(g14572),.A(g12169),.B(g9678));
  NAND2 NAND2_656(.VSS(VSS),.VDD(VDD),.Y(I14734),.A(g9732),.B(I14733));
  NAND2 NAND2_657(.VSS(VSS),.VDD(VDD),.Y(I20189),.A(g1333),.B(I20187));
  NAND2 NAND2_658(.VSS(VSS),.VDD(VDD),.Y(g21272),.A(g11268),.B(g17157));
  NAND2 NAND2_659(.VSS(VSS),.VDD(VDD),.Y(I13043),.A(g5115),.B(g5120));
  NAND2 NAND2_660(.VSS(VSS),.VDD(VDD),.Y(I14993),.A(g6527),.B(I14991));
  NAND2 NAND2_661(.VSS(VSS),.VDD(VDD),.Y(I20188),.A(g16272),.B(I20187));
  NAND3 NAND3_111(.VSS(VSS),.VDD(VDD),.Y(g13513),.A(g1351),.B(g11815),.C(g8002));
  NAND2 NAND2_662(.VSS(VSS),.VDD(VDD),.Y(g14127),.A(g11653),.B(g11435));
  NAND4 NAND4_100(.VSS(VSS),.VDD(VDD),.Y(g21462),.A(g17816),.B(g14871),.C(g17779),.D(g14829));
  NAND2 NAND2_663(.VSS(VSS),.VDD(VDD),.Y(g11961),.A(g9777),.B(g5105));
  NAND2 NAND2_664(.VSS(VSS),.VDD(VDD),.Y(g12079),.A(g1792),.B(g8195));
  NAND2 NAND2_665(.VSS(VSS),.VDD(VDD),.Y(g28860),.A(g27775),.B(g14586));
  NAND4 NAND4_101(.VSS(VSS),.VDD(VDD),.Y(g13897),.A(g3211),.B(g11217),.C(g3329),.D(g11519));
  NAND2 NAND2_666(.VSS(VSS),.VDD(VDD),.Y(I20460),.A(g17515),.B(g14187));
  NAND2 NAND2_667(.VSS(VSS),.VDD(VDD),.Y(I24383),.A(g23721),.B(g14347));
  NAND2 NAND2_668(.VSS(VSS),.VDD(VDD),.Y(g12078),.A(g8187),.B(g8093));
  NAND2 NAND2_669(.VSS(VSS),.VDD(VDD),.Y(I26071),.A(g26026),.B(I26070));
  NAND2 NAND2_670(.VSS(VSS),.VDD(VDD),.Y(I15212),.A(g10035),.B(g1714));
  NAND2 NAND2_671(.VSS(VSS),.VDD(VDD),.Y(g14956),.A(g12604),.B(g10281));
  NAND2 NAND2_672(.VSS(VSS),.VDD(VDD),.Y(I11879),.A(g4430),.B(I11877));
  NAND2 NAND2_673(.VSS(VSS),.VDD(VDD),.Y(g14889),.A(g12609),.B(g12824));
  NAND4 NAND4_102(.VSS(VSS),.VDD(VDD),.Y(g16757),.A(g13911),.B(g13886),.C(g14120),.D(g11675));
  NAND2 NAND2_674(.VSS(VSS),.VDD(VDD),.Y(I11878),.A(g4388),.B(I11877));
  NAND3 NAND3_112(.VSS(VSS),.VDD(VDD),.Y(g28987),.A(g27886),.B(g2070),.C(g7411));
  NAND3 NAND3_113(.VSS(VSS),.VDD(VDD),.Y(g25435),.A(g22432),.B(g2342),.C(g8316));
  NAND2 NAND2_675(.VSS(VSS),.VDD(VDD),.Y(I23979),.A(g23198),.B(I23978));
  NAND2 NAND2_676(.VSS(VSS),.VDD(VDD),.Y(g24989),.A(g21345),.B(g23363));
  NAND2 NAND2_677(.VSS(VSS),.VDD(VDD),.Y(g12159),.A(g8765),.B(g4864));
  NAND2 NAND2_678(.VSS(VSS),.VDD(VDD),.Y(g12125),.A(g9728),.B(g5101));
  NAND2 NAND2_679(.VSS(VSS),.VDD(VDD),.Y(I21978),.A(g19620),.B(I21976));
  NAND2 NAND2_680(.VSS(VSS),.VDD(VDD),.Y(I22974),.A(g19638),.B(I22972));
  NAND2 NAND2_681(.VSS(VSS),.VDD(VDD),.Y(I23978),.A(g23198),.B(g13670));
  NAND2 NAND2_682(.VSS(VSS),.VDD(VDD),.Y(g24988),.A(g546),.B(g23088));
  NAND2 NAND2_683(.VSS(VSS),.VDD(VDD),.Y(g24924),.A(g20007),.B(g23172));
  NAND2 NAND2_684(.VSS(VSS),.VDD(VDD),.Y(I15149),.A(g5659),.B(I15147));
  NAND2 NAND2_685(.VSS(VSS),.VDD(VDD),.Y(g21360),.A(g11510),.B(g17157));
  NAND2 NAND2_686(.VSS(VSS),.VDD(VDD),.Y(I23986),.A(g22182),.B(I23985));
  NAND2 NAND2_687(.VSS(VSS),.VDD(VDD),.Y(g27295),.A(g24776),.B(g26208));
  NAND4 NAND4_103(.VSS(VSS),.VDD(VDD),.Y(g20271),.A(g16925),.B(g14054),.C(g16657),.D(g16628));
  NAND2 NAND2_688(.VSS(VSS),.VDD(VDD),.Y(g11149),.A(g1564),.B(g7948));
  NAND2 NAND2_689(.VSS(VSS),.VDD(VDD),.Y(I15148),.A(g9864),.B(I15147));
  NAND2 NAND2_690(.VSS(VSS),.VDD(VDD),.Y(g28969),.A(g27854),.B(g8267));
  NAND2 NAND2_691(.VSS(VSS),.VDD(VDD),.Y(I26367),.A(g26400),.B(I26366));
  NAND2 NAND2_692(.VSS(VSS),.VDD(VDD),.Y(I26394),.A(g26488),.B(I26393));
  NAND2 NAND2_693(.VSS(VSS),.VDD(VDD),.Y(g12144),.A(I15003),.B(I15004));
  NAND2 NAND2_694(.VSS(VSS),.VDD(VDD),.Y(g9543),.A(g2217),.B(g2185));
  NAND4 NAND4_104(.VSS(VSS),.VDD(VDD),.Y(g13097),.A(g5204),.B(g12002),.C(g5339),.D(g9780));
  NAND2 NAND2_695(.VSS(VSS),.VDD(VDD),.Y(g10520),.A(g7195),.B(g7115));
  NAND2 NAND2_696(.VSS(VSS),.VDD(VDD),.Y(g13104),.A(g1404),.B(g10794));
  NAND2 NAND2_697(.VSS(VSS),.VDD(VDD),.Y(g12336),.A(I15175),.B(I15176));
  NAND2 NAND2_698(.VSS(VSS),.VDD(VDD),.Y(g14520),.A(g9369),.B(g12163));
  NAND2 NAND2_699(.VSS(VSS),.VDD(VDD),.Y(I14187),.A(g3470),.B(I14185));
  NAND2 NAND2_700(.VSS(VSS),.VDD(VDD),.Y(g7150),.A(g5016),.B(g5062));
  NAND2 NAND2_701(.VSS(VSS),.VDD(VDD),.Y(I25220),.A(g482),.B(I25219));
  NAND4 NAND4_105(.VSS(VSS),.VDD(VDD),.Y(g20199),.A(g16815),.B(g13968),.C(g16749),.D(g13907));
  NAND2 NAND2_702(.VSS(VSS),.VDD(VDD),.Y(g11971),.A(g8249),.B(g8302));
  NAND2 NAND2_703(.VSS(VSS),.VDD(VDD),.Y(g28870),.A(g27796),.B(g14588));
  NAND3 NAND3_114(.VSS(VSS),.VDD(VDD),.Y(g34048),.A(g33669),.B(g10583),.C(g7442));
  NAND2 NAND2_704(.VSS(VSS),.VDD(VDD),.Y(I13079),.A(g5467),.B(I13077));
  NAND2 NAND2_705(.VSS(VSS),.VDD(VDD),.Y(I13444),.A(g239),.B(I13442));
  NAND2 NAND2_706(.VSS(VSS),.VDD(VDD),.Y(I32432),.A(g34056),.B(I32431));
  NAND2 NAND2_707(.VSS(VSS),.VDD(VDD),.Y(g14546),.A(g12125),.B(g9613));
  NAND2 NAND2_708(.VSS(VSS),.VDD(VDD),.Y(g14089),.A(g11755),.B(g4717));
  NAND2 NAND2_709(.VSS(VSS),.VDD(VDD),.Y(g22688),.A(g20219),.B(g2936));
  NAND4 NAND4_106(.VSS(VSS),.VDD(VDD),.Y(g20198),.A(g16813),.B(g13958),.C(g16745),.D(g13927));
  NAND4 NAND4_107(.VSS(VSS),.VDD(VDD),.Y(g17706),.A(g3921),.B(g11255),.C(g3983),.D(g13933));
  NAND4 NAND4_108(.VSS(VSS),.VDD(VDD),.Y(g17597),.A(g3191),.B(g13700),.C(g3303),.D(g8481));
  NAND2 NAND2_710(.VSS(VSS),.VDD(VDD),.Y(I12074),.A(g996),.B(g979));
  NAND2 NAND2_711(.VSS(VSS),.VDD(VDD),.Y(I13078),.A(g5462),.B(I13077));
  NAND4 NAND4_109(.VSS(VSS),.VDD(VDD),.Y(g14088),.A(g3901),.B(g11255),.C(g4000),.D(g11631));
  NAND2 NAND2_712(.VSS(VSS),.VDD(VDD),.Y(g14024),.A(g7121),.B(g11763));
  NAND4 NAND4_110(.VSS(VSS),.VDD(VDD),.Y(g17689),.A(g6645),.B(g12137),.C(g6661),.D(g14786));
  NAND2 NAND2_713(.VSS(VSS),.VDD(VDD),.Y(I18589),.A(g14679),.B(I18587));
  NAND2 NAND2_714(.VSS(VSS),.VDD(VDD),.Y(g24528),.A(g4098),.B(g22654));
  NAND2 NAND2_715(.VSS(VSS),.VDD(VDD),.Y(g17624),.A(I18588),.B(I18589));
  NAND3 NAND3_115(.VSS(VSS),.VDD(VDD),.Y(g28867),.A(g27800),.B(g2227),.C(g2153));
  NAND2 NAND2_716(.VSS(VSS),.VDD(VDD),.Y(I18588),.A(g2370),.B(I18587));
  NAND2 NAND2_717(.VSS(VSS),.VDD(VDD),.Y(g7836),.A(g4653),.B(g4688));
  NAND2 NAND2_718(.VSS(VSS),.VDD(VDD),.Y(I20467),.A(g16663),.B(g16728));
  NAND2 NAND2_719(.VSS(VSS),.VDD(VDD),.Y(I14169),.A(g8389),.B(g3119));
  NAND2 NAND2_720(.VSS(VSS),.VDD(VDD),.Y(I14884),.A(g9500),.B(I14883));
  NAND3 NAND3_116(.VSS(VSS),.VDD(VDD),.Y(g11412),.A(g8666),.B(g6918),.C(g8697));
  NAND2 NAND2_721(.VSS(VSS),.VDD(VDD),.Y(g15702),.A(g13066),.B(g7293));
  NAND2 NAND2_722(.VSS(VSS),.VDD(VDD),.Y(g13850),.A(g11279),.B(g8396));
  NAND2 NAND2_723(.VSS(VSS),.VDD(VDD),.Y(g15904),.A(I17380),.B(I17381));
  NAND2 NAND2_724(.VSS(VSS),.VDD(VDD),.Y(g25049),.A(g21344),.B(g23462));
  NAND3 NAND3_117(.VSS(VSS),.VDD(VDD),.Y(g12289),.A(g9978),.B(g9766),.C(g9708));
  NAND2 NAND2_725(.VSS(VSS),.VDD(VDD),.Y(g14659),.A(g12646),.B(g12443));
  NAND4 NAND4_111(.VSS(VSS),.VDD(VDD),.Y(g14625),.A(g3897),.B(g11225),.C(g4031),.D(g8595));
  NAND4 NAND4_112(.VSS(VSS),.VDD(VDD),.Y(g14987),.A(g6593),.B(g12211),.C(g6692),.D(g12721));
  NAND4 NAND4_113(.VSS(VSS),.VDD(VDD),.Y(g20161),.A(g17732),.B(g17706),.C(g17670),.D(g14625));
  NAND2 NAND2_726(.VSS(VSS),.VDD(VDD),.Y(g22885),.A(g9104),.B(g20154));
  NAND2 NAND2_727(.VSS(VSS),.VDD(VDD),.Y(g12023),.A(g2453),.B(g8373));
  NAND2 NAND2_728(.VSS(VSS),.VDD(VDD),.Y(g28910),.A(g27854),.B(g14614));
  NAND4 NAND4_114(.VSS(VSS),.VDD(VDD),.Y(g13896),.A(g3227),.B(g11194),.C(g3281),.D(g11350));
  NAND2 NAND2_729(.VSS(VSS),.VDD(VDD),.Y(I23917),.A(g23975),.B(g9333));
  NAND2 NAND2_730(.VSS(VSS),.VDD(VDD),.Y(g25048),.A(g542),.B(g23088));
  NAND2 NAND2_731(.VSS(VSS),.VDD(VDD),.Y(g12224),.A(I15088),.B(I15089));
  NAND2 NAND2_732(.VSS(VSS),.VDD(VDD),.Y(g14943),.A(g7791),.B(g12622));
  NAND2 NAND2_733(.VSS(VSS),.VDD(VDD),.Y(I13336),.A(g1691),.B(I13334));
  NAND2 NAND2_734(.VSS(VSS),.VDD(VDD),.Y(g27687),.A(g25200),.B(g26714));
  NAND2 NAND2_735(.VSS(VSS),.VDD(VDD),.Y(g14968),.A(g12739),.B(g10312));
  NAND2 NAND2_736(.VSS(VSS),.VDD(VDD),.Y(g11959),.A(g8316),.B(g2342));
  NAND2 NAND2_737(.VSS(VSS),.VDD(VDD),.Y(g13627),.A(g11172),.B(g8388));
  NAND2 NAND2_738(.VSS(VSS),.VDD(VDD),.Y(I22684),.A(g11893),.B(I22683));
  NAND2 NAND2_739(.VSS(VSS),.VDD(VDD),.Y(I20167),.A(g990),.B(I20165));
  NAND2 NAND2_740(.VSS(VSS),.VDD(VDD),.Y(g14855),.A(g12700),.B(g12824));
  NAND2 NAND2_741(.VSS(VSS),.VDD(VDD),.Y(I12729),.A(g4291),.B(I12728));
  NAND4 NAND4_115(.VSS(VSS),.VDD(VDD),.Y(g13050),.A(g5543),.B(g12029),.C(g5654),.D(g9864));
  NAND4 NAND4_116(.VSS(VSS),.VDD(VDD),.Y(g13958),.A(g3610),.B(g11238),.C(g3618),.D(g11389));
  NAND2 NAND2_742(.VSS(VSS),.VDD(VDD),.Y(I12728),.A(g4291),.B(g4287));
  NAND3 NAND3_118(.VSS(VSS),.VDD(VDD),.Y(g28877),.A(g27937),.B(g7490),.C(g7431));
  NAND2 NAND2_743(.VSS(VSS),.VDD(VDD),.Y(g20068),.A(g11293),.B(g17794));
  NAND2 NAND2_744(.VSS(VSS),.VDD(VDD),.Y(I26366),.A(g26400),.B(g14211));
  NAND2 NAND2_745(.VSS(VSS),.VDD(VDD),.Y(I14531),.A(g8840),.B(I14530));
  NAND2 NAND2_746(.VSS(VSS),.VDD(VDD),.Y(g13742),.A(g11780),.B(g11283));
  NAND2 NAND2_747(.VSS(VSS),.VDD(VDD),.Y(g11944),.A(I14765),.B(I14766));
  NAND2 NAND2_748(.VSS(VSS),.VDD(VDD),.Y(g7620),.A(I12097),.B(I12098));
  NAND2 NAND2_749(.VSS(VSS),.VDD(VDD),.Y(g8010),.A(I12345),.B(I12346));
  NAND2 NAND2_750(.VSS(VSS),.VDD(VDD),.Y(I14186),.A(g8442),.B(I14185));
  NAND2 NAND2_751(.VSS(VSS),.VDD(VDD),.Y(g17287),.A(g7262),.B(g14228));
  NAND2 NAND2_752(.VSS(VSS),.VDD(VDD),.Y(g12195),.A(g2619),.B(g8381));
  NAND2 NAND2_753(.VSS(VSS),.VDD(VDD),.Y(g17596),.A(g8686),.B(g14367));
  NAND2 NAND2_754(.VSS(VSS),.VDD(VDD),.Y(g25514),.A(g12540),.B(g22498));
  NAND2 NAND2_755(.VSS(VSS),.VDD(VDD),.Y(g24792),.A(I23950),.B(I23951));
  NAND2 NAND2_756(.VSS(VSS),.VDD(VDD),.Y(g17243),.A(g7247),.B(g14212));
  NAND2 NAND2_757(.VSS(VSS),.VDD(VDD),.Y(g12525),.A(g7522),.B(g6668));
  NAND2 NAND2_758(.VSS(VSS),.VDD(VDD),.Y(g12016),.A(g1648),.B(g8093));
  NAND2 NAND2_759(.VSS(VSS),.VDD(VDD),.Y(g23281),.A(g18957),.B(g2898));
  NAND2 NAND2_760(.VSS(VSS),.VDD(VDD),.Y(g21301),.A(g11371),.B(g17157));
  NAND2 NAND2_761(.VSS(VSS),.VDD(VDD),.Y(g21377),.A(g11560),.B(g17157));
  NAND2 NAND2_762(.VSS(VSS),.VDD(VDD),.Y(g14055),.A(g11697),.B(g11763));
  NAND4 NAND4_117(.VSS(VSS),.VDD(VDD),.Y(g17773),.A(g5965),.B(g14549),.C(g5976),.D(g9935));
  NAND2 NAND2_763(.VSS(VSS),.VDD(VDD),.Y(I18485),.A(g1677),.B(g14611));
  NAND2 NAND2_764(.VSS(VSS),.VDD(VDD),.Y(g14978),.A(g12716),.B(g10491));
  NAND4 NAND4_118(.VSS(VSS),.VDD(VDD),.Y(g15780),.A(g5937),.B(g14549),.C(g6012),.D(g14701));
  NAND2 NAND2_765(.VSS(VSS),.VDD(VDD),.Y(I17475),.A(g13336),.B(I17474));
  NAND4 NAND4_119(.VSS(VSS),.VDD(VDD),.Y(g14590),.A(g3546),.B(g11207),.C(g3680),.D(g8542));
  NAND2 NAND2_766(.VSS(VSS),.VDD(VDD),.Y(g24918),.A(g136),.B(g23088));
  NAND4 NAND4_120(.VSS(VSS),.VDD(VDD),.Y(g17670),.A(g3893),.B(g13772),.C(g4005),.D(g8595));
  NAND2 NAND2_767(.VSS(VSS),.VDD(VDD),.Y(g22839),.A(g20114),.B(g2988));
  NAND2 NAND2_768(.VSS(VSS),.VDD(VDD),.Y(g23699),.A(g21012),.B(g11160));
  NAND2 NAND2_769(.VSS(VSS),.VDD(VDD),.Y(I29302),.A(g29496),.B(g12121));
  NAND2 NAND2_770(.VSS(VSS),.VDD(VDD),.Y(g25473),.A(g12437),.B(g22432));
  NAND2 NAND2_771(.VSS(VSS),.VDD(VDD),.Y(g14741),.A(g12711),.B(g10421));
  NAND2 NAND2_772(.VSS(VSS),.VDD(VDD),.Y(g27705),.A(g25237),.B(g26782));
  NAND2 NAND2_773(.VSS(VSS),.VDD(VDD),.Y(g22838),.A(g20219),.B(g2960));
  NAND4 NAND4_121(.VSS(VSS),.VDD(VDD),.Y(g17734),.A(g5272),.B(g14490),.C(g5283),.D(g9780));
  NAND2 NAND2_774(.VSS(VSS),.VDD(VDD),.Y(g28923),.A(g27775),.B(g8195));
  NAND3 NAND3_119(.VSS(VSS),.VDD(VDD),.Y(g16282),.A(g4933),.B(g13939),.C(g12088));
  NAND2 NAND2_775(.VSS(VSS),.VDD(VDD),.Y(g9442),.A(g5424),.B(g5428));
  NAND2 NAND2_776(.VSS(VSS),.VDD(VDD),.Y(g27679),.A(g25186),.B(g26685));
  NAND2 NAND2_777(.VSS(VSS),.VDD(VDD),.Y(I15129),.A(g9914),.B(I15128));
  NAND2 NAND2_778(.VSS(VSS),.VDD(VDD),.Y(g12042),.A(g9086),.B(g703));
  NAND2 NAND2_779(.VSS(VSS),.VDD(VDD),.Y(I15002),.A(g9691),.B(g1700));
  NAND2 NAND2_780(.VSS(VSS),.VDD(VDD),.Y(I26095),.A(g13539),.B(I26093));
  NAND2 NAND2_781(.VSS(VSS),.VDD(VDD),.Y(g12255),.A(g9958),.B(g6140));
  NAND2 NAND2_782(.VSS(VSS),.VDD(VDD),.Y(g11002),.A(g7475),.B(g862));
  NAND2 NAND2_783(.VSS(VSS),.VDD(VDD),.Y(I15128),.A(g9914),.B(g2527));
  NAND2 NAND2_784(.VSS(VSS),.VDD(VDD),.Y(g13057),.A(g969),.B(g11294));
  NAND2 NAND2_785(.VSS(VSS),.VDD(VDD),.Y(g14735),.A(g12739),.B(g12571));
  NAND2 NAND2_786(.VSS(VSS),.VDD(VDD),.Y(g12188),.A(g8249),.B(g1894));
  NAND2 NAND2_787(.VSS(VSS),.VDD(VDD),.Y(g12124),.A(g8741),.B(g4674));
  NAND2 NAND2_788(.VSS(VSS),.VDD(VDD),.Y(I13392),.A(g1825),.B(I13390));
  NAND3 NAND3_120(.VSS(VSS),.VDD(VDD),.Y(g11245),.A(g7636),.B(g7733),.C(g7697));
  NAND2 NAND2_789(.VSS(VSS),.VDD(VDD),.Y(I15299),.A(g10112),.B(I15298));
  NAND3 NAND3_121(.VSS(VSS),.VDD(VDD),.Y(g12460),.A(g10093),.B(g5644),.C(g5694));
  NAND3 NAND3_122(.VSS(VSS),.VDD(VDD),.Y(g12686),.A(g7097),.B(g6682),.C(g6736));
  NAND2 NAND2_790(.VSS(VSS),.VDD(VDD),.Y(I20166),.A(g16246),.B(I20165));
  NAND2 NAND2_791(.VSS(VSS),.VDD(VDD),.Y(g11323),.A(I14351),.B(I14352));
  NAND4 NAND4_122(.VSS(VSS),.VDD(VDD),.Y(g14695),.A(g5583),.B(g12029),.C(g5637),.D(g12301));
  NAND2 NAND2_792(.VSS(VSS),.VDD(VDD),.Y(g14018),.A(g10323),.B(g11483));
  NAND2 NAND2_793(.VSS(VSS),.VDD(VDD),.Y(I15298),.A(g10112),.B(g1982));
  NAND3 NAND3_123(.VSS(VSS),.VDD(VDD),.Y(g11533),.A(g6905),.B(g3639),.C(g3698));
  NAND2 NAND2_794(.VSS(VSS),.VDD(VDD),.Y(g21403),.A(g11652),.B(g17157));
  NAND2 NAND2_795(.VSS(VSS),.VDD(VDD),.Y(g20783),.A(g14616),.B(g17225));
  NAND3 NAND3_124(.VSS(VSS),.VDD(VDD),.Y(g12294),.A(g10044),.B(g7018),.C(g10090));
  NAND2 NAND2_796(.VSS(VSS),.VDD(VDD),.Y(g17618),.A(I18580),.B(I18581));
  NAND3 NAND3_125(.VSS(VSS),.VDD(VDD),.Y(g28885),.A(g27742),.B(g1668),.C(g7268));
  NAND4 NAND4_123(.VSS(VSS),.VDD(VDD),.Y(g22306),.A(g4584),.B(g4616),.C(g13202),.D(g19071));
  NAND2 NAND2_797(.VSS(VSS),.VDD(VDD),.Y(I22873),.A(g21228),.B(I22871));
  NAND2 NAND2_798(.VSS(VSS),.VDD(VDD),.Y(I11865),.A(g4434),.B(I11864));
  NAND2 NAND2_799(.VSS(VSS),.VDD(VDD),.Y(I14230),.A(g8055),.B(I14228));
  NAND4 NAND4_124(.VSS(VSS),.VDD(VDD),.Y(g17468),.A(g3215),.B(g13700),.C(g3317),.D(g8481));
  NAND2 NAND2_800(.VSS(VSS),.VDD(VDD),.Y(I21993),.A(g7670),.B(I21992));
  NAND4 NAND4_125(.VSS(VSS),.VDD(VDD),.Y(g15787),.A(g6283),.B(g14575),.C(g6358),.D(g14745));
  NAND4 NAND4_126(.VSS(VSS),.VDD(VDD),.Y(g14706),.A(g6287),.B(g12101),.C(g6369),.D(g12672));
  NAND2 NAND2_801(.VSS(VSS),.VDD(VDD),.Y(I14992),.A(g9685),.B(I14991));
  NAND4 NAND4_127(.VSS(VSS),.VDD(VDD),.Y(g21385),.A(g17736),.B(g14696),.C(g17679),.D(g14636));
  NAND2 NAND2_802(.VSS(VSS),.VDD(VDD),.Y(I14510),.A(g8721),.B(I14508));
  NAND4 NAND4_128(.VSS(VSS),.VDD(VDD),.Y(g15743),.A(g5893),.B(g14497),.C(g6005),.D(g9935));
  NAND2 NAND2_803(.VSS(VSS),.VDD(VDD),.Y(g21354),.A(g11468),.B(g17157));
  NAND2 NAND2_804(.VSS(VSS),.VDD(VDD),.Y(g14688),.A(g12604),.B(g12453));
  NAND3 NAND3_126(.VSS(VSS),.VDD(VDD),.Y(g28287),.A(g10504),.B(g26131),.C(g26973));
  NAND2 NAND2_805(.VSS(VSS),.VDD(VDD),.Y(g12915),.A(g12806),.B(g12632));
  NAND2 NAND2_806(.VSS(VSS),.VDD(VDD),.Y(I13383),.A(g269),.B(I13382));
  NAND2 NAND2_807(.VSS(VSS),.VDD(VDD),.Y(g11445),.A(g9771),.B(g3976));
  NAND2 NAND2_808(.VSS(VSS),.VDD(VDD),.Y(g14157),.A(g11715),.B(g11763));
  NAND2 NAND2_809(.VSS(VSS),.VDD(VDD),.Y(g22666),.A(g18957),.B(g2878));
  NAND4 NAND4_129(.VSS(VSS),.VDD(VDD),.Y(g13499),.A(g11479),.B(g11442),.C(g11410),.D(g11382));
  NAND2 NAND2_810(.VSS(VSS),.VDD(VDD),.Y(I13065),.A(g4308),.B(g4304));
  NAND2 NAND2_811(.VSS(VSS),.VDD(VDD),.Y(g14066),.A(g11514),.B(g11473));
  NAND4 NAND4_130(.VSS(VSS),.VDD(VDD),.Y(g13498),.A(g12577),.B(g12522),.C(g12462),.D(g12416));
  NAND2 NAND2_812(.VSS(VSS),.VDD(VDD),.Y(I15080),.A(g1968),.B(I15078));
  NAND2 NAND2_813(.VSS(VSS),.VDD(VDD),.Y(g17363),.A(g8635),.B(g14367));
  NAND3 NAND3_127(.VSS(VSS),.VDD(VDD),.Y(g28942),.A(g27858),.B(g2331),.C(g7335));
  NAND2 NAND2_814(.VSS(VSS),.VDD(VDD),.Y(g17217),.A(g7239),.B(g14194));
  NAND2 NAND2_815(.VSS(VSS),.VDD(VDD),.Y(g21190),.A(g6077),.B(g17420));
  NAND2 NAND2_816(.VSS(VSS),.VDD(VDD),.Y(g14876),.A(g12492),.B(g12443));
  NAND2 NAND2_817(.VSS(VSS),.VDD(VDD),.Y(g14885),.A(g12651),.B(g12505));
  NAND4 NAND4_131(.VSS(VSS),.VDD(VDD),.Y(g14854),.A(g5555),.B(g12093),.C(g5654),.D(g12563));
  NAND3 NAND3_128(.VSS(VSS),.VDD(VDD),.Y(g10511),.A(g4628),.B(g7202),.C(g4621));
  NAND2 NAND2_818(.VSS(VSS),.VDD(VDD),.Y(g11432),.A(g10295),.B(g8864));
  NAND2 NAND2_819(.VSS(VSS),.VDD(VDD),.Y(I23601),.A(g22360),.B(I23600));
  NAND2 NAND2_820(.VSS(VSS),.VDD(VDD),.Y(g13432),.A(g4793),.B(g10831));
  NAND2 NAND2_821(.VSS(VSS),.VDD(VDD),.Y(I14275),.A(g8218),.B(g3484));
  NAND2 NAND2_822(.VSS(VSS),.VDD(VDD),.Y(g12155),.A(g7753),.B(g7717));
  NAND4 NAND4_132(.VSS(VSS),.VDD(VDD),.Y(g12822),.A(g6978),.B(g7236),.C(g7224),.D(g7163));
  NAND2 NAND2_823(.VSS(VSS),.VDD(VDD),.Y(g15027),.A(g12667),.B(g10341));
  NAND2 NAND2_824(.VSS(VSS),.VDD(VDD),.Y(I15342),.A(g2541),.B(I15340));
  NAND2 NAND2_825(.VSS(VSS),.VDD(VDD),.Y(g28930),.A(g27833),.B(g8201));
  NAND2 NAND2_826(.VSS(VSS),.VDD(VDD),.Y(I24439),.A(g23771),.B(I24438));
  NAND2 NAND2_827(.VSS(VSS),.VDD(VDD),.Y(g28965),.A(g27882),.B(g8255));
  NAND2 NAND2_828(.VSS(VSS),.VDD(VDD),.Y(g30573),.A(g29355),.B(g19666));
  NAND2 NAND2_829(.VSS(VSS),.VDD(VDD),.Y(I24438),.A(g23771),.B(g14411));
  NAND2 NAND2_830(.VSS(VSS),.VDD(VDD),.Y(g15710),.A(g319),.B(g13385));
  NAND2 NAND2_831(.VSS(VSS),.VDD(VDD),.Y(g9715),.A(g5011),.B(g4836));
  NAND2 NAND2_832(.VSS(VSS),.VDD(VDD),.Y(g28131),.A(g27051),.B(g25838));
  NAND3 NAND3_129(.VSS(VSS),.VDD(VDD),.Y(g31509),.A(g599),.B(g29933),.C(g12323));
  NAND2 NAND2_833(.VSS(VSS),.VDD(VDD),.Y(g10916),.A(g1146),.B(g7854));
  NAND2 NAND2_834(.VSS(VSS),.VDD(VDD),.Y(I12241),.A(g1111),.B(I12240));
  NAND4 NAND4_133(.VSS(VSS),.VDD(VDD),.Y(g33933),.A(g33394),.B(g12491),.C(g12819),.D(g12796));
  NAND2 NAND2_835(.VSS(VSS),.VDD(VDD),.Y(g12589),.A(g7591),.B(g6692));
  NAND2 NAND2_836(.VSS(VSS),.VDD(VDD),.Y(g12194),.A(g8373),.B(g8273));
  NAND2 NAND2_837(.VSS(VSS),.VDD(VDD),.Y(g10550),.A(g7268),.B(g7308));
  NAND4 NAND4_134(.VSS(VSS),.VDD(VDD),.Y(g13529),.A(g11590),.B(g11544),.C(g11492),.D(g11446));
  NAND2 NAND2_838(.VSS(VSS),.VDD(VDD),.Y(I14517),.A(g10147),.B(I14516));
  NAND3 NAND3_130(.VSS(VSS),.VDD(VDD),.Y(g12588),.A(g10169),.B(g6336),.C(g6386));
  NAND2 NAND2_839(.VSS(VSS),.VDD(VDD),.Y(g27401),.A(I26094),.B(I26095));
  NAND3 NAND3_131(.VSS(VSS),.VDD(VDD),.Y(g12524),.A(g7074),.B(g7087),.C(g10212));
  NAND2 NAND2_840(.VSS(VSS),.VDD(VDD),.Y(g23659),.A(g9434),.B(g20854));
  NAND2 NAND2_841(.VSS(VSS),.VDD(VDD),.Y(g11330),.A(g9483),.B(g1193));
  NAND3 NAND3_132(.VSS(VSS),.VDD(VDD),.Y(g13528),.A(g11294),.B(g7549),.C(g1008));
  NAND2 NAND2_842(.VSS(VSS),.VDD(VDD),.Y(g13330),.A(g4664),.B(g11006));
  NAND2 NAND2_843(.VSS(VSS),.VDD(VDD),.Y(g10307),.A(I13730),.B(I13731));
  NAND2 NAND2_844(.VSS(VSS),.VDD(VDD),.Y(I15365),.A(g2675),.B(I15363));
  NAND2 NAND2_845(.VSS(VSS),.VDD(VDD),.Y(g14085),.A(g7121),.B(g11584));
  NAND4 NAND4_135(.VSS(VSS),.VDD(VDD),.Y(g17740),.A(g5945),.B(g14497),.C(g6012),.D(g12351));
  NAND2 NAND2_846(.VSS(VSS),.VDD(VDD),.Y(g13764),.A(g11252),.B(g3072));
  NAND2 NAND2_847(.VSS(VSS),.VDD(VDD),.Y(g8238),.A(I12469),.B(I12470));
  NAND4 NAND4_136(.VSS(VSS),.VDD(VDD),.Y(g14596),.A(g12196),.B(g9775),.C(g12124),.D(g9663));
  NAND2 NAND2_848(.VSS(VSS),.VDD(VDD),.Y(g12119),.A(g2351),.B(g8267));
  NAND4 NAND4_137(.VSS(VSS),.VDD(VDD),.Y(g14054),.A(g3550),.B(g11238),.C(g3649),.D(g11576));
  NAND2 NAND2_849(.VSS(VSS),.VDD(VDD),.Y(I22711),.A(g11915),.B(I22710));
  NAND3 NAND3_133(.VSS(VSS),.VDD(VDD),.Y(g7701),.A(g4859),.B(g4849),.C(g4843));
  NAND4 NAND4_138(.VSS(VSS),.VDD(VDD),.Y(g21339),.A(g15725),.B(g13084),.C(g15713),.D(g13050));
  NAND2 NAND2_850(.VSS(VSS),.VDD(VDD),.Y(g13960),.A(g11669),.B(g11537));
  NAND2 NAND2_851(.VSS(VSS),.VDD(VDD),.Y(g32057),.A(g31003),.B(g13297));
  NAND2 NAND2_852(.VSS(VSS),.VDD(VDD),.Y(g12118),.A(g8259),.B(g8150));
  NAND2 NAND2_853(.VSS(VSS),.VDD(VDD),.Y(g12022),.A(g7335),.B(g2331));
  NAND4 NAND4_139(.VSS(VSS),.VDD(VDD),.Y(g21338),.A(g15741),.B(g15734),.C(g15728),.D(g13097));
  NAND2 NAND2_854(.VSS(VSS),.VDD(VDD),.Y(I26070),.A(g26026),.B(g13517));
  NAND2 NAND2_855(.VSS(VSS),.VDD(VDD),.Y(I17474),.A(g13336),.B(g1105));
  NAND4 NAND4_140(.VSS(VSS),.VDD(VDD),.Y(g16723),.A(g3606),.B(g13730),.C(g3676),.D(g11576));
  NAND2 NAND2_856(.VSS(VSS),.VDD(VDD),.Y(g14773),.A(g12711),.B(g12581));
  NAND3 NAND3_134(.VSS(VSS),.VDD(VDD),.Y(g24544),.A(g22666),.B(g22661),.C(g22651));
  NAND2 NAND2_857(.VSS(VSS),.VDD(VDD),.Y(g13709),.A(g11755),.B(g11261));
  NAND2 NAND2_858(.VSS(VSS),.VDD(VDD),.Y(g25389),.A(g22457),.B(g12082));
  NAND2 NAND2_859(.VSS(VSS),.VDD(VDD),.Y(g12285),.A(I15122),.B(I15123));
  NAND2 NAND2_860(.VSS(VSS),.VDD(VDD),.Y(I15087),.A(g9832),.B(g2393));
  NAND2 NAND2_861(.VSS(VSS),.VDD(VDD),.Y(g14655),.A(g4743),.B(g11755));
  NAND2 NAND2_862(.VSS(VSS),.VDD(VDD),.Y(g11708),.A(g10147),.B(g10110));
  NAND2 NAND2_863(.VSS(VSS),.VDD(VDD),.Y(g13708),.A(g11200),.B(g8507));
  NAND2 NAND2_864(.VSS(VSS),.VDD(VDD),.Y(g12053),.A(g2587),.B(g8418));
  NAND2 NAND2_865(.VSS(VSS),.VDD(VDD),.Y(g16097),.A(g13319),.B(g10998));
  NAND2 NAND2_866(.VSS(VSS),.VDD(VDD),.Y(I26094),.A(g26055),.B(I26093));
  NAND2 NAND2_867(.VSS(VSS),.VDD(VDD),.Y(I24415),.A(g23751),.B(I24414));
  NAND2 NAND2_868(.VSS(VSS),.VDD(VDD),.Y(I15043),.A(g1834),.B(I15041));
  NAND2 NAND2_869(.VSS(VSS),.VDD(VDD),.Y(g13043),.A(g10521),.B(g969));
  NAND2 NAND2_870(.VSS(VSS),.VDD(VDD),.Y(g14930),.A(g12609),.B(g12515));
  NAND2 NAND2_871(.VSS(VSS),.VDD(VDD),.Y(g14993),.A(g12695),.B(g12453));
  NAND2 NAND2_872(.VSS(VSS),.VDD(VDD),.Y(I17381),.A(g1129),.B(I17379));
  NAND2 NAND2_873(.VSS(VSS),.VDD(VDD),.Y(g24678),.A(g22994),.B(g23010));
  NAND2 NAND2_874(.VSS(VSS),.VDD(VDD),.Y(g14838),.A(g12492),.B(g12405));
  NAND2 NAND2_875(.VSS(VSS),.VDD(VDD),.Y(g14965),.A(g12609),.B(g12571));
  NAND2 NAND2_876(.VSS(VSS),.VDD(VDD),.Y(g22908),.A(g9104),.B(g20175));
  NAND4 NAND4_141(.VSS(VSS),.VDD(VDD),.Y(g13069),.A(g5889),.B(g12067),.C(g6000),.D(g9935));
  NAND2 NAND2_877(.VSS(VSS),.VDD(VDD),.Y(g29702),.A(g28395),.B(g13712));
  NAND3 NAND3_135(.VSS(VSS),.VDD(VDD),.Y(g34162),.A(g785),.B(g33823),.C(g11679));
  NAND2 NAND2_878(.VSS(VSS),.VDD(VDD),.Y(g15717),.A(g10754),.B(g13092));
  NAND2 NAND2_879(.VSS(VSS),.VDD(VDD),.Y(I13401),.A(g2246),.B(g2250));
  NAND2 NAND2_880(.VSS(VSS),.VDD(VDD),.Y(g11955),.A(g8302),.B(g1917));
  NAND2 NAND2_881(.VSS(VSS),.VDD(VDD),.Y(g13955),.A(g11621),.B(g11527));
  NAND2 NAND2_882(.VSS(VSS),.VDD(VDD),.Y(g11970),.A(g1760),.B(g8241));
  NAND2 NAND2_883(.VSS(VSS),.VDD(VDD),.Y(g28410),.A(g27074),.B(g13679));
  NAND2 NAND2_884(.VSS(VSS),.VDD(VDD),.Y(g19962),.A(g11470),.B(g17794));
  NAND2 NAND2_885(.VSS(VSS),.VDD(VDD),.Y(g10618),.A(g10153),.B(g9913));
  NAND2 NAND2_886(.VSS(VSS),.VDD(VDD),.Y(I14351),.A(g8890),.B(I14350));
  NAND2 NAND2_887(.VSS(VSS),.VDD(VDD),.Y(g27693),.A(g25216),.B(g26752));
  NAND2 NAND2_888(.VSS(VSS),.VDD(VDD),.Y(I11864),.A(g4434),.B(g4401));
  NAND2 NAND2_889(.VSS(VSS),.VDD(VDD),.Y(g34220),.A(I32186),.B(I32187));
  NAND2 NAND2_890(.VSS(VSS),.VDD(VDD),.Y(g28363),.A(g27064),.B(g13593));
  NAND2 NAND2_891(.VSS(VSS),.VDD(VDD),.Y(g17568),.A(I18486),.B(I18487));
  NAND2 NAND2_892(.VSS(VSS),.VDD(VDD),.Y(g14279),.A(g12111),.B(g9246));
  NAND2 NAND2_893(.VSS(VSS),.VDD(VDD),.Y(g7887),.A(I12278),.B(I12279));
  NAND2 NAND2_894(.VSS(VSS),.VDD(VDD),.Y(I13749),.A(g4608),.B(g4584));
  NAND2 NAND2_895(.VSS(VSS),.VDD(VDD),.Y(g13886),.A(g11804),.B(g4922));
  NAND2 NAND2_896(.VSS(VSS),.VDD(VDD),.Y(g7228),.A(g6398),.B(g6444));
  NAND2 NAND2_897(.VSS(VSS),.VDD(VDD),.Y(g11994),.A(g8310),.B(g8365));
  NAND2 NAND2_898(.VSS(VSS),.VDD(VDD),.Y(g15723),.A(g10775),.B(g13104));
  NAND3 NAND3_136(.VSS(VSS),.VDD(VDD),.Y(g23978),.A(g572),.B(g21389),.C(g12323));
  NAND4 NAND4_142(.VSS(VSS),.VDD(VDD),.Y(g13967),.A(g3929),.B(g11225),.C(g3983),.D(g11419));
  NAND2 NAND2_899(.VSS(VSS),.VDD(VDD),.Y(I12345),.A(g3106),.B(I12344));
  NAND2 NAND2_900(.VSS(VSS),.VDD(VDD),.Y(I14790),.A(g6167),.B(I14788));
  NAND2 NAND2_901(.VSS(VSS),.VDD(VDD),.Y(I14516),.A(g10147),.B(g661));
  NAND2 NAND2_902(.VSS(VSS),.VDD(VDD),.Y(g23590),.A(g20682),.B(g11111));
  NAND2 NAND2_903(.VSS(VSS),.VDD(VDD),.Y(I12849),.A(g4281),.B(I12848));
  NAND2 NAND2_904(.VSS(VSS),.VDD(VDD),.Y(g12008),.A(g9932),.B(g5798));
  NAND4 NAND4_143(.VSS(VSS),.VDD(VDD),.Y(g17814),.A(g5579),.B(g14522),.C(g5673),.D(g12563));
  NAND2 NAND2_905(.VSS(VSS),.VDD(VDD),.Y(g22638),.A(g18957),.B(g2886));
  NAND2 NAND2_906(.VSS(VSS),.VDD(VDD),.Y(I12848),.A(g4281),.B(g4277));
  NAND2 NAND2_907(.VSS(VSS),.VDD(VDD),.Y(g12476),.A(g7498),.B(g6704));
  NAND3 NAND3_137(.VSS(VSS),.VDD(VDD),.Y(g13459),.A(g7479),.B(g11294),.C(g11846));
  NAND4 NAND4_144(.VSS(VSS),.VDD(VDD),.Y(g21384),.A(g17734),.B(g14686),.C(g17675),.D(g14663));
  NAND2 NAND2_908(.VSS(VSS),.VDD(VDD),.Y(I23587),.A(g4332),.B(I23585));
  NAND2 NAND2_909(.VSS(VSS),.VDD(VDD),.Y(g8889),.A(g3684),.B(g4871));
  NAND2 NAND2_910(.VSS(VSS),.VDD(VDD),.Y(g14038),.A(g11514),.B(g11435));
  NAND2 NAND2_911(.VSS(VSS),.VDD(VDD),.Y(g23067),.A(g20887),.B(g10721));
  NAND2 NAND2_912(.VSS(VSS),.VDD(VDD),.Y(g10601),.A(g896),.B(g7397));
  NAND4 NAND4_145(.VSS(VSS),.VDD(VDD),.Y(g13918),.A(g3259),.B(g11217),.C(g3267),.D(g11350));
  NAND4 NAND4_146(.VSS(VSS),.VDD(VDD),.Y(g16925),.A(g3574),.B(g13799),.C(g3668),.D(g11576));
  NAND2 NAND2_913(.VSS(VSS),.VDD(VDD),.Y(g14601),.A(g12318),.B(g6466));
  NAND2 NAND2_914(.VSS(VSS),.VDD(VDD),.Y(I18538),.A(g14642),.B(I18536));
  NAND2 NAND2_915(.VSS(VSS),.VDD(VDD),.Y(g8871),.A(I12841),.B(I12842));
  NAND2 NAND2_916(.VSS(VSS),.VDD(VDD),.Y(I15079),.A(g9827),.B(I15078));
  NAND2 NAND2_917(.VSS(VSS),.VDD(VDD),.Y(g14677),.A(I16779),.B(I16780));
  NAND2 NAND2_918(.VSS(VSS),.VDD(VDD),.Y(I12263),.A(g1448),.B(I12261));
  NAND2 NAND2_919(.VSS(VSS),.VDD(VDD),.Y(g11545),.A(I14498),.B(I14499));
  NAND3 NAND3_138(.VSS(VSS),.VDD(VDD),.Y(g11444),.A(g6905),.B(g6918),.C(g8733));
  NAND2 NAND2_920(.VSS(VSS),.VDD(VDD),.Y(g13079),.A(g1312),.B(g11336));
  NAND2 NAND2_921(.VSS(VSS),.VDD(VDD),.Y(I15078),.A(g9827),.B(g1968));
  NAND2 NAND2_922(.VSS(VSS),.VDD(VDD),.Y(g12239),.A(I15106),.B(I15107));
  NAND2 NAND2_923(.VSS(VSS),.VDD(VDD),.Y(g20201),.A(I20468),.B(I20469));
  NAND2 NAND2_924(.VSS(VSS),.VDD(VDD),.Y(g8500),.A(g3431),.B(g3423));
  NAND2 NAND2_925(.VSS(VSS),.VDD(VDD),.Y(g14937),.A(g12667),.B(g10421));
  NAND2 NAND2_926(.VSS(VSS),.VDD(VDD),.Y(g26025),.A(g22405),.B(g24631));
  NAND4 NAND4_147(.VSS(VSS),.VDD(VDD),.Y(g13086),.A(g6235),.B(g12101),.C(g6346),.D(g10003));
  NAND2 NAND2_927(.VSS(VSS),.VDD(VDD),.Y(g16681),.A(I17884),.B(I17885));
  NAND4 NAND4_148(.VSS(VSS),.VDD(VDD),.Y(g17578),.A(g5212),.B(g14399),.C(g5283),.D(g12497));
  NAND2 NAND2_928(.VSS(VSS),.VDD(VDD),.Y(g12941),.A(g7167),.B(g10537));
  NAND2 NAND2_929(.VSS(VSS),.VDD(VDD),.Y(g19795),.A(g13600),.B(g16275));
  NAND2 NAND2_930(.VSS(VSS),.VDD(VDD),.Y(g12185),.A(g9905),.B(g799));
  NAND4 NAND4_149(.VSS(VSS),.VDD(VDD),.Y(g21402),.A(g17757),.B(g14740),.C(g17716),.D(g14674));
  NAND2 NAND2_931(.VSS(VSS),.VDD(VDD),.Y(g17586),.A(g14638),.B(g14601));
  NAND2 NAND2_932(.VSS(VSS),.VDD(VDD),.Y(g11977),.A(g8373),.B(g2476));
  NAND2 NAND2_933(.VSS(VSS),.VDD(VDD),.Y(g13977),.A(g11610),.B(g11729));
  NAND2 NAND2_934(.VSS(VSS),.VDD(VDD),.Y(I14530),.A(g8840),.B(g8873));
  NAND2 NAND2_935(.VSS(VSS),.VDD(VDD),.Y(g8737),.A(I12729),.B(I12730));
  NAND2 NAND2_936(.VSS(VSS),.VDD(VDD),.Y(g15011),.A(g12716),.B(g12632));
  NAND2 NAND2_937(.VSS(VSS),.VDD(VDD),.Y(g34227),.A(I32203),.B(I32204));
  NAND2 NAND2_938(.VSS(VSS),.VDD(VDD),.Y(g14015),.A(g11658),.B(g11747));
  NAND2 NAND2_939(.VSS(VSS),.VDD(VDD),.Y(g11561),.A(I14517),.B(I14518));
  NAND2 NAND2_940(.VSS(VSS),.VDD(VDD),.Y(g25172),.A(g5052),.B(g23560));
  NAND2 NAND2_941(.VSS(VSS),.VDD(VDD),.Y(I22872),.A(g12150),.B(I22871));
  NAND2 NAND2_942(.VSS(VSS),.VDD(VDD),.Y(g25996),.A(g24601),.B(g22838));
  NAND4 NAND4_150(.VSS(VSS),.VDD(VDD),.Y(g20170),.A(g16741),.B(g13897),.C(g16687),.D(g13866));
  NAND2 NAND2_943(.VSS(VSS),.VDD(VDD),.Y(g10556),.A(g7971),.B(g8133));
  NAND2 NAND2_944(.VSS(VSS),.VDD(VDD),.Y(g13823),.A(g11313),.B(g3774));
  NAND2 NAND2_945(.VSS(VSS),.VDD(VDD),.Y(I13454),.A(g1959),.B(I13452));
  NAND2 NAND2_946(.VSS(VSS),.VDD(VDD),.Y(I21992),.A(g7670),.B(g19638));
  NAND2 NAND2_947(.VSS(VSS),.VDD(VDD),.Y(g14223),.A(g9092),.B(g11858));
  NAND2 NAND2_948(.VSS(VSS),.VDD(VDD),.Y(g17493),.A(g8659),.B(g14367));
  NAND2 NAND2_949(.VSS(VSS),.VDD(VDD),.Y(g15959),.A(I17405),.B(I17406));
  NAND4 NAND4_151(.VSS(VSS),.VDD(VDD),.Y(g27577),.A(g25019),.B(g25002),.C(g24988),.D(g25765));
  NAND2 NAND2_950(.VSS(VSS),.VDD(VDD),.Y(I15364),.A(g10182),.B(I15363));
  NAND3 NAND3_139(.VSS(VSS),.VDD(VDD),.Y(g12577),.A(g7051),.B(g5990),.C(g6044));
  NAND2 NAND2_951(.VSS(VSS),.VDD(VDD),.Y(g14110),.A(g11692),.B(g8906));
  NAND2 NAND2_952(.VSS(VSS),.VDD(VDD),.Y(g9246),.A(g847),.B(g812));
  NAND4 NAND4_152(.VSS(VSS),.VDD(VDD),.Y(g15742),.A(g5575),.B(g12093),.C(g5637),.D(g14669));
  NAND2 NAND2_953(.VSS(VSS),.VDD(VDD),.Y(I23586),.A(g22409),.B(I23585));
  NAND2 NAND2_954(.VSS(VSS),.VDD(VDD),.Y(g9203),.A(g3706),.B(g3752));
  NAND4 NAND4_153(.VSS(VSS),.VDD(VDD),.Y(g14740),.A(g5913),.B(g12129),.C(g6031),.D(g12614));
  NAND2 NAND2_955(.VSS(VSS),.VDD(VDD),.Y(I13382),.A(g269),.B(g246));
  NAND2 NAND2_956(.VSS(VSS),.VDD(VDD),.Y(I15289),.A(g6697),.B(I15287));
  NAND2 NAND2_957(.VSS(VSS),.VDD(VDD),.Y(g19358),.A(g15723),.B(g1399));
  NAND2 NAND2_958(.VSS(VSS),.VDD(VDD),.Y(I13519),.A(g2514),.B(I13518));
  NAND3 NAND3_140(.VSS(VSS),.VDD(VDD),.Y(g16299),.A(g8160),.B(g8112),.C(g13706));
  NAND3 NAND3_141(.VSS(VSS),.VDD(VDD),.Y(g31003),.A(g27163),.B(g29497),.C(g19644));
  NAND2 NAND2_959(.VSS(VSS),.VDD(VDD),.Y(g14953),.A(g12646),.B(g12405));
  NAND2 NAND2_960(.VSS(VSS),.VDD(VDD),.Y(I15288),.A(g10061),.B(I15287));
  NAND2 NAND2_961(.VSS(VSS),.VDD(VDD),.Y(I13518),.A(g2514),.B(g2518));
  NAND2 NAND2_962(.VSS(VSS),.VDD(VDD),.Y(g12083),.A(g2217),.B(g8205));
  NAND2 NAND2_963(.VSS(VSS),.VDD(VDD),.Y(I15308),.A(g2407),.B(I15306));
  NAND2 NAND2_964(.VSS(VSS),.VDD(VDD),.Y(g11224),.A(I14290),.B(I14291));
  NAND2 NAND2_965(.VSS(VSS),.VDD(VDD),.Y(g13288),.A(g10946),.B(g1442));
  NAND4 NAND4_154(.VSS(VSS),.VDD(VDD),.Y(g15730),.A(g6609),.B(g14556),.C(g6711),.D(g10061));
  NAND2 NAND2_966(.VSS(VSS),.VDD(VDD),.Y(g14800),.A(g7704),.B(g12443));
  NAND2 NAND2_967(.VSS(VSS),.VDD(VDD),.Y(I24414),.A(g23751),.B(g14382));
  NAND2 NAND2_968(.VSS(VSS),.VDD(VDD),.Y(g29046),.A(g27779),.B(g9640));
  NAND3 NAND3_142(.VSS(VSS),.VDD(VDD),.Y(g13495),.A(g1008),.B(g11786),.C(g7972));
  NAND2 NAND2_969(.VSS(VSS),.VDD(VDD),.Y(I29261),.A(g29485),.B(g12046));
  NAND2 NAND2_970(.VSS(VSS),.VDD(VDD),.Y(g24809),.A(g19965),.B(g23132));
  NAND2 NAND2_971(.VSS(VSS),.VDD(VDD),.Y(I22846),.A(g21228),.B(I22844));
  NAND2 NAND2_972(.VSS(VSS),.VDD(VDD),.Y(g24808),.A(I23986),.B(I23987));
  NAND2 NAND2_973(.VSS(VSS),.VDD(VDD),.Y(I13729),.A(g4534),.B(g4537));
  NAND2 NAND2_974(.VSS(VSS),.VDD(VDD),.Y(g10587),.A(g2421),.B(g7456));
  NAND2 NAND2_975(.VSS(VSS),.VDD(VDD),.Y(g11374),.A(g9536),.B(g1536));
  NAND2 NAND2_976(.VSS(VSS),.VDD(VDD),.Y(g28391),.A(g27064),.B(g13637));
  NAND2 NAND2_977(.VSS(VSS),.VDD(VDD),.Y(g12415),.A(g7496),.B(g5976));
  NAND2 NAND2_978(.VSS(VSS),.VDD(VDD),.Y(g21287),.A(g14616),.B(g17571));
  NAND2 NAND2_979(.VSS(VSS),.VDD(VDD),.Y(g19506),.A(g4087),.B(g15825));
  NAND2 NAND2_980(.VSS(VSS),.VDD(VDD),.Y(g10909),.A(g7304),.B(g1116));
  NAND3 NAND3_143(.VSS(VSS),.VDD(VDD),.Y(g20733),.A(g14406),.B(g17290),.C(g9509));
  NAND4 NAND4_155(.VSS(VSS),.VDD(VDD),.Y(g21307),.A(g15719),.B(g13067),.C(g15709),.D(g13040));
  NAND2 NAND2_981(.VSS(VSS),.VDD(VDD),.Y(g15002),.A(g12609),.B(g10312));
  NAND2 NAND2_982(.VSS(VSS),.VDD(VDD),.Y(I25243),.A(g490),.B(I25242));
  NAND2 NAND2_983(.VSS(VSS),.VDD(VDD),.Y(g13260),.A(g1116),.B(g10666));
  NAND2 NAND2_984(.VSS(VSS),.VDD(VDD),.Y(g14908),.A(g7812),.B(g10491));
  NAND2 NAND2_985(.VSS(VSS),.VDD(VDD),.Y(g10569),.A(g2287),.B(g7418));
  NAND2 NAND2_986(.VSS(VSS),.VDD(VDD),.Y(I22929),.A(g12223),.B(g21228));
  NAND2 NAND2_987(.VSS(VSS),.VDD(VDD),.Y(I15195),.A(g6005),.B(I15193));
  NAND2 NAND2_988(.VSS(VSS),.VDD(VDD),.Y(I17405),.A(g13378),.B(I17404));
  NAND2 NAND2_989(.VSS(VSS),.VDD(VDD),.Y(I12344),.A(g3106),.B(g3111));
  NAND4 NAND4_156(.VSS(VSS),.VDD(VDD),.Y(g14569),.A(g3195),.B(g11194),.C(g3329),.D(g8481));
  NAND2 NAND2_990(.VSS(VSS),.VDD(VDD),.Y(g11489),.A(g9661),.B(g3618));
  NAND2 NAND2_991(.VSS(VSS),.VDD(VDD),.Y(g10568),.A(g7328),.B(g7374));
  NAND2 NAND2_992(.VSS(VSS),.VDD(VDD),.Y(g25895),.A(g1259),.B(g24453));
  NAND2 NAND2_993(.VSS(VSS),.VDD(VDD),.Y(g16316),.A(g9429),.B(g13518));
  NAND2 NAND2_994(.VSS(VSS),.VDD(VDD),.Y(g11559),.A(I14509),.B(I14510));
  NAND2 NAND2_995(.VSS(VSS),.VDD(VDD),.Y(g11424),.A(g9662),.B(g4012));
  NAND2 NAND2_996(.VSS(VSS),.VDD(VDD),.Y(I13566),.A(g2652),.B(I13564));
  NAND2 NAND2_997(.VSS(VSS),.VDD(VDD),.Y(g23655),.A(I22793),.B(I22794));
  NAND2 NAND2_998(.VSS(VSS),.VDD(VDD),.Y(I29271),.A(g12050),.B(I29269));
  NAND2 NAND2_999(.VSS(VSS),.VDD(VDD),.Y(g9883),.A(g5782),.B(g5774));
  NAND2 NAND2_1000(.VSS(VSS),.VDD(VDD),.Y(g14123),.A(g10685),.B(g10928));
  NAND4 NAND4_157(.VSS(VSS),.VDD(VDD),.Y(g15737),.A(g13240),.B(g13115),.C(g7903),.D(g13210));
  NAND2 NAND2_1001(.VSS(VSS),.VDD(VDD),.Y(g14807),.A(g7738),.B(g12453));
  NAND3 NAND3_144(.VSS(VSS),.VDD(VDD),.Y(g19903),.A(g13707),.B(g16319),.C(g8227));
  NAND2 NAND2_1002(.VSS(VSS),.VDD(VDD),.Y(g12115),.A(g1926),.B(g8249));
  NAND2 NAND2_1003(.VSS(VSS),.VDD(VDD),.Y(g14974),.A(g12744),.B(g12622));
  NAND4 NAND4_158(.VSS(VSS),.VDD(VDD),.Y(g17790),.A(g6311),.B(g14575),.C(g6322),.D(g10003));
  NAND3 NAND3_145(.VSS(VSS),.VDD(VDD),.Y(g17137),.A(g13727),.B(g13511),.C(g13527));
  NAND2 NAND2_1004(.VSS(VSS),.VDD(VDD),.Y(I13139),.A(g6154),.B(g6159));
  NAND3 NAND3_146(.VSS(VSS),.VDD(VDD),.Y(g11544),.A(g8700),.B(g3990),.C(g4045));
  NAND4 NAND4_159(.VSS(VSS),.VDD(VDD),.Y(g13544),.A(g7972),.B(g10521),.C(g7549),.D(g1008));
  NAND2 NAND2_1005(.VSS(VSS),.VDD(VDD),.Y(g24570),.A(g22957),.B(g2941));
  NAND2 NAND2_1006(.VSS(VSS),.VDD(VDD),.Y(g12052),.A(g7387),.B(g2465));
  NAND2 NAND2_1007(.VSS(VSS),.VDD(VDD),.Y(g14638),.A(g9626),.B(g12361));
  NAND2 NAND2_1008(.VSS(VSS),.VDD(VDD),.Y(I15042),.A(g9752),.B(I15041));
  NAND2 NAND2_1009(.VSS(VSS),.VDD(VDD),.Y(I15255),.A(g1848),.B(I15253));
  NAND2 NAND2_1010(.VSS(VSS),.VDD(VDD),.Y(I13852),.A(g7397),.B(I13850));
  NAND2 NAND2_1011(.VSS(VSS),.VDD(VDD),.Y(g14841),.A(g12593),.B(g12443));
  NAND3 NAND3_147(.VSS(VSS),.VDD(VDD),.Y(g25385),.A(g22369),.B(g1783),.C(g8241));
  NAND2 NAND2_1012(.VSS(VSS),.VDD(VDD),.Y(g24567),.A(g22957),.B(g2917));
  NAND2 NAND2_1013(.VSS(VSS),.VDD(VDD),.Y(g11189),.A(I14248),.B(I14249));
  NAND2 NAND2_1014(.VSS(VSS),.VDD(VDD),.Y(g11679),.A(g8836),.B(g802));
  NAND2 NAND2_1015(.VSS(VSS),.VDD(VDD),.Y(I23600),.A(g22360),.B(g4322));
  NAND3 NAND3_148(.VSS(VSS),.VDD(VDD),.Y(g29778),.A(g294),.B(g28444),.C(g23204));
  NAND4 NAND4_160(.VSS(VSS),.VDD(VDD),.Y(g13124),.A(g10666),.B(g7661),.C(g979),.D(g1061));
  NAND2 NAND2_1016(.VSS(VSS),.VDD(VDD),.Y(g25888),.A(g914),.B(g24439));
  NAND2 NAND2_1017(.VSS(VSS),.VDD(VDD),.Y(g31971),.A(g30573),.B(g10511));
  NAND2 NAND2_1018(.VSS(VSS),.VDD(VDD),.Y(g23210),.A(g18957),.B(g2882));
  NAND4 NAND4_161(.VSS(VSS),.VDD(VDD),.Y(g16696),.A(g13871),.B(g13855),.C(g14682),.D(g12340));
  NAND4 NAND4_162(.VSS(VSS),.VDD(VDD),.Y(g20185),.A(g16772),.B(g13928),.C(g16723),.D(g13882));
  NAND2 NAND2_1019(.VSS(VSS),.VDD(VDD),.Y(g10578),.A(g7174),.B(g6058));
  NAND3 NAND3_149(.VSS(VSS),.VDD(VDD),.Y(g20675),.A(g14377),.B(g17246),.C(g9442));
  NAND2 NAND2_1020(.VSS(VSS),.VDD(VDD),.Y(g20092),.A(g11373),.B(g17794));
  NAND4 NAND4_163(.VSS(VSS),.VDD(VDD),.Y(g14014),.A(g3199),.B(g11217),.C(g3298),.D(g11519));
  NAND2 NAND2_1021(.VSS(VSS),.VDD(VDD),.Y(g11938),.A(g8259),.B(g2208));
  NAND2 NAND2_1022(.VSS(VSS),.VDD(VDD),.Y(g10586),.A(g7380),.B(g7418));
  NAND4 NAND4_164(.VSS(VSS),.VDD(VDD),.Y(g13093),.A(g10649),.B(g7661),.C(g979),.D(g1061));
  NAND2 NAND2_1023(.VSS(VSS),.VDD(VDD),.Y(g8873),.A(I12849),.B(I12850));
  NAND2 NAND2_1024(.VSS(VSS),.VDD(VDD),.Y(g8632),.A(g1514),.B(g1500));
  NAND2 NAND2_1025(.VSS(VSS),.VDD(VDD),.Y(g9538),.A(g1792),.B(g1760));
  NAND2 NAND2_1026(.VSS(VSS),.VDD(VDD),.Y(I20221),.A(g16272),.B(g11170));
  NAND2 NAND2_1027(.VSS(VSS),.VDD(VDD),.Y(I12240),.A(g1111),.B(g1105));
  NAND2 NAND2_1028(.VSS(VSS),.VDD(VDD),.Y(g9509),.A(g5770),.B(g5774));
  NAND2 NAND2_1029(.VSS(VSS),.VDD(VDD),.Y(g23286),.A(g6875),.B(g20887));
  NAND2 NAND2_1030(.VSS(VSS),.VDD(VDD),.Y(g25426),.A(g12371),.B(g22369));
  NAND2 NAND2_1031(.VSS(VSS),.VDD(VDD),.Y(g29672),.A(g28376),.B(g13672));
  NAND2 NAND2_1032(.VSS(VSS),.VDD(VDD),.Y(g17593),.A(I18537),.B(I18538));
  NAND2 NAND2_1033(.VSS(VSS),.VDD(VDD),.Y(g14116),.A(g11697),.B(g11584));
  NAND2 NAND2_1034(.VSS(VSS),.VDD(VDD),.Y(I32185),.A(g33665),.B(g33661));
  NAND2 NAND2_1035(.VSS(VSS),.VDD(VDD),.Y(I14509),.A(g370),.B(I14508));
  NAND2 NAND2_1036(.VSS(VSS),.VDD(VDD),.Y(g10041),.A(I13565),.B(I13566));
  NAND2 NAND2_1037(.VSS(VSS),.VDD(VDD),.Y(g14720),.A(g12593),.B(g10266));
  NAND2 NAND2_1038(.VSS(VSS),.VDD(VDD),.Y(I32518),.A(g34422),.B(I32516));
  NAND3 NAND3_150(.VSS(VSS),.VDD(VDD),.Y(g16259),.A(g4743),.B(g13908),.C(g12054));
  NAND2 NAND2_1039(.VSS(VSS),.VDD(VDD),.Y(I14508),.A(g370),.B(g8721));
  NAND3 NAND3_151(.VSS(VSS),.VDD(VDD),.Y(g16225),.A(g13544),.B(g13528),.C(g13043));
  NAND2 NAND2_1040(.VSS(VSS),.VDD(VDD),.Y(g14041),.A(g11610),.B(g11473));
  NAND2 NAND2_1041(.VSS(VSS),.VDD(VDD),.Y(g21187),.A(g14616),.B(g17364));
  NAND2 NAND2_1042(.VSS(VSS),.VDD(VDD),.Y(I22710),.A(g11915),.B(g21434));
  NAND2 NAND2_1043(.VSS(VSS),.VDD(VDD),.Y(g12207),.A(g9887),.B(g5794));
  NAND2 NAND2_1044(.VSS(VSS),.VDD(VDD),.Y(g23975),.A(I23119),.B(I23120));
  NAND2 NAND2_1045(.VSS(VSS),.VDD(VDD),.Y(g12539),.A(I15341),.B(I15342));
  NAND2 NAND2_1046(.VSS(VSS),.VDD(VDD),.Y(I24463),.A(g14437),.B(I24461));
  NAND4 NAND4_165(.VSS(VSS),.VDD(VDD),.Y(g15753),.A(g6239),.B(g14529),.C(g6351),.D(g10003));
  NAND2 NAND2_1047(.VSS(VSS),.VDD(VDD),.Y(g12538),.A(I15334),.B(I15335));
  NAND2 NAND2_1048(.VSS(VSS),.VDD(VDD),.Y(I12262),.A(g1454),.B(I12261));
  NAND2 NAND2_1049(.VSS(VSS),.VDD(VDD),.Y(I13184),.A(g6505),.B(I13182));
  NAND2 NAND2_1050(.VSS(VSS),.VDD(VDD),.Y(I14213),.A(g9295),.B(I14211));
  NAND4 NAND4_166(.VSS(VSS),.VDD(VDD),.Y(g15736),.A(g6295),.B(g14575),.C(g6373),.D(g10003));
  NAND4 NAND4_167(.VSS(VSS),.VDD(VDD),.Y(g17635),.A(g3542),.B(g13730),.C(g3654),.D(g8542));
  NAND2 NAND2_1051(.VSS(VSS),.VDD(VDD),.Y(g16069),.A(I17447),.B(I17448));
  NAND2 NAND2_1052(.VSS(VSS),.VDD(VDD),.Y(g13915),.A(g11566),.B(g11473));
  NAND2 NAND2_1053(.VSS(VSS),.VDD(VDD),.Y(I22945),.A(g9492),.B(I22944));
  NAND2 NAND2_1054(.VSS(VSS),.VDD(VDD),.Y(g14142),.A(g11715),.B(g8958));
  NAND3 NAND3_152(.VSS(VSS),.VDD(VDD),.Y(g33925),.A(g33394),.B(g4462),.C(g4467));
  NAND4 NAND4_168(.VSS(VSS),.VDD(VDD),.Y(g16657),.A(g3554),.B(g13730),.C(g3625),.D(g11576));
  NAND2 NAND2_1055(.VSS(VSS),.VDD(VDD),.Y(I14205),.A(g8508),.B(I14204));
  NAND3 NAND3_153(.VSS(VSS),.VDD(VDD),.Y(g15843),.A(g7922),.B(g7503),.C(g13264));
  NAND4 NAND4_169(.VSS(VSS),.VDD(VDD),.Y(g14517),.A(g3231),.B(g11217),.C(g3321),.D(g8481));
  NAND2 NAND2_1056(.VSS(VSS),.VDD(VDD),.Y(g24906),.A(g8743),.B(g23088));
  NAND2 NAND2_1057(.VSS(VSS),.VDD(VDD),.Y(g26714),.A(g9316),.B(g25175));
  NAND2 NAND2_1058(.VSS(VSS),.VDD(VDD),.Y(g23666),.A(g20875),.B(g11139));
  NAND2 NAND2_1059(.VSS(VSS),.VDD(VDD),.Y(I26417),.A(g26519),.B(g14247));
  NAND4 NAND4_170(.VSS(VSS),.VDD(VDD),.Y(g21363),.A(g17708),.B(g14664),.C(g17640),.D(g14598));
  NAND2 NAND2_1060(.VSS(VSS),.VDD(VDD),.Y(I32439),.A(g34227),.B(g34220));
  NAND2 NAND2_1061(.VSS(VSS),.VDD(VDD),.Y(g12100),.A(I14956),.B(I14957));
  NAND2 NAND2_1062(.VSS(VSS),.VDD(VDD),.Y(I17380),.A(g13336),.B(I17379));
  NAND2 NAND2_1063(.VSS(VSS),.VDD(VDD),.Y(g24566),.A(g22755),.B(g22713));
  NAND2 NAND2_1064(.VSS(VSS),.VDD(VDD),.Y(g22711),.A(g19581),.B(g7888));
  NAND2 NAND2_1065(.VSS(VSS),.VDD(VDD),.Y(g14130),.A(g11621),.B(g8906));
  NAND2 NAND2_1066(.VSS(VSS),.VDD(VDD),.Y(I18682),.A(g14752),.B(I18680));
  NAND2 NAND2_1067(.VSS(VSS),.VDD(VDD),.Y(g17474),.A(g14547),.B(g14521));
  NAND3 NAND3_154(.VSS(VSS),.VDD(VDD),.Y(g28516),.A(g10857),.B(g26105),.C(g27155));
  NAND2 NAND2_1068(.VSS(VSS),.VDD(VDD),.Y(g11419),.A(I14428),.B(I14429));
  NAND2 NAND2_1069(.VSS(VSS),.VDD(VDD),.Y(g29097),.A(g9700),.B(g27858));
  NAND4 NAND4_171(.VSS(VSS),.VDD(VDD),.Y(g15709),.A(g5224),.B(g14399),.C(g5327),.D(g9780));
  NAND4 NAND4_172(.VSS(VSS),.VDD(VDD),.Y(g27882),.A(g21228),.B(g25307),.C(g26424),.D(g26213));
  NAND3 NAND3_155(.VSS(VSS),.VDD(VDD),.Y(g11155),.A(g4776),.B(g7892),.C(g9030));
  NAND2 NAND2_1070(.VSS(VSS),.VDD(VDD),.Y(I14350),.A(g8890),.B(g8848));
  NAND2 NAND2_1071(.VSS(VSS),.VDD(VDD),.Y(g15708),.A(g7340),.B(g13083));
  NAND3 NAND3_156(.VSS(VSS),.VDD(VDD),.Y(g12414),.A(g7028),.B(g7041),.C(g10165));
  NAND2 NAND2_1072(.VSS(VSS),.VDD(VDD),.Y(g13822),.A(g8160),.B(g11306));
  NAND3 NAND3_157(.VSS(VSS),.VDD(VDD),.Y(g13266),.A(g12440),.B(g9920),.C(g9843));
  NAND2 NAND2_1073(.VSS(VSS),.VDD(VDD),.Y(g25527),.A(g21294),.B(g23462));
  NAND2 NAND2_1074(.VSS(VSS),.VDD(VDD),.Y(I12098),.A(g1322),.B(I12096));
  NAND2 NAND2_1075(.VSS(VSS),.VDD(VDD),.Y(g14727),.A(g12604),.B(g12505));
  NAND2 NAND2_1076(.VSS(VSS),.VDD(VDD),.Y(I12251),.A(g1124),.B(g1129));
  NAND2 NAND2_1077(.VSS(VSS),.VDD(VDD),.Y(I22717),.A(g11916),.B(g21434));
  NAND2 NAND2_1078(.VSS(VSS),.VDD(VDD),.Y(g17492),.A(g8655),.B(g14367));
  NAND2 NAND2_1079(.VSS(VSS),.VDD(VDD),.Y(I17448),.A(g956),.B(I17446));
  NAND2 NAND2_1080(.VSS(VSS),.VDD(VDD),.Y(I15167),.A(g9904),.B(I15166));
  NAND2 NAND2_1081(.VSS(VSS),.VDD(VDD),.Y(I15194),.A(g9935),.B(I15193));
  NAND2 NAND2_1082(.VSS(VSS),.VDD(VDD),.Y(I17404),.A(g13378),.B(g1472));
  NAND2 NAND2_1083(.VSS(VSS),.VDD(VDD),.Y(I31985),.A(g33648),.B(I31983));
  NAND2 NAND2_1084(.VSS(VSS),.VDD(VDD),.Y(g21186),.A(g14616),.B(g17363));
  NAND2 NAND2_1085(.VSS(VSS),.VDD(VDD),.Y(g23685),.A(I22823),.B(I22824));
  NAND2 NAND2_1086(.VSS(VSS),.VDD(VDD),.Y(g7223),.A(I11878),.B(I11879));
  NAND2 NAND2_1087(.VSS(VSS),.VDD(VDD),.Y(g14600),.A(g9564),.B(g12311));
  NAND4 NAND4_173(.VSS(VSS),.VDD(VDD),.Y(g14781),.A(g6259),.B(g12173),.C(g6377),.D(g12672));
  NAND2 NAND2_1088(.VSS(VSS),.VDD(VDD),.Y(g24576),.A(g22957),.B(g2902));
  NAND4 NAND4_174(.VSS(VSS),.VDD(VDD),.Y(g13119),.A(g6625),.B(g12211),.C(g6715),.D(g10061));
  NAND2 NAND2_1089(.VSS(VSS),.VDD(VDD),.Y(g21417),.A(g11677),.B(g17157));
  NAND2 NAND2_1090(.VSS(VSS),.VDD(VDD),.Y(g11118),.A(I14170),.B(I14171));
  NAND2 NAND2_1091(.VSS(VSS),.VDD(VDD),.Y(g12114),.A(g8241),.B(g8146));
  NAND4 NAND4_175(.VSS(VSS),.VDD(VDD),.Y(g13118),.A(g5897),.B(g12067),.C(g6031),.D(g9935));
  NAND2 NAND2_1092(.VSS(VSS),.VDD(VDD),.Y(g21334),.A(g14616),.B(g17596));
  NAND2 NAND2_1093(.VSS(VSS),.VDD(VDD),.Y(g24609),.A(g22850),.B(g22650));
  NAND2 NAND2_1094(.VSS(VSS),.VDD(VDD),.Y(g20200),.A(I20461),.B(I20462));
  NAND2 NAND2_1095(.VSS(VSS),.VDD(VDD),.Y(I29295),.A(g29495),.B(g12117));
  NAND2 NAND2_1096(.VSS(VSS),.VDD(VDD),.Y(g22663),.A(I21977),.B(I21978));
  NAND3 NAND3_158(.VSS(VSS),.VDD(VDD),.Y(g33299),.A(g608),.B(g32296),.C(g12323));
  NAND2 NAND2_1097(.VSS(VSS),.VDD(VDD),.Y(g23762),.A(I22900),.B(I22901));
  NAND2 NAND2_1098(.VSS(VSS),.VDD(VDD),.Y(I15053),.A(g2259),.B(I15051));
  NAND2 NAND2_1099(.VSS(VSS),.VDD(VDD),.Y(I15254),.A(g10078),.B(I15253));
  NAND2 NAND2_1100(.VSS(VSS),.VDD(VDD),.Y(g27141),.A(I25846),.B(I25847));
  NAND2 NAND2_1101(.VSS(VSS),.VDD(VDD),.Y(I25909),.A(g24782),.B(I25907));
  NAND2 NAND2_1102(.VSS(VSS),.VDD(VDD),.Y(g24798),.A(I23962),.B(I23963));
  NAND4 NAND4_176(.VSS(VSS),.VDD(VDD),.Y(g14422),.A(g3187),.B(g11194),.C(g3298),.D(g8481));
  NAND2 NAND2_1103(.VSS(VSS),.VDD(VDD),.Y(g24973),.A(g21272),.B(g23462));
  NAND4 NAND4_177(.VSS(VSS),.VDD(VDD),.Y(g20184),.A(g16770),.B(g13918),.C(g16719),.D(g13896));
  NAND2 NAND2_1104(.VSS(VSS),.VDD(VDD),.Y(g23909),.A(g7028),.B(g20739));
  NAND2 NAND2_1105(.VSS(VSS),.VDD(VDD),.Y(I25908),.A(g26256),.B(I25907));
  NAND2 NAND2_1106(.VSS(VSS),.VDD(VDD),.Y(g22757),.A(g20114),.B(g7891));
  NAND2 NAND2_1107(.VSS(VSS),.VDD(VDD),.Y(g12332),.A(I15167),.B(I15168));
  NAND2 NAND2_1108(.VSS(VSS),.VDD(VDD),.Y(g25019),.A(g20055),.B(g23172));
  NAND2 NAND2_1109(.VSS(VSS),.VDD(VDD),.Y(g25018),.A(g20107),.B(g23154));
  NAND2 NAND2_1110(.VSS(VSS),.VDD(VDD),.Y(I18633),.A(g2504),.B(g14713));
  NAND4 NAND4_178(.VSS(VSS),.VDD(VDD),.Y(g14542),.A(g3582),.B(g11238),.C(g3672),.D(g8542));
  NAND2 NAND2_1111(.VSS(VSS),.VDD(VDD),.Y(g14021),.A(g11697),.B(g8958));
  NAND2 NAND2_1112(.VSS(VSS),.VDD(VDD),.Y(g24934),.A(g21283),.B(g23462));
  NAND2 NAND2_1113(.VSS(VSS),.VDD(VDD),.Y(I25242),.A(g490),.B(g24744));
  NAND4 NAND4_179(.VSS(VSS),.VDD(VDD),.Y(g17757),.A(g5909),.B(g14549),.C(g6005),.D(g12614));
  NAND4 NAND4_180(.VSS(VSS),.VDD(VDD),.Y(g10726),.A(g7304),.B(g7661),.C(g979),.D(g1061));
  NAND2 NAND2_1114(.VSS(VSS),.VDD(VDD),.Y(g23747),.A(I22865),.B(I22866));
  NAND3 NAND3_159(.VSS(VSS),.VDD(VDD),.Y(g10614),.A(g9024),.B(g8977),.C(g8928));
  NAND4 NAND4_181(.VSS(VSS),.VDD(VDD),.Y(g27833),.A(g21228),.B(g25282),.C(g26424),.D(g26190));
  NAND2 NAND2_1115(.VSS(VSS),.VDD(VDD),.Y(g12049),.A(g2208),.B(g8150));
  NAND2 NAND2_1116(.VSS(VSS),.VDD(VDD),.Y(g10905),.A(g1116),.B(g7304));
  NAND2 NAND2_1117(.VSS(VSS),.VDD(VDD),.Y(I15166),.A(g9904),.B(g9823));
  NAND2 NAND2_1118(.VSS(VSS),.VDD(VDD),.Y(g14905),.A(g12785),.B(g7142));
  NAND2 NAND2_1119(.VSS(VSS),.VDD(VDD),.Y(g12048),.A(g7369),.B(g2040));
  NAND4 NAND4_182(.VSS(VSS),.VDD(VDD),.Y(g20214),.A(g16854),.B(g13993),.C(g16776),.D(g13967));
  NAND2 NAND2_1120(.VSS(VSS),.VDD(VDD),.Y(g28109),.A(g27051),.B(g25783));
  NAND2 NAND2_1121(.VSS(VSS),.VDD(VDD),.Y(g12221),.A(I15079),.B(I15080));
  NAND4 NAND4_183(.VSS(VSS),.VDD(VDD),.Y(g27613),.A(g24942),.B(g24933),.C(g25048),.D(g26871));
  NAND2 NAND2_1122(.VSS(VSS),.VDD(VDD),.Y(g11892),.A(g7777),.B(g9086));
  NAND2 NAND2_1123(.VSS(VSS),.VDD(VDD),.Y(g13892),.A(g11653),.B(g11473));
  NAND3 NAND3_160(.VSS(VSS),.VDD(VDD),.Y(g13476),.A(g7503),.B(g11336),.C(g11869));
  NAND4 NAND4_184(.VSS(VSS),.VDD(VDD),.Y(g21416),.A(g17775),.B(g14781),.C(g17744),.D(g14706));
  NAND2 NAND2_1124(.VSS(VSS),.VDD(VDD),.Y(I13141),.A(g6159),.B(I13139));
  NAND2 NAND2_1125(.VSS(VSS),.VDD(VDD),.Y(I14249),.A(g8091),.B(I14247));
  NAND2 NAND2_1126(.VSS(VSS),.VDD(VDD),.Y(I17379),.A(g13336),.B(g1129));
  NAND2 NAND2_1127(.VSS(VSS),.VDD(VDD),.Y(I17925),.A(g1478),.B(I17923));
  NAND2 NAND2_1128(.VSS(VSS),.VDD(VDD),.Y(I23949),.A(g23162),.B(g13603));
  NAND2 NAND2_1129(.VSS(VSS),.VDD(VDD),.Y(g14797),.A(g12593),.B(g12405));
  NAND3 NAND3_161(.VSS(VSS),.VDD(VDD),.Y(g27273),.A(g10504),.B(g26131),.C(g26105));
  NAND2 NAND2_1130(.VSS(VSS),.VDD(VDD),.Y(I14482),.A(g655),.B(I14480));
  NAND4 NAND4_185(.VSS(VSS),.VDD(VDD),.Y(g16687),.A(g3255),.B(g13700),.C(g3325),.D(g11519));
  NAND2 NAND2_1131(.VSS(VSS),.VDD(VDD),.Y(g13712),.A(g8984),.B(g11283));
  NAND4 NAND4_186(.VSS(VSS),.VDD(VDD),.Y(g17634),.A(g3219),.B(g11217),.C(g3281),.D(g13877));
  NAND2 NAND2_1132(.VSS(VSS),.VDD(VDD),.Y(g11914),.A(g8187),.B(g1648));
  NAND4 NAND4_187(.VSS(VSS),.VDD(VDD),.Y(g17872),.A(g6617),.B(g14602),.C(g6711),.D(g12721));
  NAND2 NAND2_1133(.VSS(VSS),.VDD(VDD),.Y(g12947),.A(g7184),.B(g10561));
  NAND2 NAND2_1134(.VSS(VSS),.VDD(VDD),.Y(I14248),.A(g1322),.B(I14247));
  NAND2 NAND2_1135(.VSS(VSS),.VDD(VDD),.Y(I22944),.A(g9492),.B(g19620));
  NAND4 NAND4_188(.VSS(VSS),.VDD(VDD),.Y(g8728),.A(g3618),.B(g3661),.C(g3632),.D(g3654));
  NAND2 NAND2_1136(.VSS(VSS),.VDD(VDD),.Y(I14204),.A(g8508),.B(g3821));
  NAND2 NAND2_1137(.VSS(VSS),.VDD(VDD),.Y(g25300),.A(g22369),.B(g12018));
  NAND3 NAND3_162(.VSS(VSS),.VDD(VDD),.Y(g27463),.A(g287),.B(g26330),.C(g23204));
  NAND4 NAND4_189(.VSS(VSS),.VDD(VDD),.Y(g13907),.A(g3941),.B(g11225),.C(g4023),.D(g11631));
  NAND2 NAND2_1138(.VSS(VSS),.VDD(VDD),.Y(g28381),.A(g27074),.B(g13621));
  NAND2 NAND2_1139(.VSS(VSS),.VDD(VDD),.Y(g29057),.A(g27800),.B(g9649));
  NAND2 NAND2_1140(.VSS(VSS),.VDD(VDD),.Y(g12463),.A(g7513),.B(g6322));
  NAND2 NAND2_1141(.VSS(VSS),.VDD(VDD),.Y(g14136),.A(g11571),.B(g8906));
  NAND2 NAND2_1142(.VSS(VSS),.VDD(VDD),.Y(g14408),.A(g6069),.B(g11924));
  NAND2 NAND2_1143(.VSS(VSS),.VDD(VDD),.Y(g12972),.A(g7209),.B(g10578));
  NAND2 NAND2_1144(.VSS(VSS),.VDD(VDD),.Y(g28174),.A(g1270),.B(g27059));
  NAND3 NAND3_163(.VSS(VSS),.VDD(VDD),.Y(g28796),.A(g27858),.B(g7418),.C(g7335));
  NAND2 NAND2_1145(.VSS(VSS),.VDD(VDD),.Y(g31753),.A(I29314),.B(I29315));
  NAND2 NAND2_1146(.VSS(VSS),.VDD(VDD),.Y(I22793),.A(g11956),.B(I22792));
  NAND3 NAND3_164(.VSS(VSS),.VDD(VDD),.Y(g16260),.A(g4888),.B(g13910),.C(g12088));
  NAND2 NAND2_1147(.VSS(VSS),.VDD(VDD),.Y(g7823),.A(I12218),.B(I12219));
  NAND3 NAND3_165(.VSS(VSS),.VDD(VDD),.Y(g28840),.A(g27858),.B(g7380),.C(g2287));
  NAND3 NAND3_166(.VSS(VSS),.VDD(VDD),.Y(g11382),.A(g8644),.B(g6895),.C(g8663));
  NAND2 NAND2_1148(.VSS(VSS),.VDD(VDD),.Y(I15176),.A(g2661),.B(I15174));
  NAND2 NAND2_1149(.VSS(VSS),.VDD(VDD),.Y(I12203),.A(g1094),.B(g1135));
  NAND3 NAND3_167(.VSS(VSS),.VDD(VDD),.Y(g19632),.A(g1413),.B(g1542),.C(g16047));
  NAND2 NAND2_1150(.VSS(VSS),.VDD(VDD),.Y(I24440),.A(g14411),.B(I24438));
  NAND2 NAND2_1151(.VSS(VSS),.VDD(VDD),.Y(g11675),.A(g8984),.B(g4912));
  NAND4 NAND4_190(.VSS(VSS),.VDD(VDD),.Y(g13176),.A(g10715),.B(g7675),.C(g1322),.D(g1404));
  NAND2 NAND2_1152(.VSS(VSS),.VDD(VDD),.Y(g13092),.A(g1061),.B(g10761));
  NAND2 NAND2_1153(.VSS(VSS),.VDD(VDD),.Y(g26269),.A(I25243),.B(I25244));
  NAND3 NAND3_168(.VSS(VSS),.VDD(VDD),.Y(g34550),.A(g626),.B(g34359),.C(g12323));
  NAND2 NAND2_1154(.VSS(VSS),.VDD(VDD),.Y(g11154),.A(I14212),.B(I14213));
  NAND2 NAND2_1155(.VSS(VSS),.VDD(VDD),.Y(g29737),.A(g28421),.B(g13779));
  NAND3 NAND3_169(.VSS(VSS),.VDD(VDD),.Y(g28522),.A(g10857),.B(g26131),.C(g27142));
  NAND2 NAND2_1156(.VSS(VSS),.VDD(VDD),.Y(g8678),.A(g376),.B(g358));
  NAND2 NAND2_1157(.VSS(VSS),.VDD(VDD),.Y(g17592),.A(I18530),.B(I18531));
  NAND3 NAND3_170(.VSS(VSS),.VDD(VDD),.Y(g16893),.A(g10685),.B(g13252),.C(g703));
  NAND2 NAND2_1158(.VSS(VSS),.VDD(VDD),.Y(g10537),.A(g7138),.B(g5366));
  NAND2 NAND2_1159(.VSS(VSS),.VDD(VDD),.Y(I14331),.A(g225),.B(I14330));
  NAND2 NAND2_1160(.VSS(VSS),.VDD(VDD),.Y(g8105),.A(g3068),.B(g3072));
  NAND2 NAND2_1161(.VSS(VSS),.VDD(VDD),.Y(I31984),.A(g33653),.B(I31983));
  NAND2 NAND2_1162(.VSS(VSS),.VDD(VDD),.Y(g16713),.A(I17924),.B(I17925));
  NAND2 NAND2_1163(.VSS(VSS),.VDD(VDD),.Y(I20462),.A(g14187),.B(I20460));
  NAND2 NAND2_1164(.VSS(VSS),.VDD(VDD),.Y(I29255),.A(g12017),.B(I29253));
  NAND2 NAND2_1165(.VSS(VSS),.VDD(VDD),.Y(I24462),.A(g23796),.B(I24461));
  NAND4 NAND4_191(.VSS(VSS),.VDD(VDD),.Y(g17820),.A(g5925),.B(g14549),.C(g6019),.D(g12614));
  NAND2 NAND2_1166(.VSS(VSS),.VDD(VDD),.Y(g31709),.A(I29285),.B(I29286));
  NAND4 NAND4_192(.VSS(VSS),.VDD(VDD),.Y(g15752),.A(g5921),.B(g12129),.C(g5983),.D(g14701));
  NAND2 NAND2_1167(.VSS(VSS),.VDD(VDD),.Y(I29270),.A(g29486),.B(I29269));
  NAND2 NAND2_1168(.VSS(VSS),.VDD(VDD),.Y(g28949),.A(g27903),.B(g14643));
  NAND2 NAND2_1169(.VSS(VSS),.VDD(VDD),.Y(I13463),.A(g2380),.B(I13462));
  NAND2 NAND2_1170(.VSS(VSS),.VDD(VDD),.Y(g31708),.A(I29278),.B(I29279));
  NAND4 NAND4_193(.VSS(VSS),.VDD(VDD),.Y(g17846),.A(g6271),.B(g14575),.C(g6365),.D(g12672));
  NAND2 NAND2_1171(.VSS(VSS),.VDD(VDD),.Y(g17396),.A(g7345),.B(g14272));
  NAND4 NAND4_194(.VSS(VSS),.VDD(VDD),.Y(g14750),.A(g6633),.B(g12137),.C(g6715),.D(g12721));
  NAND3 NAND3_171(.VSS(VSS),.VDD(VDD),.Y(g24584),.A(g22852),.B(g22836),.C(g22715));
  NAND2 NAND2_1172(.VSS(VSS),.VDD(VDD),.Y(I14212),.A(g9252),.B(I14211));
  NAND2 NAND2_1173(.VSS(VSS),.VDD(VDD),.Y(g7167),.A(g5360),.B(g5406));
  NAND2 NAND2_1174(.VSS(VSS),.VDD(VDD),.Y(g10796),.A(g7537),.B(g7523));
  NAND2 NAND2_1175(.VSS(VSS),.VDD(VDD),.Y(g20107),.A(g11404),.B(g17794));
  NAND2 NAND2_1176(.VSS(VSS),.VDD(VDD),.Y(g11906),.A(I14713),.B(I14714));
  NAND2 NAND2_1177(.VSS(VSS),.VDD(VDD),.Y(I12403),.A(g3813),.B(I12401));
  NAND2 NAND2_1178(.VSS(VSS),.VDD(VDD),.Y(g16093),.A(I17461),.B(I17462));
  NAND3 NAND3_172(.VSS(VSS),.VDD(VDD),.Y(g12344),.A(g10093),.B(g7041),.C(g10130));
  NAND3 NAND3_173(.VSS(VSS),.VDD(VDD),.Y(g13083),.A(g4392),.B(g10590),.C(g4434));
  NAND2 NAND2_1179(.VSS(VSS),.VDD(VDD),.Y(I32441),.A(g34220),.B(I32439));
  NAND2 NAND2_1180(.VSS(VSS),.VDD(VDD),.Y(g13284),.A(g10695),.B(g1157));
  NAND2 NAND2_1181(.VSS(VSS),.VDD(VDD),.Y(g7549),.A(g1018),.B(g1030));
  NAND2 NAND2_1182(.VSS(VSS),.VDD(VDD),.Y(g25341),.A(g22417),.B(g12047));
  NAND2 NAND2_1183(.VSS(VSS),.VDD(VDD),.Y(g29722),.A(g28410),.B(g13742));
  NAND2 NAND2_1184(.VSS(VSS),.VDD(VDD),.Y(g25268),.A(g21124),.B(g23692));
  NAND4 NAND4_195(.VSS(VSS),.VDD(VDD),.Y(g16875),.A(g3223),.B(g13765),.C(g3317),.D(g11519));
  NAND2 NAND2_1185(.VSS(VSS),.VDD(VDD),.Y(g7598),.A(I12075),.B(I12076));
  NAND2 NAND2_1186(.VSS(VSS),.VDD(VDD),.Y(I32758),.A(g25779),.B(I32756));
  NAND4 NAND4_196(.VSS(VSS),.VDD(VDD),.Y(g14663),.A(g5236),.B(g12002),.C(g5290),.D(g12239));
  NAND2 NAND2_1187(.VSS(VSS),.VDD(VDD),.Y(g24804),.A(g19916),.B(g23105));
  NAND3 NAND3_174(.VSS(VSS),.VDD(VDD),.Y(g24652),.A(g22712),.B(g22940),.C(g22757));
  NAND4 NAND4_197(.VSS(VSS),.VDD(VDD),.Y(g13139),.A(g6589),.B(g12137),.C(g6723),.D(g10061));
  NAND4 NAND4_198(.VSS(VSS),.VDD(VDD),.Y(g15713),.A(g5571),.B(g14425),.C(g5673),.D(g9864));
  NAND2 NAND2_1188(.VSS(VSS),.VDD(VDD),.Y(I14369),.A(g8481),.B(I14368));
  NAND2 NAND2_1189(.VSS(VSS),.VDD(VDD),.Y(g34469),.A(I32517),.B(I32518));
  NAND2 NAND2_1190(.VSS(VSS),.VDD(VDD),.Y(I15333),.A(g10152),.B(g2116));
  NAND3 NAND3_175(.VSS(VSS),.VDD(VDD),.Y(g19546),.A(g15969),.B(g10841),.C(g10884));
  NAND2 NAND2_1191(.VSS(VSS),.VDD(VDD),.Y(g8227),.A(g3770),.B(g3774));
  NAND2 NAND2_1192(.VSS(VSS),.VDD(VDD),.Y(I14368),.A(g8481),.B(g3303));
  NAND2 NAND2_1193(.VSS(VSS),.VDD(VDD),.Y(g12028),.A(I14884),.B(I14885));
  NAND2 NAND2_1194(.VSS(VSS),.VDD(VDD),.Y(g15042),.A(g12806),.B(g10491));
  NAND2 NAND2_1195(.VSS(VSS),.VDD(VDD),.Y(g21253),.A(g6423),.B(g17482));
  NAND2 NAND2_1196(.VSS(VSS),.VDD(VDD),.Y(I29277),.A(g29488),.B(g12081));
  NAND2 NAND2_1197(.VSS(VSS),.VDD(VDD),.Y(g23781),.A(I22937),.B(I22938));
  NAND2 NAND2_1198(.VSS(VSS),.VDD(VDD),.Y(g13963),.A(g11715),.B(g11584));
  NAND4 NAND4_199(.VSS(VSS),.VDD(VDD),.Y(g17640),.A(g5264),.B(g14399),.C(g5335),.D(g12497));
  NAND2 NAND2_1199(.VSS(VSS),.VDD(VDD),.Y(I14229),.A(g979),.B(I14228));
  NAND4 NAND4_200(.VSS(VSS),.VDD(VDD),.Y(g21351),.A(g15729),.B(g13098),.C(g15720),.D(g13069));
  NAND2 NAND2_1200(.VSS(VSS),.VDD(VDD),.Y(g26666),.A(g9229),.B(g25144));
  NAND2 NAND2_1201(.VSS(VSS),.VDD(VDD),.Y(I14228),.A(g979),.B(g8055));
  NAND2 NAND2_1202(.VSS(VSS),.VDD(VDD),.Y(g15030),.A(g12716),.B(g12680));
  NAND4 NAND4_201(.VSS(VSS),.VDD(VDD),.Y(g27903),.A(g21228),.B(g25316),.C(g26424),.D(g26218));
  NAND3 NAND3_176(.VSS(VSS),.VDD(VDD),.Y(g13554),.A(g11336),.B(g7582),.C(g1351));
  NAND2 NAND2_1203(.VSS(VSS),.VDD(VDD),.Y(I17924),.A(g13378),.B(I17923));
  NAND3 NAND3_177(.VSS(VSS),.VDD(VDD),.Y(g12491),.A(g7285),.B(g4462),.C(g6961));
  NAND3 NAND3_178(.VSS(VSS),.VDD(VDD),.Y(g28780),.A(g27742),.B(g7308),.C(g1636));
  NAND2 NAND2_1204(.VSS(VSS),.VDD(VDD),.Y(I22753),.A(g11937),.B(g21434));
  NAND2 NAND2_1205(.VSS(VSS),.VDD(VDD),.Y(g11312),.A(g8565),.B(g3794));
  NAND2 NAND2_1206(.VSS(VSS),.VDD(VDD),.Y(g11200),.A(g8592),.B(g3798));
  NAND2 NAND2_1207(.VSS(VSS),.VDD(VDD),.Y(g25038),.A(g21331),.B(g23363));
  NAND3 NAND3_179(.VSS(VSS),.VDD(VDD),.Y(g13115),.A(g1008),.B(g11786),.C(g11294));
  NAND2 NAND2_1208(.VSS(VSS),.VDD(VDD),.Y(I15052),.A(g9759),.B(I15051));
  NAND2 NAND2_1209(.VSS(VSS),.VDD(VDD),.Y(g14933),.A(g12700),.B(g12571));
  NAND2 NAND2_1210(.VSS(VSS),.VDD(VDD),.Y(I14925),.A(g5835),.B(I14923));
  NAND2 NAND2_1211(.VSS(VSS),.VDD(VDD),.Y(g16155),.A(I17495),.B(I17496));
  NAND2 NAND2_1212(.VSS(VSS),.VDD(VDD),.Y(g17662),.A(I18634),.B(I18635));
  NAND3 NAND3_180(.VSS(VSS),.VDD(VDD),.Y(g28820),.A(g27742),.B(g1668),.C(g1592));
  NAND2 NAND2_1213(.VSS(VSS),.VDD(VDD),.Y(I12546),.A(g194),.B(I12544));
  NAND2 NAND2_1214(.VSS(VSS),.VDD(VDD),.Y(I17461),.A(g13378),.B(I17460));
  NAND2 NAND2_1215(.VSS(VSS),.VDD(VDD),.Y(g14851),.A(g7738),.B(g12505));
  NAND2 NAND2_1216(.VSS(VSS),.VDD(VDD),.Y(g27767),.A(I26367),.B(I26368));
  NAND2 NAND2_1217(.VSS(VSS),.VDD(VDD),.Y(g9775),.A(g4831),.B(g4681));
  NAND4 NAND4_202(.VSS(VSS),.VDD(VDD),.Y(g20371),.A(g16956),.B(g14088),.C(g16694),.D(g16660));
  NAND2 NAND2_1218(.VSS(VSS),.VDD(VDD),.Y(g24951),.A(g199),.B(g23088));
  NAND2 NAND2_1219(.VSS(VSS),.VDD(VDD),.Y(g24972),.A(g19962),.B(g23172));
  NAND2 NAND2_1220(.VSS(VSS),.VDD(VDD),.Y(g12767),.A(g4467),.B(g6961));
  NAND2 NAND2_1221(.VSS(VSS),.VDD(VDD),.Y(g13798),.A(g11280),.B(g3423));
  NAND2 NAND2_1222(.VSS(VSS),.VDD(VDD),.Y(g11973),.A(g8365),.B(g2051));
  NAND2 NAND2_1223(.VSS(VSS),.VDD(VDD),.Y(g30580),.A(g29335),.B(g19666));
  NAND2 NAND2_1224(.VSS(VSS),.VDD(VDD),.Y(g29657),.A(g28363),.B(g13634));
  NAND4 NAND4_203(.VSS(VSS),.VDD(VDD),.Y(g17779),.A(g6637),.B(g14556),.C(g6704),.D(g12471));
  NAND2 NAND2_1225(.VSS(VSS),.VDD(VDD),.Y(g11674),.A(g8676),.B(g4674));
  NAND2 NAND2_1226(.VSS(VSS),.VDD(VDD),.Y(g7879),.A(I12262),.B(I12263));
  NAND2 NAND2_1227(.VSS(VSS),.VDD(VDD),.Y(g23726),.A(g9559),.B(g21140));
  NAND2 NAND2_1228(.VSS(VSS),.VDD(VDD),.Y(I20203),.A(g16246),.B(g11147));
  NAND2 NAND2_1229(.VSS(VSS),.VDD(VDD),.Y(g16524),.A(g13822),.B(g13798));
  NAND2 NAND2_1230(.VSS(VSS),.VDD(VDD),.Y(g26685),.A(g9264),.B(g25160));
  NAND2 NAND2_1231(.VSS(VSS),.VDD(VDD),.Y(I14429),.A(g4005),.B(I14427));
  NAND2 NAND2_1232(.VSS(VSS),.VDD(VDD),.Y(g14574),.A(g12256),.B(g6120));
  NAND2 NAND2_1233(.VSS(VSS),.VDD(VDD),.Y(g12191),.A(I15052),.B(I15053));
  NAND4 NAND4_204(.VSS(VSS),.VDD(VDD),.Y(g14452),.A(g3538),.B(g11207),.C(g3649),.D(g8542));
  NAND2 NAND2_1234(.VSS(VSS),.VDD(VDD),.Y(g11934),.A(g8139),.B(g8187));
  NAND2 NAND2_1235(.VSS(VSS),.VDD(VDD),.Y(g16119),.A(I17475),.B(I17476));
  NAND2 NAND2_1236(.VSS(VSS),.VDD(VDD),.Y(I14428),.A(g8595),.B(I14427));
  NAND2 NAND2_1237(.VSS(VSS),.VDD(VDD),.Y(g12521),.A(g7471),.B(g5969));
  NAND4 NAND4_205(.VSS(VSS),.VDD(VDD),.Y(g17647),.A(g5905),.B(g14497),.C(g5976),.D(g12614));
  NAND2 NAND2_1238(.VSS(VSS),.VDD(VDD),.Y(I29313),.A(g29501),.B(g12154));
  NAND2 NAND2_1239(.VSS(VSS),.VDD(VDD),.Y(g8609),.A(g1171),.B(g1157));
  NAND2 NAND2_1240(.VSS(VSS),.VDD(VDD),.Y(g19450),.A(g11471),.B(g17794));
  NAND2 NAND2_1241(.VSS(VSS),.VDD(VDD),.Y(I14765),.A(g9808),.B(I14764));
  NAND2 NAND2_1242(.VSS(VSS),.VDD(VDD),.Y(g11761),.A(I14610),.B(I14611));
  NAND2 NAND2_1243(.VSS(VSS),.VDD(VDD),.Y(g22651),.A(g20114),.B(g2873));
  NAND2 NAND2_1244(.VSS(VSS),.VDD(VDD),.Y(I29285),.A(g29489),.B(I29284));
  NAND2 NAND2_1245(.VSS(VSS),.VDD(VDD),.Y(g14051),.A(g10323),.B(g11527));
  NAND2 NAND2_1246(.VSS(VSS),.VDD(VDD),.Y(g14072),.A(g11571),.B(g11483));
  NAND4 NAND4_206(.VSS(VSS),.VDD(VDD),.Y(g16749),.A(g3957),.B(g13772),.C(g4027),.D(g11631));
  NAND2 NAND2_1247(.VSS(VSS),.VDD(VDD),.Y(g20163),.A(g16663),.B(g13938));
  NAND4 NAND4_207(.VSS(VSS),.VDD(VDD),.Y(g15782),.A(g6585),.B(g14556),.C(g6697),.D(g10061));
  NAND2 NAND2_1248(.VSS(VSS),.VDD(VDD),.Y(I29254),.A(g29482),.B(I29253));
  NAND2 NAND2_1249(.VSS(VSS),.VDD(VDD),.Y(I15214),.A(g1714),.B(I15212));
  NAND4 NAND4_208(.VSS(VSS),.VDD(VDD),.Y(g14780),.A(g6275),.B(g12101),.C(g6329),.D(g12423));
  NAND2 NAND2_1250(.VSS(VSS),.VDD(VDD),.Y(g12045),.A(g1783),.B(g8146));
  NAND3 NAND3_181(.VSS(VSS),.VDD(VDD),.Y(g10820),.A(g9985),.B(g9920),.C(g9843));
  NAND4 NAND4_209(.VSS(VSS),.VDD(VDD),.Y(g14820),.A(g6307),.B(g12173),.C(g6315),.D(g12423));
  NAND4 NAND4_210(.VSS(VSS),.VDD(VDD),.Y(g17513),.A(g3247),.B(g13765),.C(g3325),.D(g8481));
  NAND3 NAND3_182(.VSS(VSS),.VDD(VDD),.Y(g28827),.A(g27837),.B(g7362),.C(g1862));
  NAND2 NAND2_1251(.VSS(VSS),.VDD(VDD),.Y(g25531),.A(g22763),.B(g2868));
  NAND3 NAND3_183(.VSS(VSS),.VDD(VDD),.Y(g15853),.A(g14714),.B(g9417),.C(g12337));
  NAND2 NAND2_1252(.VSS(VSS),.VDD(VDD),.Y(I15241),.A(g10003),.B(g6351));
  NAND3 NAND3_184(.VSS(VSS),.VDD(VDD),.Y(g12462),.A(g7051),.B(g7064),.C(g10190));
  NAND2 NAND2_1253(.VSS(VSS),.VDD(VDD),.Y(g13241),.A(g7503),.B(g10544));
  NAND2 NAND2_1254(.VSS(VSS),.VDD(VDD),.Y(g25186),.A(g5396),.B(g23602));
  NAND2 NAND2_1255(.VSS(VSS),.VDD(VDD),.Y(g14691),.A(g12695),.B(g12505));
  NAND3 NAND3_185(.VSS(VSS),.VDD(VDD),.Y(g25953),.A(g22756),.B(g24570),.C(g22688));
  NAND2 NAND2_1256(.VSS(VSS),.VDD(VDD),.Y(g8803),.A(g128),.B(g4646));
  NAND2 NAND2_1257(.VSS(VSS),.VDD(VDD),.Y(g9954),.A(g6128),.B(g6120));
  NAND2 NAND2_1258(.VSS(VSS),.VDD(VDD),.Y(I22792),.A(g11956),.B(g21434));
  NAND2 NAND2_1259(.VSS(VSS),.VDD(VDD),.Y(I22967),.A(g21228),.B(I22965));
  NAND4 NAND4_211(.VSS(VSS),.VDD(VDD),.Y(g13100),.A(g6581),.B(g12137),.C(g6692),.D(g10061));
  NAND2 NAND2_1260(.VSS(VSS),.VDD(VDD),.Y(g23575),.A(I22711),.B(I22712));
  NAND2 NAND2_1261(.VSS(VSS),.VDD(VDD),.Y(g20173),.A(g16696),.B(g13972));
  NAND2 NAND2_1262(.VSS(VSS),.VDD(VDD),.Y(g10929),.A(g1099),.B(g7854));
  NAND2 NAND2_1263(.VSS(VSS),.VDD(VDD),.Y(g31669),.A(I29254),.B(I29255));
  NAND3 NAND3_186(.VSS(VSS),.VDD(VDD),.Y(g15864),.A(g14833),.B(g12543),.C(g12487));
  NAND2 NAND2_1264(.VSS(VSS),.VDD(VDD),.Y(g33669),.A(g33378),.B(g862));
  NAND2 NAND2_1265(.VSS(VSS),.VDD(VDD),.Y(g25334),.A(g21253),.B(g23756));
  NAND4 NAND4_212(.VSS(VSS),.VDD(VDD),.Y(g17723),.A(g6597),.B(g14556),.C(g6668),.D(g12721));
  NAND2 NAND2_1266(.VSS(VSS),.VDD(VDD),.Y(g10583),.A(g7475),.B(g862));
  NAND3 NAND3_187(.VSS(VSS),.VDD(VDD),.Y(g10928),.A(g8181),.B(g8137),.C(g417));
  NAND4 NAND4_213(.VSS(VSS),.VDD(VDD),.Y(g15748),.A(g13257),.B(g13130),.C(g7922),.D(g13241));
  NAND2 NAND2_1267(.VSS(VSS),.VDD(VDD),.Y(g21283),.A(g11291),.B(g17157));
  NAND2 NAND2_1268(.VSS(VSS),.VDD(VDD),.Y(g9912),.A(I13463),.B(I13464));
  NAND2 NAND2_1269(.VSS(VSS),.VDD(VDD),.Y(I13045),.A(g5120),.B(I13043));
  NAND4 NAND4_214(.VSS(VSS),.VDD(VDD),.Y(g20134),.A(g17572),.B(g14542),.C(g17495),.D(g14452));
  NAND4 NAND4_215(.VSS(VSS),.VDD(VDD),.Y(g13515),.A(g12628),.B(g12588),.C(g12524),.D(g12464));
  NAND4 NAND4_216(.VSS(VSS),.VDD(VDD),.Y(g13882),.A(g3590),.B(g11207),.C(g3672),.D(g11576));
  NAND2 NAND2_1270(.VSS(VSS),.VDD(VDD),.Y(g24760),.A(I23918),.B(I23919));
  NAND2 NAND2_1271(.VSS(VSS),.VDD(VDD),.Y(I23961),.A(g23184),.B(g13631));
  NAND2 NAND2_1272(.VSS(VSS),.VDD(VDD),.Y(g25216),.A(g6088),.B(g23678));
  NAND2 NAND2_1273(.VSS(VSS),.VDD(VDD),.Y(g14113),.A(g11626),.B(g11537));
  NAND2 NAND2_1274(.VSS(VSS),.VDD(VDD),.Y(I24385),.A(g14347),.B(I24383));
  NAND2 NAND2_1275(.VSS(VSS),.VDD(VDD),.Y(g15036),.A(g12780),.B(g12581));
  NAND2 NAND2_1276(.VSS(VSS),.VDD(VDD),.Y(g19597),.A(g1199),.B(g15995));
  NAND2 NAND2_1277(.VSS(VSS),.VDD(VDD),.Y(g12629),.A(g7812),.B(g7142));
  NAND2 NAND2_1278(.VSS(VSS),.VDD(VDD),.Y(I12877),.A(g4200),.B(I12876));
  NAND2 NAND2_1279(.VSS(VSS),.VDD(VDD),.Y(I13462),.A(g2380),.B(g2384));
  NAND2 NAND2_1280(.VSS(VSS),.VDD(VDD),.Y(g8847),.A(g4831),.B(g4681));
  NAND3 NAND3_188(.VSS(VSS),.VDD(VDD),.Y(g12628),.A(g7074),.B(g6336),.C(g6390));
  NAND3 NAND3_189(.VSS(VSS),.VDD(VDD),.Y(g22850),.A(g1536),.B(g19581),.C(g10699));
  NAND2 NAND2_1281(.VSS(VSS),.VDD(VDD),.Y(g11441),.A(g9599),.B(g3267));
  NAND2 NAND2_1282(.VSS(VSS),.VDD(VDD),.Y(I13140),.A(g6154),.B(I13139));
  NAND2 NAND2_1283(.VSS(VSS),.VDD(VDD),.Y(I22901),.A(g21228),.B(I22899));
  NAND3 NAND3_190(.VSS(VSS),.VDD(VDD),.Y(g28786),.A(g27837),.B(g7405),.C(g7322));
  NAND2 NAND2_1284(.VSS(VSS),.VDD(VDD),.Y(g11206),.A(I14276),.B(I14277));
  NAND3 NAND3_191(.VSS(VSS),.VDD(VDD),.Y(g16238),.A(g4698),.B(g13883),.C(g12054));
  NAND2 NAND2_1285(.VSS(VSS),.VDD(VDD),.Y(I14499),.A(g8737),.B(I14497));
  NAND2 NAND2_1286(.VSS(VSS),.VDD(VDD),.Y(g17412),.A(g14520),.B(g14489));
  NAND2 NAND2_1287(.VSS(VSS),.VDD(VDD),.Y(I18625),.A(g2079),.B(g14712));
  NAND2 NAND2_1288(.VSS(VSS),.VDD(VDD),.Y(g14768),.A(g12662),.B(g12571));
  NAND2 NAND2_1289(.VSS(VSS),.VDD(VDD),.Y(g28945),.A(g27854),.B(g8211));
  NAND4 NAND4_217(.VSS(VSS),.VDD(VDD),.Y(g14803),.A(g5208),.B(g12059),.C(g5308),.D(g12497));
  NAND2 NAND2_1290(.VSS(VSS),.VDD(VDD),.Y(I14498),.A(g9020),.B(I14497));
  NAND3 NAND3_192(.VSS(VSS),.VDD(VDD),.Y(g33679),.A(g33394),.B(g10737),.C(g10308));
  NAND2 NAND2_1291(.VSS(VSS),.VDD(VDD),.Y(g12147),.A(g8302),.B(g8201));
  NAND2 NAND2_1292(.VSS(VSS),.VDD(VDD),.Y(I12402),.A(g3808),.B(I12401));
  NAND2 NAND2_1293(.VSS(VSS),.VDD(VDD),.Y(I15107),.A(g5313),.B(I15105));
  NAND2 NAND2_1294(.VSS(VSS),.VDD(VDD),.Y(I22823),.A(g11978),.B(I22822));
  NAND2 NAND2_1295(.VSS(VSS),.VDD(VDD),.Y(I14611),.A(g8678),.B(I14609));
  NAND2 NAND2_1296(.VSS(VSS),.VDD(VDD),.Y(I14924),.A(g9558),.B(I14923));
  NAND2 NAND2_1297(.VSS(VSS),.VDD(VDD),.Y(g12370),.A(I15213),.B(I15214));
  NAND2 NAND2_1298(.VSS(VSS),.VDD(VDD),.Y(g25974),.A(g24576),.B(g22837));
  NAND4 NAND4_218(.VSS(VSS),.VDD(VDD),.Y(g17716),.A(g5957),.B(g14497),.C(g6027),.D(g12614));
  NAND2 NAND2_1299(.VSS(VSS),.VDD(VDD),.Y(g15008),.A(g12780),.B(g10341));
  NAND2 NAND2_1300(.VSS(VSS),.VDD(VDD),.Y(I23971),.A(g490),.B(I23969));
  NAND2 NAND2_1301(.VSS(VSS),.VDD(VDD),.Y(g25293),.A(g21190),.B(g23726));
  NAND2 NAND2_1302(.VSS(VSS),.VDD(VDD),.Y(g12151),.A(g8316),.B(g8211));
  NAND2 NAND2_1303(.VSS(VSS),.VDD(VDD),.Y(g19854),.A(I20222),.B(I20223));
  NAND4 NAND4_219(.VSS(VSS),.VDD(VDD),.Y(g13940),.A(g11426),.B(g8889),.C(g11707),.D(g8829));
  NAND2 NAND2_1304(.VSS(VSS),.VDD(VDD),.Y(I22966),.A(g12288),.B(I22965));
  NAND2 NAND2_1305(.VSS(VSS),.VDD(VDD),.Y(g23949),.A(g7074),.B(g21012));
  NAND2 NAND2_1306(.VSS(VSS),.VDD(VDD),.Y(g28448),.A(g23975),.B(g27377));
  NAND2 NAND2_1307(.VSS(VSS),.VDD(VDD),.Y(I15263),.A(g10081),.B(I15262));
  NAND2 NAND2_1308(.VSS(VSS),.VDD(VDD),.Y(g10552),.A(g2153),.B(g7374));
  NAND4 NAND4_220(.VSS(VSS),.VDD(VDD),.Y(g8751),.A(g3969),.B(g4012),.C(g3983),.D(g4005));
  NAND3 NAND3_193(.VSS(VSS),.VDD(VDD),.Y(g15907),.A(g14833),.B(g9417),.C(g12487));
  NAND2 NAND2_1309(.VSS(VSS),.VDD(VDD),.Y(g22681),.A(I21993),.B(I21994));
  NAND2 NAND2_1310(.VSS(VSS),.VDD(VDD),.Y(g11135),.A(I14186),.B(I14187));
  NAND2 NAND2_1311(.VSS(VSS),.VDD(VDD),.Y(I14330),.A(g225),.B(g9966));
  NAND2 NAND2_1312(.VSS(VSS),.VDD(VDD),.Y(g19916),.A(g3029),.B(g16313));
  NAND4 NAND4_221(.VSS(VSS),.VDD(VDD),.Y(g16728),.A(g13884),.B(g13870),.C(g14089),.D(g11639));
  NAND2 NAND2_1313(.VSS(VSS),.VDD(VDD),.Y(g12227),.A(g8418),.B(g8330));
  NAND2 NAND2_1314(.VSS(VSS),.VDD(VDD),.Y(I14764),.A(g9808),.B(g5821));
  NAND2 NAND2_1315(.VSS(VSS),.VDD(VDD),.Y(g11962),.A(I14789),.B(I14790));
  NAND2 NAND2_1316(.VSS(VSS),.VDD(VDD),.Y(I29284),.A(g29489),.B(g12085));
  NAND2 NAND2_1317(.VSS(VSS),.VDD(VDD),.Y(I31973),.A(g33641),.B(I31972));
  NAND2 NAND2_1318(.VSS(VSS),.VDD(VDD),.Y(I29304),.A(g12121),.B(I29302));
  NAND2 NAND2_1319(.VSS(VSS),.VDD(VDD),.Y(I18581),.A(g14678),.B(I18579));
  NAND2 NAND2_1320(.VSS(VSS),.VDD(VDD),.Y(I26051),.A(g13500),.B(I26049));
  NAND2 NAND2_1321(.VSS(VSS),.VDD(VDD),.Y(I25847),.A(g24799),.B(I25845));
  NAND2 NAND2_1322(.VSS(VSS),.VDD(VDD),.Y(I26072),.A(g13517),.B(I26070));
  NAND2 NAND2_1323(.VSS(VSS),.VDD(VDD),.Y(I11825),.A(g4593),.B(I11824));
  NAND2 NAND2_1324(.VSS(VSS),.VDD(VDD),.Y(I12876),.A(g4200),.B(g4180));
  NAND2 NAND2_1325(.VSS(VSS),.VDD(VDD),.Y(g14999),.A(g12739),.B(g12824));
  NAND3 NAND3_194(.VSS(VSS),.VDD(VDD),.Y(g16304),.A(g4765),.B(g13970),.C(g12054));
  NAND2 NAND2_1326(.VSS(VSS),.VDD(VDD),.Y(g12044),.A(g1657),.B(g8139));
  NAND2 NAND2_1327(.VSS(VSS),.VDD(VDD),.Y(I15004),.A(g1700),.B(I15002));
  NAND4 NAND4_222(.VSS(VSS),.VDD(VDD),.Y(g21509),.A(g17820),.B(g14898),.C(g17647),.D(g17608));
  NAND4 NAND4_223(.VSS(VSS),.VDD(VDD),.Y(g17765),.A(g6649),.B(g14556),.C(g6719),.D(g12721));
  NAND2 NAND2_1328(.VSS(VSS),.VDD(VDD),.Y(I14259),.A(g3133),.B(I14257));
  NAND2 NAND2_1329(.VSS(VSS),.VDD(VDD),.Y(I17495),.A(g13378),.B(I17494));
  NAND2 NAND2_1330(.VSS(VSS),.VDD(VDD),.Y(g27377),.A(g10685),.B(g25930));
  NAND4 NAND4_224(.VSS(VSS),.VDD(VDD),.Y(g24926),.A(g20172),.B(g20163),.C(g23357),.D(g13995));
  NAND2 NAND2_1331(.VSS(VSS),.VDD(VDD),.Y(g25275),.A(g22342),.B(g11991));
  NAND2 NAND2_1332(.VSS(VSS),.VDD(VDD),.Y(g12301),.A(I15148),.B(I15149));
  NAND2 NAND2_1333(.VSS(VSS),.VDD(VDD),.Y(I14258),.A(g8154),.B(I14257));
  NAND2 NAND2_1334(.VSS(VSS),.VDD(VDD),.Y(g12120),.A(g2476),.B(g8273));
  NAND4 NAND4_225(.VSS(VSS),.VDD(VDD),.Y(g27738),.A(g21228),.B(g25243),.C(g26424),.D(g26148));
  NAND2 NAND2_1335(.VSS(VSS),.VDD(VDD),.Y(I32440),.A(g34227),.B(I32439));
  NAND2 NAND2_1336(.VSS(VSS),.VDD(VDD),.Y(g25237),.A(g6434),.B(g23711));
  NAND2 NAND2_1337(.VSS(VSS),.VDD(VDD),.Y(I15106),.A(g9780),.B(I15105));
  NAND2 NAND2_1338(.VSS(VSS),.VDD(VDD),.Y(g13273),.A(g1459),.B(g10699));
  NAND2 NAND2_1339(.VSS(VSS),.VDD(VDD),.Y(g19335),.A(g15717),.B(g1056));
  NAND2 NAND2_1340(.VSS(VSS),.VDD(VDD),.Y(g10961),.A(g1442),.B(g7876));
  NAND3 NAND3_195(.VSS(VSS),.VDD(VDD),.Y(g29679),.A(g153),.B(g28353),.C(g23042));
  NAND4 NAND4_226(.VSS(VSS),.VDD(VDD),.Y(g15729),.A(g5949),.B(g14549),.C(g6027),.D(g9935));
  NAND2 NAND2_1341(.VSS(VSS),.VDD(VDD),.Y(g14505),.A(g12073),.B(g9961));
  NAND2 NAND2_1342(.VSS(VSS),.VDD(VDD),.Y(I12287),.A(g1484),.B(g1300));
  NAND2 NAND2_1343(.VSS(VSS),.VDD(VDD),.Y(I14955),.A(g9620),.B(g6181));
  NAND2 NAND2_1344(.VSS(VSS),.VDD(VDD),.Y(g19965),.A(g3380),.B(g16424));
  NAND3 NAND3_196(.VSS(VSS),.VDD(VDD),.Y(g11951),.A(g9166),.B(g847),.C(g703));
  NAND4 NAND4_227(.VSS(VSS),.VDD(VDD),.Y(g15728),.A(g5200),.B(g14399),.C(g5313),.D(g9780));
  NAND2 NAND2_1345(.VSS(VSS),.VDD(VDD),.Y(g13951),.A(g10295),.B(g11729));
  NAND2 NAND2_1346(.VSS(VSS),.VDD(VDD),.Y(I12076),.A(g979),.B(I12074));
  NAND2 NAND2_1347(.VSS(VSS),.VDD(VDD),.Y(g23047),.A(g482),.B(g20000));
  NAND2 NAND2_1348(.VSS(VSS),.VDD(VDD),.Y(g13795),.A(g11216),.B(g401));
  NAND3 NAND3_197(.VSS(VSS),.VDD(VDD),.Y(g28896),.A(g27837),.B(g1936),.C(g1862));
  NAND2 NAND2_1349(.VSS(VSS),.VDD(VDD),.Y(I14171),.A(g3119),.B(I14169));
  NAND2 NAND2_1350(.VSS(VSS),.VDD(VDD),.Y(g20871),.A(g14434),.B(g17396));
  NAND2 NAND2_1351(.VSS(VSS),.VDD(VDD),.Y(I22893),.A(g12189),.B(I22892));
  NAND2 NAND2_1352(.VSS(VSS),.VDD(VDD),.Y(I12269),.A(g1141),.B(g956));
  NAND2 NAND2_1353(.VSS(VSS),.VDD(VDD),.Y(I13044),.A(g5115),.B(I13043));
  NAND4 NAND4_228(.VSS(VSS),.VDD(VDD),.Y(g17775),.A(g6255),.B(g14575),.C(g6351),.D(g12672));
  NAND2 NAND2_1354(.VSS(VSS),.VDD(VDD),.Y(I22865),.A(g12146),.B(I22864));
  NAND2 NAND2_1355(.VSS(VSS),.VDD(VDD),.Y(g23756),.A(g9621),.B(g21206));
  NAND2 NAND2_1356(.VSS(VSS),.VDD(VDD),.Y(g14723),.A(g7704),.B(g12772));
  NAND2 NAND2_1357(.VSS(VSS),.VDD(VDD),.Y(g23780),.A(I22930),.B(I22931));
  NAND2 NAND2_1358(.VSS(VSS),.VDD(VDD),.Y(g14433),.A(g12035),.B(g9890));
  NAND2 NAND2_1359(.VSS(VSS),.VDD(VDD),.Y(I24384),.A(g23721),.B(I24383));
  NAND4 NAND4_229(.VSS(VSS),.VDD(VDD),.Y(g21350),.A(g15751),.B(g15742),.C(g15735),.D(g13108));
  NAND2 NAND2_1360(.VSS(VSS),.VDD(VDD),.Y(g16312),.A(g13580),.B(g13574));
  NAND2 NAND2_1361(.VSS(VSS),.VDD(VDD),.Y(g14104),.A(g11514),.B(g8864));
  NAND2 NAND2_1362(.VSS(VSS),.VDD(VDD),.Y(I25846),.A(g26212),.B(I25845));
  NAND2 NAND2_1363(.VSS(VSS),.VDD(VDD),.Y(g14343),.A(g11961),.B(g9670));
  NAND2 NAND2_1364(.VSS(VSS),.VDD(VDD),.Y(g10971),.A(g7867),.B(g7886));
  NAND2 NAND2_1365(.VSS(VSS),.VDD(VDD),.Y(g28958),.A(g27833),.B(g8249));
  NAND2 NAND2_1366(.VSS(VSS),.VDD(VDD),.Y(g14971),.A(g12667),.B(g12581));
  NAND4 NAND4_230(.VSS(VSS),.VDD(VDD),.Y(g16745),.A(g3594),.B(g13730),.C(g3661),.D(g11389));
  NAND2 NAND2_1367(.VSS(VSS),.VDD(VDD),.Y(g31748),.A(I29303),.B(I29304));
  NAND2 NAND2_1368(.VSS(VSS),.VDD(VDD),.Y(g26208),.A(g7975),.B(g24751));
  NAND4 NAND4_231(.VSS(VSS),.VDD(VDD),.Y(g16813),.A(g3614),.B(g13799),.C(g3625),.D(g8542));
  NAND2 NAND2_1369(.VSS(VSS),.VDD(VDD),.Y(I22938),.A(g21228),.B(I22936));
  NAND2 NAND2_1370(.VSS(VSS),.VDD(VDD),.Y(g27824),.A(I26394),.B(I26395));
  NAND2 NAND2_1371(.VSS(VSS),.VDD(VDD),.Y(g13920),.A(g11621),.B(g11483));
  NAND2 NAND2_1372(.VSS(VSS),.VDD(VDD),.Y(I17460),.A(g13378),.B(g1300));
  NAND2 NAND2_1373(.VSS(VSS),.VDD(VDD),.Y(g24591),.A(g22833),.B(g22642));
  NAND2 NAND2_1374(.VSS(VSS),.VDD(VDD),.Y(g24776),.A(g3040),.B(g23052));
  NAND2 NAND2_1375(.VSS(VSS),.VDD(VDD),.Y(I14817),.A(g9962),.B(I14816));
  NAND2 NAND2_1376(.VSS(VSS),.VDD(VDD),.Y(g25236),.A(I24415),.B(I24416));
  NAND2 NAND2_1377(.VSS(VSS),.VDD(VDD),.Y(I15121),.A(g9910),.B(g2102));
  NAND2 NAND2_1378(.VSS(VSS),.VDD(VDD),.Y(g34422),.A(I32432),.B(I32433));
  NAND3 NAND3_198(.VSS(VSS),.VDD(VDD),.Y(g28857),.A(g27779),.B(g1802),.C(g1728));
  NAND2 NAND2_1379(.VSS(VSS),.VDD(VDD),.Y(g14133),.A(g11692),.B(g11747));
  NAND2 NAND2_1380(.VSS(VSS),.VDD(VDD),.Y(I12279),.A(g1472),.B(I12277));
  NAND2 NAND2_1381(.VSS(VSS),.VDD(VDD),.Y(I14532),.A(g8873),.B(I14530));
  NAND2 NAND2_1382(.VSS(VSS),.VDD(VDD),.Y(g13121),.A(g11117),.B(g8411));
  NAND3 NAND3_199(.VSS(VSS),.VDD(VDD),.Y(g28793),.A(g27800),.B(g7328),.C(g2153));
  NAND2 NAND2_1383(.VSS(VSS),.VDD(VDD),.Y(I13403),.A(g2250),.B(I13401));
  NAND2 NAND2_1384(.VSS(VSS),.VDD(VDD),.Y(I12278),.A(g1467),.B(I12277));
  NAND2 NAND2_1385(.VSS(VSS),.VDD(VDD),.Y(g24950),.A(g19442),.B(g23154));
  NAND2 NAND2_1386(.VSS(VSS),.VDD(VDD),.Y(I12469),.A(g405),.B(I12468));
  NAND3 NAND3_200(.VSS(VSS),.VDD(VDD),.Y(g27931),.A(g25425),.B(g25381),.C(g25780));
  NAND3 NAND3_201(.VSS(VSS),.VDD(VDD),.Y(g28765),.A(g27800),.B(g7374),.C(g7280));
  NAND2 NAND2_1387(.VSS(VSS),.VDD(VDD),.Y(g7611),.A(g4057),.B(g4064));
  NAND2 NAND2_1388(.VSS(VSS),.VDD(VDD),.Y(g14011),.A(g10295),.B(g11473));
  NAND4 NAND4_232(.VSS(VSS),.VDD(VDD),.Y(g20151),.A(g17598),.B(g14570),.C(g17514),.D(g14519));
  NAND2 NAND2_1389(.VSS(VSS),.VDD(VDD),.Y(g20172),.A(g16876),.B(g8131));
  NAND2 NAND2_1390(.VSS(VSS),.VDD(VDD),.Y(I12468),.A(g405),.B(g392));
  NAND2 NAND2_1391(.VSS(VSS),.VDD(VDD),.Y(g13291),.A(g10715),.B(g1500));
  NAND3 NAND3_202(.VSS(VSS),.VDD(VDD),.Y(g11173),.A(g4966),.B(g7898),.C(g9064));
  NAND2 NAND2_1392(.VSS(VSS),.VDD(VDD),.Y(g12190),.A(g8365),.B(g8255));
  NAND2 NAND2_1393(.VSS(VSS),.VDD(VDD),.Y(g22753),.A(g1536),.B(g19632));
  NAND3 NAND3_203(.VSS(VSS),.VDD(VDD),.Y(g28504),.A(g758),.B(g27528),.C(g11679));
  NAND4 NAND4_233(.VSS(VSS),.VDD(VDD),.Y(g21357),.A(g15736),.B(g13109),.C(g15726),.D(g13086));
  NAND3 NAND3_204(.VSS(VSS),.VDD(VDD),.Y(g31009),.A(g27187),.B(g29503),.C(g19644));
  NAND2 NAND2_1394(.VSS(VSS),.VDD(VDD),.Y(g14627),.A(g12553),.B(g12772));
  NAND2 NAND2_1395(.VSS(VSS),.VDD(VDD),.Y(g23357),.A(g20201),.B(g11231));
  NAND2 NAND2_1396(.VSS(VSS),.VDD(VDD),.Y(g14959),.A(g12695),.B(g12798));
  NAND2 NAND2_1397(.VSS(VSS),.VDD(VDD),.Y(g14379),.A(g5723),.B(g11907));
  NAND2 NAND2_1398(.VSS(VSS),.VDD(VDD),.Y(g22650),.A(g7888),.B(g19581));
  NAND3 NAND3_205(.VSS(VSS),.VDD(VDD),.Y(g11134),.A(g8138),.B(g8240),.C(g8301));
  NAND2 NAND2_1399(.VSS(VSS),.VDD(VDD),.Y(g23105),.A(g8097),.B(g19887));
  NAND2 NAND2_1400(.VSS(VSS),.VDD(VDD),.Y(g13134),.A(g11134),.B(g8470));
  NAND2 NAND2_1401(.VSS(VSS),.VDD(VDD),.Y(g14378),.A(g11979),.B(g9731));
  NAND2 NAND2_1402(.VSS(VSS),.VDD(VDD),.Y(g7209),.A(g6052),.B(g6098));
  NAND2 NAND2_1403(.VSS(VSS),.VDD(VDD),.Y(g12024),.A(g8381),.B(g8418));
  NAND4 NAND4_234(.VSS(VSS),.VDD(VDD),.Y(g17650),.A(g6299),.B(g12101),.C(g6315),.D(g14745));
  NAND2 NAND2_1404(.VSS(VSS),.VDD(VDD),.Y(g10603),.A(g10077),.B(g9751));
  NAND4 NAND4_235(.VSS(VSS),.VDD(VDD),.Y(g17736),.A(g5563),.B(g14522),.C(g5659),.D(g12563));
  NAND4 NAND4_236(.VSS(VSS),.VDD(VDD),.Y(g15798),.A(g6629),.B(g14602),.C(g6704),.D(g14786));
  NAND2 NAND2_1405(.VSS(VSS),.VDD(VDD),.Y(g25021),.A(g21417),.B(g23363));
  NAND2 NAND2_1406(.VSS(VSS),.VDD(VDD),.Y(I11824),.A(g4593),.B(g4601));
  NAND2 NAND2_1407(.VSS(VSS),.VDD(VDD),.Y(g15674),.A(g921),.B(g13110));
  NAND2 NAND2_1408(.VSS(VSS),.VDD(VDD),.Y(g9310),.A(I13078),.B(I13079));
  NAND2 NAND2_1409(.VSS(VSS),.VDD(VDD),.Y(I14289),.A(g8282),.B(g3835));
  NAND3 NAND3_206(.VSS(VSS),.VDD(VDD),.Y(g28298),.A(g10533),.B(g26131),.C(g26990));
  NAND2 NAND2_1410(.VSS(VSS),.VDD(VDD),.Y(g9663),.A(g128),.B(g4646));
  NAND4 NAND4_237(.VSS(VSS),.VDD(VDD),.Y(g13927),.A(g3578),.B(g11207),.C(g3632),.D(g11389));
  NAND2 NAND2_1411(.VSS(VSS),.VDD(VDD),.Y(I17494),.A(g13378),.B(g1448));
  NAND2 NAND2_1412(.VSS(VSS),.VDD(VDD),.Y(g29118),.A(g27886),.B(g9755));
  NAND2 NAND2_1413(.VSS(VSS),.VDD(VDD),.Y(I12217),.A(g1437),.B(g1478));
  NAND4 NAND4_238(.VSS(VSS),.VDD(VDD),.Y(g14730),.A(g5615),.B(g12093),.C(g5623),.D(g12301));
  NAND2 NAND2_1414(.VSS(VSS),.VDD(VDD),.Y(g22709),.A(g1193),.B(g19611));
  NAND2 NAND2_1415(.VSS(VSS),.VDD(VDD),.Y(I22822),.A(g11978),.B(g21434));
  NAND2 NAND2_1416(.VSS(VSS),.VDD(VDD),.Y(g13240),.A(g1046),.B(g10521));
  NAND2 NAND2_1417(.VSS(VSS),.VDD(VDD),.Y(g24957),.A(g21359),.B(g23462));
  NAND2 NAND2_1418(.VSS(VSS),.VDD(VDD),.Y(g11491),.A(g9982),.B(g4000));
  NAND2 NAND2_1419(.VSS(VSS),.VDD(VDD),.Y(g12644),.A(g10233),.B(g4531));
  NAND2 NAND2_1420(.VSS(VSS),.VDD(VDD),.Y(g11903),.A(g9099),.B(g3712));
  NAND2 NAND2_1421(.VSS(VSS),.VDD(VDD),.Y(I14816),.A(g9962),.B(g6513));
  NAND2 NAND2_1422(.VSS(VSS),.VDD(VDD),.Y(I32203),.A(g33937),.B(I32202));
  NAND2 NAND2_1423(.VSS(VSS),.VDD(VDD),.Y(g23890),.A(g7004),.B(g20682));
  NAND3 NAND3_207(.VSS(VSS),.VDD(VDD),.Y(g12969),.A(g4388),.B(g7178),.C(g10476));
  NAND2 NAND2_1424(.VSS(VSS),.VDD(VDD),.Y(I13520),.A(g2518),.B(I13518));
  NAND2 NAND2_1425(.VSS(VSS),.VDD(VDD),.Y(g20645),.A(g14344),.B(g17243));
  NAND2 NAND2_1426(.VSS(VSS),.VDD(VDD),.Y(g28856),.A(g27738),.B(g8093));
  NAND2 NAND2_1427(.VSS(VSS),.VDD(VDD),.Y(g14548),.A(g12208),.B(g5774));
  NAND2 NAND2_1428(.VSS(VSS),.VDD(VDD),.Y(g17225),.A(g8612),.B(g14367));
  NAND4 NAND4_239(.VSS(VSS),.VDD(VDD),.Y(g17708),.A(g5216),.B(g14490),.C(g5313),.D(g12497));
  NAND2 NAND2_1429(.VSS(VSS),.VDD(VDD),.Y(g12197),.A(g7296),.B(g5290));
  NAND2 NAND2_1430(.VSS(VSS),.VDD(VDD),.Y(g8434),.A(g3080),.B(g3072));
  NAND3 NAND3_208(.VSS(VSS),.VDD(VDD),.Y(g28512),.A(g10857),.B(g27155),.C(g27142));
  NAND2 NAND2_1431(.VSS(VSS),.VDD(VDD),.Y(g23552),.A(I22684),.B(I22685));
  NAND2 NAND2_1432(.VSS(VSS),.VDD(VDD),.Y(g15005),.A(g12667),.B(g12622));
  NAND2 NAND2_1433(.VSS(VSS),.VDD(VDD),.Y(g14317),.A(g5033),.B(g11862));
  NAND2 NAND2_1434(.VSS(VSS),.VDD(VDD),.Y(g12411),.A(g7393),.B(g5276));
  NAND3 NAND3_209(.VSS(VSS),.VDD(VDD),.Y(g8347),.A(g4358),.B(g4349),.C(g4340));
  NAND2 NAND2_1435(.VSS(VSS),.VDD(VDD),.Y(I15262),.A(g10081),.B(g2273));
  NAND2 NAND2_1436(.VSS(VSS),.VDD(VDD),.Y(g23778),.A(I22922),.B(I22923));
  NAND2 NAND2_1437(.VSS(VSS),.VDD(VDD),.Y(g11395),.A(g9601),.B(g3983));
  NAND2 NAND2_1438(.VSS(VSS),.VDD(VDD),.Y(I13497),.A(g255),.B(g232));
  NAND2 NAND2_1439(.VSS(VSS),.VDD(VDD),.Y(g11990),.A(g9166),.B(g703));
  NAND2 NAND2_1440(.VSS(VSS),.VDD(VDD),.Y(g13990),.A(g11669),.B(g11584));
  NAND2 NAND2_1441(.VSS(VSS),.VDD(VDD),.Y(g23786),.A(I22945),.B(I22946));
  NAND2 NAND2_1442(.VSS(VSS),.VDD(VDD),.Y(I18487),.A(g14611),.B(I18485));
  NAND2 NAND2_1443(.VSS(VSS),.VDD(VDD),.Y(g13898),.A(g11621),.B(g11747));
  NAND2 NAND2_1444(.VSS(VSS),.VDD(VDD),.Y(I22864),.A(g12146),.B(g21228));
  NAND4 NAND4_240(.VSS(VSS),.VDD(VDD),.Y(g21356),.A(g15780),.B(g15752),.C(g15743),.D(g13118));
  NAND2 NAND2_1445(.VSS(VSS),.VDD(VDD),.Y(I12373),.A(g3457),.B(I12372));
  NAND4 NAND4_241(.VSS(VSS),.VDD(VDD),.Y(g14626),.A(g12232),.B(g9852),.C(g12159),.D(g9715));
  NAND3 NAND3_210(.VSS(VSS),.VDD(VDD),.Y(g24661),.A(g23210),.B(g23195),.C(g22984));
  NAND3 NAND3_211(.VSS(VSS),.VDD(VDD),.Y(g24547),.A(g22638),.B(g22643),.C(g22754));
  NAND2 NAND2_1446(.VSS(VSS),.VDD(VDD),.Y(I31972),.A(g33641),.B(g33631));
  NAND2 NAND2_1447(.VSS(VSS),.VDD(VDD),.Y(g12450),.A(g7738),.B(g10281));
  NAND3 NAND3_212(.VSS(VSS),.VDD(VDD),.Y(g10775),.A(g7960),.B(g7943),.C(g8470));
  NAND2 NAND2_1448(.VSS(VSS),.VDD(VDD),.Y(g9295),.A(I13066),.B(I13067));
  NAND2 NAND2_1449(.VSS(VSS),.VDD(VDD),.Y(g12819),.A(g9848),.B(g6961));
  NAND2 NAND2_1450(.VSS(VSS),.VDD(VDD),.Y(g12910),.A(g11002),.B(g10601));
  NAND3 NAND3_213(.VSS(VSS),.VDD(VDD),.Y(g34174),.A(g617),.B(g33851),.C(g12323));
  NAND4 NAND4_242(.VSS(VSS),.VDD(VDD),.Y(g17792),.A(g6601),.B(g14602),.C(g6697),.D(g12721));
  NAND2 NAND2_1451(.VSS(VSS),.VDD(VDD),.Y(I22900),.A(g12193),.B(I22899));
  NAND2 NAND2_1452(.VSS(VSS),.VDD(VDD),.Y(g10737),.A(g6961),.B(g9848));
  NAND2 NAND2_1453(.VSS(VSS),.VDD(VDD),.Y(g25537),.A(g22763),.B(g2873));
  NAND2 NAND2_1454(.VSS(VSS),.VDD(VDD),.Y(g12111),.A(g847),.B(g9166));
  NAND3 NAND3_214(.VSS(VSS),.VDD(VDD),.Y(g28271),.A(g10533),.B(g27004),.C(g26990));
  NAND2 NAND2_1455(.VSS(VSS),.VDD(VDD),.Y(g13861),.A(g1459),.B(g10671));
  NAND2 NAND2_1456(.VSS(VSS),.VDD(VDD),.Y(g21331),.A(g11402),.B(g17157));
  NAND4 NAND4_243(.VSS(VSS),.VDD(VDD),.Y(g13573),.A(g8002),.B(g10544),.C(g7582),.D(g1351));
  NAND2 NAND2_1457(.VSS(VSS),.VDD(VDD),.Y(g23932),.A(g7051),.B(g20875));
  NAND2 NAND2_1458(.VSS(VSS),.VDD(VDD),.Y(I14713),.A(g9671),.B(I14712));
  NAND3 NAND3_215(.VSS(VSS),.VDD(VDD),.Y(g12590),.A(g7097),.B(g7110),.C(g10229));
  NAND2 NAND2_1459(.VSS(VSS),.VDD(VDD),.Y(g33083),.A(g7805),.B(g32118));
  NAND2 NAND2_1460(.VSS(VSS),.VDD(VDD),.Y(g11389),.A(I14399),.B(I14400));
  NAND2 NAND2_1461(.VSS(VSS),.VDD(VDD),.Y(g25492),.A(g12479),.B(g22457));
  NAND2 NAND2_1462(.VSS(VSS),.VDD(VDD),.Y(g14697),.A(g12662),.B(g12824));
  NAND2 NAND2_1463(.VSS(VSS),.VDD(VDD),.Y(g9966),.A(I13498),.B(I13499));
  NAND2 NAND2_1464(.VSS(VSS),.VDD(VDD),.Y(g7184),.A(g5706),.B(g5752));
  NAND2 NAND2_1465(.VSS(VSS),.VDD(VDD),.Y(g9705),.A(g2619),.B(g2587));
  NAND2 NAND2_1466(.VSS(VSS),.VDD(VDD),.Y(I14610),.A(g8993),.B(I14609));
  NAND2 NAND2_1467(.VSS(VSS),.VDD(VDD),.Y(I26368),.A(g14211),.B(I26366));
  NAND2 NAND2_1468(.VSS(VSS),.VDD(VDD),.Y(I29263),.A(g12046),.B(I29261));
  NAND2 NAND2_1469(.VSS(VSS),.VDD(VDD),.Y(g11534),.A(g7121),.B(g8958));
  NAND2 NAND2_1470(.VSS(VSS),.VDD(VDD),.Y(I23602),.A(g4322),.B(I23600));
  NAND2 NAND2_1471(.VSS(VSS),.VDD(VDD),.Y(g20784),.A(g14616),.B(g17595));
  NAND3 NAND3_216(.VSS(VSS),.VDD(VDD),.Y(g28736),.A(g27742),.B(g7308),.C(g7252));
  NAND4 NAND4_244(.VSS(VSS),.VDD(VDD),.Y(g19265),.A(g15721),.B(g15715),.C(g13091),.D(g15710));
  NAND4 NAND4_245(.VSS(VSS),.VDD(VDD),.Y(g13098),.A(g5933),.B(g12129),.C(g6023),.D(g9935));
  NAND2 NAND2_1472(.VSS(VSS),.VDD(VDD),.Y(I20487),.A(g16696),.B(I20486));
  NAND2 NAND2_1473(.VSS(VSS),.VDD(VDD),.Y(g11251),.A(g8438),.B(g3092));
  NAND2 NAND2_1474(.VSS(VSS),.VDD(VDD),.Y(g25381),.A(g538),.B(g23088));
  NAND2 NAND2_1475(.VSS(VSS),.VDD(VDD),.Y(I23970),.A(g22202),.B(I23969));
  NAND4 NAND4_246(.VSS(VSS),.VDD(VDD),.Y(g13462),.A(g12449),.B(g12412),.C(g12342),.D(g12294));
  NAND3 NAND3_217(.VSS(VSS),.VDD(VDD),.Y(g28843),.A(g27907),.B(g7456),.C(g7387));
  NAND3 NAND3_218(.VSS(VSS),.VDD(VDD),.Y(g19510),.A(g15969),.B(g10841),.C(g10899));
  NAND2 NAND2_1476(.VSS(VSS),.VDD(VDD),.Y(g20181),.A(g13252),.B(g16846));
  NAND2 NAND2_1477(.VSS(VSS),.VDD(VDD),.Y(g12019),.A(g7322),.B(g1906));
  NAND4 NAND4_247(.VSS(VSS),.VDD(VDD),.Y(g17598),.A(g3949),.B(g13824),.C(g4027),.D(g8595));
  NAND2 NAND2_1478(.VSS(VSS),.VDD(VDD),.Y(g12196),.A(g8764),.B(g4688));
  NAND2 NAND2_1479(.VSS(VSS),.VDD(VDD),.Y(g11997),.A(g2319),.B(g8316));
  NAND2 NAND2_1480(.VSS(VSS),.VDD(VDD),.Y(I20469),.A(g16728),.B(I20467));
  NAND2 NAND2_1481(.VSS(VSS),.VDD(VDD),.Y(I21994),.A(g19638),.B(I21992));
  NAND2 NAND2_1482(.VSS(VSS),.VDD(VDD),.Y(I12242),.A(g1105),.B(I12240));
  NAND3 NAND3_219(.VSS(VSS),.VDD(VDD),.Y(g12526),.A(g10194),.B(g7110),.C(g10213));
  NAND4 NAND4_248(.VSS(VSS),.VDD(VDD),.Y(g15725),.A(g5603),.B(g14522),.C(g5681),.D(g9864));
  NAND2 NAND2_1483(.VSS(VSS),.VDD(VDD),.Y(I20468),.A(g16663),.B(I20467));
  NAND2 NAND2_1484(.VSS(VSS),.VDD(VDD),.Y(g29154),.A(g27937),.B(g9835));
  NAND4 NAND4_249(.VSS(VSS),.VDD(VDD),.Y(g21433),.A(g17792),.B(g14830),.C(g17765),.D(g14750));
  NAND2 NAND2_1485(.VSS(VSS),.VDD(VDD),.Y(I22892),.A(g12189),.B(g21228));
  NAND2 NAND2_1486(.VSS(VSS),.VDD(VDD),.Y(g19442),.A(g11431),.B(g17794));
  NAND2 NAND2_1487(.VSS(VSS),.VDD(VDD),.Y(g12402),.A(g7704),.B(g10266));
  NAND2 NAND2_1488(.VSS(VSS),.VDD(VDD),.Y(g10611),.A(g10115),.B(g9831));
  NAND2 NAND2_1489(.VSS(VSS),.VDD(VDD),.Y(I13111),.A(g5813),.B(I13109));
  NAND2 NAND2_1490(.VSS(VSS),.VDD(VDD),.Y(g13871),.A(g4955),.B(g11834));
  NAND2 NAND2_1491(.VSS(VSS),.VDD(VDD),.Y(I23919),.A(g9333),.B(I23917));
  NAND2 NAND2_1492(.VSS(VSS),.VDD(VDD),.Y(I18486),.A(g1677),.B(I18485));
  NAND3 NAND3_220(.VSS(VSS),.VDD(VDD),.Y(g28259),.A(g10504),.B(g26987),.C(g26973));
  NAND2 NAND2_1493(.VSS(VSS),.VDD(VDD),.Y(g14924),.A(g12558),.B(g12505));
  NAND2 NAND2_1494(.VSS(VSS),.VDD(VDD),.Y(I22712),.A(g21434),.B(I22710));
  NAND2 NAND2_1495(.VSS(VSS),.VDD(VDD),.Y(g17656),.A(I18626),.B(I18627));
  NAND2 NAND2_1496(.VSS(VSS),.VDD(VDD),.Y(I20187),.A(g16272),.B(g1333));
  NAND4 NAND4_250(.VSS(VSS),.VDD(VDD),.Y(g15744),.A(g6641),.B(g14602),.C(g6719),.D(g10061));
  NAND2 NAND2_1497(.VSS(VSS),.VDD(VDD),.Y(I17476),.A(g1105),.B(I17474));
  NAND2 NAND2_1498(.VSS(VSS),.VDD(VDD),.Y(I23918),.A(g23975),.B(I23917));
  NAND2 NAND2_1499(.VSS(VSS),.VDD(VDD),.Y(I18580),.A(g1945),.B(I18579));
  NAND2 NAND2_1500(.VSS(VSS),.VDD(VDD),.Y(I26050),.A(g25997),.B(I26049));
  NAND2 NAND2_1501(.VSS(VSS),.VDD(VDD),.Y(I13384),.A(g246),.B(I13382));
  NAND2 NAND2_1502(.VSS(VSS),.VDD(VDD),.Y(g12001),.A(I14854),.B(I14855));
  NAND2 NAND2_1503(.VSS(VSS),.VDD(VDD),.Y(I13067),.A(g4304),.B(I13065));
  NAND2 NAND2_1504(.VSS(VSS),.VDD(VDD),.Y(I12841),.A(g4222),.B(I12840));
  NAND2 NAND2_1505(.VSS(VSS),.VDD(VDD),.Y(I11877),.A(g4388),.B(g4430));
  NAND2 NAND2_1506(.VSS(VSS),.VDD(VDD),.Y(g10529),.A(g1592),.B(g7308));
  NAND2 NAND2_1507(.VSS(VSS),.VDD(VDD),.Y(g13628),.A(g3372),.B(g11107));
  NAND2 NAND2_1508(.VSS(VSS),.VDD(VDD),.Y(g23850),.A(g12185),.B(g19462));
  NAND2 NAND2_1509(.VSS(VSS),.VDD(VDD),.Y(g13911),.A(g11834),.B(g4917));
  NAND2 NAND2_1510(.VSS(VSS),.VDD(VDD),.Y(I18531),.A(g14640),.B(I18529));
  NAND2 NAND2_1511(.VSS(VSS),.VDD(VDD),.Y(g17364),.A(g8639),.B(g14367));
  NAND3 NAND3_221(.VSS(VSS),.VDD(VDD),.Y(g28955),.A(g27837),.B(g1936),.C(g7362));
  NAND2 NAND2_1512(.VSS(VSS),.VDD(VDD),.Y(I14277),.A(g3484),.B(I14275));
  NAND2 NAND2_1513(.VSS(VSS),.VDD(VDD),.Y(I21977),.A(g7680),.B(I21976));
  NAND4 NAND4_251(.VSS(VSS),.VDD(VDD),.Y(g14696),.A(g5567),.B(g12093),.C(g5685),.D(g12563));
  NAND2 NAND2_1514(.VSS(VSS),.VDD(VDD),.Y(I24363),.A(g23687),.B(g14320));
  NAND2 NAND2_1515(.VSS(VSS),.VDD(VDD),.Y(g8163),.A(g3419),.B(g3423));
  NAND3 NAND3_222(.VSS(VSS),.VDD(VDD),.Y(g15962),.A(g14833),.B(g9417),.C(g9340));
  NAND2 NAND2_1516(.VSS(VSS),.VDD(VDD),.Y(g14764),.A(g7738),.B(g12798));
  NAND2 NAND2_1517(.VSS(VSS),.VDD(VDD),.Y(g11591),.A(I14531),.B(I14532));
  NAND3 NAND3_223(.VSS(VSS),.VDD(VDD),.Y(g21011),.A(g14504),.B(g17399),.C(g9629));
  NAND2 NAND2_1518(.VSS(VSS),.VDD(VDD),.Y(I15147),.A(g9864),.B(g5659));
  NAND2 NAND2_1519(.VSS(VSS),.VDD(VDD),.Y(g12066),.A(I14924),.B(I14925));
  NAND2 NAND2_1520(.VSS(VSS),.VDD(VDD),.Y(I20486),.A(g16696),.B(g16757));
  NAND2 NAND2_1521(.VSS(VSS),.VDD(VDD),.Y(g24943),.A(g20068),.B(g23172));
  NAND3 NAND3_224(.VSS(VSS),.VDD(VDD),.Y(g20644),.A(g14342),.B(g17220),.C(g9372));
  NAND2 NAND2_1522(.VSS(VSS),.VDD(VDD),.Y(g27876),.A(I26418),.B(I26419));
  NAND3 NAND3_225(.VSS(VSS),.VDD(VDD),.Y(g15833),.A(g14714),.B(g12378),.C(g12337));
  NAND2 NAND2_1523(.VSS(VSS),.VDD(VDD),.Y(I13402),.A(g2246),.B(I13401));
  NAND2 NAND2_1524(.VSS(VSS),.VDD(VDD),.Y(g11355),.A(g9551),.B(g3310));
  NAND3 NAND3_226(.VSS(VSS),.VDD(VDD),.Y(g28994),.A(g27907),.B(g2495),.C(g7424));
  NAND2 NAND2_1525(.VSS(VSS),.VDD(VDD),.Y(g14868),.A(g12755),.B(g12680));
  NAND2 NAND2_1526(.VSS(VSS),.VDD(VDD),.Y(g17571),.A(g8579),.B(g14367));
  NAND2 NAND2_1527(.VSS(VSS),.VDD(VDD),.Y(I11866),.A(g4401),.B(I11864));
  NAND4 NAND4_252(.VSS(VSS),.VDD(VDD),.Y(g27854),.A(g21228),.B(g25283),.C(g26424),.D(g26195));
  NAND2 NAND2_1528(.VSS(VSS),.VDD(VDD),.Y(g25062),.A(g21403),.B(g23363));
  NAND2 NAND2_1529(.VSS(VSS),.VDD(VDD),.Y(I20223),.A(g11170),.B(I20221));
  NAND2 NAND2_1530(.VSS(VSS),.VDD(VDD),.Y(g16507),.A(g13797),.B(g13764));
  NAND2 NAND2_1531(.VSS(VSS),.VDD(VDD),.Y(g11858),.A(g9014),.B(g3010));
  NAND2 NAND2_1532(.VSS(VSS),.VDD(VDD),.Y(I14352),.A(g8848),.B(I14350));
  NAND2 NAND2_1533(.VSS(VSS),.VDD(VDD),.Y(I17883),.A(g13336),.B(g1135));
  NAND2 NAND2_1534(.VSS(VSS),.VDD(VDD),.Y(g11172),.A(g8478),.B(g3096));
  NAND3 NAND3_227(.VSS(VSS),.VDD(VDD),.Y(g12511),.A(g7028),.B(g5644),.C(g5698));
  NAND2 NAND2_1535(.VSS(VSS),.VDD(VDD),.Y(g22687),.A(g19560),.B(g7870));
  NAND2 NAND2_1536(.VSS(VSS),.VDD(VDD),.Y(g7885),.A(I12270),.B(I12271));
  NAND2 NAND2_1537(.VSS(VSS),.VDD(VDD),.Y(g11996),.A(g7280),.B(g2197));
  NAND4 NAND4_253(.VSS(VSS),.VDD(VDD),.Y(g17495),.A(g3566),.B(g13730),.C(g3668),.D(g8542));
  NAND2 NAND2_1538(.VSS(VSS),.VDD(VDD),.Y(g23379),.A(g20216),.B(g11248));
  NAND2 NAND2_1539(.VSS(VSS),.VDD(VDD),.Y(I14170),.A(g8389),.B(I14169));
  NAND2 NAND2_1540(.VSS(VSS),.VDD(VDD),.Y(I13077),.A(g5462),.B(g5467));
  NAND2 NAND2_1541(.VSS(VSS),.VDD(VDD),.Y(g23112),.A(g21024),.B(g10733));
  NAND3 NAND3_228(.VSS(VSS),.VDD(VDD),.Y(g20870),.A(g14432),.B(g17315),.C(g9567));
  NAND4 NAND4_254(.VSS(VSS),.VDD(VDD),.Y(g17816),.A(g6657),.B(g14602),.C(g6668),.D(g10061));
  NAND2 NAND2_1542(.VSS(VSS),.VDD(VDD),.Y(g14258),.A(g9203),.B(g11903));
  NAND2 NAND2_1543(.VSS(VSS),.VDD(VDD),.Y(g11394),.A(g9600),.B(g3661));
  NAND2 NAND2_1544(.VSS(VSS),.VDD(VDD),.Y(g22643),.A(g20136),.B(g18954));
  NAND2 NAND2_1545(.VSS(VSS),.VDD(VDD),.Y(g34051),.A(I31973),.B(I31974));
  NAND4 NAND4_255(.VSS(VSS),.VDD(VDD),.Y(g21386),.A(g15798),.B(g15788),.C(g15782),.D(g13139));
  NAND2 NAND2_1546(.VSS(VSS),.VDD(VDD),.Y(I18587),.A(g2370),.B(g14679));
  NAND4 NAND4_256(.VSS(VSS),.VDD(VDD),.Y(g21603),.A(g17872),.B(g14987),.C(g17723),.D(g17689));
  NAND2 NAND2_1547(.VSS(VSS),.VDD(VDD),.Y(I14853),.A(g9433),.B(g5142));
  NAND2 NAND2_1548(.VSS(VSS),.VDD(VDD),.Y(g27550),.A(g24943),.B(g25772));
  NAND2 NAND2_1549(.VSS(VSS),.VDD(VDD),.Y(g9485),.A(g1657),.B(g1624));
  NAND2 NAND2_1550(.VSS(VSS),.VDD(VDD),.Y(g14069),.A(g11653),.B(g8864));
  NAND2 NAND2_1551(.VSS(VSS),.VDD(VDD),.Y(g22668),.A(g20219),.B(g2912));
  NAND2 NAND2_1552(.VSS(VSS),.VDD(VDD),.Y(g10602),.A(g7411),.B(g7451));
  NAND3 NAND3_229(.VSS(VSS),.VDD(VDD),.Y(g11446),.A(g8700),.B(g6941),.C(g8734));
  NAND2 NAND2_1553(.VSS(VSS),.VDD(VDD),.Y(g14810),.A(g12700),.B(g10312));
  NAND2 NAND2_1554(.VSS(VSS),.VDD(VDD),.Y(g15033),.A(g12806),.B(g7142));
  NAND2 NAND2_1555(.VSS(VSS),.VDD(VDD),.Y(g12287),.A(g8381),.B(g2587));
  NAND4 NAND4_257(.VSS(VSS),.VDD(VDD),.Y(g21429),.A(g17788),.B(g14803),.C(g17578),.D(g17520));
  NAND4 NAND4_258(.VSS(VSS),.VDD(VDD),.Y(g17669),.A(g3570),.B(g11238),.C(g3632),.D(g13902));
  NAND2 NAND2_1556(.VSS(VSS),.VDD(VDD),.Y(g12307),.A(g7395),.B(g5983));
  NAND2 NAND2_1557(.VSS(VSS),.VDD(VDD),.Y(g14879),.A(g12646),.B(g10266));
  NAND2 NAND2_1558(.VSS(VSS),.VDD(VDD),.Y(I13066),.A(g4308),.B(I13065));
  NAND4 NAND4_259(.VSS(VSS),.VDD(VDD),.Y(g17668),.A(g3235),.B(g13765),.C(g3310),.D(g13877));
  NAND2 NAND2_1559(.VSS(VSS),.VDD(VDD),.Y(g23428),.A(g13945),.B(g20522));
  NAND2 NAND2_1560(.VSS(VSS),.VDD(VDD),.Y(g13058),.A(g10544),.B(g1312));
  NAND3 NAND3_230(.VSS(VSS),.VDD(VDD),.Y(g28977),.A(g27937),.B(g2629),.C(g2555));
  NAND2 NAND2_1561(.VSS(VSS),.VDD(VDD),.Y(g12431),.A(I15254),.B(I15255));
  NAND2 NAND2_1562(.VSS(VSS),.VDD(VDD),.Y(g20979),.A(g5385),.B(g17309));
  NAND3 NAND3_231(.VSS(VSS),.VDD(VDD),.Y(g28783),.A(g27779),.B(g7315),.C(g1728));
  NAND2 NAND2_1563(.VSS(VSS),.VDD(VDD),.Y(g20055),.A(g11269),.B(g17794));
  NAND4 NAND4_260(.VSS(VSS),.VDD(VDD),.Y(g20111),.A(g17513),.B(g14517),.C(g17468),.D(g14422));
  NAND2 NAND2_1564(.VSS(VSS),.VDD(VDD),.Y(g17525),.A(g14600),.B(g14574));
  NAND2 NAND2_1565(.VSS(VSS),.VDD(VDD),.Y(I13511),.A(g2093),.B(I13509));
  NAND2 NAND2_1566(.VSS(VSS),.VDD(VDD),.Y(g12341),.A(g7512),.B(g5308));
  NAND2 NAND2_1567(.VSS(VSS),.VDD(VDD),.Y(g28823),.A(g27738),.B(g14565));
  NAND2 NAND2_1568(.VSS(VSS),.VDD(VDD),.Y(I14276),.A(g8218),.B(I14275));
  NAND2 NAND2_1569(.VSS(VSS),.VDD(VDD),.Y(I21976),.A(g7680),.B(g19620));
  NAND2 NAND2_1570(.VSS(VSS),.VDD(VDD),.Y(g16291),.A(g13551),.B(g13545));
  NAND2 NAND2_1571(.VSS(VSS),.VDD(VDD),.Y(I23985),.A(g22182),.B(g482));
  NAND2 NAND2_1572(.VSS(VSS),.VDD(VDD),.Y(g13281),.A(g10916),.B(g1099));
  NAND2 NAND2_1573(.VSS(VSS),.VDD(VDD),.Y(g27670),.A(g25172),.B(g26666));
  NAND2 NAND2_1574(.VSS(VSS),.VDD(VDD),.Y(g22713),.A(g20114),.B(g2890));
  NAND2 NAND2_1575(.VSS(VSS),.VDD(VDD),.Y(g11957),.A(g8205),.B(g8259));
  NAND4 NAND4_261(.VSS(VSS),.VDD(VDD),.Y(g28336),.A(g27064),.B(g24756),.C(g27163),.D(g19644));
  NAND2 NAND2_1576(.VSS(VSS),.VDD(VDD),.Y(I32202),.A(g33937),.B(g33670));
  NAND2 NAND2_1577(.VSS(VSS),.VDD(VDD),.Y(g13739),.A(g11773),.B(g11261));
  NAND3 NAND3_232(.VSS(VSS),.VDD(VDD),.Y(g25396),.A(g22384),.B(g2208),.C(g8259));
  NAND3 NAND3_233(.VSS(VSS),.VDD(VDD),.Y(g28966),.A(g27858),.B(g2361),.C(g7380));
  NAND2 NAND2_1578(.VSS(VSS),.VDD(VDD),.Y(g14918),.A(g12646),.B(g12772));
  NAND4 NAND4_262(.VSS(VSS),.VDD(VDD),.Y(g20150),.A(g17705),.B(g17669),.C(g17635),.D(g14590));
  NAND2 NAND2_1579(.VSS(VSS),.VDD(VDD),.Y(g14079),.A(g11626),.B(g11763));
  NAND4 NAND4_263(.VSS(VSS),.VDD(VDD),.Y(g17705),.A(g3586),.B(g13799),.C(g3661),.D(g13902));
  NAND2 NAND2_1580(.VSS(VSS),.VDD(VDD),.Y(g8292),.A(g218),.B(g215));
  NAND2 NAND2_1581(.VSS(VSS),.VDD(VDD),.Y(g14599),.A(g12207),.B(g9739));
  NAND2 NAND2_1582(.VSS(VSS),.VDD(VDD),.Y(I12253),.A(g1129),.B(I12251));
  NAND4 NAND4_264(.VSS(VSS),.VDD(VDD),.Y(g17679),.A(g5611),.B(g14425),.C(g5681),.D(g12563));
  NAND2 NAND2_1583(.VSS(VSS),.VDD(VDD),.Y(g7869),.A(I12252),.B(I12253));
  NAND2 NAND2_1584(.VSS(VSS),.VDD(VDD),.Y(g10598),.A(g7191),.B(g6404));
  NAND4 NAND4_265(.VSS(VSS),.VDD(VDD),.Y(g15788),.A(g6613),.B(g12211),.C(g6675),.D(g14786));
  NAND2 NAND2_1585(.VSS(VSS),.VDD(VDD),.Y(I18579),.A(g1945),.B(g14678));
  NAND4 NAND4_266(.VSS(VSS),.VDD(VDD),.Y(g14598),.A(g5248),.B(g12002),.C(g5331),.D(g12497));
  NAND2 NAND2_1586(.VSS(VSS),.VDD(VDD),.Y(I14733),.A(g9732),.B(g5475));
  NAND2 NAND2_1587(.VSS(VSS),.VDD(VDD),.Y(g15829),.A(g4112),.B(g13831));
  NAND4 NAND4_267(.VSS(VSS),.VDD(VDD),.Y(g17686),.A(g6251),.B(g14529),.C(g6322),.D(g12672));
  NAND2 NAND2_1588(.VSS(VSS),.VDD(VDD),.Y(I12372),.A(g3457),.B(g3462));
  NAND2 NAND2_1589(.VSS(VSS),.VDD(VDD),.Y(g14817),.A(g12711),.B(g12622));
  NAND3 NAND3_234(.VSS(VSS),.VDD(VDD),.Y(g28288),.A(g10533),.B(g26105),.C(g27004));
  NAND2 NAND2_1590(.VSS(VSS),.VDD(VDD),.Y(g19913),.A(g11430),.B(g17794));
  NAND2 NAND2_1591(.VSS(VSS),.VDD(VDD),.Y(g19614),.A(g1542),.B(g16047));
  NAND2 NAND2_1592(.VSS(VSS),.VDD(VDD),.Y(g22875),.A(g20516),.B(g2980));
  NAND2 NAND2_1593(.VSS(VSS),.VDD(VDD),.Y(g25020),.A(g21377),.B(g23462));
  NAND2 NAND2_1594(.VSS(VSS),.VDD(VDD),.Y(g7442),.A(g896),.B(g890));
  NAND2 NAND2_1595(.VSS(VSS),.VDD(VDD),.Y(g24917),.A(g19913),.B(g23172));
  NAND2 NAND2_1596(.VSS(VSS),.VDD(VDD),.Y(g10561),.A(g7157),.B(g5712));
  NAND4 NAND4_268(.VSS(VSS),.VDD(VDD),.Y(g27468),.A(g24951),.B(g24932),.C(g24925),.D(g26852));
  NAND2 NAND2_1597(.VSS(VSS),.VDD(VDD),.Y(I22921),.A(g14677),.B(g21284));
  NAND2 NAND2_1598(.VSS(VSS),.VDD(VDD),.Y(g27306),.A(g24787),.B(g26235));
  NAND2 NAND2_1599(.VSS(VSS),.VDD(VDD),.Y(g19530),.A(g15829),.B(g10841));
  NAND2 NAND2_1600(.VSS(VSS),.VDD(VDD),.Y(g12286),.A(I15129),.B(I15130));
  NAND2 NAND2_1601(.VSS(VSS),.VDD(VDD),.Y(g14656),.A(g12553),.B(g12405));
  NAND2 NAND2_1602(.VSS(VSS),.VDD(VDD),.Y(g9177),.A(g3355),.B(g3401));
  NAND2 NAND2_1603(.VSS(VSS),.VDD(VDD),.Y(g22837),.A(g20219),.B(g2907));
  NAND2 NAND2_1604(.VSS(VSS),.VDD(VDD),.Y(g12306),.A(g7394),.B(g5666));
  NAND2 NAND2_1605(.VSS(VSS),.VDD(VDD),.Y(I26461),.A(g14306),.B(I26459));
  NAND2 NAND2_1606(.VSS(VSS),.VDD(VDD),.Y(I24416),.A(g14382),.B(I24414));
  NAND4 NAND4_269(.VSS(VSS),.VDD(VDD),.Y(g16604),.A(g3251),.B(g11194),.C(g3267),.D(g13877));
  NAND2 NAND2_1607(.VSS(VSS),.VDD(VDD),.Y(I22799),.A(g11960),.B(g21434));
  NAND4 NAND4_270(.VSS(VSS),.VDD(VDD),.Y(g13551),.A(g11812),.B(g7479),.C(g7903),.D(g10521));
  NAND2 NAND2_1608(.VSS(VSS),.VDD(VDD),.Y(g10336),.A(I13750),.B(I13751));
  NAND2 NAND2_1609(.VSS(VSS),.VDD(VDD),.Y(g28976),.A(g27903),.B(g8273));
  NAND2 NAND2_1610(.VSS(VSS),.VDD(VDD),.Y(I14712),.A(g9671),.B(g5128));
  NAND2 NAND2_1611(.VSS(VSS),.VDD(VDD),.Y(I13335),.A(g1687),.B(I13334));
  NAND4 NAND4_271(.VSS(VSS),.VDD(VDD),.Y(g16770),.A(g3263),.B(g13765),.C(g3274),.D(g8481));
  NAND2 NAND2_1612(.VSS(VSS),.VDD(VDD),.Y(g8561),.A(g3782),.B(g3774));
  NAND2 NAND2_1613(.VSS(VSS),.VDD(VDD),.Y(I22973),.A(g9657),.B(I22972));
  NAND2 NAND2_1614(.VSS(VSS),.VDD(VDD),.Y(g26248),.A(I25220),.B(I25221));
  NAND2 NAND2_1615(.VSS(VSS),.VDD(VDD),.Y(g12187),.A(I15042),.B(I15043));
  NAND2 NAND2_1616(.VSS(VSS),.VDD(VDD),.Y(I29262),.A(g29485),.B(I29261));
  NAND3 NAND3_235(.VSS(VSS),.VDD(VDD),.Y(g11490),.A(g8666),.B(g3639),.C(g3694));
  NAND2 NAND2_1617(.VSS(VSS),.VDD(VDD),.Y(I26393),.A(g26488),.B(g14227));
//
  NOR2 NOR2_0(.VSS(VSS),.VDD(VDD),.Y(g30249),.A(g5297),.B(g28982));
  NOR2 NOR2_1(.VSS(VSS),.VDD(VDD),.Y(g33141),.A(g32099),.B(g8400));
  NOR2 NOR2_2(.VSS(VSS),.VDD(VDD),.Y(g13824),.A(g8623),.B(g11702));
  NOR2 NOR2_3(.VSS(VSS),.VDD(VDD),.Y(g27479),.A(g9056),.B(g26616));
  NOR2 NOR2_4(.VSS(VSS),.VDD(VDD),.Y(g12479),.A(g2028),.B(g8310));
  NOR2 NOR2_5(.VSS(VSS),.VDD(VDD),.Y(g20854),.A(g5381),.B(g17243));
  NOR2 NOR2_6(.VSS(VSS),.VDD(VDD),.Y(g33135),.A(g32090),.B(g8350));
  NOR4 NOR4_0(.VSS(VSS),.VDD(VDD),.Y(g7675),.A(g1554),.B(g1559),.C(g1564),.D(g1548));
  NOR4 NOR4_1(.VSS(VSS),.VDD(VDD),.Y(g12486),.A(g9055),.B(g9013),.C(g8957),.D(g8905));
  NOR2 NOR2_7(.VSS(VSS),.VDD(VDD),.Y(g9694),.A(g1936),.B(g1862));
  NOR2 NOR2_8(.VSS(VSS),.VDD(VDD),.Y(g8906),.A(g3530),.B(g3522));
  NOR2 NOR2_9(.VSS(VSS),.VDD(VDD),.Y(g14816),.A(g10166),.B(g12252));
  NOR2 NOR2_10(.VSS(VSS),.VDD(VDD),.Y(g12223),.A(g2051),.B(g8365));
  NOR2 NOR2_11(.VSS(VSS),.VDD(VDD),.Y(g14687),.A(g5352),.B(g12166));
  NOR2 NOR2_12(.VSS(VSS),.VDD(VDD),.Y(g14752),.A(g12540),.B(g10040));
  NOR2 NOR2_13(.VSS(VSS),.VDD(VDD),.Y(g16272),.A(g13580),.B(g11189));
  NOR2 NOR2_14(.VSS(VSS),.VDD(VDD),.Y(g22524),.A(g19720),.B(g1361));
  NOR2 NOR2_15(.VSS(VSS),.VDD(VDD),.Y(g25778),.A(g25459),.B(g25420));
  NOR2 NOR2_16(.VSS(VSS),.VDD(VDD),.Y(g26212),.A(g23837),.B(g25408));
  NOR2 NOR2_17(.VSS(VSS),.VDD(VDD),.Y(g17194),.A(g11039),.B(g13480));
  NOR2 NOR2_18(.VSS(VSS),.VDD(VDD),.Y(g14392),.A(g12114),.B(g9537));
  NOR2 NOR2_19(.VSS(VSS),.VDD(VDD),.Y(g13700),.A(g3288),.B(g11615));
  NOR2 NOR2_20(.VSS(VSS),.VDD(VDD),.Y(g11658),.A(g8021),.B(g3506));
  NOR2 NOR2_21(.VSS(VSS),.VDD(VDD),.Y(g15718),.A(g13858),.B(g11330));
  NOR3 NOR3_0(.VSS(VSS),.VDD(VDD),.Y(g10488),.A(g4616),.B(g7133),.C(g10336));
  NOR3 NOR3_1(.VSS(VSS),.VDD(VDD),.Y(g29107),.A(g6203),.B(g7791),.C(g26977));
  NOR3 NOR3_2(.VSS(VSS),.VDD(VDD),.Y(g10893),.A(g1189),.B(g7715),.C(g7749));
  NOR2 NOR2_22(.VSS(VSS),.VDD(VDD),.Y(g25932),.A(g7680),.B(g24528));
  NOR2 NOR2_23(.VSS(VSS),.VDD(VDD),.Y(g29141),.A(g9374),.B(g27999));
  NOR2 NOR2_24(.VSS(VSS),.VDD(VDD),.Y(g14713),.A(g12483),.B(g9974));
  NOR2 NOR2_25(.VSS(VSS),.VDD(VDD),.Y(g31507),.A(g9064),.B(g29556));
  NOR2 NOR2_26(.VSS(VSS),.VDD(VDD),.Y(g15099),.A(g13191),.B(g12869));
  NOR2 NOR2_27(.VSS(VSS),.VDD(VDD),.Y(g11527),.A(g8165),.B(g8114));
  NOR3 NOR3_3(.VSS(VSS),.VDD(VDD),.Y(g32715),.A(g31327),.B(I30261),.C(I30262));
  NOR2 NOR2_28(.VSS(VSS),.VDD(VDD),.Y(g15098),.A(g13191),.B(g6927));
  NOR2 NOR2_29(.VSS(VSS),.VDD(VDD),.Y(g30148),.A(g28799),.B(g7335));
  NOR2 NOR2_30(.VSS(VSS),.VDD(VDD),.Y(g23602),.A(g9672),.B(g20979));
  NOR2 NOR2_31(.VSS(VSS),.VDD(VDD),.Y(g28470),.A(g8021),.B(g27617));
  NOR2 NOR2_32(.VSS(VSS),.VDD(VDD),.Y(g16220),.A(g13499),.B(g4939));
  NOR2 NOR2_33(.VSS(VSS),.VDD(VDD),.Y(g14679),.A(g12437),.B(g9911));
  NOR2 NOR2_34(.VSS(VSS),.VDD(VDD),.Y(g23955),.A(g2823),.B(g18890));
  NOR2 NOR2_35(.VSS(VSS),.VDD(VDD),.Y(g33163),.A(g32099),.B(g7809));
  NOR2 NOR2_36(.VSS(VSS),.VDD(VDD),.Y(g24619),.A(g23554),.B(g23581));
  NOR2 NOR2_37(.VSS(VSS),.VDD(VDD),.Y(g14188),.A(g9162),.B(g12259));
  NOR2 NOR2_38(.VSS(VSS),.VDD(VDD),.Y(g14124),.A(g8830),.B(g11083));
  NOR2 NOR2_39(.VSS(VSS),.VDD(VDD),.Y(g14678),.A(g12432),.B(g9907));
  NOR2 NOR2_40(.VSS(VSS),.VDD(VDD),.Y(g16246),.A(g13551),.B(g11169));
  NOR2 NOR2_41(.VSS(VSS),.VDD(VDD),.Y(g12117),.A(g10113),.B(g9755));
  NOR2 NOR2_42(.VSS(VSS),.VDD(VDD),.Y(g29361),.A(g7553),.B(g28174));
  NOR2 NOR2_43(.VSS(VSS),.VDD(VDD),.Y(g15140),.A(g12887),.B(g13680));
  NOR2 NOR2_44(.VSS(VSS),.VDD(VDD),.Y(g14093),.A(g8833),.B(g11083));
  NOR2 NOR2_45(.VSS(VSS),.VDD(VDD),.Y(g15061),.A(g6815),.B(g13394));
  NOR3 NOR3_4(.VSS(VSS),.VDD(VDD),.Y(g13910),.A(g4899),.B(g4975),.C(g11173));
  NOR2 NOR2_46(.VSS(VSS),.VDD(VDD),.Y(g13202),.A(g8347),.B(g10511));
  NOR2 NOR2_47(.VSS(VSS),.VDD(VDD),.Y(g12123),.A(g6856),.B(g2748));
  NOR2 NOR2_48(.VSS(VSS),.VDD(VDD),.Y(g27772),.A(g7297),.B(g25839));
  NOR2 NOR2_49(.VSS(VSS),.VDD(VDD),.Y(g12772),.A(g5188),.B(g9300));
  NOR2 NOR2_50(.VSS(VSS),.VDD(VDD),.Y(g31121),.A(g4776),.B(g29540));
  NOR2 NOR2_51(.VSS(VSS),.VDD(VDD),.Y(g23918),.A(g2799),.B(g21382));
  NOR2 NOR2_52(.VSS(VSS),.VDD(VDD),.Y(g15162),.A(g13809),.B(g12904));
  NOR2 NOR2_53(.VSS(VSS),.VDD(VDD),.Y(g11384),.A(g8538),.B(g8540));
  NOR2 NOR2_54(.VSS(VSS),.VDD(VDD),.Y(g23079),.A(g8390),.B(g19965));
  NOR2 NOR2_55(.VSS(VSS),.VDD(VDD),.Y(g29106),.A(g9451),.B(g28020));
  NOR2 NOR2_56(.VSS(VSS),.VDD(VDD),.Y(g13094),.A(g7487),.B(g10762));
  NOR2 NOR2_57(.VSS(VSS),.VDD(VDD),.Y(g26603),.A(g24908),.B(g24900));
  NOR3 NOR3_5(.VSS(VSS),.VDD(VDD),.Y(g29033),.A(g5511),.B(g7738),.C(g28010));
  NOR2 NOR2_58(.VSS(VSS),.VDD(VDD),.Y(g15628),.A(g11907),.B(g14228));
  NOR3 NOR3_6(.VSS(VSS),.VDD(VDD),.Y(g32520),.A(g31554),.B(I30054),.C(I30055));
  NOR2 NOR2_59(.VSS(VSS),.VDD(VDD),.Y(g17239),.A(g11119),.B(g13518));
  NOR3 NOR3_7(.VSS(VSS),.VDD(VDD),.Y(g31134),.A(g8033),.B(g29679),.C(g24732));
  NOR2 NOR2_60(.VSS(VSS),.VDD(VDD),.Y(g33134),.A(g7686),.B(g32057));
  NOR2 NOR2_61(.VSS(VSS),.VDD(VDD),.Y(g16227),.A(g1554),.B(g13574));
  NOR2 NOR2_62(.VSS(VSS),.VDD(VDD),.Y(g27007),.A(g5706),.B(g25821));
  NOR2 NOR2_63(.VSS(VSS),.VDD(VDD),.Y(g31506),.A(g4793),.B(g29540));
  NOR2 NOR2_64(.VSS(VSS),.VDD(VDD),.Y(g15071),.A(g6831),.B(g13416));
  NOR2 NOR2_65(.VSS(VSS),.VDD(VDD),.Y(g15147),.A(g13716),.B(g12892));
  NOR3 NOR3_8(.VSS(VSS),.VDD(VDD),.Y(g15754),.A(g341),.B(g7440),.C(g13385));
  NOR2 NOR2_66(.VSS(VSS),.VDD(VDD),.Y(g14037),.A(g8748),.B(g11083));
  NOR2 NOR2_67(.VSS(VSS),.VDD(VDD),.Y(g15825),.A(g7666),.B(g13217));
  NOR2 NOR2_68(.VSS(VSS),.VDD(VDD),.Y(g16044),.A(g10961),.B(g13861));
  NOR2 NOR2_69(.VSS(VSS),.VDD(VDD),.Y(g27720),.A(g9253),.B(g25791));
  NOR2 NOR2_70(.VSS(VSS),.VDD(VDD),.Y(g14419),.A(g12152),.B(g9546));
  NOR2 NOR2_71(.VSS(VSS),.VDD(VDD),.Y(g29012),.A(g5863),.B(g28020));
  NOR2 NOR2_72(.VSS(VSS),.VDD(VDD),.Y(g15151),.A(g13745),.B(g7027));
  NOR2 NOR2_73(.VSS(VSS),.VDD(VDD),.Y(g14418),.A(g12151),.B(g9594));
  NOR2 NOR2_74(.VSS(VSS),.VDD(VDD),.Y(g10266),.A(g5188),.B(g5180));
  NOR2 NOR2_75(.VSS(VSS),.VDD(VDD),.Y(g25958),.A(g7779),.B(g24609));
  NOR3 NOR3_9(.VSS(VSS),.VDD(VDD),.Y(g32296),.A(g9044),.B(g31509),.C(g12259));
  NOR2 NOR2_76(.VSS(VSS),.VDD(VDD),.Y(g31491),.A(g8938),.B(g29725));
  NOR2 NOR2_77(.VSS(VSS),.VDD(VDD),.Y(g11280),.A(g8647),.B(g3408));
  NOR2 NOR2_78(.VSS(VSS),.VDD(VDD),.Y(g25944),.A(g7716),.B(g24591));
  NOR2 NOR2_79(.VSS(VSS),.VDD(VDD),.Y(g29359),.A(g7528),.B(g28167));
  NOR2 NOR2_80(.VSS(VSS),.VDD(VDD),.Y(g12806),.A(g9472),.B(g9407));
  NOR2 NOR2_81(.VSS(VSS),.VDD(VDD),.Y(g14194),.A(g5029),.B(g10515));
  NOR2 NOR2_82(.VSS(VSS),.VDD(VDD),.Y(g19413),.A(g17151),.B(g14221));
  NOR3 NOR3_10(.VSS(VSS),.VDD(VDD),.Y(g24953),.A(g10262),.B(g23978),.C(g12259));
  NOR2 NOR2_83(.VSS(VSS),.VDD(VDD),.Y(g15059),.A(g12839),.B(g13350));
  NOR2 NOR2_84(.VSS(VSS),.VDD(VDD),.Y(g26298),.A(g8297),.B(g24825));
  NOR2 NOR2_85(.VSS(VSS),.VDD(VDD),.Y(g30129),.A(g28739),.B(g14537));
  NOR2 NOR2_86(.VSS(VSS),.VDD(VDD),.Y(g15058),.A(g12838),.B(g13350));
  NOR3 NOR3_11(.VSS(VSS),.VDD(VDD),.Y(g11231),.A(g7928),.B(g4801),.C(g4793));
  NOR2 NOR2_87(.VSS(VSS),.VDD(VDD),.Y(g17284),.A(g9253),.B(g14317));
  NOR2 NOR2_88(.VSS(VSS),.VDD(VDD),.Y(g12193),.A(g2342),.B(g8316));
  NOR2 NOR2_89(.VSS(VSS),.VDD(VDD),.Y(g11885),.A(g7153),.B(g7167));
  NOR3 NOR3_12(.VSS(VSS),.VDD(VDD),.Y(g29173),.A(g9259),.B(g27999),.C(g7704));
  NOR2 NOR2_90(.VSS(VSS),.VDD(VDD),.Y(g14313),.A(g12016),.B(g9250));
  NOR2 NOR2_91(.VSS(VSS),.VDD(VDD),.Y(g28476),.A(g27627),.B(g26547));
  NOR2 NOR2_92(.VSS(VSS),.VDD(VDD),.Y(g16226),.A(g8052),.B(g13545));
  NOR2 NOR2_93(.VSS(VSS),.VDD(VDD),.Y(g11763),.A(g3881),.B(g8172));
  NOR2 NOR2_94(.VSS(VSS),.VDD(VDD),.Y(g25504),.A(g22550),.B(g7222));
  NOR2 NOR2_95(.VSS(VSS),.VDD(VDD),.Y(g15120),.A(g12873),.B(g13605));
  NOR3 NOR3_13(.VSS(VSS),.VDD(VDD),.Y(g32910),.A(g31327),.B(I30468),.C(I30469));
  NOR2 NOR2_96(.VSS(VSS),.VDD(VDD),.Y(g25317),.A(g9766),.B(g23782));
  NOR2 NOR2_97(.VSS(VSS),.VDD(VDD),.Y(g10808),.A(g8509),.B(g7611));
  NOR2 NOR2_98(.VSS(VSS),.VDD(VDD),.Y(g15146),.A(g13716),.B(g7003));
  NOR2 NOR2_99(.VSS(VSS),.VDD(VDD),.Y(g14036),.A(g8725),.B(g11083));
  NOR2 NOR2_100(.VSS(VSS),.VDD(VDD),.Y(g34737),.A(g34706),.B(g30003));
  NOR2 NOR2_101(.VSS(VSS),.VDD(VDD),.Y(g12437),.A(g2319),.B(g8267));
  NOR2 NOR2_102(.VSS(VSS),.VDD(VDD),.Y(g27703),.A(g9607),.B(g25791));
  NOR2 NOR2_103(.VSS(VSS),.VDD(VDD),.Y(g20000),.A(g13661),.B(g16264));
  NOR2 NOR2_104(.VSS(VSS),.VDD(VDD),.Y(g13480),.A(g3017),.B(g11858));
  NOR2 NOR2_105(.VSS(VSS),.VDD(VDD),.Y(g14642),.A(g12374),.B(g9829));
  NOR2 NOR2_106(.VSS(VSS),.VDD(VDD),.Y(g12347),.A(g9321),.B(g9274));
  NOR2 NOR2_107(.VSS(VSS),.VDD(VDD),.Y(g14064),.A(g9214),.B(g12259));
  NOR2 NOR2_108(.VSS(VSS),.VDD(VDD),.Y(g13076),.A(g7443),.B(g10741));
  NOR2 NOR2_109(.VSS(VSS),.VDD(VDD),.Y(g33098),.A(g31997),.B(g4616));
  NOR3 NOR3_14(.VSS(VSS),.VDD(VDD),.Y(g28519),.A(g8011),.B(g27602),.C(g10295));
  NOR4 NOR4_2(.VSS(VSS),.VDD(VDD),.Y(g12821),.A(g7132),.B(g10223),.C(g7149),.D(g10261));
  NOR2 NOR2_110(.VSS(VSS),.VDD(VDD),.Y(g27063),.A(g26485),.B(g26516));
  NOR2 NOR2_111(.VSS(VSS),.VDD(VDD),.Y(g24751),.A(g3034),.B(g23105));
  NOR2 NOR2_112(.VSS(VSS),.VDD(VDD),.Y(g29903),.A(g6928),.B(g28484));
  NOR2 NOR2_113(.VSS(VSS),.VDD(VDD),.Y(g11773),.A(g8883),.B(g4785));
  NOR2 NOR2_114(.VSS(VSS),.VDD(VDD),.Y(g27516),.A(g9180),.B(g26657));
  NOR2 NOR2_115(.VSS(VSS),.VDD(VDD),.Y(g33140),.A(g7693),.B(g32072));
  NOR2 NOR2_116(.VSS(VSS),.VDD(VDD),.Y(g13341),.A(g7863),.B(g10762));
  NOR2 NOR2_117(.VSS(VSS),.VDD(VDD),.Y(g12137),.A(g6682),.B(g7097));
  NOR2 NOR2_118(.VSS(VSS),.VDD(VDD),.Y(g13670),.A(g8123),.B(g10756));
  NOR3 NOR3_15(.VSS(VSS),.VDD(VDD),.Y(g10555),.A(g7227),.B(g4601),.C(g4608));
  NOR2 NOR2_119(.VSS(VSS),.VDD(VDD),.Y(g20841),.A(g17847),.B(g12027));
  NOR3 NOR3_16(.VSS(VSS),.VDD(VDD),.Y(g23042),.A(g16581),.B(g19462),.C(g10685));
  NOR2 NOR2_120(.VSS(VSS),.VDD(VDD),.Y(g14712),.A(g12479),.B(g9971));
  NOR2 NOR2_121(.VSS(VSS),.VDD(VDD),.Y(g13335),.A(g7851),.B(g10741));
  NOR2 NOR2_122(.VSS(VSS),.VDD(VDD),.Y(g19890),.A(g16987),.B(g8058));
  NOR2 NOR2_123(.VSS(VSS),.VDD(VDD),.Y(g14914),.A(g12822),.B(g12797));
  NOR2 NOR2_124(.VSS(VSS),.VDD(VDD),.Y(g24391),.A(g22190),.B(g14645));
  NOR2 NOR2_125(.VSS(VSS),.VDD(VDD),.Y(g15127),.A(g12879),.B(g13605));
  NOR2 NOR2_126(.VSS(VSS),.VDD(VDD),.Y(g30271),.A(g7041),.B(g29008));
  NOR2 NOR2_127(.VSS(VSS),.VDD(VDD),.Y(g23124),.A(g8443),.B(g20011));
  NOR2 NOR2_128(.VSS(VSS),.VDD(VDD),.Y(g23678),.A(g9809),.B(g21190));
  NOR2 NOR2_129(.VSS(VSS),.VDD(VDD),.Y(g16024),.A(g14216),.B(g11890));
  NOR2 NOR2_130(.VSS(VSS),.VDD(VDD),.Y(g12208),.A(g10096),.B(g5759));
  NOR2 NOR2_131(.VSS(VSS),.VDD(VDD),.Y(g33447),.A(g31978),.B(g7643));
  NOR2 NOR2_132(.VSS(VSS),.VDD(VDD),.Y(g26330),.A(g8631),.B(g24825));
  NOR2 NOR2_133(.VSS(VSS),.VDD(VDD),.Y(g23686),.A(g2767),.B(g21066));
  NOR2 NOR2_134(.VSS(VSS),.VDD(VDD),.Y(g20014),.A(g17096),.B(g11244));
  NOR2 NOR2_135(.VSS(VSS),.VDD(VDD),.Y(g33162),.A(g4859),.B(g32072));
  NOR2 NOR2_136(.VSS(VSS),.VDD(VDD),.Y(g29898),.A(g6895),.B(g28458));
  NOR2 NOR2_137(.VSS(VSS),.VDD(VDD),.Y(g12453),.A(g9444),.B(g5527));
  NOR2 NOR2_138(.VSS(VSS),.VDD(VDD),.Y(g15095),.A(g13177),.B(g12866));
  NOR2 NOR2_139(.VSS(VSS),.VDD(VDD),.Y(g29191),.A(g7738),.B(g28010));
  NOR2 NOR2_140(.VSS(VSS),.VDD(VDD),.Y(g19778),.A(g16268),.B(g1061));
  NOR2 NOR2_141(.VSS(VSS),.VDD(VDD),.Y(g11618),.A(g8114),.B(g8070));
  NOR2 NOR2_142(.VSS(VSS),.VDD(VDD),.Y(g14382),.A(g9390),.B(g11139));
  NOR2 NOR2_143(.VSS(VSS),.VDD(VDD),.Y(g14176),.A(g9044),.B(g12259));
  NOR2 NOR2_144(.VSS(VSS),.VDD(VDD),.Y(g14092),.A(g8774),.B(g11083));
  NOR2 NOR2_145(.VSS(VSS),.VDD(VDD),.Y(g19999),.A(g16232),.B(g13742));
  NOR2 NOR2_146(.VSS(VSS),.VDD(VDD),.Y(g22400),.A(g19345),.B(g15718));
  NOR2 NOR2_147(.VSS(VSS),.VDD(VDD),.Y(g20720),.A(g17847),.B(g9299));
  NOR3 NOR3_17(.VSS(VSS),.VDD(VDD),.Y(g11469),.A(g650),.B(g9903),.C(g645));
  NOR2 NOR2_148(.VSS(VSS),.VDD(VDD),.Y(g12593),.A(g9234),.B(g5164));
  NOR2 NOR2_149(.VSS(VSS),.VDD(VDD),.Y(g12346),.A(g9931),.B(g9933));
  NOR3 NOR3_18(.VSS(VSS),.VDD(VDD),.Y(g24720),.A(g1322),.B(g23051),.C(g19793));
  NOR2 NOR2_150(.VSS(VSS),.VDD(VDD),.Y(g11039),.A(g9056),.B(g9092));
  NOR2 NOR2_151(.VSS(VSS),.VDD(VDD),.Y(g11306),.A(g3412),.B(g8647));
  NOR2 NOR2_152(.VSS(VSS),.VDD(VDD),.Y(g30132),.A(g28789),.B(g7362));
  NOR2 NOR2_153(.VSS(VSS),.VDD(VDD),.Y(g22539),.A(g1030),.B(g19699));
  NOR2 NOR2_154(.VSS(VSS),.VDD(VDD),.Y(g8958),.A(g3881),.B(g3873));
  NOR2 NOR2_155(.VSS(VSS),.VDD(VDD),.Y(g33147),.A(g32090),.B(g7788));
  NOR2 NOR2_156(.VSS(VSS),.VDD(VDD),.Y(g9061),.A(g3401),.B(g3361));
  NOR2 NOR2_157(.VSS(VSS),.VDD(VDD),.Y(g19932),.A(g3376),.B(g16296));
  NOR2 NOR2_158(.VSS(VSS),.VDD(VDD),.Y(g25887),.A(g24984),.B(g11706));
  NOR2 NOR2_159(.VSS(VSS),.VDD(VDD),.Y(g15089),.A(g13144),.B(g12861));
  NOR2 NOR2_160(.VSS(VSS),.VDD(VDD),.Y(g15088),.A(g13144),.B(g6874));
  NOR3 NOR3_19(.VSS(VSS),.VDD(VDD),.Y(g13937),.A(g8883),.B(g4785),.C(g11155));
  NOR3 NOR3_20(.VSS(VSS),.VDD(VDD),.Y(g21277),.A(g9417),.B(g9340),.C(g17467));
  NOR2 NOR2_161(.VSS(VSS),.VDD(VDD),.Y(g29032),.A(g9300),.B(g27999));
  NOR2 NOR2_162(.VSS(VSS),.VDD(VDD),.Y(g15126),.A(g12878),.B(g13605));
  NOR2 NOR2_163(.VSS(VSS),.VDD(VDD),.Y(g11666),.A(g8172),.B(g8125));
  NOR2 NOR2_164(.VSS(VSS),.VDD(VDD),.Y(g16581),.A(g13756),.B(g8086));
  NOR2 NOR2_165(.VSS(VSS),.VDD(VDD),.Y(g11363),.A(g8626),.B(g8751));
  NOR2 NOR2_166(.VSS(VSS),.VDD(VDD),.Y(g11217),.A(g8531),.B(g6875));
  NOR2 NOR2_167(.VSS(VSS),.VDD(VDD),.Y(g31318),.A(g4785),.B(g29697));
  NOR2 NOR2_168(.VSS(VSS),.VDD(VDD),.Y(g12711),.A(g6209),.B(g9326));
  NOR3 NOR3_21(.VSS(VSS),.VDD(VDD),.Y(g8177),.A(g4966),.B(g4991),.C(g4983));
  NOR2 NOR2_169(.VSS(VSS),.VDD(VDD),.Y(g30171),.A(g28880),.B(g7431));
  NOR2 NOR2_170(.VSS(VSS),.VDD(VDD),.Y(g17515),.A(g13221),.B(g10828));
  NOR2 NOR2_171(.VSS(VSS),.VDD(VDD),.Y(g15060),.A(g13350),.B(g6814));
  NOR3 NOR3_22(.VSS(VSS),.VDD(VDD),.Y(g12492),.A(g7704),.B(g5170),.C(g5164));
  NOR2 NOR2_172(.VSS(VSS),.VDD(VDD),.Y(g26545),.A(g24881),.B(g24855));
  NOR2 NOR2_173(.VSS(VSS),.VDD(VDD),.Y(g27982),.A(g7212),.B(g25856));
  NOR2 NOR2_174(.VSS(VSS),.VDD(VDD),.Y(g27381),.A(g8075),.B(g26657));
  NOR2 NOR2_175(.VSS(VSS),.VDD(VDD),.Y(g14415),.A(g12147),.B(g9590));
  NOR2 NOR2_176(.VSS(VSS),.VDD(VDD),.Y(g13110),.A(g7841),.B(g10741));
  NOR3 NOR3_23(.VSS(VSS),.VDD(VDD),.Y(g26598),.A(g8990),.B(g13756),.C(g24732));
  NOR2 NOR2_177(.VSS(VSS),.VDD(VDD),.Y(g33146),.A(g4669),.B(g32057));
  NOR2 NOR2_178(.VSS(VSS),.VDD(VDD),.Y(g29071),.A(g5873),.B(g28020));
  NOR2 NOR2_179(.VSS(VSS),.VDD(VDD),.Y(g29370),.A(g28585),.B(g28599));
  NOR2 NOR2_180(.VSS(VSS),.VDD(VDD),.Y(g33427),.A(g10278),.B(g31950));
  NOR2 NOR2_181(.VSS(VSS),.VDD(VDD),.Y(g22399),.A(g1367),.B(g19720));
  NOR2 NOR2_182(.VSS(VSS),.VDD(VDD),.Y(g10312),.A(g5881),.B(g5873));
  NOR2 NOR2_183(.VSS(VSS),.VDD(VDD),.Y(g15055),.A(g6808),.B(g13350));
  NOR2 NOR2_184(.VSS(VSS),.VDD(VDD),.Y(g15070),.A(g6829),.B(g13416));
  NOR2 NOR2_185(.VSS(VSS),.VDD(VDD),.Y(g30159),.A(g28799),.B(g14589));
  NOR2 NOR2_186(.VSS(VSS),.VDD(VDD),.Y(g23560),.A(g9607),.B(g20838));
  NOR2 NOR2_187(.VSS(VSS),.VDD(VDD),.Y(g12483),.A(g2453),.B(g8324));
  NOR2 NOR2_188(.VSS(VSS),.VDD(VDD),.Y(g11216),.A(g7998),.B(g8037));
  NOR2 NOR2_189(.VSS(VSS),.VDD(VDD),.Y(g10799),.A(g347),.B(g7541));
  NOR2 NOR2_190(.VSS(VSS),.VDD(VDD),.Y(g12553),.A(g5170),.B(g9206));
  NOR2 NOR2_191(.VSS(VSS),.VDD(VDD),.Y(g23642),.A(g9733),.B(g21124));
  NOR2 NOR2_192(.VSS(VSS),.VDD(VDD),.Y(g15067),.A(g12842),.B(g13394));
  NOR2 NOR2_193(.VSS(VSS),.VDD(VDD),.Y(g15094),.A(g13177),.B(g12865));
  NOR2 NOR2_194(.VSS(VSS),.VDD(VDD),.Y(g30144),.A(g28789),.B(g7322));
  NOR2 NOR2_195(.VSS(VSS),.VDD(VDD),.Y(g24453),.A(g7446),.B(g22325));
  NOR2 NOR2_196(.VSS(VSS),.VDD(VDD),.Y(g15150),.A(g12895),.B(g13745));
  NOR2 NOR2_197(.VSS(VSS),.VDD(VDD),.Y(g31127),.A(g4966),.B(g29556));
  NOR3 NOR3_24(.VSS(VSS),.VDD(VDD),.Y(g13908),.A(g4709),.B(g8796),.C(g11155));
  NOR2 NOR2_198(.VSS(VSS),.VDD(VDD),.Y(g12252),.A(g9995),.B(g10185));
  NOR2 NOR2_199(.VSS(VSS),.VDD(VDD),.Y(g26309),.A(g8575),.B(g24825));
  NOR2 NOR2_200(.VSS(VSS),.VDD(VDD),.Y(g11747),.A(g3530),.B(g8114));
  NOR2 NOR2_201(.VSS(VSS),.VDD(VDD),.Y(g13568),.A(g8046),.B(g12527));
  NOR2 NOR2_202(.VSS(VSS),.VDD(VDD),.Y(g16066),.A(g10929),.B(g13307));
  NOR2 NOR2_203(.VSS(VSS),.VDD(VDD),.Y(g16231),.A(g13515),.B(g4771));
  NOR2 NOR2_204(.VSS(VSS),.VDD(VDD),.Y(g33103),.A(g32176),.B(g31212));
  NOR2 NOR2_205(.VSS(VSS),.VDD(VDD),.Y(g19793),.A(g16292),.B(g1404));
  NOR2 NOR2_206(.VSS(VSS),.VDD(VDD),.Y(g33095),.A(g31997),.B(g7236));
  NOR2 NOR2_207(.VSS(VSS),.VDD(VDD),.Y(g12847),.A(g6838),.B(g10430));
  NOR2 NOR2_208(.VSS(VSS),.VDD(VDD),.Y(g25144),.A(g5046),.B(g23623));
  NOR2 NOR2_209(.VSS(VSS),.VDD(VDD),.Y(g13772),.A(g3990),.B(g11702));
  NOR2 NOR2_210(.VSS(VSS),.VDD(VDD),.Y(g28515),.A(g3881),.B(g27635));
  NOR2 NOR2_211(.VSS(VSS),.VDD(VDD),.Y(g28414),.A(g27467),.B(g26347));
  NOR2 NOR2_212(.VSS(VSS),.VDD(VDD),.Y(g30288),.A(g7087),.B(g29073));
  NOR2 NOR2_213(.VSS(VSS),.VDD(VDD),.Y(g26976),.A(g5016),.B(g25791));
  NOR2 NOR2_214(.VSS(VSS),.VDD(VDD),.Y(g29146),.A(g6565),.B(g26994));
  NOR2 NOR2_215(.VSS(VSS),.VDD(VDD),.Y(g12851),.A(g6846),.B(g10430));
  NOR2 NOR2_216(.VSS(VSS),.VDD(VDD),.Y(g14539),.A(g11977),.B(g9833));
  NOR2 NOR2_217(.VSS(VSS),.VDD(VDD),.Y(g9649),.A(g2227),.B(g2153));
  NOR2 NOR2_218(.VSS(VSS),.VDD(VDD),.Y(g14538),.A(g11973),.B(g9828));
  NOR2 NOR2_219(.VSS(VSS),.VDD(VDD),.Y(g28584),.A(g7121),.B(g27635));
  NOR2 NOR2_220(.VSS(VSS),.VDD(VDD),.Y(g16287),.A(g13622),.B(g11144));
  NOR2 NOR2_221(.VSS(VSS),.VDD(VDD),.Y(g33089),.A(g31978),.B(g4322));
  NOR2 NOR2_222(.VSS(VSS),.VDD(VDD),.Y(g15102),.A(g14591),.B(g6954));
  NOR2 NOR2_223(.VSS(VSS),.VDD(VDD),.Y(g15157),.A(g13782),.B(g12900));
  NOR2 NOR2_224(.VSS(VSS),.VDD(VDD),.Y(g33088),.A(g31997),.B(g7224));
  NOR2 NOR2_225(.VSS(VSS),.VDD(VDD),.Y(g22514),.A(g19699),.B(g1018));
  NOR2 NOR2_226(.VSS(VSS),.VDD(VDD),.Y(g12311),.A(g6109),.B(g10136));
  NOR2 NOR2_227(.VSS(VSS),.VDD(VDD),.Y(g15066),.A(g12841),.B(g13394));
  NOR2 NOR2_228(.VSS(VSS),.VDD(VDD),.Y(g24575),.A(g23498),.B(g23514));
  NOR2 NOR2_229(.VSS(VSS),.VDD(VDD),.Y(g30260),.A(g7018),.B(g28982));
  NOR2 NOR2_230(.VSS(VSS),.VDD(VDD),.Y(g23883),.A(g2779),.B(g21067));
  NOR2 NOR2_231(.VSS(VSS),.VDD(VDD),.Y(g26865),.A(g25328),.B(g25290));
  NOR2 NOR2_232(.VSS(VSS),.VDD(VDD),.Y(g31126),.A(g7928),.B(g29540));
  NOR2 NOR2_233(.VSS(VSS),.VDD(VDD),.Y(g16268),.A(g7913),.B(g13121));
  NOR2 NOR2_234(.VSS(VSS),.VDD(VDD),.Y(g12780),.A(g9402),.B(g9326));
  NOR2 NOR2_235(.VSS(VSS),.VDD(VDD),.Y(g14515),.A(g12225),.B(g9761));
  NOR2 NOR2_236(.VSS(VSS),.VDD(VDD),.Y(g14414),.A(g12145),.B(g9639));
  NOR2 NOR2_237(.VSS(VSS),.VDD(VDD),.Y(g11493),.A(g8964),.B(g8967));
  NOR2 NOR2_238(.VSS(VSS),.VDD(VDD),.Y(g25954),.A(g7750),.B(g24591));
  NOR2 NOR2_239(.VSS(VSS),.VDD(VDD),.Y(g23729),.A(g17482),.B(g21206));
  NOR2 NOR2_240(.VSS(VSS),.VDD(VDD),.Y(g20982),.A(g17929),.B(g12065));
  NOR2 NOR2_241(.VSS(VSS),.VDD(VDD),.Y(g19880),.A(g16201),.B(g13634));
  NOR2 NOR2_242(.VSS(VSS),.VDD(VDD),.Y(g27731),.A(g9229),.B(g25791));
  NOR2 NOR2_243(.VSS(VSS),.VDD(VDD),.Y(g12846),.A(g6837),.B(g10430));
  NOR2 NOR2_244(.VSS(VSS),.VDD(VDD),.Y(g22535),.A(g19699),.B(g1030));
  NOR2 NOR2_245(.VSS(VSS),.VDD(VDD),.Y(g13806),.A(g11245),.B(g4076));
  NOR2 NOR2_246(.VSS(VSS),.VDD(VDD),.Y(g29889),.A(g6905),.B(g28471));
  NOR2 NOR2_247(.VSS(VSS),.VDD(VDD),.Y(g26686),.A(g23678),.B(g25189));
  NOR2 NOR2_248(.VSS(VSS),.VDD(VDD),.Y(g13517),.A(g8541),.B(g12692));
  NOR2 NOR2_249(.VSS(VSS),.VDD(VDD),.Y(g20390),.A(g17182),.B(g14257));
  NOR2 NOR2_250(.VSS(VSS),.VDD(VDD),.Y(g29181),.A(g6573),.B(g26994));
  NOR2 NOR2_251(.VSS(VSS),.VDD(VDD),.Y(g21284),.A(g16646),.B(g9690));
  NOR2 NOR2_252(.VSS(VSS),.VDD(VDD),.Y(g26267),.A(g8033),.B(g24732));
  NOR2 NOR2_253(.VSS(VSS),.VDD(VDD),.Y(g12405),.A(g9374),.B(g5180));
  NOR2 NOR2_254(.VSS(VSS),.VDD(VDD),.Y(g16210),.A(g13479),.B(g4894));
  NOR2 NOR2_255(.VSS(VSS),.VDD(VDD),.Y(g15054),.A(g12837),.B(g13350));
  NOR2 NOR2_256(.VSS(VSS),.VDD(VDD),.Y(g27046),.A(g7544),.B(g25888));
  NOR2 NOR2_257(.VSS(VSS),.VDD(VDD),.Y(g15156),.A(g13782),.B(g7050));
  NOR2 NOR2_258(.VSS(VSS),.VDD(VDD),.Y(g30294),.A(g7110),.B(g29110));
  NOR2 NOR2_259(.VSS(VSS),.VDD(VDD),.Y(g12046),.A(g10036),.B(g9640));
  NOR2 NOR2_260(.VSS(VSS),.VDD(VDD),.Y(g14399),.A(g5297),.B(g12598));
  NOR2 NOR2_261(.VSS(VSS),.VDD(VDD),.Y(g11006),.A(g7686),.B(g7836));
  NOR2 NOR2_262(.VSS(VSS),.VDD(VDD),.Y(g12113),.A(g1648),.B(g8187));
  NOR2 NOR2_263(.VSS(VSS),.VDD(VDD),.Y(g28106),.A(g7812),.B(g26994));
  NOR2 NOR2_264(.VSS(VSS),.VDD(VDD),.Y(g25189),.A(g6082),.B(g23726));
  NOR2 NOR2_265(.VSS(VSS),.VDD(VDD),.Y(g27827),.A(g9456),.B(g25839));
  NOR2 NOR2_266(.VSS(VSS),.VDD(VDD),.Y(g9586),.A(g1668),.B(g1592));
  NOR2 NOR2_267(.VSS(VSS),.VDD(VDD),.Y(g19887),.A(g3025),.B(g16275));
  NOR2 NOR2_268(.VSS(VSS),.VDD(VDD),.Y(g29497),.A(g22763),.B(g28241));
  NOR2 NOR2_269(.VSS(VSS),.VDD(VDD),.Y(g27769),.A(g9434),.B(g25805));
  NOR2 NOR2_270(.VSS(VSS),.VDD(VDD),.Y(g15131),.A(g12881),.B(g13638));
  NOR2 NOR2_271(.VSS(VSS),.VDD(VDD),.Y(g27768),.A(g9264),.B(g25805));
  NOR2 NOR2_272(.VSS(VSS),.VDD(VDD),.Y(g30160),.A(g28846),.B(g7387));
  NOR2 NOR2_273(.VSS(VSS),.VDD(VDD),.Y(g33094),.A(g31950),.B(g4639));
  NOR2 NOR2_274(.VSS(VSS),.VDD(VDD),.Y(g14361),.A(g12079),.B(g9413));
  NOR2 NOR2_275(.VSS(VSS),.VDD(VDD),.Y(g20183),.A(g17152),.B(g14222));
  NOR2 NOR2_276(.VSS(VSS),.VDD(VDD),.Y(g28514),.A(g8165),.B(g27617));
  NOR2 NOR2_277(.VSS(VSS),.VDD(VDD),.Y(g22491),.A(g1361),.B(g19720));
  NOR2 NOR2_278(.VSS(VSS),.VDD(VDD),.Y(g16479),.A(g14719),.B(g12490));
  NOR2 NOR2_279(.VSS(VSS),.VDD(VDD),.Y(g27027),.A(g26398),.B(g26484));
  NOR2 NOR2_280(.VSS(VSS),.VDD(VDD),.Y(g24508),.A(g23577),.B(g23618));
  NOR2 NOR2_281(.VSS(VSS),.VDD(VDD),.Y(g23052),.A(g8334),.B(g19916));
  NOR2 NOR2_282(.VSS(VSS),.VDD(VDD),.Y(g12662),.A(g5863),.B(g9274));
  NOR2 NOR2_283(.VSS(VSS),.VDD(VDD),.Y(g25160),.A(g5390),.B(g23659));
  NOR2 NOR2_284(.VSS(VSS),.VDD(VDD),.Y(g12249),.A(g5763),.B(g10096));
  NOR2 NOR2_285(.VSS(VSS),.VDD(VDD),.Y(g11834),.A(g8938),.B(g8822));
  NOR2 NOR2_286(.VSS(VSS),.VDD(VDD),.Y(g12204),.A(g9927),.B(g10160));
  NOR2 NOR2_287(.VSS(VSS),.VDD(VDD),.Y(g15143),.A(g6998),.B(g13680));
  NOR2 NOR2_288(.VSS(VSS),.VDD(VDD),.Y(g30170),.A(g28846),.B(g14615));
  NOR2 NOR2_289(.VSS(VSS),.VDD(VDD),.Y(g29503),.A(g22763),.B(g28250));
  NOR2 NOR2_290(.VSS(VSS),.VDD(VDD),.Y(g14033),.A(g8808),.B(g12259));
  NOR2 NOR2_291(.VSS(VSS),.VDD(VDD),.Y(g12081),.A(g10079),.B(g9694));
  NOR2 NOR2_292(.VSS(VSS),.VDD(VDD),.Y(g13021),.A(g7544),.B(g10741));
  NOR2 NOR2_293(.VSS(VSS),.VDD(VDD),.Y(g22521),.A(g1036),.B(g19699));
  NOR2 NOR2_294(.VSS(VSS),.VDD(VDD),.Y(g27647),.A(g3004),.B(g26616));
  NOR2 NOR2_295(.VSS(VSS),.VDD(VDD),.Y(g11913),.A(g7197),.B(g9166));
  NOR2 NOR2_296(.VSS(VSS),.VDD(VDD),.Y(g13913),.A(g8859),.B(g11083));
  NOR2 NOR2_297(.VSS(VSS),.VDD(VDD),.Y(g27356),.A(g9429),.B(g26657));
  NOR2 NOR2_298(.VSS(VSS),.VDD(VDD),.Y(g7601),.A(g1322),.B(g1333));
  NOR2 NOR2_299(.VSS(VSS),.VDD(VDD),.Y(g15168),.A(g13835),.B(g12909));
  NOR2 NOR2_300(.VSS(VSS),.VDD(VDD),.Y(g27826),.A(g9501),.B(g25821));
  NOR2 NOR2_301(.VSS(VSS),.VDD(VDD),.Y(g29910),.A(g3990),.B(g28484));
  NOR3 NOR3_25(.VSS(VSS),.VDD(VDD),.Y(g11607),.A(g8848),.B(g8993),.C(g376));
  NOR2 NOR2_302(.VSS(VSS),.VDD(VDD),.Y(g14514),.A(g11959),.B(g9760));
  NOR2 NOR2_303(.VSS(VSS),.VDD(VDD),.Y(g11346),.A(g7980),.B(g7964));
  NOR3 NOR3_26(.VSS(VSS),.VDD(VDD),.Y(g29070),.A(g5857),.B(g7766),.C(g28020));
  NOR2 NOR2_304(.VSS(VSS),.VDD(VDD),.Y(g12651),.A(g9269),.B(g5511));
  NOR2 NOR2_305(.VSS(VSS),.VDD(VDD),.Y(g10421),.A(g6227),.B(g9518));
  NOR2 NOR2_306(.VSS(VSS),.VDD(VDD),.Y(g30119),.A(g28761),.B(g7315));
  NOR2 NOR2_307(.VSS(VSS),.VDD(VDD),.Y(g14163),.A(g8997),.B(g12259));
  NOR2 NOR2_308(.VSS(VSS),.VDD(VDD),.Y(g11797),.A(g8883),.B(g8796));
  NOR2 NOR2_309(.VSS(VSS),.VDD(VDD),.Y(g19919),.A(g16987),.B(g11205));
  NOR2 NOR2_310(.VSS(VSS),.VDD(VDD),.Y(g30276),.A(g7074),.B(g29073));
  NOR2 NOR2_311(.VSS(VSS),.VDD(VDD),.Y(g30285),.A(g7097),.B(g29110));
  NOR2 NOR2_312(.VSS(VSS),.VDD(VDD),.Y(g19444),.A(g17192),.B(g14295));
  NOR2 NOR2_313(.VSS(VSS),.VDD(VDD),.Y(g12505),.A(g9444),.B(g9381));
  NOR2 NOR2_314(.VSS(VSS),.VDD(VDD),.Y(g27717),.A(g9492),.B(g26745));
  NOR2 NOR2_315(.VSS(VSS),.VDD(VDD),.Y(g9100),.A(g3752),.B(g3712));
  NOR2 NOR2_316(.VSS(VSS),.VDD(VDD),.Y(g12026),.A(g9417),.B(g9340));
  NOR2 NOR2_317(.VSS(VSS),.VDD(VDD),.Y(g8984),.A(g4899),.B(g4975));
  NOR2 NOR2_318(.VSS(VSS),.VDD(VDD),.Y(g14121),.A(g8891),.B(g12259));
  NOR2 NOR2_319(.VSS(VSS),.VDD(VDD),.Y(g25022),.A(g714),.B(g23324));
  NOR2 NOR2_320(.VSS(VSS),.VDD(VDD),.Y(g11891),.A(g812),.B(g9166));
  NOR2 NOR2_321(.VSS(VSS),.VDD(VDD),.Y(g16242),.A(g13529),.B(g4961));
  NOR2 NOR2_322(.VSS(VSS),.VDD(VDD),.Y(g28491),.A(g8114),.B(g27617));
  NOR2 NOR2_323(.VSS(VSS),.VDD(VDD),.Y(g33085),.A(g31978),.B(g4311));
  NOR2 NOR2_324(.VSS(VSS),.VDD(VDD),.Y(g14291),.A(g9839),.B(g12155));
  NOR2 NOR2_325(.VSS(VSS),.VDD(VDD),.Y(g11537),.A(g8229),.B(g3873));
  NOR2 NOR2_326(.VSS(VSS),.VDD(VDD),.Y(g27343),.A(g8005),.B(g26616));
  NOR2 NOR2_327(.VSS(VSS),.VDD(VDD),.Y(g28981),.A(g9234),.B(g27999));
  NOR2 NOR2_328(.VSS(VSS),.VDD(VDD),.Y(g29077),.A(g6555),.B(g26994));
  NOR2 NOR2_329(.VSS(VSS),.VDD(VDD),.Y(g12646),.A(g9234),.B(g9206));
  NOR3 NOR3_27(.VSS(VSS),.VDD(VDD),.Y(g11283),.A(g7953),.B(g4991),.C(g9064));
  NOR2 NOR2_330(.VSS(VSS),.VDD(VDD),.Y(g10760),.A(g1046),.B(g7479));
  NOR2 NOR2_331(.VSS(VSS),.VDD(VDD),.Y(g11303),.A(g8497),.B(g8500));
  NOR2 NOR2_332(.VSS(VSS),.VDD(VDD),.Y(g31942),.A(g8977),.B(g30583));
  NOR2 NOR2_333(.VSS(VSS),.VDD(VDD),.Y(g27368),.A(g8119),.B(g26657));
  NOR2 NOR2_334(.VSS(VSS),.VDD(VDD),.Y(g21206),.A(g6419),.B(g17396));
  NOR2 NOR2_335(.VSS(VSS),.VDD(VDD),.Y(g12850),.A(g10430),.B(g6845));
  NOR2 NOR2_336(.VSS(VSS),.VDD(VDD),.Y(g13796),.A(g9158),.B(g12527));
  NOR2 NOR2_337(.VSS(VSS),.VDD(VDD),.Y(g28521),.A(g27649),.B(g26604));
  NOR2 NOR2_338(.VSS(VSS),.VDD(VDD),.Y(g31965),.A(g30583),.B(g4358));
  NOR2 NOR2_339(.VSS(VSS),.VDD(VDD),.Y(g33131),.A(g4659),.B(g32057));
  NOR4 NOR4_3(.VSS(VSS),.VDD(VDD),.Y(g12228),.A(g10222),.B(g10206),.C(g10184),.D(g10335));
  NOR2 NOR2_340(.VSS(VSS),.VDD(VDD),.Y(g10649),.A(g1183),.B(g8407));
  NOR3 NOR3_28(.VSS(VSS),.VDD(VDD),.Y(g12716),.A(g7812),.B(g6555),.C(g6549));
  NOR2 NOR2_341(.VSS(VSS),.VDD(VDD),.Y(g15123),.A(g6975),.B(g13605));
  NOR2 NOR2_342(.VSS(VSS),.VDD(VDD),.Y(g10491),.A(g6573),.B(g9576));
  NOR2 NOR2_343(.VSS(VSS),.VDD(VDD),.Y(g20027),.A(g16242),.B(g13779));
  NOR2 NOR2_344(.VSS(VSS),.VDD(VDD),.Y(g21652),.A(g17619),.B(g17663));
  NOR2 NOR2_345(.VSS(VSS),.VDD(VDD),.Y(g27379),.A(g8492),.B(g26636));
  NOR2 NOR2_346(.VSS(VSS),.VDD(VDD),.Y(g11483),.A(g8165),.B(g3522));
  NOR2 NOR2_347(.VSS(VSS),.VDD(VDD),.Y(g31469),.A(g8822),.B(g29725));
  NOR2 NOR2_348(.VSS(VSS),.VDD(VDD),.Y(g11862),.A(g7134),.B(g7150));
  NOR2 NOR2_349(.VSS(VSS),.VDD(VDD),.Y(g12050),.A(g10038),.B(g9649));
  NOR2 NOR2_350(.VSS(VSS),.VDD(VDD),.Y(g24779),.A(g3736),.B(g23167));
  NOR2 NOR2_351(.VSS(VSS),.VDD(VDD),.Y(g16237),.A(g8088),.B(g13574));
  NOR3 NOR3_29(.VSS(VSS),.VDD(VDD),.Y(g29916),.A(g8681),.B(g28504),.C(g11083));
  NOR2 NOR2_352(.VSS(VSS),.VDD(VDD),.Y(g23135),.A(g16476),.B(g19981));
  NOR2 NOR2_353(.VSS(VSS),.VDD(VDD),.Y(g15992),.A(g10929),.B(g13846));
  NOR2 NOR2_354(.VSS(VSS),.VDD(VDD),.Y(g28462),.A(g3512),.B(g27617));
  NOR2 NOR2_355(.VSS(VSS),.VDD(VDD),.Y(g13326),.A(g10929),.B(g10905));
  NOR2 NOR2_356(.VSS(VSS),.VDD(VDD),.Y(g14767),.A(g10130),.B(g12204));
  NOR2 NOR2_357(.VSS(VSS),.VDD(VDD),.Y(g14395),.A(g12118),.B(g9542));
  NOR2 NOR2_358(.VSS(VSS),.VDD(VDD),.Y(g17420),.A(g9456),.B(g14408));
  NOR2 NOR2_359(.VSS(VSS),.VDD(VDD),.Y(g10899),.A(g4064),.B(g8451));
  NOR2 NOR2_360(.VSS(VSS),.VDD(VDD),.Y(g22540),.A(g19720),.B(g1373));
  NOR2 NOR2_361(.VSS(VSS),.VDD(VDD),.Y(g11252),.A(g8620),.B(g3057));
  NOR2 NOR2_362(.VSS(VSS),.VDD(VDD),.Y(g11621),.A(g3512),.B(g7985));
  NOR2 NOR2_363(.VSS(VSS),.VDD(VDD),.Y(g15578),.A(g7216),.B(g14279));
  NOR2 NOR2_364(.VSS(VSS),.VDD(VDD),.Y(g20998),.A(g18065),.B(g9450));
  NOR2 NOR2_365(.VSS(VSS),.VDD(VDD),.Y(g33143),.A(g32293),.B(g31518));
  NOR4 NOR4_4(.VSS(VSS),.VDD(VDD),.Y(g7661),.A(g1211),.B(g1216),.C(g1221),.D(g1205));
  NOR2 NOR2_366(.VSS(VSS),.VDD(VDD),.Y(g29180),.A(g9569),.B(g26977));
  NOR2 NOR2_367(.VSS(VSS),.VDD(VDD),.Y(g14247),.A(g9934),.B(g10869));
  NOR2 NOR2_368(.VSS(VSS),.VDD(VDD),.Y(g13872),.A(g8745),.B(g11083));
  NOR2 NOR2_369(.VSS(VSS),.VDD(VDD),.Y(g25501),.A(g23918),.B(g14645));
  NOR2 NOR2_370(.VSS(VSS),.VDD(VDD),.Y(g20717),.A(g5037),.B(g17217));
  NOR2 NOR2_371(.VSS(VSS),.VDD(VDD),.Y(g14272),.A(g6411),.B(g10598));
  NOR2 NOR2_372(.VSS(VSS),.VDD(VDD),.Y(g12129),.A(g9992),.B(g7051));
  NOR2 NOR2_373(.VSS(VSS),.VDD(VDD),.Y(g12002),.A(g5297),.B(g7004));
  NOR3 NOR3_30(.VSS(VSS),.VDD(VDD),.Y(g11213),.A(g4776),.B(g7892),.C(g9030));
  NOR2 NOR2_374(.VSS(VSS),.VDD(VDD),.Y(g15142),.A(g13680),.B(g12889));
  NOR2 NOR2_375(.VSS(VSS),.VDD(VDD),.Y(g33084),.A(g31978),.B(g7655));
  NOR2 NOR2_376(.VSS(VSS),.VDD(VDD),.Y(g20149),.A(g17091),.B(g14185));
  NOR2 NOR2_377(.VSS(VSS),.VDD(VDD),.Y(g26609),.A(g146),.B(g24732));
  NOR2 NOR2_378(.VSS(VSS),.VDD(VDD),.Y(g15130),.A(g13638),.B(g6985));
  NOR2 NOR2_379(.VSS(VSS),.VDD(VDD),.Y(g24148),.A(g19268),.B(g19338));
  NOR2 NOR2_380(.VSS(VSS),.VDD(VDD),.Y(g15165),.A(g12907),.B(g13835));
  NOR2 NOR2_381(.VSS(VSS),.VDD(VDD),.Y(g31373),.A(g4975),.B(g29725));
  NOR2 NOR2_382(.VSS(VSS),.VDD(VDD),.Y(g11780),.A(g4899),.B(g8822));
  NOR2 NOR2_383(.VSS(VSS),.VDD(VDD),.Y(g14360),.A(g12078),.B(g9484));
  NOR2 NOR2_384(.VSS(VSS),.VDD(VDD),.Y(g9835),.A(g2629),.B(g2555));
  NOR2 NOR2_385(.VSS(VSS),.VDD(VDD),.Y(g14447),.A(g11938),.B(g9698));
  NOR2 NOR2_386(.VSS(VSS),.VDD(VDD),.Y(g12856),.A(g10430),.B(g6855));
  NOR2 NOR2_387(.VSS(VSS),.VDD(VDD),.Y(g29187),.A(g7704),.B(g27999));
  NOR3 NOR3_31(.VSS(VSS),.VDD(VDD),.Y(g11846),.A(g7635),.B(g7518),.C(g7548));
  NOR2 NOR2_388(.VSS(VSS),.VDD(VDD),.Y(g16209),.A(g13478),.B(g4749));
  NOR2 NOR2_389(.VSS(VSS),.VDD(VDD),.Y(g14911),.A(g10213),.B(g12364));
  NOR2 NOR2_390(.VSS(VSS),.VDD(VDD),.Y(g27499),.A(g9095),.B(g26636));
  NOR3 NOR3_32(.VSS(VSS),.VDD(VDD),.Y(g28540),.A(g8125),.B(g27635),.C(g7121));
  NOR2 NOR2_391(.VSS(VSS),.VDD(VDD),.Y(g15372),.A(g817),.B(g14279));
  NOR2 NOR2_392(.VSS(VSS),.VDD(VDD),.Y(g14754),.A(g12821),.B(g2988));
  NOR2 NOR2_393(.VSS(VSS),.VDD(VDD),.Y(g27722),.A(g7247),.B(g25805));
  NOR2 NOR2_394(.VSS(VSS),.VDD(VDD),.Y(g31117),.A(g4991),.B(g29556));
  NOR2 NOR2_395(.VSS(VSS),.VDD(VDD),.Y(g27924),.A(g9946),.B(g25839));
  NOR2 NOR2_396(.VSS(VSS),.VDD(VDD),.Y(g33117),.A(g31261),.B(g32205));
  NOR2 NOR2_397(.VSS(VSS),.VDD(VDD),.Y(g22190),.A(g2827),.B(g18949));
  NOR2 NOR2_398(.VSS(VSS),.VDD(VDD),.Y(g8720),.A(g358),.B(g365));
  NOR2 NOR2_399(.VSS(VSS),.VDD(VDD),.Y(g15063),.A(g6818),.B(g13394));
  NOR2 NOR2_400(.VSS(VSS),.VDD(VDD),.Y(g30934),.A(g29836),.B(g29850));
  NOR2 NOR2_401(.VSS(VSS),.VDD(VDD),.Y(g19984),.A(g17096),.B(g8171));
  NOR2 NOR2_402(.VSS(VSS),.VDD(VDD),.Y(g15137),.A(g6992),.B(g13680));
  NOR2 NOR2_403(.VSS(VSS),.VDD(VDD),.Y(g12432),.A(g1894),.B(g8249));
  NOR2 NOR2_404(.VSS(VSS),.VDD(VDD),.Y(g24959),.A(g8858),.B(g23324));
  NOR2 NOR2_405(.VSS(VSS),.VDD(VDD),.Y(g17190),.A(g723),.B(g14279));
  NOR2 NOR2_406(.VSS(VSS),.VDD(VDD),.Y(g14394),.A(g12116),.B(g9414));
  NOR2 NOR2_407(.VSS(VSS),.VDD(VDD),.Y(g14367),.A(g9547),.B(g12289));
  NOR2 NOR2_408(.VSS(VSS),.VDD(VDD),.Y(g16292),.A(g7943),.B(g13134));
  NOR2 NOR2_409(.VSS(VSS),.VDD(VDD),.Y(g11357),.A(g8558),.B(g8561));
  NOR3 NOR3_33(.VSS(VSS),.VDD(VDD),.Y(g29179),.A(g9311),.B(g28010),.C(g7738));
  NOR2 NOR2_410(.VSS(VSS),.VDD(VDD),.Y(g14420),.A(g12153),.B(g9490));
  NOR2 NOR2_411(.VSS(VSS),.VDD(VDD),.Y(g12198),.A(g9797),.B(g9800));
  NOR2 NOR2_412(.VSS(VSS),.VDD(VDD),.Y(g19853),.A(g15746),.B(g1052));
  NOR3 NOR3_34(.VSS(VSS),.VDD(VDD),.Y(g27528),.A(g8770),.B(g26352),.C(g11083));
  NOR2 NOR2_413(.VSS(VSS),.VDD(VDD),.Y(g10318),.A(g25),.B(g22));
  NOR2 NOR2_414(.VSS(VSS),.VDD(VDD),.Y(g14446),.A(g12190),.B(g9644));
  NOR2 NOR2_415(.VSS(VSS),.VDD(VDD),.Y(g14227),.A(g9863),.B(g10838));
  NOR2 NOR2_416(.VSS(VSS),.VDD(VDD),.Y(g20857),.A(g17929),.B(g9380));
  NOR2 NOR2_417(.VSS(VSS),.VDD(VDD),.Y(g27960),.A(g7134),.B(g25791));
  NOR2 NOR2_418(.VSS(VSS),.VDD(VDD),.Y(g14540),.A(g12287),.B(g9834));
  NOR2 NOR2_419(.VSS(VSS),.VDD(VDD),.Y(g19401),.A(g17193),.B(g14296));
  NOR2 NOR2_420(.VSS(VSS),.VDD(VDD),.Y(g17700),.A(g14792),.B(g12983));
  NOR2 NOR2_421(.VSS(VSS),.VDD(VDD),.Y(g17625),.A(g14541),.B(g12123));
  NOR2 NOR2_422(.VSS(VSS),.VDD(VDD),.Y(g15073),.A(g12844),.B(g13416));
  NOR3 NOR3_35(.VSS(VSS),.VDD(VDD),.Y(g28481),.A(g3506),.B(g10323),.C(g27617));
  NOR2 NOR2_423(.VSS(VSS),.VDD(VDD),.Y(g10281),.A(g5535),.B(g5527));
  NOR2 NOR2_424(.VSS(VSS),.VDD(VDD),.Y(g15122),.A(g6959),.B(g13605));
  NOR2 NOR2_425(.VSS(VSS),.VDD(VDD),.Y(g26515),.A(g24843),.B(g24822));
  NOR2 NOR2_426(.VSS(VSS),.VDD(VDD),.Y(g12708),.A(g9518),.B(g9462));
  NOR2 NOR2_427(.VSS(VSS),.VDD(VDD),.Y(g25005),.A(g6811),.B(g23324));
  NOR2 NOR2_428(.VSS(VSS),.VDD(VDD),.Y(g10699),.A(g8526),.B(g1514));
  NOR2 NOR2_429(.VSS(VSS),.VDD(VDD),.Y(g15153),.A(g13745),.B(g12897));
  NOR2 NOR2_430(.VSS(VSS),.VDD(VDD),.Y(g31116),.A(g7892),.B(g29540));
  NOR3 NOR3_36(.VSS(VSS),.VDD(VDD),.Y(g11248),.A(g7953),.B(g4991),.C(g4983));
  NOR3 NOR3_37(.VSS(VSS),.VDD(VDD),.Y(g32780),.A(g31327),.B(I30330),.C(I30331));
  NOR2 NOR2_431(.VSS(VSS),.VDD(VDD),.Y(g15136),.A(g13680),.B(g12885));
  NOR2 NOR2_432(.VSS(VSS),.VDD(VDD),.Y(g29908),.A(g6918),.B(g28471));
  NOR2 NOR2_433(.VSS(VSS),.VDD(VDD),.Y(g27879),.A(g9523),.B(g25856));
  NOR2 NOR2_434(.VSS(VSS),.VDD(VDD),.Y(g22450),.A(g19345),.B(g15724));
  NOR3 NOR3_38(.VSS(VSS),.VDD(VDD),.Y(g12970),.A(g10555),.B(g10510),.C(g10488));
  NOR2 NOR2_435(.VSS(VSS),.VDD(VDD),.Y(g27878),.A(g9559),.B(g25839));
  NOR2 NOR2_436(.VSS(VSS),.VDD(VDD),.Y(g27337),.A(g8334),.B(g26616));
  NOR2 NOR2_437(.VSS(VSS),.VDD(VDD),.Y(g15164),.A(g13835),.B(g12906));
  NOR2 NOR2_438(.VSS(VSS),.VDD(VDD),.Y(g11945),.A(g7212),.B(g7228));
  NOR2 NOR2_439(.VSS(VSS),.VDD(VDD),.Y(g11999),.A(g9654),.B(g7423));
  NOR2 NOR2_440(.VSS(VSS),.VDD(VDD),.Y(g10715),.A(g8526),.B(g8466));
  NOR3 NOR3_39(.VSS(VSS),.VDD(VDD),.Y(g21389),.A(g10143),.B(g17748),.C(g12259));
  NOR2 NOR2_441(.VSS(VSS),.VDD(VDD),.Y(g20995),.A(g5727),.B(g17287));
  NOR2 NOR2_442(.VSS(VSS),.VDD(VDD),.Y(g28520),.A(g8229),.B(g27635));
  NOR2 NOR2_443(.VSS(VSS),.VDD(VDD),.Y(g25407),.A(g23871),.B(g14645));
  NOR2 NOR2_444(.VSS(VSS),.VDD(VDD),.Y(g27010),.A(g6052),.B(g25839));
  NOR2 NOR2_445(.VSS(VSS),.VDD(VDD),.Y(g11932),.A(g843),.B(g9166));
  NOR2 NOR2_446(.VSS(VSS),.VDD(VDD),.Y(g33130),.A(g32265),.B(g31497));
  NOR2 NOR2_447(.VSS(VSS),.VDD(VDD),.Y(g11448),.A(g4191),.B(g8790));
  NOR2 NOR2_448(.VSS(VSS),.VDD(VDD),.Y(g14490),.A(g9853),.B(g12598));
  NOR2 NOR2_449(.VSS(VSS),.VDD(VDD),.Y(g19907),.A(g16210),.B(g13676));
  NOR2 NOR2_450(.VSS(VSS),.VDD(VDD),.Y(g21140),.A(g6073),.B(g17312));
  NOR2 NOR2_451(.VSS(VSS),.VDD(VDD),.Y(g15091),.A(g13177),.B(g12863));
  NOR2 NOR2_452(.VSS(VSS),.VDD(VDD),.Y(g33437),.A(g31997),.B(g10275));
  NOR2 NOR2_453(.VSS(VSS),.VDD(VDD),.Y(g29007),.A(g9269),.B(g28010));
  NOR2 NOR2_454(.VSS(VSS),.VDD(VDD),.Y(g10671),.A(g1526),.B(g8466));
  NOR2 NOR2_455(.VSS(VSS),.VDD(VDD),.Y(g14181),.A(g9083),.B(g12259));
  NOR2 NOR2_456(.VSS(VSS),.VDD(VDD),.Y(g23871),.A(g2811),.B(g21348));
  NOR2 NOR2_457(.VSS(VSS),.VDD(VDD),.Y(g27353),.A(g8097),.B(g26616));
  NOR2 NOR2_458(.VSS(VSS),.VDD(VDD),.Y(g16183),.A(g9223),.B(g13545));
  NOR2 NOR2_459(.VSS(VSS),.VDD(VDD),.Y(g27823),.A(g9792),.B(g25805));
  NOR4 NOR4_5(.VSS(VSS),.VDD(VDD),.Y(g11148),.A(g8052),.B(g9197),.C(g9174),.D(g9050));
  NOR2 NOR2_460(.VSS(VSS),.VDD(VDD),.Y(g12680),.A(g9631),.B(g9576));
  NOR2 NOR2_461(.VSS(VSS),.VDD(VDD),.Y(g19935),.A(g17062),.B(g8113));
  NOR2 NOR2_462(.VSS(VSS),.VDD(VDD),.Y(g31372),.A(g8796),.B(g29697));
  NOR2 NOR2_463(.VSS(VSS),.VDD(VDD),.Y(g25141),.A(g22228),.B(g10334));
  NOR2 NOR2_464(.VSS(VSS),.VDD(VDD),.Y(g33175),.A(g32099),.B(g7828));
  NOR2 NOR2_465(.VSS(VSS),.VDD(VDD),.Y(g24145),.A(g19402),.B(g19422));
  NOR2 NOR2_466(.VSS(VSS),.VDD(VDD),.Y(g27966),.A(g7153),.B(g25805));
  NOR3 NOR3_40(.VSS(VSS),.VDD(VDD),.Y(g13971),.A(g8938),.B(g4975),.C(g11173));
  NOR2 NOR2_467(.VSS(VSS),.VDD(VDD),.Y(g29035),.A(g9321),.B(g28020));
  NOR2 NOR2_468(.VSS(VSS),.VDD(VDD),.Y(g14211),.A(g9779),.B(g10823));
  NOR2 NOR2_469(.VSS(VSS),.VDD(VDD),.Y(g27364),.A(g8426),.B(g26616));
  NOR2 NOR2_470(.VSS(VSS),.VDD(VDD),.Y(g33137),.A(g4849),.B(g32072));
  NOR2 NOR2_471(.VSS(VSS),.VDD(VDD),.Y(g12017),.A(g9969),.B(g9586));
  NOR2 NOR2_472(.VSS(VSS),.VDD(VDD),.Y(g12364),.A(g10102),.B(g10224));
  NOR2 NOR2_473(.VSS(VSS),.VDD(VDD),.Y(g30613),.A(g4507),.B(g29365));
  NOR2 NOR2_474(.VSS(VSS),.VDD(VDD),.Y(g29142),.A(g5535),.B(g28010));
  NOR2 NOR2_475(.VSS(VSS),.VDD(VDD),.Y(g14497),.A(g5990),.B(g12705));
  NOR2 NOR2_476(.VSS(VSS),.VDD(VDD),.Y(g30273),.A(g5990),.B(g29036));
  NOR2 NOR2_477(.VSS(VSS),.VDD(VDD),.Y(g30106),.A(g28739),.B(g7268));
  NOR2 NOR2_478(.VSS(VSS),.VDD(VDD),.Y(g12288),.A(g2610),.B(g8418));
  NOR3 NOR3_41(.VSS(VSS),.VDD(VDD),.Y(g29193),.A(g9529),.B(g26994),.C(g7812));
  NOR2 NOR2_479(.VSS(VSS),.VDD(VDD),.Y(g19906),.A(g16209),.B(g13672));
  NOR2 NOR2_480(.VSS(VSS),.VDD(VDD),.Y(g12571),.A(g9511),.B(g9451));
  NOR2 NOR2_481(.VSS(VSS),.VDD(VDD),.Y(g12308),.A(g9951),.B(g9954));
  NOR2 NOR2_482(.VSS(VSS),.VDD(VDD),.Y(g25004),.A(g676),.B(g23324));
  NOR2 NOR2_483(.VSS(VSS),.VDD(VDD),.Y(g28496),.A(g3179),.B(g27602));
  NOR2 NOR2_484(.VSS(VSS),.VDD(VDD),.Y(g29165),.A(g5881),.B(g28020));
  NOR2 NOR2_485(.VSS(VSS),.VDD(VDD),.Y(g14339),.A(g12289),.B(g2735));
  NOR2 NOR2_486(.VSS(VSS),.VDD(VDD),.Y(g16072),.A(g10961),.B(g13273));
  NOR2 NOR2_487(.VSS(VSS),.VDD(VDD),.Y(g10338),.A(g5062),.B(g5022));
  NOR2 NOR2_488(.VSS(VSS),.VDD(VDD),.Y(g15062),.A(g6817),.B(g13394));
  NOR2 NOR2_489(.VSS(VSS),.VDD(VDD),.Y(g28986),.A(g5517),.B(g28010));
  NOR2 NOR2_490(.VSS(VSS),.VDD(VDD),.Y(g29006),.A(g5180),.B(g27999));
  NOR2 NOR2_491(.VSS(VSS),.VDD(VDD),.Y(g25947),.A(g1199),.B(g24591));
  NOR2 NOR2_492(.VSS(VSS),.VDD(VDD),.Y(g15508),.A(g10320),.B(g14279));
  NOR2 NOR2_493(.VSS(VSS),.VDD(VDD),.Y(g13959),.A(g3698),.B(g11309));
  NOR2 NOR2_494(.VSS(VSS),.VDD(VDD),.Y(g27954),.A(g10014),.B(g25856));
  NOR2 NOR2_495(.VSS(VSS),.VDD(VDD),.Y(g12752),.A(g9576),.B(g9529));
  NOR2 NOR2_496(.VSS(VSS),.VDD(VDD),.Y(g11958),.A(g9543),.B(g7327));
  NOR2 NOR2_497(.VSS(VSS),.VDD(VDD),.Y(g12374),.A(g2185),.B(g8205));
  NOR2 NOR2_498(.VSS(VSS),.VDD(VDD),.Y(g13378),.A(g11374),.B(g11017));
  NOR2 NOR2_499(.VSS(VSS),.VDD(VDD),.Y(g14411),.A(g9460),.B(g11160));
  NOR2 NOR2_500(.VSS(VSS),.VDD(VDD),.Y(g13603),.A(g8009),.B(g10721));
  NOR2 NOR2_501(.VSS(VSS),.VDD(VDD),.Y(g13944),.A(g10262),.B(g12259));
  NOR2 NOR2_502(.VSS(VSS),.VDD(VDD),.Y(g14867),.A(g10191),.B(g12314));
  NOR2 NOR2_503(.VSS(VSS),.VDD(VDD),.Y(g14450),.A(g12195),.B(g9598));
  NOR2 NOR2_504(.VSS(VSS),.VDD(VDD),.Y(g29175),.A(g6227),.B(g26977));
  NOR2 NOR2_505(.VSS(VSS),.VDD(VDD),.Y(g10819),.A(g7479),.B(g1041));
  NOR2 NOR2_506(.VSS(VSS),.VDD(VDD),.Y(g13730),.A(g3639),.B(g11663));
  NOR3 NOR3_42(.VSS(VSS),.VDD(VDD),.Y(g34359),.A(g9162),.B(g34174),.C(g12259));
  NOR2 NOR2_507(.VSS(VSS),.VDD(VDD),.Y(g14707),.A(g10143),.B(g12259));
  NOR2 NOR2_508(.VSS(VSS),.VDD(VDD),.Y(g28457),.A(g7980),.B(g27602));
  NOR3 NOR3_43(.VSS(VSS),.VDD(VDD),.Y(g32212),.A(g8859),.B(g31262),.C(g11083));
  NOR3 NOR3_44(.VSS(VSS),.VDD(VDD),.Y(g12558),.A(g7738),.B(g5517),.C(g5511));
  NOR2 NOR2_509(.VSS(VSS),.VDD(VDD),.Y(g13765),.A(g8531),.B(g11615));
  NOR2 NOR2_510(.VSS(VSS),.VDD(VDD),.Y(g15051),.A(g6801),.B(g13350));
  NOR2 NOR2_511(.VSS(VSS),.VDD(VDD),.Y(g15072),.A(g13416),.B(g12843));
  NOR2 NOR2_512(.VSS(VSS),.VDD(VDD),.Y(g7192),.A(g6444),.B(g6404));
  NOR2 NOR2_513(.VSS(VSS),.VDD(VDD),.Y(g29873),.A(g6875),.B(g28458));
  NOR2 NOR2_514(.VSS(VSS),.VDD(VDD),.Y(g17180),.A(g1559),.B(g13574));
  NOR3 NOR3_45(.VSS(VSS),.VDD(VDD),.Y(g22993),.A(g1322),.B(g16292),.C(g19873));
  NOR2 NOR2_515(.VSS(VSS),.VDD(VDD),.Y(g14094),.A(g8770),.B(g11083));
  NOR2 NOR2_516(.VSS(VSS),.VDD(VDD),.Y(g15152),.A(g13745),.B(g12896));
  NOR2 NOR2_517(.VSS(VSS),.VDD(VDD),.Y(g33109),.A(g31997),.B(g4584));
  NOR2 NOR2_518(.VSS(VSS),.VDD(VDD),.Y(g12189),.A(g1917),.B(g8302));
  NOR2 NOR2_519(.VSS(VSS),.VDD(VDD),.Y(g13129),.A(g7553),.B(g10762));
  NOR2 NOR2_520(.VSS(VSS),.VDD(VDD),.Y(g10801),.A(g1041),.B(g7479));
  NOR2 NOR2_521(.VSS(VSS),.VDD(VDD),.Y(g17694),.A(g12435),.B(g12955));
  NOR2 NOR2_522(.VSS(VSS),.VDD(VDD),.Y(g33108),.A(g32183),.B(g31228));
  NOR2 NOR2_523(.VSS(VSS),.VDD(VDD),.Y(g30134),.A(g28768),.B(g7280));
  NOR3 NOR3_46(.VSS(VSS),.VDD(VDD),.Y(g11626),.A(g7121),.B(g3863),.C(g3857));
  NOR2 NOR2_524(.VSS(VSS),.VDD(VDD),.Y(g10695),.A(g8462),.B(g8407));
  NOR2 NOR2_525(.VSS(VSS),.VDD(VDD),.Y(g27093),.A(g26712),.B(g26749));
  NOR2 NOR2_526(.VSS(VSS),.VDD(VDD),.Y(g17619),.A(g10179),.B(g12955));
  NOR2 NOR2_527(.VSS(VSS),.VDD(VDD),.Y(g12093),.A(g9924),.B(g7028));
  NOR2 NOR2_528(.VSS(VSS),.VDD(VDD),.Y(g26649),.A(g9037),.B(g24732));
  NOR2 NOR2_529(.VSS(VSS),.VDD(VDD),.Y(g27875),.A(g9875),.B(g25821));
  NOR2 NOR2_530(.VSS(VSS),.VDD(VDD),.Y(g33174),.A(g8714),.B(g32072));
  NOR3 NOR3_47(.VSS(VSS),.VDD(VDD),.Y(g11232),.A(g4966),.B(g7898),.C(g9064));
  NOR2 NOR2_531(.VSS(VSS),.VDD(VDD),.Y(g29034),.A(g5527),.B(g28010));
  NOR2 NOR2_532(.VSS(VSS),.VDD(VDD),.Y(g19400),.A(g17139),.B(g14206));
  NOR2 NOR2_533(.VSS(VSS),.VDD(VDD),.Y(g21127),.A(g18065),.B(g12099));
  NOR2 NOR2_534(.VSS(VSS),.VDD(VDD),.Y(g11697),.A(g8080),.B(g3857));
  NOR2 NOR2_535(.VSS(VSS),.VDD(VDD),.Y(g11995),.A(g9645),.B(g7410));
  NOR2 NOR2_536(.VSS(VSS),.VDD(VDD),.Y(g16027),.A(g10929),.B(g13260));
  NOR3 NOR3_48(.VSS(VSS),.VDD(VDD),.Y(g11261),.A(g7928),.B(g4801),.C(g9030));
  NOR2 NOR2_537(.VSS(VSS),.VDD(VDD),.Y(g14001),.A(g739),.B(g11083));
  NOR2 NOR2_538(.VSS(VSS),.VDD(VDD),.Y(g30240),.A(g7004),.B(g28982));
  NOR4 NOR4_6(.VSS(VSS),.VDD(VDD),.Y(g24631),.A(g20516),.B(g20436),.C(g20219),.D(g22957));
  NOR2 NOR2_539(.VSS(VSS),.VDD(VDD),.Y(g12160),.A(g9721),.B(g9724));
  NOR2 NOR2_540(.VSS(VSS),.VDD(VDD),.Y(g13512),.A(g9077),.B(g12527));
  NOR2 NOR2_541(.VSS(VSS),.VDD(VDD),.Y(g28480),.A(g8059),.B(g27602));
  NOR4 NOR4_7(.VSS(VSS),.VDD(VDD),.Y(g23956),.A(g18957),.B(g18918),.C(g20136),.D(g20114));
  NOR2 NOR2_542(.VSS(VSS),.VDD(VDD),.Y(g8933),.A(g4709),.B(g4785));
  NOR2 NOR2_543(.VSS(VSS),.VDD(VDD),.Y(g31483),.A(g4899),.B(g29725));
  NOR2 NOR2_544(.VSS(VSS),.VDD(VDD),.Y(g13831),.A(g11245),.B(g7666));
  NOR2 NOR2_545(.VSS(VSS),.VDD(VDD),.Y(g12201),.A(g5417),.B(g10047));
  NOR2 NOR2_546(.VSS(VSS),.VDD(VDD),.Y(g29164),.A(g9444),.B(g28010));
  NOR2 NOR2_547(.VSS(VSS),.VDD(VDD),.Y(g12467),.A(g9472),.B(g9407));
  NOR2 NOR2_548(.VSS(VSS),.VDD(VDD),.Y(g30262),.A(g5644),.B(g29008));
  NOR2 NOR2_549(.VSS(VSS),.VDD(VDD),.Y(g13989),.A(g8697),.B(g11309));
  NOR2 NOR2_550(.VSS(VSS),.VDD(VDD),.Y(g13056),.A(g7400),.B(g10741));
  NOR2 NOR2_551(.VSS(VSS),.VDD(VDD),.Y(g16090),.A(g10961),.B(g13315));
  NOR2 NOR2_552(.VSS(VSS),.VDD(VDD),.Y(g26573),.A(g24897),.B(g24884));
  NOR2 NOR2_553(.VSS(VSS),.VDD(VDD),.Y(g11924),.A(g7187),.B(g7209));
  NOR2 NOR2_554(.VSS(VSS),.VDD(VDD),.Y(g29109),.A(g9472),.B(g26994));
  NOR2 NOR2_555(.VSS(VSS),.VDD(VDD),.Y(g27352),.A(g7975),.B(g26616));
  NOR2 NOR2_556(.VSS(VSS),.VDD(VDD),.Y(g26247),.A(g7995),.B(g24732));
  NOR2 NOR2_557(.VSS(VSS),.VDD(VDD),.Y(g7781),.A(g4064),.B(g4057));
  NOR2 NOR2_558(.VSS(VSS),.VDD(VDD),.Y(g12419),.A(g9402),.B(g9326));
  NOR2 NOR2_559(.VSS(VSS),.VDD(VDD),.Y(g25770),.A(g25417),.B(g25377));
  NOR2 NOR2_560(.VSS(VSS),.VDD(VDD),.Y(g29108),.A(g6219),.B(g26977));
  NOR2 NOR2_561(.VSS(VSS),.VDD(VDD),.Y(g24976),.A(g671),.B(g23324));
  NOR2 NOR2_562(.VSS(VSS),.VDD(VDD),.Y(g12418),.A(g9999),.B(g10001));
  NOR2 NOR2_563(.VSS(VSS),.VDD(VDD),.Y(g12170),.A(g10047),.B(g5413));
  NOR2 NOR2_564(.VSS(VSS),.VDD(VDD),.Y(g26098),.A(g9073),.B(g24732));
  NOR2 NOR2_565(.VSS(VSS),.VDD(VDD),.Y(g23024),.A(g7936),.B(g19407));
  NOR2 NOR2_566(.VSS(VSS),.VDD(VDD),.Y(g13342),.A(g10961),.B(g10935));
  NOR2 NOR2_567(.VSS(VSS),.VDD(VDD),.Y(g13031),.A(g7301),.B(g10741));
  NOR2 NOR2_568(.VSS(VSS),.VDD(VDD),.Y(g12853),.A(g6848),.B(g10430));
  NOR3 NOR3_49(.VSS(VSS),.VDD(VDD),.Y(g33851),.A(g8854),.B(g33299),.C(g12259));
  NOR2 NOR2_569(.VSS(VSS),.VDD(VDD),.Y(g29174),.A(g9511),.B(g28020));
  NOR3 NOR3_50(.VSS(VSS),.VDD(VDD),.Y(g21250),.A(g9417),.B(g9340),.C(g17494));
  NOR2 NOR2_570(.VSS(VSS),.VDD(VDD),.Y(g21658),.A(g17694),.B(g17727));
  NOR2 NOR2_571(.VSS(VSS),.VDD(VDD),.Y(g22654),.A(g7733),.B(g19506));
  NOR2 NOR2_572(.VSS(VSS),.VDD(VDD),.Y(g25521),.A(g23955),.B(g14645));
  NOR3 NOR3_51(.VSS(VSS),.VDD(VDD),.Y(g11869),.A(g7649),.B(g7534),.C(g7581));
  NOR2 NOR2_573(.VSS(VSS),.VDD(VDD),.Y(g15647),.A(g11924),.B(g14248));
  NOR2 NOR2_574(.VSS(VSS),.VDD(VDD),.Y(g28469),.A(g3171),.B(g27602));
  NOR2 NOR2_575(.VSS(VSS),.VDD(VDD),.Y(g15090),.A(g13144),.B(g12862));
  NOR3 NOR3_52(.VSS(VSS),.VDD(VDD),.Y(g28468),.A(g3155),.B(g10295),.C(g27602));
  NOR2 NOR2_576(.VSS(VSS),.VDD(VDD),.Y(g10341),.A(g6227),.B(g6219));
  NOR2 NOR2_577(.VSS(VSS),.VDD(VDD),.Y(g25247),.A(g23763),.B(g14645));
  NOR2 NOR2_578(.VSS(VSS),.VDD(VDD),.Y(g27704),.A(g7239),.B(g25791));
  NOR2 NOR2_579(.VSS(VSS),.VDD(VDD),.Y(g11225),.A(g3990),.B(g6928));
  NOR2 NOR2_580(.VSS(VSS),.VDD(VDD),.Y(g26162),.A(g23052),.B(g24751));
  NOR3 NOR3_53(.VSS(VSS),.VDD(VDD),.Y(g16646),.A(g13437),.B(g11020),.C(g11372));
  NOR2 NOR2_581(.VSS(VSS),.VDD(VDD),.Y(g12466),.A(g10057),.B(g10059));
  NOR2 NOR2_582(.VSS(VSS),.VDD(VDD),.Y(g25777),.A(g25482),.B(g25456));
  NOR2 NOR2_583(.VSS(VSS),.VDD(VDD),.Y(g14335),.A(g12045),.B(g9283));
  NOR2 NOR2_584(.VSS(VSS),.VDD(VDD),.Y(g12101),.A(g6336),.B(g7074));
  NOR2 NOR2_585(.VSS(VSS),.VDD(VDD),.Y(g26628),.A(g8990),.B(g24732));
  NOR2 NOR2_586(.VSS(VSS),.VDD(VDD),.Y(g29040),.A(g6209),.B(g26977));
  NOR2 NOR2_587(.VSS(VSS),.VDD(VDD),.Y(g30162),.A(g28880),.B(g7462));
  NOR2 NOR2_588(.VSS(VSS),.VDD(VDD),.Y(g8864),.A(g3179),.B(g3171));
  NOR2 NOR2_589(.VSS(VSS),.VDD(VDD),.Y(g24383),.A(g22409),.B(g22360));
  NOR2 NOR2_590(.VSS(VSS),.VDD(VDD),.Y(g27733),.A(g9305),.B(g25805));
  NOR3 NOR3_54(.VSS(VSS),.VDD(VDD),.Y(g13970),.A(g8883),.B(g8796),.C(g11155));
  NOR4 NOR4_8(.VSS(VSS),.VDD(VDD),.Y(g11171),.A(g8088),.B(g9226),.C(g9200),.D(g9091));
  NOR3 NOR3_55(.VSS(VSS),.VDD(VDD),.Y(g29183),.A(g9392),.B(g28020),.C(g7766));
  NOR3 NOR3_56(.VSS(VSS),.VDD(VDD),.Y(g24875),.A(g8725),.B(g23850),.C(g11083));
  NOR2 NOR2_591(.VSS(VSS),.VDD(VDD),.Y(g12166),.A(g9856),.B(g10124));
  NOR3 NOR3_57(.VSS(VSS),.VDD(VDD),.Y(g14278),.A(g562),.B(g12259),.C(g9217));
  NOR2 NOR2_592(.VSS(VSS),.VDD(VDD),.Y(g13994),.A(g4049),.B(g11363));
  NOR2 NOR2_593(.VSS(VSS),.VDD(VDD),.Y(g15149),.A(g13745),.B(g12894));
  NOR2 NOR2_594(.VSS(VSS),.VDD(VDD),.Y(g25447),.A(g23883),.B(g14645));
  NOR2 NOR2_595(.VSS(VSS),.VDD(VDD),.Y(g14306),.A(g10060),.B(g10887));
  NOR3 NOR3_58(.VSS(VSS),.VDD(VDD),.Y(g29933),.A(g8808),.B(g28500),.C(g12259));
  NOR2 NOR2_596(.VSS(VSS),.VDD(VDD),.Y(g15148),.A(g13716),.B(g12893));
  NOR2 NOR2_597(.VSS(VSS),.VDD(VDD),.Y(g15097),.A(g12868),.B(g13191));
  NOR2 NOR2_598(.VSS(VSS),.VDD(VDD),.Y(g30147),.A(g28768),.B(g14567));
  NOR2 NOR2_599(.VSS(VSS),.VDD(VDD),.Y(g13919),.A(g3347),.B(g11276));
  NOR2 NOR2_600(.VSS(VSS),.VDD(VDD),.Y(g9755),.A(g2070),.B(g1996));
  NOR2 NOR2_601(.VSS(VSS),.VDD(VDD),.Y(g13078),.A(g7446),.B(g10762));
  NOR2 NOR2_602(.VSS(VSS),.VDD(VDD),.Y(g23695),.A(g17420),.B(g21140));
  NOR2 NOR2_603(.VSS(VSS),.VDD(VDD),.Y(g19951),.A(g16219),.B(g13709));
  NOR3 NOR3_59(.VSS(VSS),.VDD(VDD),.Y(g25776),.A(g7166),.B(g24380),.C(g24369));
  NOR2 NOR2_604(.VSS(VSS),.VDD(VDD),.Y(g25785),.A(g25488),.B(g25462));
  NOR2 NOR2_605(.VSS(VSS),.VDD(VDD),.Y(g10884),.A(g7650),.B(g8451));
  NOR2 NOR2_606(.VSS(VSS),.VDD(VDD),.Y(g27382),.A(g8219),.B(g26657));
  NOR2 NOR2_607(.VSS(VSS),.VDD(VDD),.Y(g28953),.A(g5170),.B(g27999));
  NOR2 NOR2_608(.VSS(VSS),.VDD(VDD),.Y(g24494),.A(g23513),.B(g23532));
  NOR2 NOR2_609(.VSS(VSS),.VDD(VDD),.Y(g15133),.A(g12883),.B(g13638));
  NOR3 NOR3_60(.VSS(VSS),.VDD(VDD),.Y(g32650),.A(g31579),.B(I30192),.C(I30193));
  NOR2 NOR2_610(.VSS(VSS),.VDD(VDD),.Y(g13125),.A(g7863),.B(g10762));
  NOR2 NOR2_611(.VSS(VSS),.VDD(VDD),.Y(g10666),.A(g8462),.B(g1171));
  NOR2 NOR2_612(.VSS(VSS),.VDD(VDD),.Y(g25950),.A(g1070),.B(g24591));
  NOR2 NOR2_613(.VSS(VSS),.VDD(VDD),.Y(g7142),.A(g6573),.B(g6565));
  NOR2 NOR2_614(.VSS(VSS),.VDD(VDD),.Y(g12154),.A(g10155),.B(g9835));
  NOR2 NOR2_615(.VSS(VSS),.VDD(VDD),.Y(g29072),.A(g9402),.B(g26977));
  NOR4 NOR4_9(.VSS(VSS),.VDD(VDD),.Y(g9602),.A(g4688),.B(g4681),.C(g4674),.D(g4646));
  NOR2 NOR2_616(.VSS(VSS),.VDD(VDD),.Y(g14556),.A(g6682),.B(g12790));
  NOR2 NOR2_617(.VSS(VSS),.VDD(VDD),.Y(g26645),.A(g23602),.B(g25160));
  NOR2 NOR2_618(.VSS(VSS),.VDD(VDD),.Y(g13336),.A(g11330),.B(g11011));
  NOR2 NOR2_619(.VSS(VSS),.VDD(VDD),.Y(g21256),.A(g15483),.B(g12179));
  NOR3 NOR3_61(.VSS(VSS),.VDD(VDD),.Y(g22983),.A(g979),.B(g16268),.C(g19853));
  NOR2 NOR2_620(.VSS(VSS),.VDD(VDD),.Y(g9015),.A(g3050),.B(g3010));
  NOR2 NOR2_621(.VSS(VSS),.VDD(VDD),.Y(g15050),.A(g12834),.B(g13350));
  NOR2 NOR2_622(.VSS(VSS),.VDD(VDD),.Y(g12729),.A(g1657),.B(g8139));
  NOR2 NOR2_623(.VSS(VSS),.VDD(VDD),.Y(g13631),.A(g8068),.B(g10733));
  NOR2 NOR2_624(.VSS(VSS),.VDD(VDD),.Y(g10922),.A(g7650),.B(g4057));
  NOR2 NOR2_625(.VSS(VSS),.VDD(VDD),.Y(g25446),.A(g23686),.B(g14645));
  NOR2 NOR2_626(.VSS(VSS),.VDD(VDD),.Y(g22517),.A(g19720),.B(g1345));
  NOR4 NOR4_10(.VSS(VSS),.VDD(VDD),.Y(g10179),.A(g2098),.B(g1964),.C(g1830),.D(g1696));
  NOR4 NOR4_11(.VSS(VSS),.VDD(VDD),.Y(g9664),.A(g4878),.B(g4871),.C(g4864),.D(g4836));
  NOR2 NOR2_627(.VSS(VSS),.VDD(VDD),.Y(g15096),.A(g13191),.B(g12867));
  NOR2 NOR2_628(.VSS(VSS),.VDD(VDD),.Y(g30146),.A(g28833),.B(g7411));
  NOR2 NOR2_629(.VSS(VSS),.VDD(VDD),.Y(g25540),.A(g22409),.B(g22360));
  NOR2 NOR2_630(.VSS(VSS),.VDD(VDD),.Y(g14178),.A(g8899),.B(g11083));
  NOR2 NOR2_631(.VSS(VSS),.VDD(VDD),.Y(g31482),.A(g8883),.B(g29697));
  NOR2 NOR2_632(.VSS(VSS),.VDD(VDD),.Y(g30290),.A(g6682),.B(g29110));
  NOR2 NOR2_633(.VSS(VSS),.VDD(VDD),.Y(g28568),.A(g10323),.B(g27617));
  NOR2 NOR2_634(.VSS(VSS),.VDD(VDD),.Y(g25203),.A(g6428),.B(g23756));
  NOR2 NOR2_635(.VSS(VSS),.VDD(VDD),.Y(g11309),.A(g8587),.B(g8728));
  NOR3 NOR3_62(.VSS(VSS),.VDD(VDD),.Y(g11571),.A(g10323),.B(g3512),.C(g3506));
  NOR2 NOR2_636(.VSS(VSS),.VDD(VDD),.Y(g22523),.A(g1345),.B(g19720));
  NOR2 NOR2_637(.VSS(VSS),.VDD(VDD),.Y(g14417),.A(g12149),.B(g9648));
  NOR2 NOR2_638(.VSS(VSS),.VDD(VDD),.Y(g12622),.A(g9569),.B(g9518));
  NOR2 NOR2_639(.VSS(VSS),.VDD(VDD),.Y(g26715),.A(g23711),.B(g25203));
  NOR2 NOR2_640(.VSS(VSS),.VDD(VDD),.Y(g23763),.A(g2795),.B(g21276));
  NOR2 NOR2_641(.VSS(VSS),.VDD(VDD),.Y(g14334),.A(g12044),.B(g9337));
  NOR2 NOR2_642(.VSS(VSS),.VDD(VDD),.Y(g16232),.A(g13516),.B(g4950));
  NOR2 NOR2_643(.VSS(VSS),.VDD(VDD),.Y(g11976),.A(g9595),.B(g7379));
  NOR2 NOR2_644(.VSS(VSS),.VDD(VDD),.Y(g33090),.A(g31997),.B(g4593));
  NOR3 NOR3_63(.VSS(VSS),.VDD(VDD),.Y(g31233),.A(g8522),.B(g29778),.C(g24825));
  NOR2 NOR2_645(.VSS(VSS),.VDD(VDD),.Y(g17727),.A(g12486),.B(g12983));
  NOR2 NOR2_646(.VSS(VSS),.VDD(VDD),.Y(g11954),.A(g9538),.B(g7314));
  NOR2 NOR2_647(.VSS(VSS),.VDD(VDD),.Y(g13954),.A(g8663),.B(g11276));
  NOR2 NOR2_648(.VSS(VSS),.VDD(VDD),.Y(g28510),.A(g3530),.B(g27617));
  NOR2 NOR2_649(.VSS(VSS),.VDD(VDD),.Y(g12333),.A(g1624),.B(g8139));
  NOR2 NOR2_650(.VSS(VSS),.VDD(VDD),.Y(g26297),.A(g8519),.B(g24825));
  NOR2 NOR2_651(.VSS(VSS),.VDD(VDD),.Y(g15129),.A(g6984),.B(g13638));
  NOR2 NOR2_652(.VSS(VSS),.VDD(VDD),.Y(g12852),.A(g6847),.B(g10430));
  NOR2 NOR2_653(.VSS(VSS),.VDD(VDD),.Y(g15057),.A(g6810),.B(g13350));
  NOR2 NOR2_654(.VSS(VSS),.VDD(VDD),.Y(g11669),.A(g3863),.B(g8026));
  NOR2 NOR2_655(.VSS(VSS),.VDD(VDD),.Y(g15128),.A(g13638),.B(g12880));
  NOR2 NOR2_656(.VSS(VSS),.VDD(VDD),.Y(g14000),.A(g8766),.B(g12259));
  NOR2 NOR2_657(.VSS(VSS),.VDD(VDD),.Y(g33449),.A(g10311),.B(g31950));
  NOR2 NOR2_658(.VSS(VSS),.VDD(VDD),.Y(g33448),.A(g7785),.B(g31950));
  NOR2 NOR2_659(.VSS(VSS),.VDD(VDD),.Y(g14568),.A(g12000),.B(g9915));
  NOR2 NOR2_660(.VSS(VSS),.VDD(VDD),.Y(g17175),.A(g1216),.B(g13545));
  NOR2 NOR2_661(.VSS(VSS),.VDD(VDD),.Y(g10123),.A(g4294),.B(g4297));
  NOR2 NOR2_662(.VSS(VSS),.VDD(VDD),.Y(g21655),.A(g17657),.B(g17700));
  NOR3 NOR3_64(.VSS(VSS),.VDD(VDD),.Y(g34354),.A(g9003),.B(g34162),.C(g11083));
  NOR3 NOR3_65(.VSS(VSS),.VDD(VDD),.Y(g12609),.A(g7766),.B(g5863),.C(g5857));
  NOR4 NOR4_12(.VSS(VSS),.VDD(VDD),.Y(g14751),.A(g10622),.B(g10617),.C(g10609),.D(g10603));
  NOR2 NOR2_663(.VSS(VSS),.VDD(VDD),.Y(g14772),.A(g6044),.B(g12252));
  NOR2 NOR2_664(.VSS(VSS),.VDD(VDD),.Y(g8182),.A(g405),.B(g392));
  NOR2 NOR2_665(.VSS(VSS),.VDD(VDD),.Y(g28493),.A(g3873),.B(g27635));
  NOR2 NOR2_666(.VSS(VSS),.VDD(VDD),.Y(g26546),.A(g24858),.B(g24846));
  NOR2 NOR2_667(.VSS(VSS),.VDD(VDD),.Y(g19981),.A(g3727),.B(g16316));
  NOR2 NOR2_668(.VSS(VSS),.VDD(VDD),.Y(g28340),.A(g27439),.B(g26339));
  NOR2 NOR2_669(.VSS(VSS),.VDD(VDD),.Y(g14416),.A(g12148),.B(g9541));
  NOR2 NOR2_670(.VSS(VSS),.VDD(VDD),.Y(g11610),.A(g7980),.B(g3155));
  NOR2 NOR2_671(.VSS(VSS),.VDD(VDD),.Y(g25784),.A(g25507),.B(g25485));
  NOR2 NOR2_672(.VSS(VSS),.VDD(VDD),.Y(g27973),.A(g7187),.B(g25839));
  NOR2 NOR2_673(.VSS(VSS),.VDD(VDD),.Y(g33148),.A(g4854),.B(g32072));
  NOR2 NOR2_674(.VSS(VSS),.VDD(VDD),.Y(g25956),.A(g1413),.B(g24609));
  NOR2 NOR2_675(.VSS(VSS),.VDD(VDD),.Y(g11255),.A(g8623),.B(g6928));
  NOR2 NOR2_676(.VSS(VSS),.VDD(VDD),.Y(g33097),.A(g31950),.B(g4628));
  NOR2 NOR2_677(.VSS(VSS),.VDD(VDD),.Y(g14391),.A(g12112),.B(g9585));
  NOR2 NOR2_678(.VSS(VSS),.VDD(VDD),.Y(g12798),.A(g5535),.B(g9381));
  NOR3 NOR3_66(.VSS(VSS),.VDD(VDD),.Y(g10510),.A(g7183),.B(g4593),.C(g4584));
  NOR2 NOR2_679(.VSS(VSS),.VDD(VDD),.Y(g11270),.A(g8431),.B(g8434));
  NOR2 NOR2_680(.VSS(VSS),.VDD(VDD),.Y(g16198),.A(g9247),.B(g13574));
  NOR2 NOR2_681(.VSS(VSS),.VDD(VDD),.Y(g7352),.A(g1526),.B(g1514));
  NOR2 NOR2_682(.VSS(VSS),.VDD(VDD),.Y(g26625),.A(g23560),.B(g25144));
  NOR2 NOR2_683(.VSS(VSS),.VDD(VDD),.Y(g27732),.A(g9364),.B(g25791));
  NOR3 NOR3_67(.VSS(VSS),.VDD(VDD),.Y(g13939),.A(g4899),.B(g8822),.C(g11173));
  NOR2 NOR2_684(.VSS(VSS),.VDD(VDD),.Y(g32017),.A(g31504),.B(g23475));
  NOR2 NOR2_685(.VSS(VSS),.VDD(VDD),.Y(g26296),.A(g8287),.B(g24732));
  NOR2 NOR2_686(.VSS(VSS),.VDD(VDD),.Y(g26338),.A(g8458),.B(g24825));
  NOR2 NOR2_687(.VSS(VSS),.VDD(VDD),.Y(g15056),.A(g6809),.B(g13350));
  NOR2 NOR2_688(.VSS(VSS),.VDD(VDD),.Y(g27400),.A(g8553),.B(g26657));
  NOR2 NOR2_689(.VSS(VSS),.VDD(VDD),.Y(g10615),.A(g1636),.B(g7308));
  NOR2 NOR2_690(.VSS(VSS),.VDD(VDD),.Y(g31133),.A(g7953),.B(g29556));
  NOR2 NOR2_691(.VSS(VSS),.VDD(VDD),.Y(g33133),.A(g32278),.B(g31503));
  NOR2 NOR2_692(.VSS(VSS),.VDD(VDD),.Y(g28475),.A(g3863),.B(g27635));
  NOR2 NOR2_693(.VSS(VSS),.VDD(VDD),.Y(g21143),.A(g15348),.B(g9517));
  NOR2 NOR2_694(.VSS(VSS),.VDD(VDD),.Y(g19388),.A(g17181),.B(g14256));
  NOR2 NOR2_695(.VSS(VSS),.VDD(VDD),.Y(g15145),.A(g12891),.B(g13716));
  NOR2 NOR2_696(.VSS(VSS),.VDD(VDD),.Y(g24439),.A(g7400),.B(g22312));
  NOR2 NOR2_697(.VSS(VSS),.VDD(VDD),.Y(g9700),.A(g2361),.B(g2287));
  NOR2 NOR2_698(.VSS(VSS),.VDD(VDD),.Y(g11201),.A(g4125),.B(g7765));
  NOR2 NOR2_699(.VSS(VSS),.VDD(VDD),.Y(g33112),.A(g31240),.B(g32194));
  NOR2 NOR2_700(.VSS(VSS),.VDD(VDD),.Y(g27771),.A(g9809),.B(g25839));
  NOR2 NOR2_701(.VSS(VSS),.VDD(VDD),.Y(g19140),.A(g7939),.B(g15695));
  NOR2 NOR2_702(.VSS(VSS),.VDD(VDD),.Y(g19997),.A(g16231),.B(g13739));
  NOR2 NOR2_703(.VSS(VSS),.VDD(VDD),.Y(g15132),.A(g12882),.B(g13638));
  NOR2 NOR2_704(.VSS(VSS),.VDD(VDD),.Y(g12235),.A(g9234),.B(g9206));
  NOR2 NOR2_705(.VSS(VSS),.VDD(VDD),.Y(g33096),.A(g31997),.B(g4608));
  NOR2 NOR2_706(.VSS(VSS),.VDD(VDD),.Y(g14362),.A(g12080),.B(g9338));
  NOR2 NOR2_707(.VSS(VSS),.VDD(VDD),.Y(g22537),.A(g19720),.B(g1367));
  NOR2 NOR2_708(.VSS(VSS),.VDD(VDD),.Y(g15161),.A(g13809),.B(g7073));
  NOR2 NOR2_709(.VSS(VSS),.VDD(VDD),.Y(g14165),.A(g8951),.B(g11083));
  NOR2 NOR2_710(.VSS(VSS),.VDD(VDD),.Y(g29104),.A(g5188),.B(g27999));
  NOR2 NOR2_711(.VSS(VSS),.VDD(VDD),.Y(g12515),.A(g9511),.B(g5873));
  NOR2 NOR2_712(.VSS(VSS),.VDD(VDD),.Y(g15087),.A(g12860),.B(g13144));
  NOR2 NOR2_713(.VSS(VSS),.VDD(VDD),.Y(g32424),.A(g8721),.B(g31294));
  NOR2 NOR2_714(.VSS(VSS),.VDD(VDD),.Y(g34496),.A(g34370),.B(g27648));
  NOR2 NOR2_715(.VSS(VSS),.VDD(VDD),.Y(g14437),.A(g9527),.B(g11178));
  NOR2 NOR2_716(.VSS(VSS),.VDD(VDD),.Y(g11194),.A(g3288),.B(g6875));
  NOR2 NOR2_717(.VSS(VSS),.VDD(VDD),.Y(g15069),.A(g6828),.B(g13416));
  NOR2 NOR2_718(.VSS(VSS),.VDD(VDD),.Y(g14347),.A(g9309),.B(g11123));
  NOR3 NOR3_68(.VSS(VSS),.VDD(VDD),.Y(g14253),.A(g10032),.B(g12259),.C(g9217));
  NOR2 NOR2_719(.VSS(VSS),.VDD(VDD),.Y(g15068),.A(g6826),.B(g13416));
  NOR2 NOR2_720(.VSS(VSS),.VDD(VDD),.Y(g17174),.A(g9194),.B(g14279));
  NOR2 NOR2_721(.VSS(VSS),.VDD(VDD),.Y(g34067),.A(g33859),.B(g11772));
  NOR2 NOR2_722(.VSS(VSS),.VDD(VDD),.Y(g11119),.A(g9180),.B(g9203));
  NOR2 NOR2_723(.VSS(VSS),.VDD(VDD),.Y(g30150),.A(g28846),.B(g7424));
  NOR2 NOR2_724(.VSS(VSS),.VDD(VDD),.Y(g33129),.A(g8630),.B(g32072));
  NOR2 NOR2_725(.VSS(VSS),.VDD(VDD),.Y(g10821),.A(g7503),.B(g1384));
  NOR4 NOR4_13(.VSS(VSS),.VDD(VDD),.Y(g12435),.A(g9012),.B(g8956),.C(g8904),.D(g8863));
  NOR2 NOR2_726(.VSS(VSS),.VDD(VDD),.Y(g33128),.A(g4653),.B(g32057));
  NOR2 NOR2_727(.VSS(VSS),.VDD(VDD),.Y(g14821),.A(g6390),.B(g12314));
  NOR2 NOR2_728(.VSS(VSS),.VDD(VDD),.Y(g22522),.A(g19699),.B(g1024));
  NOR2 NOR2_729(.VSS(VSS),.VDD(VDD),.Y(g11313),.A(g8669),.B(g3759));
  NOR2 NOR2_730(.VSS(VSS),.VDD(VDD),.Y(g27345),.A(g9360),.B(g26636));
  NOR2 NOR2_731(.VSS(VSS),.VDD(VDD),.Y(g12744),.A(g9402),.B(g6203));
  NOR2 NOR2_732(.VSS(VSS),.VDD(VDD),.Y(g14516),.A(g12227),.B(g9704));
  NOR2 NOR2_733(.VSS(VSS),.VDD(VDD),.Y(g11276),.A(g8534),.B(g8691));
  NOR2 NOR2_734(.VSS(VSS),.VDD(VDD),.Y(g12849),.A(g6840),.B(g10430));
  NOR2 NOR2_735(.VSS(VSS),.VDD(VDD),.Y(g17663),.A(g10205),.B(g12983));
  NOR2 NOR2_736(.VSS(VSS),.VDD(VDD),.Y(g12848),.A(g6839),.B(g10430));
  NOR2 NOR2_737(.VSS(VSS),.VDD(VDD),.Y(g27652),.A(g3355),.B(g26636));
  NOR2 NOR2_738(.VSS(VSS),.VDD(VDD),.Y(g26256),.A(g23873),.B(g25479));
  NOR2 NOR2_739(.VSS(VSS),.VDD(VDD),.Y(g22536),.A(g1379),.B(g19720));
  NOR2 NOR2_740(.VSS(VSS),.VDD(VDD),.Y(g15086),.A(g13144),.B(g12859));
  NOR2 NOR2_741(.VSS(VSS),.VDD(VDD),.Y(g12361),.A(g6455),.B(g10172));
  NOR2 NOR2_742(.VSS(VSS),.VDD(VDD),.Y(g14726),.A(g10090),.B(g12166));
  NOR2 NOR2_743(.VSS(VSS),.VDD(VDD),.Y(g30280),.A(g7064),.B(g29036));
  NOR3 NOR3_69(.VSS(VSS),.VDD(VDD),.Y(g32455),.A(g31566),.B(I29985),.C(I29986));
  NOR2 NOR2_744(.VSS(VSS),.VDD(VDD),.Y(g15159),.A(g13809),.B(g12902));
  NOR2 NOR2_745(.VSS(VSS),.VDD(VDD),.Y(g16288),.A(g13794),.B(g417));
  NOR2 NOR2_746(.VSS(VSS),.VDD(VDD),.Y(g14320),.A(g9257),.B(g11111));
  NOR2 NOR2_747(.VSS(VSS),.VDD(VDD),.Y(g15158),.A(g13782),.B(g12901));
  NOR2 NOR2_748(.VSS(VSS),.VDD(VDD),.Y(g30157),.A(g28833),.B(g7369));
  NOR2 NOR2_749(.VSS(VSS),.VDD(VDD),.Y(g14122),.A(g8895),.B(g12259));
  NOR2 NOR2_750(.VSS(VSS),.VDD(VDD),.Y(g15144),.A(g13716),.B(g12890));
  NOR2 NOR2_751(.VSS(VSS),.VDD(VDD),.Y(g31498),.A(g9030),.B(g29540));
  NOR3 NOR3_70(.VSS(VSS),.VDD(VDD),.Y(g28492),.A(g3857),.B(g7121),.C(g27635));
  NOR3 NOR3_71(.VSS(VSS),.VDD(VDD),.Y(g8086),.A(g168),.B(g174),.C(g182));
  NOR2 NOR2_752(.VSS(VSS),.VDD(VDD),.Y(g11907),.A(g7170),.B(g7184));
  NOR2 NOR2_753(.VSS(VSS),.VDD(VDD),.Y(g33432),.A(g31997),.B(g6978));
  NOR2 NOR2_754(.VSS(VSS),.VDD(VDD),.Y(g26314),.A(g24808),.B(g24802));
  NOR2 NOR2_755(.VSS(VSS),.VDD(VDD),.Y(g12371),.A(g1760),.B(g8195));
  NOR2 NOR2_756(.VSS(VSS),.VDD(VDD),.Y(g23835),.A(g2791),.B(g21303));
  NOR2 NOR2_757(.VSS(VSS),.VDD(VDD),.Y(g11238),.A(g8584),.B(g6905));
  NOR2 NOR2_758(.VSS(VSS),.VDD(VDD),.Y(g17213),.A(g11107),.B(g13501));
  NOR2 NOR2_759(.VSS(VSS),.VDD(VDD),.Y(g12234),.A(g9776),.B(g9778));
  NOR2 NOR2_760(.VSS(VSS),.VDD(VDD),.Y(g23586),.A(g17284),.B(g20717));
  NOR2 NOR2_761(.VSS(VSS),.VDD(VDD),.Y(g33145),.A(g8677),.B(g32072));
  NOR2 NOR2_762(.VSS(VSS),.VDD(VDD),.Y(g14164),.A(g9000),.B(g12259));
  NOR3 NOR3_72(.VSS(VSS),.VDD(VDD),.Y(g11185),.A(g8038),.B(g8183),.C(g6804));
  NOR2 NOR2_763(.VSS(VSS),.VDD(VDD),.Y(g13518),.A(g3719),.B(g11903));
  NOR2 NOR2_764(.VSS(VSS),.VDD(VDD),.Y(g16488),.A(g13697),.B(g13656));
  NOR2 NOR2_765(.VSS(VSS),.VDD(VDD),.Y(g16424),.A(g8064),.B(g13628));
  NOR2 NOR2_766(.VSS(VSS),.VDD(VDD),.Y(g26268),.A(g283),.B(g24825));
  NOR2 NOR2_767(.VSS(VSS),.VDD(VDD),.Y(g14575),.A(g10050),.B(g12749));
  NOR2 NOR2_768(.VSS(VSS),.VDD(VDD),.Y(g11935),.A(g9485),.B(g7267));
  NOR3 NOR3_73(.VSS(VSS),.VDD(VDD),.Y(g8131),.A(g4776),.B(g4801),.C(g4793));
  NOR2 NOR2_769(.VSS(VSS),.VDD(VDD),.Y(g27012),.A(g6398),.B(g25856));
  NOR3 NOR3_74(.VSS(VSS),.VDD(VDD),.Y(g13883),.A(g4709),.B(g4785),.C(g11155));
  NOR2 NOR2_770(.VSS(VSS),.VDD(VDD),.Y(g33132),.A(g4843),.B(g32072));
  NOR2 NOR2_771(.VSS(VSS),.VDD(VDD),.Y(g12163),.A(g5073),.B(g9989));
  NOR2 NOR2_772(.VSS(VSS),.VDD(VDD),.Y(g28483),.A(g8080),.B(g27635));
  NOR2 NOR2_773(.VSS(VSS),.VDD(VDD),.Y(g26993),.A(g5360),.B(g25805));
  NOR2 NOR2_774(.VSS(VSS),.VDD(VDD),.Y(g33161),.A(g32090),.B(g7806));
  NOR2 NOR2_775(.VSS(VSS),.VDD(VDD),.Y(g26667),.A(g23642),.B(g25175));
  NOR2 NOR2_776(.VSS(VSS),.VDD(VDD),.Y(g30156),.A(g28789),.B(g14587));
  NOR2 NOR2_777(.VSS(VSS),.VDD(VDD),.Y(g11729),.A(g3179),.B(g8059));
  NOR2 NOR2_778(.VSS(VSS),.VDD(VDD),.Y(g13501),.A(g3368),.B(g11881));
  NOR2 NOR2_779(.VSS(VSS),.VDD(VDD),.Y(g27829),.A(g7345),.B(g25856));
  NOR2 NOR2_780(.VSS(VSS),.VDD(VDD),.Y(g14091),.A(g8854),.B(g12259));
  NOR2 NOR2_781(.VSS(VSS),.VDD(VDD),.Y(g27828),.A(g9892),.B(g25856));
  NOR3 NOR3_75(.VSS(VSS),.VDD(VDD),.Y(g22405),.A(g18957),.B(g20136),.C(g20114));
  NOR2 NOR2_782(.VSS(VSS),.VDD(VDD),.Y(g15669),.A(g11945),.B(g14272));
  NOR2 NOR2_783(.VSS(VSS),.VDD(VDD),.Y(g12358),.A(g10019),.B(g10022));
  NOR2 NOR2_784(.VSS(VSS),.VDD(VDD),.Y(g27344),.A(g8390),.B(g26636));
  NOR2 NOR2_785(.VSS(VSS),.VDD(VDD),.Y(g12121),.A(g10117),.B(g9762));
  NOR2 NOR2_786(.VSS(VSS),.VDD(VDD),.Y(g21193),.A(g15348),.B(g12135));
  NOR2 NOR2_787(.VSS(VSS),.VDD(VDD),.Y(g22929),.A(g19773),.B(g12970));
  NOR2 NOR2_788(.VSS(VSS),.VDD(VDD),.Y(g31068),.A(g4801),.B(g29540));
  NOR2 NOR2_789(.VSS(VSS),.VDD(VDD),.Y(g11566),.A(g3161),.B(g7964));
  NOR2 NOR2_790(.VSS(VSS),.VDD(VDD),.Y(g13622),.A(g278),.B(g11166));
  NOR2 NOR2_791(.VSS(VSS),.VDD(VDD),.Y(g31970),.A(g9024),.B(g30583));
  NOR2 NOR2_792(.VSS(VSS),.VDD(VDD),.Y(g12173),.A(g10050),.B(g7074));
  NOR2 NOR2_793(.VSS(VSS),.VDD(VDD),.Y(g28509),.A(g8107),.B(g27602));
  NOR2 NOR2_794(.VSS(VSS),.VDD(VDD),.Y(g16219),.A(g13498),.B(g4760));
  NOR2 NOR2_795(.VSS(VSS),.VDD(VDD),.Y(g14522),.A(g9924),.B(g12656));
  NOR2 NOR2_796(.VSS(VSS),.VDD(VDD),.Y(g11653),.A(g7980),.B(g7964));
  NOR2 NOR2_797(.VSS(VSS),.VDD(VDD),.Y(g22357),.A(g1024),.B(g19699));
  NOR3 NOR3_76(.VSS(VSS),.VDD(VDD),.Y(g29145),.A(g6549),.B(g7812),.C(g26994));
  NOR2 NOR2_798(.VSS(VSS),.VDD(VDD),.Y(g12029),.A(g5644),.B(g7028));
  NOR2 NOR2_799(.VSS(VSS),.VDD(VDD),.Y(g10862),.A(g7701),.B(g7840));
  NOR2 NOR2_800(.VSS(VSS),.VDD(VDD),.Y(g11415),.A(g8080),.B(g8026));
  NOR2 NOR2_801(.VSS(VSS),.VDD(VDD),.Y(g29198),.A(g7766),.B(g28020));
  NOR2 NOR2_802(.VSS(VSS),.VDD(VDD),.Y(g13852),.A(g11320),.B(g8347));
  NOR2 NOR2_803(.VSS(VSS),.VDD(VDD),.Y(g30601),.A(g16279),.B(g29718));
  NOR2 NOR2_804(.VSS(VSS),.VDD(VDD),.Y(g28452),.A(g3161),.B(g27602));
  NOR2 NOR2_805(.VSS(VSS),.VDD(VDD),.Y(g27927),.A(g9621),.B(g25856));
  NOR2 NOR2_806(.VSS(VSS),.VDD(VDD),.Y(g16201),.A(g13462),.B(g4704));
  NOR2 NOR2_807(.VSS(VSS),.VDD(VDD),.Y(g15093),.A(g13177),.B(g6904));
  NOR2 NOR2_808(.VSS(VSS),.VDD(VDD),.Y(g30143),.A(g28761),.B(g14566));
  NOR2 NOR2_809(.VSS(VSS),.VDD(VDD),.Y(g23063),.A(g16313),.B(g19887));
  NOR2 NOR2_810(.VSS(VSS),.VDD(VDD),.Y(g15065),.A(g13394),.B(g12840));
  NOR2 NOR2_811(.VSS(VSS),.VDD(VDD),.Y(g30169),.A(g28833),.B(g14613));
  NOR2 NOR2_812(.VSS(VSS),.VDD(VDD),.Y(g14397),.A(g12120),.B(g9416));
  NOR2 NOR2_813(.VSS(VSS),.VDD(VDD),.Y(g12604),.A(g5517),.B(g9239));
  NOR2 NOR2_814(.VSS(VSS),.VDD(VDD),.Y(g27770),.A(g9386),.B(g25821));
  NOR2 NOR2_815(.VSS(VSS),.VDD(VDD),.Y(g19338),.A(g16031),.B(g1306));
  NOR2 NOR2_816(.VSS(VSS),.VDD(VDD),.Y(g12755),.A(g6555),.B(g9407));
  NOR2 NOR2_817(.VSS(VSS),.VDD(VDD),.Y(g33125),.A(g8606),.B(g32057));
  NOR2 NOR2_818(.VSS(VSS),.VDD(VDD),.Y(g21209),.A(g15483),.B(g9575));
  NOR2 NOR2_819(.VSS(VSS),.VDD(VDD),.Y(g14872),.A(g6736),.B(g12364));
  NOR2 NOR2_820(.VSS(VSS),.VDD(VDD),.Y(g19968),.A(g17062),.B(g11223));
  NOR2 NOR2_821(.VSS(VSS),.VDD(VDD),.Y(g23208),.A(g20035),.B(g16324));
  NOR2 NOR2_822(.VSS(VSS),.VDD(VDD),.Y(g15160),.A(g12903),.B(g13809));
  NOR2 NOR2_823(.VSS(VSS),.VDD(VDD),.Y(g13799),.A(g8584),.B(g11663));
  NOR2 NOR2_824(.VSS(VSS),.VDD(VDD),.Y(g17482),.A(g9523),.B(g14434));
  NOR2 NOR2_825(.VSS(VSS),.VDD(VDD),.Y(g33144),.A(g4664),.B(g32057));
  NOR3 NOR3_77(.VSS(VSS),.VDD(VDD),.Y(g33823),.A(g8774),.B(g33306),.C(g11083));
  NOR2 NOR2_826(.VSS(VSS),.VDD(VDD),.Y(g20234),.A(g17140),.B(g14207));
  NOR2 NOR2_827(.VSS(VSS),.VDD(VDD),.Y(g29069),.A(g9381),.B(g28010));
  NOR2 NOR2_828(.VSS(VSS),.VDD(VDD),.Y(g11184),.A(g513),.B(g9040));
  NOR2 NOR2_829(.VSS(VSS),.VDD(VDD),.Y(g7158),.A(g5752),.B(g5712));
  NOR4 NOR4_14(.VSS(VSS),.VDD(VDD),.Y(g10205),.A(g2657),.B(g2523),.C(g2389),.D(g2255));
  NOR2 NOR2_830(.VSS(VSS),.VDD(VDD),.Y(g24514),.A(g23619),.B(g23657));
  NOR2 NOR2_831(.VSS(VSS),.VDD(VDD),.Y(g30922),.A(g16662),.B(g29810));
  NOR2 NOR2_832(.VSS(VSS),.VDD(VDD),.Y(g29886),.A(g3288),.B(g28458));
  NOR2 NOR2_833(.VSS(VSS),.VDD(VDD),.Y(g11692),.A(g8021),.B(g7985));
  NOR2 NOR2_834(.VSS(VSS),.VDD(VDD),.Y(g16313),.A(g8005),.B(g13600));
  NOR2 NOR2_835(.VSS(VSS),.VDD(VDD),.Y(g27926),.A(g9467),.B(g25856));
  NOR2 NOR2_836(.VSS(VSS),.VDD(VDD),.Y(g13013),.A(g7957),.B(g10762));
  NOR2 NOR2_837(.VSS(VSS),.VDD(VDD),.Y(g19070),.A(g16957),.B(g11720));
  NOR2 NOR2_838(.VSS(VSS),.VDD(VDD),.Y(g22513),.A(g1002),.B(g19699));
  NOR2 NOR2_839(.VSS(VSS),.VDD(VDD),.Y(g15155),.A(g12899),.B(g13782));
  NOR2 NOR2_840(.VSS(VSS),.VDD(VDD),.Y(g11207),.A(g3639),.B(g6905));
  NOR2 NOR2_841(.VSS(VSS),.VDD(VDD),.Y(g15170),.A(g7118),.B(g14279));
  NOR2 NOR2_842(.VSS(VSS),.VDD(VDD),.Y(g22448),.A(g1018),.B(g19699));
  NOR2 NOR2_843(.VSS(VSS),.VDD(VDD),.Y(g13539),.A(g8594),.B(g12735));
  NOR2 NOR2_844(.VSS(VSS),.VDD(VDD),.Y(g13005),.A(g7939),.B(g10762));
  NOR2 NOR2_845(.VSS(VSS),.VDD(VDD),.Y(g25321),.A(g23835),.B(g14645));
  NOR2 NOR2_846(.VSS(VSS),.VDD(VDD),.Y(g14396),.A(g12119),.B(g9489));
  NOR2 NOR2_847(.VSS(VSS),.VDD(VDD),.Y(g14731),.A(g5698),.B(g12204));
  NOR2 NOR2_848(.VSS(VSS),.VDD(VDD),.Y(g15167),.A(g13835),.B(g12908));
  NOR2 NOR2_849(.VSS(VSS),.VDD(VDD),.Y(g14413),.A(g11914),.B(g9638));
  NOR2 NOR2_850(.VSS(VSS),.VDD(VDD),.Y(g28803),.A(g27730),.B(g22763));
  NOR2 NOR2_851(.VSS(VSS),.VDD(VDD),.Y(g11771),.A(g8921),.B(g4185));
  NOR2 NOR2_852(.VSS(VSS),.VDD(VDD),.Y(g25800),.A(g25518),.B(g25510));
  NOR2 NOR2_853(.VSS(VSS),.VDD(VDD),.Y(g27766),.A(g9716),.B(g25791));
  NOR2 NOR2_854(.VSS(VSS),.VDD(VDD),.Y(g23711),.A(g9892),.B(g21253));
  NOR2 NOR2_855(.VSS(VSS),.VDD(VDD),.Y(g30117),.A(g28739),.B(g7252));
  NOR2 NOR2_856(.VSS(VSS),.VDD(VDD),.Y(g29144),.A(g9518),.B(g26977));
  NOR2 NOR2_857(.VSS(VSS),.VDD(VDD),.Y(g19402),.A(g15979),.B(g13133));
  NOR2 NOR2_858(.VSS(VSS),.VDD(VDD),.Y(g23108),.A(g16424),.B(g19932));
  NOR2 NOR2_859(.VSS(VSS),.VDD(VDD),.Y(g17148),.A(g827),.B(g14279));
  NOR2 NOR2_860(.VSS(VSS),.VDD(VDD),.Y(g11414),.A(g8591),.B(g8593));
  NOR2 NOR2_861(.VSS(VSS),.VDD(VDD),.Y(g16476),.A(g8119),.B(g13667));
  NOR3 NOR3_78(.VSS(VSS),.VDD(VDD),.Y(g32585),.A(g31542),.B(I30123),.C(I30124));
  NOR2 NOR2_862(.VSS(VSS),.VDD(VDD),.Y(g15053),.A(g12836),.B(g13350));
  NOR2 NOR2_863(.VSS(VSS),.VDD(VDD),.Y(g28482),.A(g3522),.B(g27617));
  NOR2 NOR2_864(.VSS(VSS),.VDD(VDD),.Y(g30123),.A(g28768),.B(g7328));
  NOR3 NOR3_79(.VSS(VSS),.VDD(VDD),.Y(g27629),.A(g8891),.B(g26382),.C(g12259));
  NOR2 NOR2_865(.VSS(VSS),.VDD(VDD),.Y(g28552),.A(g10295),.B(g27602));
  NOR2 NOR2_866(.VSS(VSS),.VDD(VDD),.Y(g15101),.A(g12871),.B(g14591));
  NOR2 NOR2_867(.VSS(VSS),.VDD(VDD),.Y(g12246),.A(g9880),.B(g9883));
  NOR2 NOR2_868(.VSS(VSS),.VDD(VDD),.Y(g11584),.A(g8229),.B(g8172));
  NOR2 NOR2_869(.VSS(VSS),.VDD(VDD),.Y(g30265),.A(g7051),.B(g29036));
  NOR2 NOR2_870(.VSS(VSS),.VDD(VDD),.Y(g14640),.A(g12371),.B(g9824));
  NOR2 NOR2_871(.VSS(VSS),.VDD(VDD),.Y(g15064),.A(g6820),.B(g13394));
  NOR2 NOR2_872(.VSS(VSS),.VDD(VDD),.Y(g10803),.A(g1384),.B(g7503));
  NOR2 NOR2_873(.VSS(VSS),.VDD(VDD),.Y(g12591),.A(g504),.B(g9040));
  NOR2 NOR2_874(.VSS(VSS),.VDD(VDD),.Y(g12785),.A(g9472),.B(g6549));
  NOR2 NOR2_875(.VSS(VSS),.VDD(VDD),.Y(g27355),.A(g8443),.B(g26657));
  NOR2 NOR2_876(.VSS(VSS),.VDD(VDD),.Y(g13114),.A(g7528),.B(g10741));
  NOR2 NOR2_877(.VSS(VSS),.VDD(VDD),.Y(g27825),.A(g9316),.B(g25821));
  NOR2 NOR2_878(.VSS(VSS),.VDD(VDD),.Y(g11435),.A(g8107),.B(g3171));
  NOR2 NOR2_879(.VSS(VSS),.VDD(VDD),.Y(g11107),.A(g9095),.B(g9177));
  NOR2 NOR2_880(.VSS(VSS),.VDD(VDD),.Y(g15166),.A(g13835),.B(g7096));
  NOR2 NOR2_881(.VSS(VSS),.VDD(VDD),.Y(g12858),.A(g10365),.B(g10430));
  NOR2 NOR2_882(.VSS(VSS),.VDD(VDD),.Y(g11345),.A(g8477),.B(g8479));
  NOR2 NOR2_883(.VSS(VSS),.VDD(VDD),.Y(g33093),.A(g31997),.B(g4601));
  NOR2 NOR2_884(.VSS(VSS),.VDD(VDD),.Y(g31294),.A(g11326),.B(g29660));
  NOR2 NOR2_885(.VSS(VSS),.VDD(VDD),.Y(g11940),.A(g2712),.B(g10084));
  NOR2 NOR2_886(.VSS(VSS),.VDD(VDD),.Y(g27367),.A(g8155),.B(g26636));
  NOR2 NOR2_887(.VSS(VSS),.VDD(VDD),.Y(g14027),.A(g8734),.B(g11363));
  NOR2 NOR2_888(.VSS(VSS),.VDD(VDD),.Y(g11804),.A(g8938),.B(g4975));
  NOR2 NOR2_889(.VSS(VSS),.VDD(VDD),.Y(g15570),.A(g822),.B(g14279));
  NOR2 NOR2_890(.VSS(VSS),.VDD(VDD),.Y(g14248),.A(g6065),.B(g10578));
  NOR2 NOR2_891(.VSS(VSS),.VDD(VDD),.Y(g16215),.A(g1211),.B(g13545));
  NOR2 NOR2_892(.VSS(VSS),.VDD(VDD),.Y(g24990),.A(g8898),.B(g23324));
  NOR2 NOR2_893(.VSS(VSS),.VDD(VDD),.Y(g14003),.A(g9003),.B(g11083));
  NOR2 NOR2_894(.VSS(VSS),.VDD(VDD),.Y(g15074),.A(g12845),.B(g13416));
  NOR2 NOR2_895(.VSS(VSS),.VDD(VDD),.Y(g12318),.A(g10172),.B(g6451));
  NOR2 NOR2_896(.VSS(VSS),.VDD(VDD),.Y(g27059),.A(g7577),.B(g25895));
  NOR3 NOR3_80(.VSS(VSS),.VDD(VDD),.Y(g15594),.A(g10614),.B(g13026),.C(g7285));
  NOR2 NOR2_897(.VSS(VSS),.VDD(VDD),.Y(g12059),.A(g9853),.B(g7004));
  NOR2 NOR2_898(.VSS(VSS),.VDD(VDD),.Y(g12025),.A(g9705),.B(g7461));
  NOR2 NOR2_899(.VSS(VSS),.VDD(VDD),.Y(g33160),.A(g8672),.B(g32057));
  NOR2 NOR2_900(.VSS(VSS),.VDD(VDD),.Y(g12540),.A(g2587),.B(g8381));
  NOR2 NOR2_901(.VSS(VSS),.VDD(VDD),.Y(g13500),.A(g8480),.B(g12641));
  NOR2 NOR2_902(.VSS(VSS),.VDD(VDD),.Y(g15092),.A(g12864),.B(g13177));
  NOR2 NOR2_903(.VSS(VSS),.VDD(VDD),.Y(g28149),.A(g27598),.B(g27612));
  NOR2 NOR2_904(.VSS(VSS),.VDD(VDD),.Y(g15154),.A(g13782),.B(g12898));
  NOR2 NOR2_905(.VSS(VSS),.VDD(VDD),.Y(g21062),.A(g9547),.B(g17297));
  NOR2 NOR2_906(.VSS(VSS),.VDD(VDD),.Y(g14090),.A(g8851),.B(g12259));
  NOR2 NOR2_907(.VSS(VSS),.VDD(VDD),.Y(g13004),.A(g7933),.B(g10741));
  NOR2 NOR2_908(.VSS(VSS),.VDD(VDD),.Y(g33075),.A(g31997),.B(g7163));
  NOR2 NOR2_909(.VSS(VSS),.VDD(VDD),.Y(g19268),.A(g15979),.B(g962));
  NOR3 NOR3_81(.VSS(VSS),.VDD(VDD),.Y(g12377),.A(g6856),.B(g2748),.C(g9708));
  NOR2 NOR2_910(.VSS(VSS),.VDD(VDD),.Y(g12739),.A(g9321),.B(g9274));
  NOR2 NOR2_911(.VSS(VSS),.VDD(VDD),.Y(g30130),.A(g28761),.B(g7275));
  NOR3 NOR3_82(.VSS(VSS),.VDD(VDD),.Y(g24701),.A(g979),.B(g23024),.C(g19778));
  NOR2 NOR2_912(.VSS(VSS),.VDD(VDD),.Y(g12146),.A(g1783),.B(g8241));
  NOR2 NOR2_913(.VSS(VSS),.VDD(VDD),.Y(g12645),.A(g4467),.B(g6961));
  NOR2 NOR2_914(.VSS(VSS),.VDD(VDD),.Y(g13947),.A(g8948),.B(g11083));
  NOR2 NOR2_915(.VSS(VSS),.VDD(VDD),.Y(g11273),.A(g3061),.B(g8620));
  NOR2 NOR2_916(.VSS(VSS),.VDD(VDD),.Y(g14513),.A(g12222),.B(g9754));
  NOR3 NOR3_83(.VSS(VSS),.VDD(VDD),.Y(g29705),.A(g28399),.B(g8284),.C(g8404));
  NOR2 NOR2_917(.VSS(VSS),.VDD(VDD),.Y(g14449),.A(g12194),.B(g9653));
  NOR3 NOR3_84(.VSS(VSS),.VDD(VDD),.Y(g29189),.A(g9462),.B(g26977),.C(g7791));
  NOR2 NOR2_918(.VSS(VSS),.VDD(VDD),.Y(g33419),.A(g31978),.B(g7627));
  NOR2 NOR2_919(.VSS(VSS),.VDD(VDD),.Y(g14448),.A(g12192),.B(g9699));
  NOR2 NOR2_920(.VSS(VSS),.VDD(VDD),.Y(g11972),.A(g9591),.B(g7361));
  NOR2 NOR2_921(.VSS(VSS),.VDD(VDD),.Y(g27366),.A(g8016),.B(g26636));
  NOR2 NOR2_922(.VSS(VSS),.VDD(VDD),.Y(g7567),.A(g979),.B(g990));
  NOR2 NOR2_923(.VSS(VSS),.VDD(VDD),.Y(g14212),.A(g5373),.B(g10537));
  NOR2 NOR2_924(.VSS(VSS),.VDD(VDD),.Y(g12632),.A(g9631),.B(g6565));
  NOR2 NOR2_925(.VSS(VSS),.VDD(VDD),.Y(g24766),.A(g3385),.B(g23132));
  NOR2 NOR2_926(.VSS(VSS),.VDD(VDD),.Y(g23051),.A(g7960),.B(g19427));
  NOR3 NOR3_85(.VSS(VSS),.VDD(VDD),.Y(g34703),.A(g8899),.B(g34545),.C(g11083));
  NOR3 NOR3_86(.VSS(VSS),.VDD(VDD),.Y(g11514),.A(g10295),.B(g3161),.C(g3155));
  NOR2 NOR2_927(.VSS(VSS),.VDD(VDD),.Y(g12226),.A(g2476),.B(g8373));
  NOR2 NOR2_928(.VSS(VSS),.VDD(VDD),.Y(g31119),.A(g7898),.B(g29556));
  NOR2 NOR2_929(.VSS(VSS),.VDD(VDD),.Y(g26873),.A(g25374),.B(g25331));
  NOR2 NOR2_930(.VSS(VSS),.VDD(VDD),.Y(g11012),.A(g7693),.B(g7846));
  NOR2 NOR2_931(.VSS(VSS),.VDD(VDD),.Y(g15139),.A(g12886),.B(g13680));
  NOR2 NOR2_932(.VSS(VSS),.VDD(VDD),.Y(g26209),.A(g23124),.B(g24779));
  NOR2 NOR2_933(.VSS(VSS),.VDD(VDD),.Y(g15138),.A(g13680),.B(g6993));
  NOR2 NOR2_934(.VSS(VSS),.VDD(VDD),.Y(g11473),.A(g8107),.B(g8059));
  NOR2 NOR2_935(.VSS(VSS),.VDD(VDD),.Y(g29915),.A(g6941),.B(g28484));
  NOR2 NOR2_936(.VSS(VSS),.VDD(VDD),.Y(g27354),.A(g8064),.B(g26636));
  NOR2 NOR2_937(.VSS(VSS),.VDD(VDD),.Y(g12297),.A(g9269),.B(g9239));
  NOR2 NOR2_938(.VSS(VSS),.VDD(VDD),.Y(g13325),.A(g7841),.B(g10741));
  NOR2 NOR2_939(.VSS(VSS),.VDD(VDD),.Y(g12980),.A(g7909),.B(g10741));
  NOR2 NOR2_940(.VSS(VSS),.VDD(VDD),.Y(g12824),.A(g5881),.B(g9451));
  NOR2 NOR2_941(.VSS(VSS),.VDD(VDD),.Y(g25952),.A(g1542),.B(g24609));
  NOR2 NOR2_942(.VSS(VSS),.VDD(VDD),.Y(g13946),.A(g8651),.B(g11083));
  NOR2 NOR2_943(.VSS(VSS),.VDD(VDD),.Y(g25175),.A(g5736),.B(g23692));
  NOR2 NOR2_944(.VSS(VSS),.VDD(VDD),.Y(g14228),.A(g5719),.B(g10561));
  NOR2 NOR2_945(.VSS(VSS),.VDD(VDD),.Y(g15585),.A(g11862),.B(g14194));
  NOR2 NOR2_946(.VSS(VSS),.VDD(VDD),.Y(g26346),.A(g8522),.B(g24825));
  NOR2 NOR2_947(.VSS(VSS),.VDD(VDD),.Y(g15608),.A(g11885),.B(g14212));
  NOR2 NOR2_948(.VSS(VSS),.VDD(VDD),.Y(g15052),.A(g12835),.B(g13350));
  NOR2 NOR2_949(.VSS(VSS),.VDD(VDD),.Y(g12211),.A(g10099),.B(g7097));
  NOR2 NOR2_950(.VSS(VSS),.VDD(VDD),.Y(g31008),.A(g30004),.B(g30026));
  NOR2 NOR2_951(.VSS(VSS),.VDD(VDD),.Y(g31476),.A(g4709),.B(g29697));
  NOR2 NOR2_952(.VSS(VSS),.VDD(VDD),.Y(g29167),.A(g9576),.B(g26994));
  NOR2 NOR2_953(.VSS(VSS),.VDD(VDD),.Y(g17198),.A(g9282),.B(g14279));
  NOR2 NOR2_954(.VSS(VSS),.VDD(VDD),.Y(g27659),.A(g3706),.B(g26657));
  NOR2 NOR2_955(.VSS(VSS),.VDD(VDD),.Y(g17393),.A(g9386),.B(g14379));
  NOR2 NOR2_956(.VSS(VSS),.VDD(VDD),.Y(g12700),.A(g9321),.B(g5857));
  NOR2 NOR2_957(.VSS(VSS),.VDD(VDD),.Y(g12659),.A(g9451),.B(g9392));
  NOR2 NOR2_958(.VSS(VSS),.VDD(VDD),.Y(g12126),.A(g9989),.B(g5069));
  NOR2 NOR2_959(.VSS(VSS),.VDD(VDD),.Y(g30136),.A(g28799),.B(g7380));
  NOR2 NOR2_960(.VSS(VSS),.VDD(VDD),.Y(g19953),.A(g16220),.B(g13712));
  NOR2 NOR2_961(.VSS(VSS),.VDD(VDD),.Y(g10793),.A(g1389),.B(g7503));
  NOR2 NOR2_962(.VSS(VSS),.VDD(VDD),.Y(g14793),.A(g2988),.B(g12228));
  NOR2 NOR2_963(.VSS(VSS),.VDD(VDD),.Y(g27338),.A(g9291),.B(g26616));
  NOR2 NOR2_964(.VSS(VSS),.VDD(VDD),.Y(g12296),.A(g9860),.B(g9862));
  NOR2 NOR2_965(.VSS(VSS),.VDD(VDD),.Y(g9762),.A(g2495),.B(g2421));
  NOR2 NOR2_966(.VSS(VSS),.VDD(VDD),.Y(g23662),.A(g17393),.B(g20995));
  NOR2 NOR2_967(.VSS(VSS),.VDD(VDD),.Y(g27969),.A(g7170),.B(g25821));
  NOR2 NOR2_968(.VSS(VSS),.VDD(VDD),.Y(g14549),.A(g9992),.B(g12705));
  NOR2 NOR2_969(.VSS(VSS),.VDD(VDD),.Y(g11755),.A(g4709),.B(g8796));
  NOR2 NOR2_970(.VSS(VSS),.VDD(VDD),.Y(g29900),.A(g3639),.B(g28471));
  NOR2 NOR2_971(.VSS(VSS),.VDD(VDD),.Y(g33092),.A(g31978),.B(g4332));
  NOR2 NOR2_972(.VSS(VSS),.VDD(VDD),.Y(g11563),.A(g8059),.B(g8011));
  NOR2 NOR2_973(.VSS(VSS),.VDD(VDD),.Y(g12855),.A(g10430),.B(g6854));
  NOR2 NOR2_974(.VSS(VSS),.VDD(VDD),.Y(g31935),.A(g30583),.B(g4349));
  NOR3 NOR3_87(.VSS(VSS),.VDD(VDD),.Y(g23204),.A(g10685),.B(g19462),.C(g16488));
  NOR2 NOR2_975(.VSS(VSS),.VDD(VDD),.Y(g14002),.A(g8681),.B(g11083));
  NOR2 NOR2_976(.VSS(VSS),.VDD(VDD),.Y(g17657),.A(g14751),.B(g12955));
  NOR3 NOR3_88(.VSS(VSS),.VDD(VDD),.Y(g11191),.A(g4776),.B(g4801),.C(g9030));
  NOR2 NOR2_977(.VSS(VSS),.VDD(VDD),.Y(g28498),.A(g8172),.B(g27635));
  NOR2 NOR2_978(.VSS(VSS),.VDD(VDD),.Y(g15100),.A(g13191),.B(g12870));
  NOR2 NOR2_979(.VSS(VSS),.VDD(VDD),.Y(g12581),.A(g9569),.B(g6219));
  NOR2 NOR2_980(.VSS(VSS),.VDD(VDD),.Y(g33439),.A(g31950),.B(g4633));
  NOR2 NOR2_981(.VSS(VSS),.VDD(VDD),.Y(g7175),.A(g6098),.B(g6058));
  NOR2 NOR2_982(.VSS(VSS),.VDD(VDD),.Y(g33438),.A(g31950),.B(g4621));
  NOR2 NOR2_983(.VSS(VSS),.VDD(VDD),.Y(g7139),.A(g5406),.B(g5366));
  NOR2 NOR2_984(.VSS(VSS),.VDD(VDD),.Y(g22545),.A(g1373),.B(g19720));
  NOR3 NOR3_89(.VSS(VSS),.VDD(VDD),.Y(g28031),.A(g21209),.B(I26522),.C(I26523));
  NOR2 NOR2_985(.VSS(VSS),.VDD(VDD),.Y(g12067),.A(g5990),.B(g7051));
  NOR2 NOR2_986(.VSS(VSS),.VDD(VDD),.Y(g14512),.A(g11955),.B(g9753));
  NOR2 NOR2_987(.VSS(VSS),.VDD(VDD),.Y(g27735),.A(g7262),.B(g25821));
  NOR2 NOR2_988(.VSS(VSS),.VDD(VDD),.Y(g27877),.A(g9397),.B(g25839));
  NOR3 NOR3_90(.VSS(VSS),.VDD(VDD),.Y(g28529),.A(g8070),.B(g27617),.C(g10323));
  NOR2 NOR2_989(.VSS(VSS),.VDD(VDD),.Y(g12150),.A(g2208),.B(g8259));
  NOR2 NOR2_990(.VSS(VSS),.VDD(VDD),.Y(g33139),.A(g8650),.B(g32057));
  NOR2 NOR2_991(.VSS(VSS),.VDD(VDD),.Y(g10831),.A(g7690),.B(g7827));
  NOR2 NOR2_992(.VSS(VSS),.VDD(VDD),.Y(g13032),.A(g7577),.B(g10762));
  NOR2 NOR2_993(.VSS(VSS),.VDD(VDD),.Y(g33138),.A(g32287),.B(g31514));
  NOR2 NOR2_994(.VSS(VSS),.VDD(VDD),.Y(g14445),.A(g12188),.B(g9693));
  NOR2 NOR2_995(.VSS(VSS),.VDD(VDD),.Y(g12695),.A(g9269),.B(g9239));
  NOR3 NOR3_91(.VSS(VSS),.VDD(VDD),.Y(g29675),.A(g28380),.B(g8236),.C(g8354));
  NOR2 NOR2_996(.VSS(VSS),.VDD(VDD),.Y(g26183),.A(g23079),.B(g24766));
  NOR2 NOR2_997(.VSS(VSS),.VDD(VDD),.Y(g30252),.A(g7028),.B(g29008));
  NOR2 NOR2_998(.VSS(VSS),.VDD(VDD),.Y(g7304),.A(g1183),.B(g1171));
  NOR2 NOR2_999(.VSS(VSS),.VDD(VDD),.Y(g14611),.A(g12333),.B(g9749));
  NOR2 NOR2_1000(.VSS(VSS),.VDD(VDD),.Y(g7499),.A(g333),.B(g355));
  NOR3 NOR3_92(.VSS(VSS),.VDD(VDD),.Y(g14988),.A(g10816),.B(g10812),.C(g10805));
  NOR2 NOR2_1001(.VSS(VSS),.VDD(VDD),.Y(g11360),.A(g3763),.B(g8669));
  NOR2 NOR2_1002(.VSS(VSS),.VDD(VDD),.Y(g26872),.A(g25411),.B(g25371));
  NOR2 NOR2_1003(.VSS(VSS),.VDD(VDD),.Y(g14271),.A(g10002),.B(g10874));
  NOR2 NOR2_1004(.VSS(VSS),.VDD(VDD),.Y(g30183),.A(g28880),.B(g14644));
  NOR2 NOR2_1005(.VSS(VSS),.VDD(VDD),.Y(g19430),.A(g17150),.B(g14220));
  NOR2 NOR2_1006(.VSS(VSS),.VDD(VDD),.Y(g15141),.A(g12888),.B(g13680));
  NOR2 NOR2_1007(.VSS(VSS),.VDD(VDD),.Y(g14145),.A(g8945),.B(g12259));
  NOR2 NOR2_1008(.VSS(VSS),.VDD(VDD),.Y(g12256),.A(g10136),.B(g6105));
  NOR2 NOR2_1009(.VSS(VSS),.VDD(VDD),.Y(g25948),.A(g7752),.B(g24609));
  NOR2 NOR2_1010(.VSS(VSS),.VDD(VDD),.Y(g24497),.A(g23533),.B(g23553));
  NOR2 NOR2_1011(.VSS(VSS),.VDD(VDD),.Y(g14529),.A(g6336),.B(g12749));
  NOR2 NOR2_1012(.VSS(VSS),.VDD(VDD),.Y(g27102),.A(g26750),.B(g26779));
  NOR2 NOR2_1013(.VSS(VSS),.VDD(VDD),.Y(g15135),.A(g6990),.B(g13638));
  NOR2 NOR2_1014(.VSS(VSS),.VDD(VDD),.Y(g26574),.A(g24887),.B(g24861));
  NOR2 NOR2_1015(.VSS(VSS),.VDD(VDD),.Y(g14393),.A(g12115),.B(g9488));
  NOR2 NOR2_1016(.VSS(VSS),.VDD(VDD),.Y(g14365),.A(g12084),.B(g9339));
  NOR3 NOR3_93(.VSS(VSS),.VDD(VDD),.Y(g32845),.A(g30673),.B(I30399),.C(I30400));
  NOR2 NOR2_1017(.VSS(VSS),.VDD(VDD),.Y(g17309),.A(g9305),.B(g14344));
  NOR2 NOR2_1018(.VSS(VSS),.VDD(VDD),.Y(g15049),.A(g13350),.B(g6799));
  NOR2 NOR2_1019(.VSS(VSS),.VDD(VDD),.Y(g11950),.A(g9220),.B(g9166));
  NOR2 NOR2_1020(.VSS(VSS),.VDD(VDD),.Y(g10709),.A(g7499),.B(g351));
  NOR3 NOR3_94(.VSS(VSS),.VDD(VDD),.Y(g27511),.A(g22137),.B(g26866),.C(g20277));
  NOR2 NOR2_1021(.VSS(VSS),.VDD(VDD),.Y(g12854),.A(g6849),.B(g10430));
  NOR2 NOR2_1022(.VSS(VSS),.VDD(VDD),.Y(g28425),.A(g27493),.B(g26351));
  NOR4 NOR4_15(.VSS(VSS),.VDD(VDD),.Y(g34912),.A(g34883),.B(g20277),.C(g20242),.D(g21370));
  NOR3 NOR3_95(.VSS(VSS),.VDD(VDD),.Y(g25851),.A(g4311),.B(g24380),.C(g24369));
  NOR3 NOR3_96(.VSS(VSS),.VDD(VDD),.Y(g13996),.A(g8938),.B(g8822),.C(g11173));
  NOR3 NOR3_97(.VSS(VSS),.VDD(VDD),.Y(g28444),.A(g8575),.B(g27463),.C(g24825));
  NOR2 NOR2_1023(.VSS(VSS),.VDD(VDD),.Y(g15106),.A(g12872),.B(g10430));
  NOR2 NOR2_1024(.VSS(VSS),.VDD(VDD),.Y(g17954),.A(g832),.B(g14279));
  NOR2 NOR2_1025(.VSS(VSS),.VDD(VDD),.Y(g12550),.A(g9300),.B(g9259));
  NOR2 NOR2_1026(.VSS(VSS),.VDD(VDD),.Y(g12314),.A(g10053),.B(g10207));
  NOR2 NOR2_1027(.VSS(VSS),.VDD(VDD),.Y(g14602),.A(g10099),.B(g12790));
  NOR2 NOR2_1028(.VSS(VSS),.VDD(VDD),.Y(g27721),.A(g9672),.B(g25805));
  NOR2 NOR2_1029(.VSS(VSS),.VDD(VDD),.Y(g12085),.A(g10082),.B(g9700));
  NOR2 NOR2_1030(.VSS(VSS),.VDD(VDD),.Y(g22488),.A(g19699),.B(g1002));
  NOR2 NOR2_1031(.VSS(VSS),.VDD(VDD),.Y(g14337),.A(g12049),.B(g9284));
  NOR3 NOR3_98(.VSS(VSS),.VDD(VDD),.Y(g11203),.A(g4966),.B(g4991),.C(g9064));
  NOR2 NOR2_1032(.VSS(VSS),.VDD(VDD),.Y(g13044),.A(g7349),.B(g10762));
  NOR4 NOR4_16(.VSS(VSS),.VDD(VDD),.Y(g14792),.A(g10653),.B(g10623),.C(g10618),.D(g10611));
  NOR3 NOR3_99(.VSS(VSS),.VDD(VDD),.Y(g28353),.A(g9073),.B(g27654),.C(g24732));
  NOR2 NOR2_1033(.VSS(VSS),.VDD(VDD),.Y(g29200),.A(g7791),.B(g26977));
  NOR2 NOR2_1034(.VSS(VSS),.VDD(VDD),.Y(g9640),.A(g1802),.B(g1728));
  NOR2 NOR2_1035(.VSS(VSS),.VDD(VDD),.Y(g19063),.A(g7909),.B(g15674));
  NOR2 NOR2_1036(.VSS(VSS),.VDD(VDD),.Y(g33100),.A(g32172),.B(g31188));
  NOR2 NOR2_1037(.VSS(VSS),.VDD(VDD),.Y(g13377),.A(g7873),.B(g10762));
  NOR2 NOR2_1038(.VSS(VSS),.VDD(VDD),.Y(g14425),.A(g5644),.B(g12656));
  NOR2 NOR2_1039(.VSS(VSS),.VDD(VDD),.Y(g27734),.A(g9733),.B(g25821));
  NOR2 NOR2_1040(.VSS(VSS),.VDD(VDD),.Y(g15163),.A(g13809),.B(g12905));
  NOR2 NOR2_1041(.VSS(VSS),.VDD(VDD),.Y(g30929),.A(g29803),.B(g29835));
  NOR2 NOR2_1042(.VSS(VSS),.VDD(VDD),.Y(g19873),.A(g15755),.B(g1395));
  NOR3 NOR3_100(.VSS(VSS),.VDD(VDD),.Y(g10918),.A(g1532),.B(g7751),.C(g7778));
  NOR2 NOR2_1043(.VSS(VSS),.VDD(VDD),.Y(g19422),.A(g16031),.B(g13141));
  NOR2 NOR2_1044(.VSS(VSS),.VDD(VDD),.Y(g14444),.A(g11936),.B(g9692));
  NOR3 NOR3_101(.VSS(VSS),.VDD(VDD),.Y(g12667),.A(g7791),.B(g6209),.C(g6203));
  NOR3 NOR3_102(.VSS(VSS),.VDD(VDD),.Y(g19209),.A(g12971),.B(g15614),.C(g11320));
  NOR3 NOR3_103(.VSS(VSS),.VDD(VDD),.Y(g13698),.A(g528),.B(g12527),.C(g11185));
  NOR2 NOR2_1045(.VSS(VSS),.VDD(VDD),.Y(g31515),.A(g4983),.B(g29556));
  NOR2 NOR2_1046(.VSS(VSS),.VDD(VDD),.Y(g29184),.A(g9631),.B(g26994));
  NOR2 NOR2_1047(.VSS(VSS),.VDD(VDD),.Y(g23626),.A(g17309),.B(g20854));
  NOR2 NOR2_1048(.VSS(VSS),.VDD(VDD),.Y(g15724),.A(g13858),.B(g11374));
  NOR2 NOR2_1049(.VSS(VSS),.VDD(VDD),.Y(g24018),.A(I23162),.B(I23163));
  NOR2 NOR2_1050(.VSS(VSS),.VDD(VDD),.Y(g30282),.A(g6336),.B(g29073));
  NOR2 NOR2_1051(.VSS(VSS),.VDD(VDD),.Y(g19453),.A(g17199),.B(g14316));
  NOR2 NOR2_1052(.VSS(VSS),.VDD(VDD),.Y(g15121),.A(g12874),.B(g13605));
  NOR2 NOR2_1053(.VSS(VSS),.VDD(VDD),.Y(g12443),.A(g9374),.B(g9300));
  NOR2 NOR2_1054(.VSS(VSS),.VDD(VDD),.Y(g19436),.A(g17176),.B(g14233));
  NOR2 NOR2_1055(.VSS(VSS),.VDD(VDD),.Y(g13661),.A(g528),.B(g11185));
  NOR2 NOR2_1056(.VSS(VSS),.VDD(VDD),.Y(g11715),.A(g8080),.B(g8026));
  NOR3 NOR3_104(.VSS(VSS),.VDD(VDD),.Y(g29005),.A(g5164),.B(g7704),.C(g27999));
  NOR2 NOR2_1057(.VSS(VSS),.VDD(VDD),.Y(g33107),.A(g32180),.B(g31223));
  NOR2 NOR2_1058(.VSS(VSS),.VDD(VDD),.Y(g12601),.A(g9381),.B(g9311));
  NOR2 NOR2_1059(.VSS(VSS),.VDD(VDD),.Y(g15134),.A(g13638),.B(g12884));
  NOR2 NOR2_1060(.VSS(VSS),.VDD(VDD),.Y(g14364),.A(g12083),.B(g9415));
  NOR2 NOR2_1061(.VSS(VSS),.VDD(VDD),.Y(g25769),.A(g25453),.B(g25414));
  NOR2 NOR2_1062(.VSS(VSS),.VDD(VDD),.Y(g11385),.A(g8021),.B(g7985));

endmodule