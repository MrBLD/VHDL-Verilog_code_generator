module s1320(g723,g6269,g7729,g7287,g4370,g6425,g702,g7292,g962,g4657,g7425,g1724,g634,g9310,g7285,g5684,g648,g8234,VDD,g1234,g5143,g9128,g1798,g3860,g756,g453,g6849,g8219,g6909,g7732,g7295,g5678,g6212,g1871,g7293,g9204,g2888,g7063,g752,g722,g3077,g753,g1810,g2844,g6207,g534,g7298,g1017,g291,g3829,g1804,g49,g3859,g6675,g9305,g7730,g206,g6850,g7103,g4660,g7731,g785,g8661,g4371,g1006,g694,g1080,g1016,g7291,g7283,g3096,g1824,g4664,g4655,g4661,g7294,g6236,g5682,g9297,g9280,g7508,g1894,g8872,g7286,g8958,g7505,g9299,g6223,g1783,g4267,g754,g9378,g9314,g1944,g6895,g3191,g6648,g1829,g7514,g8663,g1553,g4373,g635,g645,g1817,g647,g7474,g7506,g7289,g43,g941,g7288,g6653,g4316,g1554,g7423,g690,g7424,g757,g1000,g8216,g5164,g5571,g1015,g1911,g7504,g3159,g751,g372,g7290,g1246,g7048,g5729,g9132,g4663,g9308,g7507,g9312,g8218,g781,g3130,g5669,g2662,g7284,g594,g8217,VSS,g1008,g1870,g755,g698,CLOCK,g633,g4372,g5687);
input g723,g752,g722,g754,g751,g702,g753,g962,g634,g49,g1553,g648,g635,VDD,g645,g647,g1234,g756,g781,g694,g43,g941,g1080,VSS,g1016,g1554,g1008,g690,g755,g698,CLOCK,g633,g1000,g757;
output g6269,g7729,g7287,g4370,g6425,g7292,g4657,g7425,g1724,g9310,g7285,g5684,g8234,g5143,g9128,g1798,g3860,g453,g6849,g8219,g6909,g7732,g7295,g5678,g6212,g1871,g7293,g9204,g2888,g7063,g3077,g1810,g2844,g6207,g534,g7298,g1017,g291,g3829,g1804,g3859,g6675,g9305,g7730,g206,g6850,g7103,g4660,g7731,g785,g8661,g4371,g1006,g7291,g7283,g3096,g1824,g4664,g4655,g4661,g7294,g6236,g5682,g9297,g9280,g7508,g1894,g8872,g7286,g8958,g7505,g9299,g6223,g1783,g4267,g9378,g9314,g1944,g6895,g3191,g6648,g1829,g7514,g8663,g4373,g1817,g7474,g7506,g7289,g7288,g6653,g4316,g7423,g7424,g8216,g5164,g5571,g1015,g1911,g7504,g3159,g372,g7290,g1246,g7048,g5729,g9132,g4663,g9308,g7507,g9312,g8218,g3130,g5669,g2662,g7284,g594,g8217,g1870,g4372,g5687;

  wire g998,g954,g9070,g6367,g7021,g4181,I11638,g9219,g7535,g98,g2896,I11696,g9113,I10834,g3462,I5942,g7071,I15263,I7478,g3964,g3993,g8464,g4908,I9573,g8812,I6998,I12158,I13376,g6462,g4746,g4810,g6264,g4313,g7593,I13320,g556,I12370,I13054,I8480,g5253,g1864,g6103,g9238,I15112,I10313,I5692,g4407,g9177,g4392,g2652,g9088,I6853,g4792,g6070,I14492,I15285,g5750,g5550,g2497,g6704,g7695,g543,g606,I14637,I15225,g1176,g3931,g758,g5121,I13478,I6003,I13088,g8792,g7164,I12927,g9182,g7632,I9059,I7504,I7517,g7719,g9319,g7992,I13794,g7119,I10320,I7568,g8639,g4891,g6604,g7113,I10678,I15082,I7512,g2905,I7688,I12776,I9745,g6997,I7618,g4585,g8076,g2895,g4622,I10062,g100,I11515,g7129,g901,g2768,g1375,g3880,I9597,I13284,I15102,I8904,g1643,g1960,g1576,g3995,I15040,g6782,I6103,g9137,g2887,g270,g8776,I14142,g2039,g7142,g2645,g2903,g5079,g8851,I11701,g7537,I8775,I8461,I11115,I12033,I6078,I5667,I14257,g1586,g7319,g6055,g6342,I11170,g7042,g6706,I12451,g6387,g2514,g7242,I15041,g7749,g6713,g9372,g1037,I5515,I15589,I5555,I10409,g456,g5345,g1416,g9361,I9271,I13570,g8832,g2651,g7090,g1597,I10256,g6979,I14009,g7337,g3890,g2916,g3219,I6198,g9011,g3700,g2330,I9278,g4305,g2923,g3761,I12229,g5412,g560,g1745,g5786,I13293,g4424,g1578,g6254,I7107,I7626,I7702,g4098,I8436,g4312,I14015,g5521,g5753,g6739,I8472,g6073,g5236,g7513,g3061,g5335,g8239,I11004,I6471,I7978,g4360,I8751,g3805,g6708,g5598,g8279,I7353,g6774,g6182,g1378,g2650,g4258,I8218,I12062,g4795,I5766,g9317,g6489,I7995,g8863,g6517,I6574,I7140,g3,I9525,I10277,I11227,I11494,g6890,I14996,I6239,g4517,g5104,I5812,g4801,I8925,I15065,I7792,g5511,g9003,g4131,g8267,I5401,I13707,I5598,g6554,I14448,g7754,I13388,g5052,I8730,g6837,g8758,g2206,g4414,g8686,I9148,g7598,g8174,g1975,g2970,g1276,I15897,g4841,g3778,g3919,I15651,I10758,g8889,I8064,g4114,I15222,I10078,g182,g8276,I6959,I5562,g2256,I6741,g5145,I12080,g6709,I15985,g5310,g4400,g8013,g4364,I14374,g4363,I10360,g1390,g1240,g8915,g7887,I13347,g4707,g5484,g2490,I7931,I8877,g4721,g4800,I15933,I6815,g8154,I10744,g7101,g1225,g5493,I7156,g7548,g4662,g2674,I12328,g6135,g5169,g7753,g2547,I14712,I13438,g2699,I15229,g1244,g1205,g2927,g4580,I7964,I9493,g9039,I7036,g8886,g8795,g9031,I8072,g5037,g4673,g2360,I7588,g5395,g6177,g1114,g8301,g3666,I7302,I6440,g4589,g9239,g6224,I11659,g9126,I7386,g7066,g4399,g4492,g1214,I12226,g5148,I5599,I10154,g7779,I12065,I12577,I15400,g6601,g3997,g6647,g7082,g4362,I8071,g3840,g8072,g6949,I6860,I5901,I10393,g1197,I13595,g587,g553,g4272,I13122,g6027,g6466,I6220,I8607,I15577,g6796,g5022,g9234,g6327,I12173,g4685,I10072,g4631,I10451,I14370,g812,g3753,I10144,g5116,g724,g13,I13903,I8432,I12316,g8460,I6012,I9947,I11206,g4836,g8262,g7536,I7752,g5364,g6403,g7196,g1665,g4719,g3095,g8300,g9025,I9636,I15720,I13617,I11758,g4242,I13822,I10847,g4560,I7186,g8808,g9362,I14403,I10705,I12523,g8331,g7273,g8981,g7269,I9383,I11116,g3935,g3085,g1571,g2208,g5088,I13487,g5642,g7700,I11725,I12996,g3500,I13271,g3858,g8363,g1537,I8709,I11272,I9534,g113,g2283,g4445,g2995,I9350,I10196,g6520,g8087,I16180,g8306,I8523,g1025,g478,I13583,I10565,g2128,I6051,g5697,I8328,g3225,g6056,g5284,g2242,g252,g2904,g5683,g5467,g6572,g2246,g775,g999,g7259,g7190,I6814,I10356,g11,I14166,g3963,g6418,g1399,I10649,I14285,g6416,g2177,g3561,I12779,I9310,g5751,g2149,g436,g765,g3937,g5662,g6923,g8852,I14857,g4785,I11156,g5167,g1308,I12564,g1868,I9837,g9054,I7804,g8691,g3750,I7811,g1541,I11485,I16138,g3911,g5009,g3577,I6757,I15814,I10439,g2393,I7928,I14739,g1562,g9002,g5089,I15726,g6859,I15909,g5278,g6966,g1646,I11109,I12629,g5291,g8510,g9214,g1409,g8736,I12598,I7148,I9774,g8315,I6075,I15881,g9112,I13396,g8861,g6380,g435,I16006,g5246,I5706,g4613,g8754,g4051,I8658,g4246,g7243,g6357,g3578,I5709,g6600,I13801,g1977,g6990,g5068,g5154,I13213,g3869,g7751,g4626,I10292,I15741,I10298,I14844,I8766,g7217,g4658,g9143,I12376,g3512,g7741,g8280,I15705,g741,I10538,g6715,I6733,I8053,g1364,g8772,g8701,g7317,g6676,g6366,g5157,g7007,I9935,g8919,I12400,g1393,I8618,g1918,g1676,g4690,g1886,I13825,g4832,I11479,g6371,g8089,g4552,g3640,I5577,g4647,g8238,g2890,I10675,g5057,g246,I14932,I6925,g3641,g5475,g6424,g9010,g7127,g9159,g5149,g7344,g9038,g1935,g4229,I9535,g5610,I13003,I15830,g7712,g5814,I10901,g7610,I9081,g2386,g5800,I15604,g1787,g3908,g4448,g1575,I12295,I8502,g7067,I8865,I15842,g642,I12454,g5802,I16165,g77,g9101,I12460,g6362,g1958,g5626,I8255,g2920,I14061,I10080,g1126,I13638,I13764,I10243,g6593,g5587,I5471,g2821,g8362,I14457,g6287,I6676,g9099,I7558,g4676,I10998,g7256,g4525,g4900,g4539,g4182,g4422,g4228,g4220,g4646,g1382,g2267,g4352,I14187,I14801,I15583,I6428,I7277,g4905,I9681,I5365,I13281,g3918,g625,g6438,g4739,I6774,g7466,I16154,g9072,I15625,g6415,I5657,g5690,g5813,I13547,g4320,I14001,g3491,g5784,g7340,g1779,g7527,g1318,g4048,g8266,I9624,g83,g3560,g109,g6130,g4111,I9177,I5923,g5401,g8199,g7615,I8108,g4526,I7885,g4540,I10790,g5025,g6695,g8759,I13927,g3949,g9369,g4888,g1195,I5559,I7118,I16173,g4268,I10166,g7102,g4227,I6233,g114,g2404,g8073,g9386,g8093,g6337,g6992,g6285,g1805,g5463,g4884,I8529,I8215,I13758,g5644,g5514,g8970,g5760,g3079,I8793,g3870,g9208,g1772,I13502,g1327,I9963,g3654,I12924,g8976,I14175,I9515,g5234,I11135,I10350,g604,g4559,g1776,I8589,I13350,I8115,g1816,g6069,g2325,g1253,g7775,g7134,I14046,I7778,g6323,g6892,g7276,g5069,g7517,g8882,I15262,I7838,I10204,I13335,g9102,g8483,g1923,I16161,I15007,I11308,g859,I13359,I14623,g4328,g7094,I12712,I8935,I13332,I14442,g3528,g4907,g5758,g4202,g7522,I12832,I10574,g4074,I8581,I11747,I13663,I12170,g9291,I11958,I12421,I5600,g9258,g7061,g2933,g5343,g2312,I7575,I12217,g2647,g1725,g7777,I11549,g8146,I12391,g2014,g6196,I11525,I5383,I11191,g6221,I9158,g6119,I12424,g8545,g5817,g6887,g5061,g7265,g2924,g303,g3844,g5054,g6673,g4254,I13362,I9502,g7092,g2392,I11867,I14088,g4456,g8977,g5576,g1887,g2383,g7583,g6651,g2477,g9044,g2992,I7308,g6215,I6134,g2051,g8753,g7717,I6457,g2309,I11335,g2329,g4590,g1186,I7539,g1348,g8583,I8446,g6209,g8648,g4001,g2926,g774,g8152,g4793,g6515,g5627,g7742,I7486,g5599,I15522,g9247,I7262,I7180,g6918,g8605,g2104,I6904,g4283,g4016,I8109,g4353,I12635,g1806,g4052,g6743,g4871,g7309,I12948,g2044,g9212,I7101,g7829,g1226,I11353,I10552,g2057,g4469,g3492,g4082,g4609,g5653,I5374,I6087,I7332,g5210,I10981,g4538,I15274,I6036,g4870,g6198,g8734,g8689,I6112,g3499,I11627,g6661,g6228,g6412,I6669,g9142,g6983,g6559,g6015,g6074,g7503,I7347,g1254,g5917,g3904,I14127,I10626,g973,g3078,g6193,g6652,g5713,g825,g6111,g5190,I11880,I14816,I12385,g4236,g9381,g8702,g7083,g4603,I9363,g121,g1585,I11037,g778,g3967,I10491,I13422,I13057,g513,g5046,g1243,g7202,g6496,g8995,I10125,g9019,g3798,I14807,g8802,g6266,g7405,I8998,I12538,g8263,g6841,I6015,g9210,g8543,g766,I8665,g6429,g6158,I10953,g4936,g1211,g3779,g7299,I11164,g5126,g8667,I13509,g8683,I15863,g1815,g521,g7592,g4276,g665,g8228,g7733,g1154,g6242,I8264,g6741,I8772,I10336,g4088,I10569,g4302,g6336,I14231,g7188,g9322,I6864,I8354,g7585,g4134,I5751,g1781,g9118,g6639,I14067,g4553,g6273,g4476,I14199,g7160,g4712,g6751,I12466,g9158,g4308,I5682,I12268,I15937,I13669,g216,I11034,I5975,g6781,g4385,I12247,I11371,g6664,I11437,g6325,I12187,g8290,I11079,I8268,g2780,I9116,g4032,I7551,g8875,I6305,g5767,g7144,I7233,g6769,g30,g3857,g5971,g4096,g6912,g5608,g8931,g1415,g4387,g3925,g8858,g4013,g5163,g4915,g632,g6616,I13305,g8307,g6395,g5085,g5101,I11835,g2265,g9379,g8295,g2573,g5746,g4901,g7024,I11425,I8040,g395,g3555,g6019,I15580,g348,g6088,g2793,g5265,g6855,g3525,I14424,g4623,g5221,I14413,g9357,g5570,g5203,g1799,I8874,g6714,g8988,g8230,I5646,I11821,I6826,I14904,I15519,g6632,g4524,I15484,g2239,g3505,g5432,g1199,I11803,g4490,g7356,g3842,I9463,I5894,I15315,g3984,I8895,g3991,I10479,g6332,g3951,g622,g6976,g4179,g6800,I13587,g4612,I15507,I14959,g7049,I12514,I6258,I8058,g6947,g2626,g9052,g5028,g597,g4050,g2209,I8357,I11165,g8755,I6834,g8608,I15423,g6117,g5178,I11497,g1372,g3314,g4303,g1961,g7532,g7041,g2989,g1695,g408,g2605,I14058,I11488,g1477,I6232,g7107,g4571,I14780,I12301,g8628,I9769,g8738,g8951,I15616,g4575,g4038,g7239,g8957,g6457,I8243,g7282,g3952,g1311,I5478,g4724,g7519,g2229,I16046,I7087,g8681,g2480,I8326,g612,g7018,g8857,g28,I13740,g7147,I15953,g1566,I10810,g7745,g2487,g6752,g5189,g5152,g4078,I10448,g4319,I11890,I12111,g9311,g3956,g2900,g6156,g7429,I11929,g7209,g7157,I11796,g1987,g4654,I10295,g4917,g5821,I15918,I13314,I15824,g1185,I12499,I15113,I14294,g6283,g6640,g8066,I9570,g6952,g6898,g5938,g9148,g4813,g5055,I8814,I15433,g3567,g6426,g2308,I8739,I15803,g4700,I11122,I11380,g6065,g7058,g953,I6680,g4962,g6822,I8537,g7079,g5490,I15251,I15672,g7791,g443,I11964,g8265,g7676,g4687,I15075,g94,g2324,g4744,g4351,I8245,g6038,g7151,g5704,g3929,g2769,I6820,g611,I12205,g7633,I15501,g5515,g6319,g5397,I5855,g1687,I6949,g4710,g1792,I11299,g1663,g8684,g6589,I15574,I10259,g8773,g7114,g2827,I6060,g8229,g7040,g2986,I10889,g3866,g874,g6761,g4689,g8820,g2833,I11981,g8319,I11149,g5299,g213,g7436,I7987,g8983,I9615,I15717,I13734,g6595,I11773,g8718,I13912,I15043,g5840,I12418,I13490,g5830,I15165,I10780,g6621,g2671,g6312,g6888,g8268,I6341,g609,I13599,g4922,g6275,g7528,g3865,I7953,I13444,g4621,I5407,g6566,g6470,g1098,g4006,I5410,g4806,g4464,I9785,I10681,g9282,g5824,I10289,I10361,g8270,I13588,g5988,g5053,g7833,g1748,g6299,g7780,g2470,g4572,g7308,g6087,I8835,g4421,g4486,I14214,g4969,I15340,I13858,g6818,g5147,g4101,g3980,g3693,g3259,I8543,g5559,g4287,g4430,I7179,I10488,I8980,I7278,g6962,g4873,g8787,I14139,g6013,g3898,g118,I14838,g7470,g9244,I8315,g9021,g5578,I10882,I5413,g2326,I7480,I6431,g1685,g6625,g8641,g7296,I11751,g7115,I9419,g6138,g2454,g6334,g4396,I13308,I8932,g3913,g1690,I12951,g1189,g6975,g3846,g300,I10826,I15708,g6180,I10702,g5204,g4437,g7607,g6392,g5071,g8703,g7783,g9279,g6295,g6716,g8704,g5108,I11858,g9363,g6920,g9248,I8477,g7520,g4197,g339,g8814,g1872,I10639,g2271,I16148,I16020,g2353,I9103,g4010,I15631,g9300,I8140,g518,g1808,I13869,g2957,g9097,g2105,I15702,I15613,I10694,I8202,g6278,I8471,g7937,g2909,g5207,g7826,g5334,I6839,g5438,I12915,g4624,g9111,I8449,g134,I11591,g92,g834,g6391,I15417,I9182,g62,g4146,g3938,I7635,I10874,I12696,I15510,I16023,g4130,g374,g5588,I16142,g7335,g1564,g5064,I11550,g6033,g4123,I11851,g8296,I12052,I11458,g5367,g8153,I7956,g6195,g7652,g7653,I12481,g6028,I15888,g2825,I15205,I14342,g773,g8902,g6204,I9222,g8880,g6361,I5763,g8181,g5443,g5317,g3429,g6658,g3086,g9096,g1462,g2709,I14725,g8751,I14260,I15169,g9,g3886,g3921,g6175,I6813,I15231,g8443,I15072,g1814,I5960,I5847,I7365,g8585,g7123,g7497,g6315,I11740,g2367,g2623,I10442,g7702,g6147,g1192,g4124,g3754,g1737,g4960,I14677,g8722,g8899,g6737,g3855,g6244,I14291,I12271,g1146,g8652,I11622,g48,g3502,I15184,g1744,g535,g5783,g4814,g5435,I6784,g8807,g5969,I14662,g677,g4958,g7757,g4829,g8905,I11158,I15533,g8940,I6887,g631,I10919,g6524,g6904,g9029,I8006,g7324,g1750,I10128,I13894,g7245,I11401,I12517,I9752,g7834,g6258,g8078,g3260,I8938,I5989,g8581,I7899,g5474,g9013,I6024,g1220,g7983,I14305,g9092,g1454,g2348,g979,g8173,I11305,I7255,I13373,g7654,g6230,g9133,I13106,g6995,I5984,g5716,I12646,g5492,g1795,I15178,g3784,I7870,I15052,g378,g4443,g9343,I15232,g906,I9910,g4608,g4080,g458,I13850,g125,I12597,g9327,g6803,I14055,g1658,I12025,g8198,g6624,I6242,g5844,g9255,I7269,g3944,I15950,g8336,g1782,g3920,I8660,g6974,g4097,g6373,g4026,g7037,g943,g4465,I15051,I6172,g9275,I11991,I13807,g5747,g7625,g6645,I7545,I12484,g3957,g6577,g1357,g8864,g8382,I13341,g3050,g4666,I10796,g1580,g3590,I15762,g623,g1007,g4033,g6994,I6072,g1649,I9233,g8090,I5389,g2327,I10300,g7495,I12202,g5568,g9105,I12993,g7253,g9022,g2359,I13541,I11884,g1853,g3338,I11239,g5005,g1387,g8835,g9026,g3966,g267,g6901,I16176,g7174,g6733,g4059,g3811,g6646,g1652,g2868,I13610,g9356,g8644,g1573,I8504,g3677,I13267,g2914,g6181,I11078,g9370,g5031,g2298,g2556,g9123,g2724,g2,I12725,g9211,g2655,I14531,g2712,g8441,g2843,g2969,g6879,I5831,g7498,I12906,I7738,I8363,g8998,I9132,I8956,g1130,I10807,g5688,g8155,I9057,I11936,g7578,g9049,g8846,g146,I9301,g5761,I7576,g476,g4022,g6538,g8092,g7509,I6894,g3013,I7882,g2314,g2352,g4895,g7411,g1005,I8254,g4436,g2664,I13979,I16151,g3875,g6106,g4037,g4263,g6109,g1231,g8340,I11018,I9845,g5001,g1310,I7706,g6146,g6488,g2616,I10516,I11656,I6302,I15388,g2979,g446,g1428,g180,g3838,I13419,I13885,g8804,g762,I16145,I7947,I8296,g7838,I5565,g4116,I12038,g7687,g2286,g8844,g4541,g8179,I15527,I5545,g4693,I12502,I6939,I7492,I7232,g4412,g1757,g5918,I6434,g4927,g6306,g7434,g8065,g4125,g7467,g8629,I10605,g7433,g9094,I14786,g4564,I11994,g375,g8231,g6321,g1896,g5592,I8613,g2361,g3933,I11136,g7582,g7614,I9089,g7554,I14674,I8637,I7417,g5781,g187,g8757,I12355,I10343,g8801,g8894,I6597,g9174,I15943,I8437,I8020,g6363,g1424,I13676,g6343,g1292,g5179,g3732,g7471,g4359,I10397,I7651,g9220,I9234,g9306,g4697,g9060,g1742,g6161,I11407,g951,g2922,I13533,g7496,I11389,g5093,g4089,g9198,g3002,I13639,g7320,g6172,g6844,g390,I6561,g3094,g7515,I12986,g6183,I10856,g7832,g8948,g714,g5693,g8222,g6698,g8273,I10643,g1812,g4638,I15230,g3972,g5596,g7604,g7132,g429,g6687,g7095,I15495,g9063,g5822,g1339,g8982,g8849,I9987,g1638,g5763,g2222,g3498,I11832,I12280,I13215,I9111,g5035,I8551,g4652,g6951,g211,g4636,I7150,g4288,g4601,g2347,g5565,I7422,g7001,I12154,I5428,I13635,g4265,g5525,g9161,I9684,I12403,I15062,g9233,I15765,I7595,g6793,I7380,I14264,g5099,g1395,I11662,g7683,g3614,g4020,g6490,I14804,I15956,I10433,I10454,g7274,g6408,g7227,g1826,g3871,g1379,g6218,I6192,g3970,g2275,g595,I12877,I9994,I14709,g4668,g6229,g3941,g5625,I6805,I11616,I15054,I11787,I11025,I11491,g8256,g6005,g4928,g9261,g7736,I9579,g1385,I14388,g4547,g5606,g8643,I7041,g1955,I9520,I7453,I11556,I10924,g8291,g4736,g3226,g7234,I8308,I8859,g9047,g4732,g6798,I12930,g7627,g6279,g7413,I15657,g1029,I10973,g8272,g8609,g162,g7553,g2510,g2323,g7697,g9048,g1252,g8017,g1149,I14234,I10867,g940,g2818,g1354,I9630,g6308,g6463,I11110,g6104,I13261,g3906,I6425,g2891,g1681,I7844,I8273,I12669,g3075,I14643,g8656,g7170,I10506,g142,I11522,g2944,g6915,g459,g9067,g5623,I10541,g1069,I11395,I14273,g4532,I8418,I12244,I13574,I14097,I10743,I7758,g8769,g173,I14079,I15962,g4081,g1549,g7275,I15298,I14942,g2902,I15696,g6406,I12592,g5699,g6179,g2889,g8855,g6289,g7441,g4463,g1778,g8008,g3768,I5512,g4036,I9425,g7750,g6297,g3706,g1819,g5823,g2074,I13425,I11443,I10708,g6257,g1312,g3934,g746,I14759,g8784,g1322,g8285,I9460,g6281,g5212,I12742,I13921,I14467,I8594,I8237,I7939,g6953,g2633,g7518,I15971,g4103,I14695,g7098,I7172,g9389,g8811,g6035,g4961,g6672,g1257,I6446,g55,g7511,g5529,g8777,I8823,g9199,I6274,g8128,g4651,g6662,g7765,g7587,g5741,g317,g179,g3926,g3316,g4335,I15053,g6905,I8005,g7159,g7772,I11939,g7480,I5386,I11151,I9633,g6643,I15974,g557,g9053,I12575,g8677,I13338,I15880,g2007,g4956,g6916,I15635,g1726,I9594,g93,g3982,g6776,g3996,I11790,g8634,g689,g9162,I15965,g4796,g7228,g2893,I12852,g6160,g3770,I13737,g7516,I11144,g6805,I12942,g7367,g3659,g3899,I10157,g3612,g2240,g465,I11707,g6856,I13882,g7770,g3540,I10315,I12891,I12496,g8631,g2282,g6170,g8442,g2262,g9191,I11377,g4252,I6267,g9334,I12550,g8360,g7725,g4411,g7169,I8483,g3527,I10224,g771,g8711,g261,I13589,g41,g9230,g626,I15308,g7226,g9036,I5772,g6133,I8787,g5127,g8341,g9034,g5481,g7445,g9366,I6831,g4741,g4425,g2016,g5091,g6105,g5518,g652,I8612,g6359,I12265,g8665,I7749,I7788,I13323,g6052,I13622,g8960,g4121,I13773,I15147,g2554,g8651,g5082,g1030,g1377,I13962,g8693,I6463,g855,I8455,g3978,g2389,g2906,I12737,g4677,g4378,g8791,g3519,I11843,g7254,I5911,g5314,g5160,g314,g7766,I11177,g3657,I14005,g8833,I7126,g6611,g4619,g6967,I11704,I14831,g6439,I15638,g3187,g4882,g4543,g888,g8748,I6273,g1857,I13066,I14338,I14245,g8709,g6414,I11729,I11793,I7548,I13524,g6833,g1863,g4327,I12933,I8052,I11757,g4475,g5648,I10421,g7260,g8922,I10535,g2866,g8974,g6778,I13244,g6188,g3910,g3617,I5969,I11920,g5787,g1499,I11186,g6724,I8288,I12003,I12903,I14416,I5715,g2268,g8524,I15848,g8715,g580,g4358,I10142,g629,g3739,I10739,I12463,g4653,g6934,g6054,g2334,I15898,g3862,g8892,g1319,g3083,I9760,g8710,I13628,g5643,g6505,g9185,g6145,I16055,g6617,g2660,I15073,g4417,g7574,I7526,g4035,I11172,g4200,I6636,g7538,I10334,g3851,g4483,g2873,g7145,I9209,g7360,g3633,I6018,g7302,g6945,I11278,g3084,g4632,g6305,g4839,I13631,I6422,g8845,I7149,g3780,g6963,g4642,g1974,g8873,g8015,g4903,g4376,g5006,g8311,I14202,g6683,I15405,g23,g7054,g5633,g8236,g610,I14100,g1304,g4511,I11080,I14052,g789,g1878,g1371,g1707,g2106,I13469,g730,g6004,g4119,g768,I9243,g6265,g2878,I5939,g8059,I9235,g4285,g4563,I8282,I7667,I16100,g7176,g3233,g3656,g8666,g8921,g6112,g1245,I11680,g8898,g6398,I15592,I14106,g4748,I7683,I9567,g1363,g1866,g792,g9109,I6057,I13605,I10804,I9993,g1800,g6397,I11641,g4885,g1084,g530,g5214,g7355,I14427,g1877,g6944,g6037,g6939,I6254,I15202,g4634,g1934,g5228,g1202,g2401,g80,g5151,g5013,g7303,I8642,g8664,g5765,g2945,I12493,I6916,I15475,g8818,g145,I13816,g7177,g6858,g7240,I8392,g3877,g628,g5478,I14969,g7588,I11732,I14789,I15978,g8339,g9209,g5176,I6118,g2584,g9062,g6075,g8768,g4869,g2972,I10457,I12684,g6978,g5789,g4812,g7580,g4266,g6474,g8287,g2394,g6036,g2397,I8029,g5124,g3604,g7015,g6511,g6696,g8329,g1329,g293,I13017,g4633,g4190,g8658,g6163,g8669,I13701,g5759,g4616,g8972,g4696,g9129,g3390,g5552,g7350,g5165,g6320,g7904,I13403,I8588,g8912,g5201,I13035,g1701,I13140,g2214,I7599,g1637,g5402,I10380,g1396,g1266,g5607,g7347,g6862,g4923,g5546,g1860,g5000,g5259,g7426,g9076,g3960,g6780,I11718,g8640,g432,g8381,g2954,I7104,g7755,g5081,g2363,I13770,I6354,g6471,I6800,g9183,g3008,g3999,g5512,I6121,g7186,g4924,g6294,g9330,g214,g2659,g617,g8563,g1194,g8942,I14238,g9203,g2371,g8067,g9201,g7225,I10522,g7836,g9200,I12475,I13099,g7233,g3831,g6925,g6091,g8770,g6154,g2862,I12277,I7888,g5032,g8939,g3712,g3258,g9093,I12415,g4107,g9035,g6330,g1832,g6996,g1753,g8172,g6787,g4044,g6816,g4592,g1545,g3012,g7205,g2644,g6622,g6758,g7149,g4695,g2555,I12409,g6606,I5868,I8180,g5440,g4824,g6523,g6686,g6688,g1751,g6121,g1682,g8907,g8706,g1784,g3049,g7529,g8933,g8668,g6948,g8523,g4497,I8143,I15334,g4963,I9064,I10786,g6318,g4606,I8808,I13241,I10071,I7317,g7740,g4656,I14288,g2976,I13189,g588,g9304,g4738,g8771,g46,I11686,g5970,I14267,I11942,I7781,g1367,I15239,I7368,g1376,g4069,g7087,g8385,g8799,I15175,g7422,I7864,g969,g7106,g4105,g7551,g3466,g6853,I10143,I15290,g891,I10646,g6873,I10485,I8412,g3948,g6775,g6459,g7563,I10842,g3517,g9004,g3557,g7222,I6686,g8303,g5137,g1431,g2235,I13698,I11974,g3642,I9196,g7267,g9350,g2479,g235,g4275,I5926,g6692,I7115,g1325,g3802,g4930,I13451,g5205,I15504,g3691,I7362,I6102,g1879,I14839,g5752,g4380,g8632,g5362,I15855,g6794,I9938,g5458,g8867,I12180,g4110,I14463,g4743,g4394,g1402,g4567,I6090,g8778,g6291,g3093,I6096,g2384,g5074,g2349,g4025,g2424,g6399,g1572,I11374,I8957,I10460,g6801,g6812,I10387,I15291,g2345,g5208,I8583,g6900,I9484,g7705,g2533,g6860,g7715,g8790,g5141,I9041,I9070,I6509,g4883,I8977,I5957,I9907,g2863,g9218,I15530,g1844,g7104,g9315,g5539,g6580,g1193,g4912,I6963,I7564,g3912,I8517,I11203,g1773,g9388,g1326,I8133,g6009,g4357,g6018,g3533,I8452,I6148,g7586,g393,g6861,g8293,g2043,g5040,I13060,g4176,g6011,I5997,g1780,g7589,g5437,I11933,g1590,I10403,g6630,g6390,I6186,g2794,g2774,I10151,I12232,I13051,g7761,I14378,g579,g2901,I6856,g6760,g1908,g6263,g4811,I9499,g1674,I9794,g4196,g5472,I14109,I8166,g3649,I9162,I16052,g3358,g5216,g3947,g4147,g4216,g313,I8817,g8337,I10627,g9015,g6937,g6928,g9313,g4921,I9558,g2943,I15571,g8016,g384,g1600,I6257,g2224,g7591,I12757,g7693,g3539,g8284,I11320,I5872,I7755,g4094,g2752,g3589,I7338,g1830,g4823,I15940,g8992,g9125,I13713,g6819,g7759,g4453,g4296,g8562,I8520,I10225,g2939,I13302,g4244,g7550,g4232,g5073,g5113,g5396,I13231,g1204,g6409,I6064,I14325,I14941,g6322,g2310,g2495,g1156,I8853,I9892,I15085,g4186,I13258,g24,g5117,g6249,I15899,g2837,g5302,g5023,g5112,I7658,g2973,g2925,g8323,g9316,g9240,g929,I12508,g489,g8836,g602,g1794,g591,I11827,g6809,g6197,g2215,I13692,g8879,g7064,g1196,g7837,I9171,g3313,g1758,I11028,g7,I12181,I10274,g1421,I13496,g4245,g4454,I9443,I9834,g6164,I14246,g9179,g6251,g8042,g6003,g8767,g5726,I10463,g6745,g7688,I9021,I8536,g3506,I11341,I8132,g2932,g7156,I16119,g4053,g8785,I8339,g945,g4021,I14279,g3819,g7235,I12319,g5769,I11575,g4808,g566,g6956,g4640,I15492,I8119,g7336,g200,g1813,g1948,I6323,g4799,g4513,I8820,I11251,g486,I12349,g7039,g6040,g1760,g8334,g9193,g5029,g6789,I6054,g3903,g5076,g6813,I11917,g2162,I6270,g1555,g601,g8775,g6891,g4554,I11163,g5649,g6050,g2520,I6251,I15190,I8844,g5114,g3897,I15924,I14436,g2949,I15990,g4913,g5264,I6911,g5487,I12643,g3922,I10836,g9222,g772,I11143,g5192,g7116,g2221,g5072,g4314,I10946,g4916,I5371,g6594,g6256,g4273,I11562,g8225,g7301,I11467,g699,g1983,g6437,g8440,g9146,g212,g9205,g4153,g202,g4704,g8859,g1158,g1926,g6635,I8769,I8907,g4611,g137,g8911,I9142,g9104,g4635,g7416,g3124,I6695,g3264,g8638,g4583,I10250,g6211,I11117,g6871,g7323,I7540,g7601,I13072,g2539,g1889,I14157,g7599,g8971,g5159,I8784,g5701,g6927,g8997,g2351,g4253,g4627,I7856,I5954,I8910,I8001,I13416,I10848,I8057,g5285,I12649,g1568,g7139,g5845,g6447,g4030,g3979,I6170,g2880,g5698,g479,I8105,g7763,I7157,g9082,I9561,g5171,g1581,g5725,I16107,I6764,I9675,I13134,I7800,I10247,g4225,g7626,g2546,g7721,I14178,g6046,g2548,I12124,I10223,g5517,g4573,g6293,I13031,g3873,g6571,g1680,g7016,g4684,g4444,g8069,I15020,I15240,g3530,g2270,g8969,g5768,g5187,I9827,g2654,I7648,g5150,I15839,I11014,g5036,I6776,g6062,g5059,I9531,g8131,I6104,I12015,g970,I5636,I13565,g1775,g9016,g2460,g831,I10494,g2637,I13544,g3883,g6238,g6872,g2816,g2743,I6723,I12999,g4918,I9954,g5668,g2343,I16058,g9339,I7423,g287,I6522,g5007,I10327,g6482,g5468,g7716,g5736,g7428,g2096,g8622,g222,I12976,I7617,g3787,g4931,g1768,g8176,I11242,I14318,g8328,g5696,g2291,g1092,I12307,g7345,I13837,g6326,g3959,g3743,g4581,I7377,g4503,I5605,g1519,g9144,I7859,g4219,g4317,g7762,I5609,g1087,g1673,g972,g8947,g7315,g5581,g7494,g2452,I15010,I7520,g32,g2100,I7195,g5222,I6133,g8493,g8837,g7255,g896,g7162,g6060,I12373,I16061,g6731,g5674,I10868,g6884,g1153,g1807,g5041,g8944,I8573,I14244,I10198,I5839,g681,g7420,g1736,I16072,g5740,I7443,I11069,g5583,I6657,I14042,g2223,g5156,g5094,I7655,g1582,g8721,g5547,I8962,g1679,g5689,g533,g6432,g2145,g6155,g5015,g2832,g6755,g4957,g417,g6834,g950,g7003,g6370,g3192,I10011,g9298,g1924,g278,g984,g9307,g875,g6885,g8457,I13023,I14064,g9055,g3822,I9145,g2677,g210,I9591,I14112,g6232,g8403,g3939,g6284,g6674,I5419,I6703,g4361,g6452,I14219,g5708,g5874,g7602,g9178,g6984,g1856,g4535,I13562,g6542,I10469,g8946,I7241,g5764,g2629,I10268,I15172,g8705,g4079,g5220,g6628,g6227,g4092,I9018,g7552,g2292,g1565,I8760,I12520,g3131,I6163,g4598,I11184,g510,I7807,g5452,g2783,I9407,I15211,g4369,g258,g2380,I9123,g4733,g936,I12286,I7981,g3680,g1324,g3882,g7014,I9466,g2665,g7263,I7145,g3988,g3893,g7210,g255,g2929,I13888,g1321,I11368,I7069,g2615,g5232,g8749,g9320,I13786,I15032,I14828,g6764,I15429,g86,I7216,I8486,g9085,g9213,g7597,I8244,g6369,g8333,g5818,g4787,g3529,g7595,I6956,g5193,g8943,I12059,I13897,I6033,I10472,g6783,I7762,g58,g5737,g1288,g4825,I6416,I15071,g1897,g2368,g4747,g9050,I7293,I10982,I11722,g6460,I11984,g1045,I9612,I11759,I12412,I14680,g8309,I7436,g4835,g4566,g1504,g8984,I11470,g4579,I10862,I11245,g3310,g7606,g5058,g4015,I8097,g1803,I12490,g7122,g2622,g3808,I9918,g3705,I7296,I11841,g5469,I14822,I8850,g6627,g2892,g3930,g183,g2313,g5482,g7546,I14193,g2253,g3692,g6597,g8906,I15759,g4521,I13353,g8760,I15862,g4904,g6311,g6552,g8611,g4122,g9294,g9124,I11824,g4332,g8938,I7676,g5287,g6444,g6866,g9140,I8945,g5700,g6267,I6130,I11344,g596,g8986,g6153,I8745,g234,g8930,g480,g6867,g477,g8823,I10597,g3867,g2810,g2761,g4239,g8949,g3900,g296,g1270,I6924,g815,I12085,I7662,g4502,I15833,g6205,g4919,g237,g2934,I6454,g7221,I11266,I13731,g6941,g4142,g2225,g7714,I14489,g4545,I7044,g7744,I8327,I9585,I5654,g9014,g4000,I10555,g4408,g1774,I13435,g6377,I8011,I10377,g3879,I12274,I14397,I13277,g7704,g4398,I14753,g8029,g5312,g658,I12813,g9202,g5566,g9221,g576,g411,g1370,g4879,g761,g6562,g6840,I13672,g9331,g2232,g5639,I10937,g7782,g5021,I15030,g6839,g605,g4084,I9099,g7009,I12367,g8383,g4379,I7680,g457,I13329,I16033,g7658,I11926,g7311,I15675,g6032,g6681,g507,I13048,g9068,I13997,g5065,g1398,g5558,I6333,g3605,I8552,g2522,I11197,g8779,g4306,I12117,g3635,g4745,g6581,g6744,g8685,I6460,I8394,g3548,g3562,g3962,g2689,I10558,I9446,g7549,I12176,g7603,I13749,I8781,g8380,g1122,I16036,g7163,g3965,g5811,g9353,g7764,g583,g7342,I9747,g6991,I9382,g7252,g1439,I12436,g5551,g1134,I7329,g321,I11233,I12897,g2344,g6435,I14381,g8330,g8909,g4163,I7902,g2091,g4027,I14169,I8209,g3992,g7487,I6124,I10079,g7758,g6379,g6006,g3849,g6456,g5624,I10384,g8980,I9678,g6699,I10532,I10172,g7446,g7488,g4315,I14251,I6540,g4968,I10770,g4159,g6717,g9333,I15199,g377,I13865,g7442,g2919,I10690,g616,g5894,g405,I7905,g4734,g5107,I9645,g8774,g275,I7867,g4692,g9075,I14130,I16090,g8989,g3503,g4577,g1952,g7100,g3587,g95,g2911,g944,g8297,g5790,I6532,g6659,I13828,I16135,I11806,g8305,I10427,g6763,g2202,g6137,g5717,g6446,I15693,g8458,g5123,g3650,g6237,g6178,I8547,g6203,g4100,g8584,g2273,g8741,g4118,g5617,I15565,g7738,g6510,g3190,g4343,g6274,g7316,I14227,I14208,g3563,g5807,g6186,g4193,I12953,I9170,g2982,g6372,g8377,I7323,g5460,I12529,I9657,I15543,I15241,I6905,I11998,I15254,I15770,I6758,I7445,I9242,I5757,g4735,g2234,g3943,g4185,I11955,g5706,g7539,I14070,g7068,g1738,I15732,I7723,I7421,g5613,g6970,g6472,g7120,g8679,g7611,g6848,g7110,g5199,g7361,g6277,I15228,g8660,I8338,I15849,g8856,g7711,g2540,g423,I6553,I8715,g8806,g7305,I7691,g6881,I6248,g2884,g5166,g3969,g6115,g1704,I9788,I11838,g1472,g1855,g5661,g6728,g9237,g6300,I12912,g8782,g108,I11586,g4249,I9955,g4892,g2966,g2245,I11398,I10519,g249,I7908,I5897,g3924,g9340,g8789,g852,g5542,g5243,g6051,I13012,g9355,g4366,g4887,I10908,I13161,I11461,g8888,I8868,I15426,g2233,I13613,g1368,g2015,g1435,g5785,g7722,g1280,I13484,g9349,g7330,g1667,g6917,I11142,g4742,g6742,g6210,I15882,g5096,g495,I8401,I15265,g3981,g1811,g2365,g7631,g5427,g7455,I15218,I14276,g8764,I10001,g2840,g9323,g7117,g7270,g8862,g3958,I12346,g4678,I8014,I9672,g504,I13695,g471,g4108,g3769,g1360,g819,g7178,g4091,I13378,g1392,g5686,g9360,g6618,g4226,I15553,I8847,I15776,I14743,g6136,I9692,g4395,I13600,I9325,g7182,g9216,g7594,g8731,g952,g6002,g1670,g7363,I6770,g1049,g8630,g8324,I8024,g8260,I10073,I12406,g8338,g8819,g4129,I10773,g8312,I6587,g527,g2672,g6048,g5444,g6382,g2883,I15017,g2985,g1467,g6838,g8321,I9768,I14657,g8332,I5754,g7088,g2502,g7349,I7629,g9188,g3853,I10745,I7082,I7505,g7790,g7187,g5654,g1945,g7112,g7739,g5516,g3520,g7307,g6376,g9071,g4493,g7010,g4604,I11455,I10849,g7510,I15681,I7400,g6469,g5197,g3188,g47,I11855,g9045,g7246,I9139,g5448,g2038,g2938,g7547,g201,I11506,g3029,g2453,g767,g4072,g6889,g2331,I14763,g9354,g1011,g4126,I12690,g6010,g7192,g3018,I6217,I12753,g2829,g5024,g8405,I7602,g3884,I6109,g1603,I7538,g5868,g6353,g8233,I6065,g2092,g8,I12193,g7359,g6799,g7034,I8164,g4297,I10430,I10766,g74,I7640,I13649,g4355,g7351,g4438,I12397,g1756,g4501,g6718,g3891,g7406,g6697,g8903,g8796,g3812,g6893,I8582,I9618,I9948,g1980,g7596,g2478,g3014,g1828,I14810,g8936,I8805,g2137,I9381,I15645,g5657,g695,I11428,I15536,g371,g7699,g8482,g8816,I9440,g8325,g6804,I14732,g9281,g1827,g7920,g4298,g5403,g141,g7756,g122,g6842,g7566,I12457,g4713,g4728,I10322,g1272,g6150,I8922,g3062,g630,g8378,g7334,I5781,I10952,g2184,g103,g3582,g6509,g8934,I8802,I8826,g6792,I9360,I16084,g3495,g6810,I15193,g1167,g1567,I13214,I8736,g1383,I11209,g1904,g4344,g1034,g6348,I11800,I13407,g5030,g8694,g3998,g8653,g5709,g3994,I15086,g1910,g3953,g9260,I14282,g7657,I9151,g3790,g7502,I10046,I14420,g1683,I6309,I9600,g6753,g1913,g402,g8091,I6740,g5039,g4880,g2877,I13209,g7031,I10466,g6478,I6917,I7950,g8987,g3946,g5672,g6120,g563,g1809,g45,g3028,g6851,g7784,g2471,I14603,I11323,I8496,g2238,g6282,g4017,I5817,I8428,I5356,g2734,g8544,g1217,g1852,g7417,I14687,I7086,g5491,g2879,I15324,I8413,g8147,g4455,I10390,g4706,g7326,g6458,g6972,I12763,I11971,g6682,I10321,I12909,g6999,g1777,g624,g2134,I12433,g2867,g5939,I7371,I12442,g7198,g6506,g7329,g1317,g2886,g6938,g9217,I11338,g6847,I13045,I15586,I14082,I14933,g7366,I11449,g8891,g3674,g8719,g4003,I7712,g3895,g7026,g8625,g7581,g1494,g7512,g2264,g6797,I11215,g3287,g1964,g3847,g6910,g8294,g2706,g4409,g4375,g8670,I7389,I8829,I14315,g8726,g4840,g9024,g1065,I6877,g1260,g5638,I9547,g5749,g10,g1430,I11066,I10197,I7305,g9273,g2375,g8955,I12088,g3076,I12022,g9157,g355,I6081,g5122,I9666,g655,g2506,g4595,g5742,g9110,g6824,g9278,g6094,I8190,g4482,g710,g1307,I6468,I9071,I8892,g2807,I13924,g926,I10509,g8713,g6508,g9241,g6483,I11257,g7070,g6473,g207,g8654,g2496,g8645,I15033,g4569,g6356,I7592,I12304,I7437,g5309,g1230,I7609,g6870,g8361,I11648,g6001,g5034,g6565,I11102,g4112,g1300,g1577,g3835,g5439,g6655,g4507,g3522,I15252,g7207,g1801,g5480,g5872,g8877,g6906,I14366,g6815,I11248,g8314,I12983,I11311,I8841,I6578,g5313,g9352,g9058,I12138,g8780,g2509,I11230,g6253,I13447,g1203,g8887,g9151,g6043,g9127,I11001,g8624,g8920,g2366,I11416,I13112,I10299,I15084,g7556,I8559,g1429,g4056,g782,g8675,I13499,g685,g5522,I10503,I14085,I14952,g8511,g5060,g7033,g1110,g2959,I8721,g7008,I11894,g6116,I6135,g8803,I7973,I15420,I12250,g6134,g6310,g8815,g2635,g7418,g6396,g5470,g9285,g4433,g5557,g172,I10625,g9095,g6108,g4168,g3783,I12888,g4023,I8659,g3928,g8950,I15273,g4789,g8040,g8890,g1616,g1012,I12511,g8421,g5083,I8727,g9116,g4231,g6843,g2870,g6344,g4403,I7797,g7682,g7165,g2625,g976,g6596,g7105,I6499,g7059,I13234,g1200,g3950,g6467,g4255,g7608,g7710,g1061,g5043,I5933,g8462,I10307,g4452,g4837,I6663,I13819,g7155,I16129,g6786,g1831,I7011,g5077,g38,I15498,g7136,g5180,g318,I13915,g2746,I7198,I9347,g6707,g2340,I10169,I12771,g6142,g1916,I7967,g7281,g6225,g6877,g4434,g9028,g1837,g7111,g4783,I7616,I10855,g5231,g6428,g8928,g9373,I14031,g769,g4139,g7038,g1247,g3976,I11332,g8953,I10366,g8075,g1384,g4354,I8063,g1313,I5732,g8082,g6445,g6465,g4256,g2824,g5562,g3652,g8728,g7437,g5593,I5432,g7143,g4702,g1524,I15711,I5542,g5569,g890,g6169,g31,g1345,g6599,g2174,g6875,I5398,g6235,g6262,I8635,g6612,g4011,I13653,I5879,I5519,g345,g3568,I16168,I11446,g1912,g4280,I12659,g6039,g9189,I13577,g7223,I15068,g1847,g7019,g8908,I5936,g5062,I14925,g2207,g4665,g2787,g4393,g6932,I7567,g6298,I15641,I9136,g27,g5494,I5506,g1579,g8965,g8606,g6823,g6125,g5087,g1155,g4629,g6971,I13506,g7266,g9087,g8316,I13876,g7691,g5433,I12965,g9181,g3511,I12958,g5217,I14980,g4166,g1584,g4681,g2621,I11350,g6605,g8994,g7524,g8745,I15791,g8512,g8881,I10280,I14964,I12292,g3848,g615,g8542,I9005,g5471,I15003,I8417,I5883,I12675,g8941,g6933,g8809,I7268,g1077,g4175,I15297,I14974,g6339,g6386,g2996,g8619,g5707,g9196,I12196,g4729,g2379,g6720,g2728,I7279,g4008,I9606,g9089,g6341,g5756,g6836,I6590,g5585,I5568,I7079,g6280,I13193,g6585,I10305,I15516,g5757,I7769,g5016,g5808,g8659,I10038,I12361,g5066,g4586,g4802,g3902,I13039,I11137,g8868,g8657,g2703,I6451,I9217,I6294,g7475,I14184,g5685,I14148,I10180,g2781,I15889,I12151,g1408,g6864,g7463,I8120,g6722,I10009,g4659,g4628,g6486,g315,g387,g7029,g6631,g4356,g3722,I6608,I12179,g4881,g4926,g1556,g5595,I11900,I13580,g6433,g7727,g5828,g6968,g7542,g7735,g7045,g9145,g5718,I6084,g6498,g9207,g6159,g4224,g2913,I9999,g5735,g2648,I9691,I12131,I8989,g8081,g351,I6006,I12687,g9346,g1041,g454,g5809,g7792,g7277,I7581,g2517,g8917,g5796,I6538,g786,g397,g158,g8838,g7771,g1869,g1752,g7776,g3521,g9367,g8895,I9539,I10028,g9083,I10253,g8602,g4615,g6351,I14025,I14136,g4104,g6475,g1909,g186,g5723,g5594,I11781,g4838,g5142,I8089,g7089,I12894,g9328,g5048,I8763,I9819,g7321,I9964,g5,g4264,g9084,g7224,g3091,g8876,I8351,g4342,g1746,g2971,g4740,g2764,g7698,g2947,g5049,g9023,g7208,g8798,I15391,I13767,I12968,I5359,I6115,g8762,g4388,g7521,g3047,I10980,g5286,g3222,g5477,g3735,I13250,g7056,g5209,g7109,g6384,g3531,g6578,I13118,I5521,g5254,g1919,g5363,I15699,g1509,g5086,I12448,g8910,I8511,g1148,g3315,I6066,I7632,g1967,I7452,I12008,g6768,g4557,g4701,g4639,g7724,g498,g7272,I7716,I5620,g9017,g8952,I8460,g7236,I15110,g6381,g1102,g1820,g6143,g6139,g8964,g2346,g6024,g6389,g5524,g6176,g4494,I6259,g4274,g3843,I6166,g5233,I11912,g7138,g7338,I15568,I12298,I6564,g2148,g4898,I15729,g7332,g8761,g5710,g6807,I6788,g2942,g5090,g3973,g7313,g3653,g5843,g8223,I15044,I15811,I12214,g5748,I15261,g5541,g4591,g8937,g6360,g2395,g840,g1842,g5219,I13787,g4649,g2782,I14771,I5789,g7333,g5835,I6437,g4031,I14430,g138,g5513,g6712,g6477,g7435,I9044,g5132,g5806,I10761,g8979,g3549,I8015,g6185,g6960,g608,I11410,g7357,g8080,I5368,g2285,g6762,I11302,g9371,I6326,g1843,I9476,I11043,I9603,I6376,g5230,I13299,g1405,g5033,g8991,I8643,g843,g3914,I11677,I10899,I8033,g544,g8805,g4670,g8744,I5416,g468,I10236,g6831,g309,g8968,g4614,I11961,I7029,g8407,g6638,g8800,g7449,g6303,g5269,I13755,g7006,I7561,I8754,g6614,I14754,g9321,g7557,g7306,g7268,I11864,g8690,g8275,g6732,I6202,g2501,I6849,g4542,g4250,g3238,g7080,I8000,g6464,g7810,I11614,I14813,g8283,g9215,g2940,I14133,I15019,I15850,I11897,g1073,I11710,g4584,I5920,I6160,I8127,g2180,I15595,g1147,I8898,g5100,g8359,I13196,I11809,I14646,g4368,g6555,g8612,g4536,g414,g6929,g7044,I14349,I15864,I15181,I6843,g4128,I7214,I10890,g7789,g2557,g5572,g9057,g8041,g7206,g5174,g356,g5680,g7023,I11365,g6553,I14485,I13761,g4777,g8281,g4605,g5739,g6152,I7533,I6443,g1888,I9025,I15411,g6168,g7768,g3221,g4610,g3556,g8610,g205,I13463,g4420,g7773,g7579,g2646,I8742,g4587,I10993,I15784,g5095,g6588,I10801,g3936,g6902,I10716,g2804,I11645,I5689,g2885,g3801,g7199,g9107,g4868,g129,g6629,g7713,g6586,g3872,I7139,I12223,g1698,g8317,g6167,I7290,g5195,g3887,g8327,I9194,g3983,I12632,I14330,I14439,I6752,I10094,I12044,g6288,g8304,g4830,I9202,g3465,g4568,g7499,g8151,g3603,g6736,g3541,g3850,I14121,g3940,I13719,g3777,I6474,g8932,g4127,I13704,g1163,g3830,g5070,g9139,I14792,g7339,g6730,g3854,g4117,g4132,g9359,g7541,g6911,g324,g5793,g3955,I10614,g6090,g4576,g2841,g5462,I7878,g5590,I7925,g5106,I15098,I11178,I7239,g5681,g3927,g1284,g7491,g4561,I7610,I5649,I13956,g9345,I7270,g661,g6059,g7331,I13797,I10271,g4935,g6958,g3579,g3723,g5526,g8635,g6657,I11778,g6068,g3968,g5238,g5425,g2263,g362,g9335,I11948,g7173,I12334,g706,g1166,g6845,I10190,I16017,g5453,g3977,g5825,I12571,g6957,g4333,g9223,g6955,g8896,g963,g6049,I5679,I8261,I11386,g7564,I12394,g4781,I10923,g7325,g6383,I12678,g4259,g4382,g1661,g5128,I11284,I12866,g4546,I16009,I15109,g5519,I12262,g2372,g990,g5846,g2963,g6649,I13413,g6345,g573,g5755,g6058,g3876,g7748,g5105,I15747,g5144,I10412,g837,I15031,g6656,g8626,g4158,I10286,g9100,I11362,g8647,I6791,g7050,g7870,g6829,g7743,g3915,I11683,g6365,I9261,g4087,g4120,g1563,g6440,I6759,g6913,g281,g3917,g4257,g5191,g9270,I6923,I8568,I11669,g7062,I12445,I14990,g6358,I11008,g9138,g9066,g3746,I6245,g297,g6385,I13365,g5772,I14951,g1394,g6314,g6693,g7523,g6907,g2960,g8175,I12128,g7180,g455,I13157,g7297,I8994,g6719,g4821,I12051,g8156,g2374,g8038,g6148,g5839,g8725,I14484,I13290,g8655,g7137,g8853,I10160,g5743,g4049,g6411,I10400,g7500,g6936,g8439,g3485,I9985,I11200,I15414,g703,I12364,g7787,I7138,g2931,I12068,g5140,g2276,g4286,g4620,g7774,I14028,g3524,I14035,I12551,g7689,g5294,g3716,I15539,g1797,g7692,g5679,I13472,g7443,I9621,I8277,I7938,I9038,I13383,g7966,g6507,I9422,g5658,g7193,g5258,g4192,g5611,I9979,g5162,g4311,g9302,g399,g6525,g6089,g1588,I7085,I8078,g6729,I10359,g6969,I8617,g6317,g599,g3878,g949,I9651,g7230,I7010,I12325,g5008,I15283,I15018,g2373,I13879,g5138,I6646,g4133,I7510,g6071,g3232,g8929,I5422,I12939,g3080,g7257,g6407,g3942,I11736,I15074,I10789,I6872,I15408,g5235,g2680,g5002,g6582,g8985,I10820,I15753,I6652,I13356,g5445,I13686,I12672,g6516,g5200,g6852,g2385,g4699,g6903,g3961,g104,g7559,g6497,g1686,g4057,I13103,g2700,I9396,g6346,g948,g3825,g6767,I12722,g598,I11326,I12854,I9582,g2614,g7028,I9126,g3588,I12532,g4426,g7022,g6461,I5908,g7181,I6716,g9077,g6141,I5676,g5268,g7696,g764,I8986,g7211,I12091,g2663,g1373,g1942,g8463,g5724,g4784,g4794,I12053,I15099,g536,I13873,g4914,g2354,g3630,g8235,g8978,g2642,I9076,I7454,g6785,g7318,g5812,I15250,I8150,g6012,g5705,g2376,I10482,g1157,I7095,g6501,g8830,g6025,I13028,I8799,I9344,g9332,I9609,g1269,g8455,g9236,I14985,g4235,I8796,g9018,g99,g4007,g6846,g4109,I5852,g5738,g6252,I12011,g8286,I5475,g8783,g2288,g1675,I11874,I15648,I9372,I10907,g6590,g4910,I7204,g516,g8178,g9114,g5172,g4593,g9091,g5109,I13800,g3818,g8925,g184,I11031,g1732,I9069,g5239,g2315,g4500,g6615,g4135,g3398,g6735,g600,g5115,I13728,g4959,g3679,I9050,g2661,g7835,g607,g8967,I9687,I10819,g2936,g8975,g6417,g2937,I10497,I15329,g5799,g9186,g8874,I6941,g1743,g7017,g6352,I12918,I6021,g2161,I12952,g4617,g6502,I14019,g6863,I6795,I13109,g5266,I8966,I12760,g2962,g1,I10933,g1569,g126,I12639,g7251,g168,g2293,g8730,I9823,g294,g4172,g4067,g5428,g5227,g1528,g7679,g4083,g8918,I6996,I5978,g6493,g6721,I6189,g8326,g8620,g9348,I10415,I15773,g5652,I10262,g6394,I10265,I8253,I7311,g2630,g8840,g3158,g6806,I5392,I7335,I11293,g4294,g7605,g3052,g4473,g4686,g7526,I14094,I9009,g4667,g2185,g8259,g6368,I14795,g8220,I9826,g5202,g1786,g7708,g2287,I10940,I5664,g9033,g7590,I13092,g8406,g9206,g4718,g1336,I7383,g4791,I13466,g4504,g4937,I8569,I10969,I10019,I14445,g7167,g4071,g6255,g1917,g2643,g8177,I8718,I6223,I7211,g3909,g540,g6144,g474,g3861,g2396,g9309,g5605,g7723,g5063,g1865,g3547,g6613,g2618,g1825,I8790,g3339,I7461,g4558,I7531,I14073,g9120,g9272,g6187,I6936,g3894,g9380,g4085,I14151,g584,I6195,g2634,g7247,I11870,g4397,g2170,I13369,g6375,g8541,g2686,I16049,g6710,g828,g7248,g8916,g6567,g1351,g9160,g8150,I5696,I5914,g2498,I5520,g7855,g1583,I14825,g3074,g4523,I7098,g236,g4389,g6041,g5459,g3011,I6203,g6598,g6171,g6194,g7121,I15723,g3532,I10965,g6107,I8883,g6302,g7686,g1118,g1229,g4028,I13126,g6184,g5418,g1004,g2295,I13659,I9588,g4199,I15264,g7244,I10925,g6556,g3974,g5820,g7421,I11383,I6539,g6404,g809,g231,g426,g5732,g8739,g6131,g7171,I5718,I7344,g3509,I12164,g2381,I15601,g1018,I8856,g4820,g5832,g7215,I7466,I7911,g3852,g2485,I12768,g3832,I8724,g8825,g2872,g4599,g4334,g5257,g7354,g4070,g8269,g6874,g7993,I8706,g4427,g6876,g5479,I13441,g9171,I13834,g4099,g5466,g2131,g68,I7554,g5798,g3892,g1570,I16043,g2457,g1718,g1941,g7158,I11842,g4737,g4872,g4055,g5483,I15817,I9166,g3583,g6347,g1432,I12101,g1159,I9986,I7479,I14118,g4350,g1854,g6243,g1933,I14683,I9195,g1655,g3916,I5395,I13553,g3523,g7216,I8172,g1481,g2274,I8757,g1389,g8257,g6950,I6337,I5945,g8732,g8074,I10369,I9277,I10177,I7158,I7167,I5535,I11124,g7152,I11744,g492,g8318,g3497,g8839,g2521,I11569,I15921,I14196,g4435,I15738,g7279,g4578,g4565,I15546,g1296,g2532,g233,I8605,g2784,g4047,g6896,g42,g8680,g7146,I12439,g8274,g7575,I12259,g2020,I14454,g4054,g4514,g6007,I8832,g4451,g5538,g3868,I12526,g6304,g6220,g1711,g130,I15042,I5377,g4645,I10525,g1694,g1380,g2640,I8034,g5616,g5671,I8528,g2894,I10783,g9288,I15275,I9953,g8513,g2269,g3237,g5842,g619,g3841,g6173,g5026,g3591,g8264,I13900,g2908,g7262,g8604,I14460,g9009,I6523,g420,g5745,I12945,I9416,g6734,g398,I8871,g4106,g4270,g4271,g5184,I11473,I10815,g8282,g7560,I15014,g4243,I11123,g4198,I11607,I6997,I12322,I13397,g6420,g2328,I13861,I7009,g7534,I7746,g7191,I9333,I10017,I5775,g7328,g8700,g2226,g1838,g2486,I13228,I11559,g9351,g7678,I8560,I14728,g4187,g9337,g6931,I15912,g7057,g4920,g1097,g9168,I5747,I6358,I11095,g883,g1789,g6290,g5042,g2316,g6122,I8838,g8302,I14012,I7523,I8090,g2562,I15660,g9338,g5826,g4878,I11150,I12190,I7584,I7320,g1486,g9227,g2777,I10888,I5380,I12544,I14049,I12989,g8062,g8404,I5425,g6766,g6825,I9181,g9081,g1793,g5801,g8793,I16126,I7731,I8558,g1739,I15242,g8884,I11287,g7827,g4423,g2377,g2958,g760,g6791,I11464,I6419,g7310,g3864,g7027,I8593,I11764,g4630,I9276,g215,I10906,g1678,I14400,g5731,g4607,g7793,g7030,g1664,g8636,g7530,I5981,g5173,g4911,g9197,g5260,g5589,I6868,g2364,I11275,g6725,g2767,g5645,g4527,g6063,I8606,g5987,g3496,g8781,g5956,I13802,g33,I5353,I7240,g4381,I16158,I10976,g4300,g12,g4809,I12135,g6174,g4309,g4068,g7183,I8041,g185,g4556,I13746,I7487,g3655,g6324,g3461,g1867,I9828,g3774,g6919,I14573,I11652,I14224,I10791,I11171,g4788,I12031,I8299,g5119,g5434,I10818,I8094,g5027,I14410,g5722,I11848,I13785,g8901,g174,g8012,g7069,I8538,g4894,g3526,g359,g8737,g3945,g8299,g1514,I13685,I15887,I8916,I8205,g6083,g5305,I15152,I8224,I6171,I6844,I8431,g8699,I8333,g8014,I13137,g7767,g738,g7232,g8865,g3128,g6239,I11987,g6,I10579,g5067,g6610,g9192,I9660,g8009,g7565,g7035,g4522,I10873,I13016,g6307,g2881,g2795,I8952,g6772,I13002,g7189,g2955,g8633,g959,g232,I11094,I15160,g8077,g9277,I15684,g8735,g1770,g1223,g6573,I12313,g8752,g2921,g3932,g4899,g9005,g6865,g3631,g1796,I13238,g5591,I15836,g8707,I13075,g9271,I11212,g7825,g8649,I7112,I14163,g6777,I7460,g7460,g7951,g5019,g1198,g8935,g8145,g7558,I10582,g4477,g7055,I15243,I10010,g6759,I5865,g649,I6143,g475,I12161,g6216,g5442,g7769,I13457,g4365,g8750,g2882,I12853,g1374,I9782,I11086,I14205,I13813,I10418,g7448,I12041,g5196,g6868,g2362,I13395,I12310,g3048,g6093,g7781,g4041,I12881,I14406,g7543,g8278,g9135,g4024,I14181,g8847,I12017,I8456,I11157,g6817,g4618,g6401,I14039,I10854,g1925,g8674,g9006,I13018,g6354,g6166,g9375,g1895,g6633,I7611,I7164,I7326,I12748,I15690,g2551,I12708,g4644,g2770,I6208,I9889,I7068,g4594,g6045,g2210,g8627,g2157,g9358,g110,g2941,g4831,g1320,g8335,g4925,g4474,g603,g3665,I14783,g8481,g354,g452,g365,g4295,g3678,g7212,g1460,g7220,g7081,g4641,g7362,g1821,g2965,g6129,g6820,g795,g6770,g3771,g37,g9147,g7454,I12552,g8743,g1333,g5092,g9065,I6209,g7314,I12108,g5673,I12241,g4512,g863,I12337,g4798,I14614,g7013,g2845,I11185,g7175,I9369,I15292,I10512,g8322,I8084,g4,I7392,I8165,g8039,g9131,I12016,g1876,g2511,I5621,g7241,g6790,g4201,g3051,g6998,g613,I6127,I7314,g3546,g5241,g9012,I7532,g1589,g7150,g9267,I14103,I6750,I14819,g5586,g7141,I12869,g1759,I9058,I11317,I12340,g6504,g9252,I14848,g6878,g9347,g6726,g4602,g6301,I11101,I13527,g5125,I14496,g5311,g6355,I13776,g1412,I14433,I15029,g6008,g6020,I11413,g4625,I15845,I12098,g4180,g3644,I15478,g1267,I8373,I11596,g8860,g1823,g228,g5603,I10314,g5129,I9477,I12141,g6857,g3684,g5984,g9001,I12576,I14115,g4669,g8973,I10061,g6826,g2458,I10060,g5597,g6313,I12586,g1235,g7126,g333,g4410,g6756,g1922,g6642,g8094,I12352,g6757,I12681,g5223,g2898,I7697,I13287,I7174,g4391,I10335,g4062,g7501,g462,g6021,I9512,g6400,g6286,I9767,I14334,g394,I15819,I10545,g4230,g5045,I12885,I6673,g6338,g3229,g8797,I16132,g6773,g1976,I9496,I11254,I10900,I9627,g6914,I6048,I13831,g1138,I15562,g1733,g7492,I14798,g6869,g2692,g8870,g1970,I11260,I9152,I11503,g7414,g7238,g4694,g9103,g7412,I6900,g5056,g6634,I7728,I12235,g5245,g9154,g9180,g6246,I15666,g8831,g5255,g4065,g9165,g6431,g8697,g618,g3611,g6309,g7264,g7486,I12541,I7215,g7439,I14468,I10776,g181,g1400,g5244,g1833,I6317,g5242,I16026,g290,g8954,g2956,g8258,g5563,I15083,g8456,g7078,I12478,g7002,g7544,g7231,g5218,I7356,I14270,g4066,g5473,g5177,g6886,g8961,I15714,g9329,I15663,g7694,I5507,I14479,g1182,I10445,I13220,g7118,g3658,g9303,g1403,g7726,I8778,g7358,I7428,I14473,I12256,g6607,I15607,g4807,g6684,g1671,g8060,g669,g4797,g1728,g822,g5579,I11875,I9053,g5555,I5842,g273,g995,g4727,g6044,g6641,g6924,I7341,g6514,g8712,g8271,I14160,g3863,g3836,g8826,g1444,I7734,g4491,I9929,g6946,g6935,I13725,g5240,g6468,g7562,g6448,I12973,g7131,g2627,I12833,g5754,g6165,g4889,g8676,g8927,I8161,g4377,g5344,g3632,g3874,g2953,I10353,g5582,g8637,I11666,g9115,g4570,g6795,I9330,g4472,g1898,g9374,g7447,g1611,g4528,g8662,I10406,g7086,I6571,I12652,g6705,I7569,g6118,g89,I13666,g7576,I7061,g6245,I15253,g6602,g6702,I11296,g6202,g5937,g3542,g4597,g8308,I8574,I12289,g8088,g2727,g4562,g4160,g6828,g4826,I13679,g6064,I13264,I13710,I14091,I6946,g8810,g8893,I8913,g5520,I15276,g4600,g9078,g887,g4304,I8490,g5118,g4095,g306,I10548,g7348,g9000,g6765,g9007,g8966,g7760,g6481,I7944,g9226,I13326,g6449,g1397,I13410,g8261,I13144,I13515,I12505,g4705,g8813,g7525,g8292,I8971,g4703,g8742,g4238,g6430,I11392,I15382,g3834,g8061,g1587,g955,I13909,g2183,g4282,g6980,I11714,I8121,I6629,I8340,g9090,I12079,I12871,I7430,g3092,g5256,g4582,g1771,I6201,g5871,I12900,I15857,g8237,g8924,I15101,g3985,g4237,g8613,g8642,g20,g3071,g7609,I13656,g8289,g3907,g8298,I12829,g105,g7099,g1749,I14767,g5810,I8291,g6014,I12936,g3901,g7531,I13640,g7036,I10193,I12220,g1785,g4019,g8817,I6739,g1224,I11752,I8046,g6427,I9543,I11978,g7540,I7444,g8724,g2721,I11476,g8727,g5734,I8546,g4720,g4279,g2474,g3230,I11047,g8603,I8512,g4804,g6388,g4367,g1708,I7459,g1688,g5744,I9250,g6882,g4637,g6092,I11482,I11633,g4929,g8962,I9642,g2834,g6422,I13164,g4374,g1459,g5436,g539,g8788,g2695,g4191,g4954,I14668,g9037,g8678,g6671,I12472,g2213,g1250,g7677,I9746,I13042,g5762,g9130,g336,g8963,g5050,I7064,I8079,g8990,I7053,I8901,g225,I8510,g3220,I9654,g9064,g2638,I5435,I15385,g8623,g5168,g2798,g636,g4549,g6296,g6034,g799,g2294,g6854,g7415,g5621,g8904,I8177,I12834,I11967,g2918,g759,g2403,g5577,I15394,g1834,g2912,I9366,I12283,I12961,g1271,I11951,g2350,I10987,I14851,g6213,g8822,g52,g9098,g3767,I8940,g2649,g5714,g9344,I11096,g2402,I9840,I11512,g8885,g1142,I7468,g6711,g7197,I11103,I14837,g2636,g4588,g5139,g5153,g1386,g1513,g5712,I9183,g8070,g1391,g889,I11908,g368,I12558,g4014,g5600,g5873,I11419,g8733,g2628,I10347,I16040,I7937,I12567,I13518,I10866,g6835,g5545,I11873,g7681,g6543,g8695,I7485,g5237,g6821,g6226,g7450,g8842,g9251,I6952,g1268,g1727,g7459,I11434,I16103,g5198,g5051,g933,g5488,g2505,g9184,I5619,I11281,I10930,g763,g5604,I13203,I7775,g5548,I10283,g7479,g6268,g9195,g627,I12382,g4938,I12826,g5540,g501,I8712,I8748,g6022,g2528,g8786,I10752,g4299,I14766,g5185,g1532,g8923,g2871,g2525,g4113,g6694,g8650,g1201,I11011,I11347,g8956,g9119,I8028,g2307,g316,I9258,g7483,g4009,g4680,I10949,g7108,I5552,I10992,g5441,g621,I7970,g3885,I11055,I10186,g4413,I8928,g567,g6189,g5615,I11224,g4090,g9030,I8974,I6728,I7850,I7875,g7616,g7032,I10018,g6689,I9084,g4819,g4349,I10835,g6830,g5183,g4115,g7140,I7893,I5861,I8880,g4004,I12253,g449,I10475,g5797,I11021,I8400,g7555,g6680,g6880,g6700,I15856,g2259,I9457,I12238,g6541,g1662,g1949,I6229,g2382,I9576,I14298,g4073,g6487,g6814,I15272,g6206,g7304,I11090,I15818,I9505,I12596,g6214,I11693,g4457,I14472,g4077,g8716,I8636,g718,g2378,g5733,g6784,g5188,g5417,g4650,I10328,I9980,g6703,I8491,g2332,g8913,g2484,g7577,g7718,g5014,g8729,g4145,g6292,I9974,I9946,g6740,I6234,I15628,I8524,g5080,g1689,g2897,g8313,g8926,g1160,g312,g5670,I11452,I7429,g5158,g4648,g7533,g8708,g8342,g5161,g240,g2961,g8582,g2617,g8829,g7444,g5573,g3896,I11440,g330,I13646,I9107,g3516,g2237,g5665,g6350,g7280,g7093,I7359,I15379,I6842,g2917,g9042,g6591,g4955,I16183,g8878,g9276,g381,g6231,I13854,I13432,g5897,I13891,g9046,g4902,I12806,g3613,g8765,g4893,g1366,g437,I7287,I9884,g6930,g7148,I9528,I11290,I15337,I6099,g6217,I11359,I8495,g1404,g5182,g6123,I12430,g7060,g6157,g1450,I6878,g4076,g9043,g2241,g4150,g6788,g4058,I11533,g6827,g7322,g4529,I15894,I9001,g4154,g8883,I10032,g327,g871,g8717,g8740,I10329,g1929,g6026,g4886,g1014,I7814,g8221,g6378,g614,I15735,g4933,g7828,g6140,g8673,g5556,g7680,g6623,I13559,I8811,g1461,I14451,g4876,g2006,g8824,g7091,I11945,g8843,I5616,g4093,g1666,g4877,g4307,I8862,g3845,g8438,g2230,g6637,g6434,g7133,g6574,g2290,I7959,I5889,g6413,g9027,g7261,g9376,g9122,I9669,g3629,g2236,g7124,g3986,g3160,g550,I6029,I16122,g154,I15196,g5831,I10092,g2284,g5564,I6643,g2641,g7703,I5362,I15871,I8193,I8151,g1769,g6660,g6393,g373,I10608,I14480,g9073,g2333,g1672,g264,g9187,I15610,I11269,g2653,I6214,g985,g295,g3764,g2790,g7300,g6333,I11923,g5833,I9095,I13716,g1901,I11861,g5795,g6738,g8996,I5404,g8384,g7493,g7737,I6348,g9235,I7129,I6906,g6410,I12199,g6162,g3574,I7498,I13428,g5181,g8841,I11576,g3038,g4890,g8688,g6441,g4029,I6970,g5461,g7584,I5948,I8983,I13454,g4691,g7353,g8834,g5489,g3340,g6754,g7734,g9008,g2306,g5632,g6587,I12167,g9301,I15111,g274,I10617,g1263,g7905,I6291,g2467,g5711,g9059,I7511,g5175,g9134,g4643,I9791,g7168,g8320,g8379,g3721,I10561,g1443,I14834,g5020,g4779,I15930,g7327,I15619,I5548,g547,I12487,I12839,g9056,g8672,I7919,g2631,I13475,g1558,g5766,g5782,g6644,g1328,g8900,g1106,g4018,I12609,I8045,g3286,g6883,g8720,g8897,g5788,I5795,g6329,g2216,g3815,g6110,g3097,g9032,g219,g1170,I10207,g7025,g2673,I8886,g691,I13687,g2311,I13344,I5966,g4934,g4169,g7271,I9978,g5537,I6093,I6157,g3518,g8827,g8461,I9804,I13722,g9377,g6132,g7440,g6402,g9108,g6270,g2632,I15208,g3019,I15481,g6723,I7891,I10436,g8310,g5523,g5819,g6961,g9385,g4155,g6374,g5084,g8687,g3905,g26,I7672,g517,I7765,I13311,g7166,g3675,g25,g639,I12331,g1388,g4012,I8186,I10592,g5213,g6436,g911,I8679,I12145,g8564,g6316,g866,I7574,I12547,I8919,g803,g6098,g4786,g4005,I13063,I10528,I12655,g4548,I6286,g7788,I14190,g21,g3602,g4489,I12427,I7173,I6178,g878,g3341,I7187,g8018,g6977,g5170,I12731,I12208,I12717,g6701,g7709,g6503,g4466,g3889,I13550,g570,g2826,g2935,g7438,g6832,I11050,I13247,g1381,g1190,g8763,g8063,I14145,g4803,g7811,g9079,I11314,g2481,g3545,g9384,I13918,I10991,g5780,g4688,I8678,g6663,g7237,I11903,g3129,g1818,g5224,I7892,I6009,I6711,I6183,I12782,I10954,I6500,I7785,g5622,I7070,I8157,I8503,I10183,I8360,g2494,I15915,g4310,I12810,I9393,g3839,g8607,I10875,g6677,g9020,I8680,g29,I6275,g195,g3989,I13084,g1236,g6331,g971,I9850,I13743,g7545,g196,g4537,g3651,g2543,g8869,g3634,g7047,g8226,I11574,g3285,I5697,I15021,I14777,g1557,I14772,g2624,g7364,g5827,I8470,g4251,g4932,g9117,g1574,g5580,g5609,g7172,g4714,I14722,g6364,g1330,g1401,I12921,I11887,g1907,I13779,g8914,I13147,I10373,I14076,I8225,g150,g7000,I8101,g7125,g3681,g6072,I6524,g8696,I12078,g5017,I6517,g5206,I14718,g8821,g4780,g8671,I8114,g6405,I11404,I14302,I12582,I14211,I8240,I10962,g9387,g1207,I11551,g5575,I9648,g6208,g6569,g7258,g1369,g4167,g1943,I13131,g7346,g8068,g3707,g1788,g3648,g3757,I7473,g1849,g6097,g5215,g6124,g4822,I11672,I6876,g6897,g8079,g4390,g3833,I7132,g7352,g2915,g6201,I5633,g1684,I9029,I11060,g8288,g6811,g7065,g2876,I16116,I13377,I13460,g6102,g9190,g117,g8766,g8866,g1053,g9061,I5695,g9074,g483,I13493,g2052,I11218,I15756,g6727,I14970,g1081,I11194,g2999,g921,g1323,g8854,I11221,I8889,I13317,I11689,g5836,I14495,g3888,I9153,g7229,g6023,I5528,g7343,g3430,g9274,g2011,I13009,g6101,g4906,g2928,I15622,g5044,g1721,I15947,g2842,I12343,g6802,g6993,g7600,I15557,g2828,g5120,g22,g5834,g8828,g3189,g2698,I12358,g6894,I12211,g1013,g7020,g8227,g7561,I11750,I7181,I5670,g6808,I5466,I8233,I9129,I9693,g2930,g1938,g8180,g1179,g846,I6151,g5047,g6771,I15959,g6349,g8871,g3971,g199,g6076,I11040,g2266,g5794,I6039,g4510,g8514,g1714,g2817,g8459,g5560,g6922,I15678,I9241,g5612,g44,g6053,I15284,g6335,I12032,g2231,g5075,I14311,g3639,g7746,g5841,g190,I13512,g6626,g2899,g2751,I9047,g7427,g5730,g849,g6190,g2561,I11615,g3694,g5618,I6767,I11132,g734,I9034,g2869,g4301,g9086,I8196,g1206,g8692,I10040,g2683,I10424,I8939,I10914,I13930,I15187,I6045,g6940,g7747,g3647,g4386,I5505,g7077,g1715,g1639,g4544,I7467,I6000,g7043,g6340,g1173,g3359,g6926,g6259,g6047,g3488,g7476,I10587,g4805,g4867,I15982,g376,I11818,g9383,I7994,g8848,g3504,g1959,g4909,g6042,g9136,g1612,g1309,g8959,I12870,g292,I11422,I13274,g1228,g7752,g9141,g4574,g8277,I5801,g8621,g1822,g6654,g2907,g2946,g5584,g9121,g7179,I7605,g3954,g8232,I15598,g2595,I13843,g3856,g1227,g8850,I10135,I13537,g2289,g4698,g6423,g5426,g6328,g6568,I8565,g6964,g4318,I6775,g7046,I11603,g673,g7128,I13782,g4596,I8134,g5628,I15100,g5211,I12148,I10093,I13846,g4790,g4679,g2801,g727,g1251,g7690,I7644,g8945,g8723,I11108,g5018,I8393,I5531,g1848,g7161,g5847,g4555,I12666,g6419,g4284,g6779,g9368,g3082,I7832,g5779,g6222,I6371,I10000,I5972,g5267,g8747,g5829,I9014,I6615,g5719,I9549,g440,I6974,I10684,g3081,g5229,I8955,g1342,g2910,g6603,I14758,I12535,g9069,I9639,I5963,g9051,g966,g7720,g4086,I9341,I12379,g4194,g2668,g7135,g7432,g5186,I11431,g3676,g4384,g3760,I13752,I7503,g3513,I15513,g620,g4776,g5916,g6061,g3923,g5549,I8733,I6501,I8152,I8949,g7365,I13906,g2205,I9336,g7184,g9259,I7350,I12388,g3515,I9548,g16,I11179,g6973,g524,I12702,g5476,g8993,g8999,g4034,I6154,g6685,g4281,g7185,g7312,g1489,g7728,g7341,I10687,g6921,I15927,g284,I11236,I14960,g8224,g4782,g6250,I12699,g9080,g3728,g65,I13173,I13296,g5677,g7096,I14124,g5194,g8794,g2272,g342,I10719,g9382,g7628,I9663,I9965,g7195,g4138,g9106,g6636,I13940,g646,g3975,g8111,g8756,g1747,I10306,g1191,g2407,I12980,I10039,I7374,I11815,I15654,g4778,I7299,I14154,g3881,I10896,I7438,I10829,g6095,g5146,g3231,I7623,I15669,g6965,I14022,g1057,g6959,I13810,g9194,I11329,g7456,g6908,I8019,I6930,g2639,g806,g4269,g9318,I9992,g3828,I13152,g6057,I15550,I13185,g4002,g6219,g6096,g5078,I14172,g5567,g1365,g7778,g942,g6570,g5574,g6149,g8698,g4383,g6650,g2952,g6151,g5614,g2948,g1677,I13225,g3643,I9555,g3514,g4102,g8682,g3510,I13004,I6226,I6368,g2536,g2073,g7701,g8071,I10500,g133,g2964,I9169,g3837,g8746,I12120,I14474,I6363,g6421,I15055,I13199,g243,I6940,g4711,I13255,I7922,g4195,I14747,g3573,g1021,g71,I7495,I6751,g9336,I12561,g2459,g5298,I9564,g3987,I12469,g6592,I11500,g4341,I11129,I6918,g916,g6899,I13481,g1802,g5561,g4462,g7634,g3610,g7130,g7278,I6299,I13682,g396,g6579,I7188,g7194,g6276,g7419,I11263,g9324,I6042,g5805,g5715,g4075,g8064,I9475,g5384,g9264,g7097,I14394,I13598,I7847,g770,g8714,g5038,g3990,g1033,g6476,g8646,g5155,I15687,g6954,g3501,g5261,g5631,g8386,I11356;
//# 31 inputs
//# 121 outputs
//# 669 D-type flipflops
//# 5378 inverters
//# 2573 gates (1114 ANDs + 849 NANDs + 512 ORs + 98 NORs)
//
//
//
  MSFF DFF_0(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g31),.DATA(g6302));
  MSFF DFF_1(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g30),.DATA(g6301));
  MSFF DFF_2(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g29),.DATA(g6300));
  MSFF DFF_3(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g28),.DATA(g6298));
  MSFF DFF_4(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g27),.DATA(g6297));
  MSFF DFF_5(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g26),.DATA(g6296));
  MSFF DFF_6(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g25),.DATA(g6295));
  MSFF DFF_7(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g24),.DATA(g6294));
  MSFF DFF_8(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g23),.DATA(g6293));
  MSFF DFF_9(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g22),.DATA(g6292));
  MSFF DFF_10(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g12),.DATA(g8662));
  MSFF DFF_11(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g11),.DATA(g6290));
  MSFF DFF_12(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g9),.DATA(g6288));
  MSFF DFF_13(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g8),.DATA(g9376));
  MSFF DFF_14(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g7),.DATA(g9375));
  MSFF DFF_15(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6),.DATA(g9374));
  MSFF DFF_16(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5),.DATA(g9373));
  MSFF DFF_17(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4),.DATA(g9372));
  MSFF DFF_18(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2),.DATA(g9361));
  MSFF DFF_19(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3),.DATA(g9360));
  MSFF DFF_20(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g48),.DATA(g9362));
  MSFF DFF_21(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g21),.DATA(g6299));
  MSFF DFF_22(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g10),.DATA(g6291));
  MSFF DFF_23(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1),.DATA(g6289));
  MSFF DFF_24(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g47),.DATA(g9389));
  MSFF DFF_25(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g46),.DATA(g8955));
  MSFF DFF_26(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g45),.DATA(g6308));
  MSFF DFF_27(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g44),.DATA(g6307));
  MSFF DFF_28(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g42),.DATA(g6306));
  MSFF DFF_29(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g41),.DATA(g6305));
  MSFF DFF_30(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g37),.DATA(g6304));
  MSFF DFF_31(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g32),.DATA(g6303));
  MSFF DFF_32(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1207),.DATA(g5173));
  MSFF DFF_33(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1211),.DATA(g5174));
  MSFF DFF_34(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1214),.DATA(g5736));
  MSFF DFF_35(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1217),.DATA(g6377));
  MSFF DFF_36(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1220),.DATA(g6378));
  MSFF DFF_37(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1223),.DATA(g6379));
  MSFF DFF_38(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1224),.DATA(g6857));
  MSFF DFF_39(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1225),.DATA(g6858));
  MSFF DFF_40(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1226),.DATA(g6859));
  MSFF DFF_41(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1227),.DATA(g7108));
  MSFF DFF_42(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1228),.DATA(g7109));
  MSFF DFF_43(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1229),.DATA(g7110));
  MSFF DFF_44(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1230),.DATA(g7300));
  MSFF DFF_45(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1240),.DATA(g1235));
  MSFF DFF_46(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1236),.DATA(g1240));
  MSFF DFF_47(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1231),.DATA(g1236));
  MSFF DFF_48(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1244),.DATA(g2659));
  MSFF DFF_49(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1245),.DATA(g1244));
  MSFF DFF_50(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1243),.DATA(g2660));
  MSFF DFF_51(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1272),.DATA(g6383));
  MSFF DFF_52(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1276),.DATA(g6384));
  MSFF DFF_53(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1280),.DATA(g7112));
  MSFF DFF_54(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1284),.DATA(g7301));
  MSFF DFF_55(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1288),.DATA(g7527));
  MSFF DFF_56(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1292),.DATA(g7302));
  MSFF DFF_57(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1300),.DATA(g7303));
  MSFF DFF_58(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1296),.DATA(g7304));
  MSFF DFF_59(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1253),.DATA(g5741));
  MSFF DFF_60(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1308),.DATA(g6385));
  MSFF DFF_61(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1309),.DATA(g1308));
  MSFF DFF_62(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1310),.DATA(g1309));
  MSFF DFF_63(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1311),.DATA(g1310));
  MSFF DFF_64(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1312),.DATA(g1311));
  MSFF DFF_65(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1304),.DATA(g1312));
  MSFF DFF_66(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1307),.DATA(g3858));
  MSFF DFF_67(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1330),.DATA(g6862));
  MSFF DFF_68(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1333),.DATA(g6863));
  MSFF DFF_69(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1336),.DATA(g6864));
  MSFF DFF_70(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1339),.DATA(g6865));
  MSFF DFF_71(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1342),.DATA(g7119));
  MSFF DFF_72(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1345),.DATA(g7528));
  MSFF DFF_73(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1348),.DATA(g7529));
  MSFF DFF_74(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1351),.DATA(g7530));
  MSFF DFF_75(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1354),.DATA(g7768));
  MSFF DFF_76(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1357),.DATA(g8675));
  MSFF DFF_77(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1360),.DATA(g8676));
  MSFF DFF_78(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1190),.DATA(g8677));
  MSFF DFF_79(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1191),.DATA(g6373));
  MSFF DFF_80(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1192),.DATA(g1191));
  MSFF DFF_81(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1193),.DATA(g1192));
  MSFF DFF_82(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1194),.DATA(g1193));
  MSFF DFF_83(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1195),.DATA(g6374));
  MSFF DFF_84(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1196),.DATA(g1195));
  MSFF DFF_85(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1197),.DATA(g1196));
  MSFF DFF_86(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1198),.DATA(g1197));
  MSFF DFF_87(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1199),.DATA(g6375));
  MSFF DFF_88(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1200),.DATA(g1199));
  MSFF DFF_89(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1201),.DATA(g1200));
  MSFF DFF_90(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1202),.DATA(g1201));
  MSFF DFF_91(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1203),.DATA(g6376));
  MSFF DFF_92(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1204),.DATA(g1203));
  MSFF DFF_93(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1205),.DATA(g1204));
  MSFF DFF_94(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1206),.DATA(g1205));
  MSFF DFF_95(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1252),.DATA(g2661));
  MSFF DFF_96(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1250),.DATA(g7111));
  MSFF DFF_97(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1251),.DATA(g6860));
  MSFF DFF_98(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1247),.DATA(g6380));
  MSFF DFF_99(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1254),.DATA(g6381));
  MSFF DFF_100(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1266),.DATA(g5739));
  MSFF DFF_101(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1260),.DATA(g6382));
  MSFF DFF_102(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1257),.DATA(g5738));
  MSFF DFF_103(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1263),.DATA(g5737));
  MSFF DFF_104(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1267),.DATA(g4656));
  MSFF DFF_105(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1268),.DATA(g5175));
  MSFF DFF_106(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1269),.DATA(g5740));
  MSFF DFF_107(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1271),.DATA(g5176));
  MSFF DFF_108(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1270),.DATA(g1271));
  MSFF DFF_109(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g172),.DATA(g1270));
  MSFF DFF_110(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1313),.DATA(g5742));
  MSFF DFF_111(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1317),.DATA(g5743));
  MSFF DFF_112(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1318),.DATA(g6861));
  MSFF DFF_113(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1319),.DATA(g7113));
  MSFF DFF_114(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1320),.DATA(g7114));
  MSFF DFF_115(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1321),.DATA(g7115));
  MSFF DFF_116(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1322),.DATA(g7116));
  MSFF DFF_117(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1323),.DATA(g7117));
  MSFF DFF_118(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1324),.DATA(g7118));
  MSFF DFF_119(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1325),.DATA(g7305));
  MSFF DFF_120(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1326),.DATA(g7306));
  MSFF DFF_121(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1327),.DATA(g7307));
  MSFF DFF_122(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1328),.DATA(g7309));
  MSFF DFF_123(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g13),.DATA(g7308));
  MSFF DFF_124(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1329),.DATA(g2663));
  MSFF DFF_125(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g20),.DATA(g6386));
  MSFF DFF_126(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1366),.DATA(g6866));
  MSFF DFF_127(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1364),.DATA(g6878));
  MSFF DFF_128(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1370),.DATA(g6876));
  MSFF DFF_129(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1368),.DATA(g6874));
  MSFF DFF_130(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1374),.DATA(g6872));
  MSFF DFF_131(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1372),.DATA(g6870));
  MSFF DFF_132(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1375),.DATA(g6869));
  MSFF DFF_133(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1365),.DATA(g6867));
  MSFF DFF_134(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1363),.DATA(g6877));
  MSFF DFF_135(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1369),.DATA(g6875));
  MSFF DFF_136(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1367),.DATA(g6873));
  MSFF DFF_137(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1373),.DATA(g6871));
  MSFF DFF_138(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1371),.DATA(g6868));
  MSFF DFF_139(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1389),.DATA(g4658));
  MSFF DFF_140(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1379),.DATA(g6879));
  MSFF DFF_141(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1377),.DATA(g6891));
  MSFF DFF_142(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1383),.DATA(g6889));
  MSFF DFF_143(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1381),.DATA(g6887));
  MSFF DFF_144(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1387),.DATA(g6885));
  MSFF DFF_145(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1385),.DATA(g6883));
  MSFF DFF_146(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1388),.DATA(g6882));
  MSFF DFF_147(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1378),.DATA(g6880));
  MSFF DFF_148(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1376),.DATA(g6890));
  MSFF DFF_149(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1382),.DATA(g6888));
  MSFF DFF_150(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1380),.DATA(g6886));
  MSFF DFF_151(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1386),.DATA(g6884));
  MSFF DFF_152(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1384),.DATA(g6881));
  MSFF DFF_153(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1390),.DATA(g4659));
  MSFF DFF_154(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1391),.DATA(g1390));
  MSFF DFF_155(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1392),.DATA(g6387));
  MSFF DFF_156(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1393),.DATA(g2664));
  MSFF DFF_157(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1395),.DATA(g1393));
  MSFF DFF_158(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1394),.DATA(g6388));
  MSFF DFF_159(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1396),.DATA(g4662));
  MSFF DFF_160(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1398),.DATA(g1396));
  MSFF DFF_161(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1397),.DATA(g6389));
  MSFF DFF_162(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1399),.DATA(g3861));
  MSFF DFF_163(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1401),.DATA(g1399));
  MSFF DFF_164(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1400),.DATA(g6390));
  MSFF DFF_165(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1402),.DATA(g6391));
  MSFF DFF_166(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1403),.DATA(g1402));
  MSFF DFF_167(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1404),.DATA(g1403));
  MSFF DFF_168(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g16),.DATA(g1404));
  MSFF DFF_169(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1189),.DATA(g6392));
  MSFF DFF_170(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1412),.DATA(g5745));
  MSFF DFF_171(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1415),.DATA(g5180));
  MSFF DFF_172(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1409),.DATA(g5178));
  MSFF DFF_173(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1416),.DATA(g4665));
  MSFF DFF_174(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1421),.DATA(g5179));
  MSFF DFF_175(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1405),.DATA(g5744));
  MSFF DFF_176(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1408),.DATA(g5177));
  MSFF DFF_177(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1429),.DATA(g2671));
  MSFF DFF_178(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1428),.DATA(g2672));
  MSFF DFF_179(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1431),.DATA(g2673));
  MSFF DFF_180(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1430),.DATA(g4666));
  MSFF DFF_181(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1424),.DATA(g3862));
  MSFF DFF_182(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1524),.DATA(g6393));
  MSFF DFF_183(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1513),.DATA(g1524));
  MSFF DFF_184(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1486),.DATA(g8226));
  MSFF DFF_185(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1481),.DATA(g7769));
  MSFF DFF_186(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1489),.DATA(g7770));
  MSFF DFF_187(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1494),.DATA(g7771));
  MSFF DFF_188(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1499),.DATA(g7772));
  MSFF DFF_189(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1504),.DATA(g7773));
  MSFF DFF_190(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1509),.DATA(g7774));
  MSFF DFF_191(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1514),.DATA(g7775));
  MSFF DFF_192(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1519),.DATA(g8227));
  MSFF DFF_193(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1462),.DATA(g8678));
  MSFF DFF_194(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1467),.DATA(g8875));
  MSFF DFF_195(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1472),.DATA(g8960));
  MSFF DFF_196(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1477),.DATA(g9036));
  MSFF DFF_197(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g727),.DATA(g8228));
  MSFF DFF_198(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1532),.DATA(g7781));
  MSFF DFF_199(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1528),.DATA(g7776));
  MSFF DFF_200(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1537),.DATA(g7777));
  MSFF DFF_201(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1541),.DATA(g7778));
  MSFF DFF_202(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1545),.DATA(g7779));
  MSFF DFF_203(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1549),.DATA(g7780));
  MSFF DFF_204(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1435),.DATA(g5181));
  MSFF DFF_205(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1439),.DATA(g5182));
  MSFF DFF_206(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1432),.DATA(g5183));
  MSFF DFF_207(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1443),.DATA(g4667));
  MSFF DFF_208(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g33),.DATA(g5184));
  MSFF DFF_209(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g38),.DATA(g5746));
  MSFF DFF_210(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1461),.DATA(g4669));
  MSFF DFF_211(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1444),.DATA(g5185));
  MSFF DFF_212(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1450),.DATA(g5186));
  MSFF DFF_213(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1454),.DATA(g5187));
  MSFF DFF_214(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1459),.DATA(g3863));
  MSFF DFF_215(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1460),.DATA(g4668));
  MSFF DFF_216(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g979),.DATA(g7104));
  MSFF DFF_217(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g966),.DATA(g8223));
  MSFF DFF_218(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g969),.DATA(g966));
  MSFF DFF_219(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g963),.DATA(g7764));
  MSFF DFF_220(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g970),.DATA(g963));
  MSFF DFF_221(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g971),.DATA(g5171));
  MSFF DFF_222(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g972),.DATA(g2653));
  MSFF DFF_223(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g973),.DATA(g8672));
  MSFF DFF_224(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g976),.DATA(g8864));
  MSFF DFF_225(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g984),.DATA(g9133));
  MSFF DFF_226(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g985),.DATA(g7515));
  MSFF DFF_227(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g990),.DATA(g7516));
  MSFF DFF_228(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g995),.DATA(g7517));
  MSFF DFF_229(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1004),.DATA(g7105));
  MSFF DFF_230(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1005),.DATA(g1004));
  MSFF DFF_231(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g998),.DATA(g1005));
  MSFF DFF_232(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g999),.DATA(g8865));
  MSFF DFF_233(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1007),.DATA(g8867));
  MSFF DFF_234(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1012),.DATA(g6851));
  MSFF DFF_235(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1014),.DATA(g1012));
  MSFF DFF_236(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1013),.DATA(g1014));
  MSFF DFF_237(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1029),.DATA(g2654));
  MSFF DFF_238(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1018),.DATA(g8869));
  MSFF DFF_239(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1021),.DATA(g8870));
  MSFF DFF_240(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1025),.DATA(g8871));
  MSFF DFF_241(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1033),.DATA(g9034));
  MSFF DFF_242(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1034),.DATA(g8957));
  MSFF DFF_243(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1030),.DATA(g7518));
  MSFF DFF_244(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1081),.DATA(g6852));
  MSFF DFF_245(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1156),.DATA(g1081));
  MSFF DFF_246(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1157),.DATA(g1156));
  MSFF DFF_247(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1159),.DATA(g1157));
  MSFF DFF_248(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1158),.DATA(g1159));
  MSFF DFF_249(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1084),.DATA(g7106));
  MSFF DFF_250(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1146),.DATA(g1612));
  MSFF DFF_251(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1147),.DATA(g1146));
  MSFF DFF_252(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1148),.DATA(g1147));
  MSFF DFF_253(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1087),.DATA(g6853));
  MSFF DFF_254(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1098),.DATA(g6854));
  MSFF DFF_255(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1102),.DATA(g6855));
  MSFF DFF_256(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1106),.DATA(g7107));
  MSFF DFF_257(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1110),.DATA(g7299));
  MSFF DFF_258(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1114),.DATA(g7521));
  MSFF DFF_259(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1118),.DATA(g7766));
  MSFF DFF_260(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1122),.DATA(g8225));
  MSFF DFF_261(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1126),.DATA(g8674));
  MSFF DFF_262(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1142),.DATA(g8874));
  MSFF DFF_263(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1173),.DATA(g7526));
  MSFF DFF_264(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1170),.DATA(g1173));
  MSFF DFF_265(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1167),.DATA(g1170));
  MSFF DFF_266(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1166),.DATA(g1167));
  MSFF DFF_267(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1077),.DATA(g7767));
  MSFF DFF_268(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1153),.DATA(g6856));
  MSFF DFF_269(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1154),.DATA(g1153));
  MSFF DFF_270(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1155),.DATA(g1154));
  MSFF DFF_271(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1185),.DATA(g1155));
  MSFF DFF_272(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1097),.DATA(g1185));
  MSFF DFF_273(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1092),.DATA(g7520));
  MSFF DFF_274(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1130),.DATA(g7522));
  MSFF DFF_275(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1134),.DATA(g7523));
  MSFF DFF_276(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1138),.DATA(g7524));
  MSFF DFF_277(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1149),.DATA(g7525));
  MSFF DFF_278(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1037),.DATA(g7519));
  MSFF DFF_279(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1041),.DATA(g7765));
  MSFF DFF_280(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1045),.DATA(g8224));
  MSFF DFF_281(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1049),.DATA(g8673));
  MSFF DFF_282(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1053),.DATA(g8873));
  MSFF DFF_283(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1057),.DATA(g8959));
  MSFF DFF_284(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1061),.DATA(g9035));
  MSFF DFF_285(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1065),.DATA(g9117));
  MSFF DFF_286(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1069),.DATA(g9134));
  MSFF DFF_287(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1073),.DATA(g9145));
  MSFF DFF_288(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1163),.DATA(g2655));
  MSFF DFF_289(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1160),.DATA(g1163));
  MSFF DFF_290(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1182),.DATA(g1160));
  MSFF DFF_291(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1186),.DATA(g1182));
  MSFF DFF_292(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1179),.DATA(g1186));
  MSFF DFF_293(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1176),.DATA(g5172));
  MSFF DFF_294(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g68),.DATA(g6774));
  MSFF DFF_295(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g71),.DATA(g6775));
  MSFF DFF_296(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g74),.DATA(g6776));
  MSFF DFF_297(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g77),.DATA(g6777));
  MSFF DFF_298(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g80),.DATA(g6778));
  MSFF DFF_299(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g83),.DATA(g6779));
  MSFF DFF_300(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g86),.DATA(g6780));
  MSFF DFF_301(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g52),.DATA(g6781));
  MSFF DFF_302(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g55),.DATA(g7733));
  MSFF DFF_303(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g62),.DATA(g7509));
  MSFF DFF_304(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g58),.DATA(g7734));
  MSFF DFF_305(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g65),.DATA(g4598));
  MSFF DFF_306(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g199),.DATA(g3832));
  MSFF DFF_307(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g200),.DATA(g199));
  MSFF DFF_308(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g201),.DATA(g200));
  MSFF DFF_309(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g190),.DATA(g201));
  MSFF DFF_310(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g195),.DATA(g3831));
  MSFF DFF_311(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g196),.DATA(g5731));
  MSFF DFF_312(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g179),.DATA(g5159));
  MSFF DFF_313(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g186),.DATA(g3830));
  MSFF DFF_314(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g187),.DATA(g5730));
  MSFF DFF_315(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g180),.DATA(g5158));
  MSFF DFF_316(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g205),.DATA(g3835));
  MSFF DFF_317(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g202),.DATA(g5732));
  MSFF DFF_318(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g181),.DATA(g5160));
  MSFF DFF_319(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g210),.DATA(g3834));
  MSFF DFF_320(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g207),.DATA(g5733));
  MSFF DFF_321(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g182),.DATA(g5161));
  MSFF DFF_322(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g146),.DATA(g7735));
  MSFF DFF_323(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g173),.DATA(g7736));
  MSFF DFF_324(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g150),.DATA(g7738));
  MSFF DFF_325(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g174),.DATA(g7737));
  MSFF DFF_326(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g154),.DATA(g7739));
  MSFF DFF_327(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g158),.DATA(g7740));
  MSFF DFF_328(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g162),.DATA(g7741));
  MSFF DFF_329(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g168),.DATA(g7742));
  MSFF DFF_330(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g183),.DATA(g6309));
  MSFF DFF_331(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g184),.DATA(g6310));
  MSFF DFF_332(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g185),.DATA(g4599));
  MSFF DFF_333(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g92),.DATA(g6794));
  MSFF DFF_334(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g89),.DATA(g92));
  MSFF DFF_335(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g93),.DATA(g5145));
  MSFF DFF_336(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g94),.DATA(g6782));
  MSFF DFF_337(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g95),.DATA(g94));
  MSFF DFF_338(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g98),.DATA(g5146));
  MSFF DFF_339(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g99),.DATA(g6783));
  MSFF DFF_340(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g100),.DATA(g99));
  MSFF DFF_341(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g103),.DATA(g5157));
  MSFF DFF_342(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g104),.DATA(g6784));
  MSFF DFF_343(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g105),.DATA(g104));
  MSFF DFF_344(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g108),.DATA(g5147));
  MSFF DFF_345(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g109),.DATA(g6785));
  MSFF DFF_346(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g110),.DATA(g109));
  MSFF DFF_347(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g113),.DATA(g5148));
  MSFF DFF_348(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g114),.DATA(g6786));
  MSFF DFF_349(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g117),.DATA(g5153));
  MSFF DFF_350(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g118),.DATA(g6787));
  MSFF DFF_351(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g121),.DATA(g5154));
  MSFF DFF_352(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g122),.DATA(g6788));
  MSFF DFF_353(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g125),.DATA(g5155));
  MSFF DFF_354(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g126),.DATA(g6789));
  MSFF DFF_355(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g129),.DATA(g5156));
  MSFF DFF_356(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g130),.DATA(g6790));
  MSFF DFF_357(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g133),.DATA(g5149));
  MSFF DFF_358(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g134),.DATA(g6791));
  MSFF DFF_359(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g137),.DATA(g5150));
  MSFF DFF_360(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g138),.DATA(g6792));
  MSFF DFF_361(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g141),.DATA(g5151));
  MSFF DFF_362(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g142),.DATA(g6793));
  MSFF DFF_363(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g145),.DATA(g5152));
  MSFF DFF_364(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g287),.DATA(g3836));
  MSFF DFF_365(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g290),.DATA(g287));
  MSFF DFF_366(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g255),.DATA(g9087));
  MSFF DFF_367(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g258),.DATA(g9088));
  MSFF DFF_368(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g261),.DATA(g9089));
  MSFF DFF_369(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g264),.DATA(g9090));
  MSFF DFF_370(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g267),.DATA(g9091));
  MSFF DFF_371(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g270),.DATA(g9092));
  MSFF DFF_372(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g281),.DATA(g9085));
  MSFF DFF_373(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g284),.DATA(g9086));
  MSFF DFF_374(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g211),.DATA(g4600));
  MSFF DFF_375(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g216),.DATA(g6311));
  MSFF DFF_376(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g212),.DATA(g4601));
  MSFF DFF_377(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g219),.DATA(g6312));
  MSFF DFF_378(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g213),.DATA(g4602));
  MSFF DFF_379(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g222),.DATA(g6313));
  MSFF DFF_380(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g214),.DATA(g4603));
  MSFF DFF_381(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g225),.DATA(g6314));
  MSFF DFF_382(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g215),.DATA(g4604));
  MSFF DFF_383(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g228),.DATA(g6315));
  MSFF DFF_384(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g231),.DATA(g4605));
  MSFF DFF_385(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g237),.DATA(g6316));
  MSFF DFF_386(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g232),.DATA(g4606));
  MSFF DFF_387(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g240),.DATA(g6317));
  MSFF DFF_388(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g233),.DATA(g4607));
  MSFF DFF_389(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g243),.DATA(g6318));
  MSFF DFF_390(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g234),.DATA(g4608));
  MSFF DFF_391(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g246),.DATA(g6319));
  MSFF DFF_392(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g235),.DATA(g4609));
  MSFF DFF_393(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g249),.DATA(g6320));
  MSFF DFF_394(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g236),.DATA(g4610));
  MSFF DFF_395(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g252),.DATA(g6321));
  MSFF DFF_396(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g273),.DATA(g4611));
  MSFF DFF_397(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g275),.DATA(g6322));
  MSFF DFF_398(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g274),.DATA(g4612));
  MSFF DFF_399(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g278),.DATA(g6323));
  MSFF DFF_400(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g368),.DATA(g3838));
  MSFF DFF_401(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g371),.DATA(g368));
  MSFF DFF_402(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g336),.DATA(g9095));
  MSFF DFF_403(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g339),.DATA(g9096));
  MSFF DFF_404(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g342),.DATA(g9097));
  MSFF DFF_405(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g345),.DATA(g9098));
  MSFF DFF_406(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g348),.DATA(g9099));
  MSFF DFF_407(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g351),.DATA(g9100));
  MSFF DFF_408(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g362),.DATA(g9093));
  MSFF DFF_409(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g365),.DATA(g9094));
  MSFF DFF_410(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g292),.DATA(g4613));
  MSFF DFF_411(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g297),.DATA(g6324));
  MSFF DFF_412(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g293),.DATA(g4614));
  MSFF DFF_413(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g300),.DATA(g6325));
  MSFF DFF_414(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g294),.DATA(g4615));
  MSFF DFF_415(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g303),.DATA(g6326));
  MSFF DFF_416(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g295),.DATA(g4616));
  MSFF DFF_417(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g306),.DATA(g6327));
  MSFF DFF_418(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g296),.DATA(g4617));
  MSFF DFF_419(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g309),.DATA(g6328));
  MSFF DFF_420(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g312),.DATA(g4618));
  MSFF DFF_421(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g318),.DATA(g6329));
  MSFF DFF_422(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g313),.DATA(g4619));
  MSFF DFF_423(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g321),.DATA(g6330));
  MSFF DFF_424(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g314),.DATA(g4620));
  MSFF DFF_425(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g324),.DATA(g6331));
  MSFF DFF_426(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g315),.DATA(g4621));
  MSFF DFF_427(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g327),.DATA(g6332));
  MSFF DFF_428(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g316),.DATA(g4622));
  MSFF DFF_429(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g330),.DATA(g6333));
  MSFF DFF_430(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g317),.DATA(g4623));
  MSFF DFF_431(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g333),.DATA(g6334));
  MSFF DFF_432(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g354),.DATA(g4624));
  MSFF DFF_433(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g356),.DATA(g6335));
  MSFF DFF_434(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g355),.DATA(g4625));
  MSFF DFF_435(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g359),.DATA(g6336));
  MSFF DFF_436(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g449),.DATA(g3840));
  MSFF DFF_437(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g452),.DATA(g449));
  MSFF DFF_438(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g417),.DATA(g9103));
  MSFF DFF_439(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g420),.DATA(g9104));
  MSFF DFF_440(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g423),.DATA(g9105));
  MSFF DFF_441(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g426),.DATA(g9106));
  MSFF DFF_442(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g429),.DATA(g9107));
  MSFF DFF_443(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g432),.DATA(g9108));
  MSFF DFF_444(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g443),.DATA(g9101));
  MSFF DFF_445(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g446),.DATA(g9102));
  MSFF DFF_446(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g373),.DATA(g4626));
  MSFF DFF_447(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g378),.DATA(g6337));
  MSFF DFF_448(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g374),.DATA(g4627));
  MSFF DFF_449(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g381),.DATA(g6338));
  MSFF DFF_450(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g375),.DATA(g4628));
  MSFF DFF_451(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g384),.DATA(g6339));
  MSFF DFF_452(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g376),.DATA(g4629));
  MSFF DFF_453(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g387),.DATA(g6340));
  MSFF DFF_454(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g377),.DATA(g4630));
  MSFF DFF_455(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g390),.DATA(g6341));
  MSFF DFF_456(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g393),.DATA(g4631));
  MSFF DFF_457(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g399),.DATA(g6342));
  MSFF DFF_458(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g394),.DATA(g4632));
  MSFF DFF_459(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g402),.DATA(g6343));
  MSFF DFF_460(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g395),.DATA(g4633));
  MSFF DFF_461(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g405),.DATA(g6344));
  MSFF DFF_462(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g396),.DATA(g4634));
  MSFF DFF_463(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g408),.DATA(g6345));
  MSFF DFF_464(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g397),.DATA(g4635));
  MSFF DFF_465(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g411),.DATA(g6346));
  MSFF DFF_466(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g398),.DATA(g4636));
  MSFF DFF_467(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g414),.DATA(g6347));
  MSFF DFF_468(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g435),.DATA(g4637));
  MSFF DFF_469(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g437),.DATA(g6348));
  MSFF DFF_470(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g436),.DATA(g4638));
  MSFF DFF_471(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g440),.DATA(g6349));
  MSFF DFF_472(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g530),.DATA(g3842));
  MSFF DFF_473(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g533),.DATA(g530));
  MSFF DFF_474(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g498),.DATA(g9111));
  MSFF DFF_475(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g501),.DATA(g9112));
  MSFF DFF_476(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g504),.DATA(g9113));
  MSFF DFF_477(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g507),.DATA(g9114));
  MSFF DFF_478(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g510),.DATA(g9115));
  MSFF DFF_479(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g513),.DATA(g9116));
  MSFF DFF_480(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g524),.DATA(g9109));
  MSFF DFF_481(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g527),.DATA(g9110));
  MSFF DFF_482(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g454),.DATA(g4639));
  MSFF DFF_483(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g459),.DATA(g6350));
  MSFF DFF_484(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g455),.DATA(g4640));
  MSFF DFF_485(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g462),.DATA(g6351));
  MSFF DFF_486(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g456),.DATA(g4641));
  MSFF DFF_487(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g465),.DATA(g6352));
  MSFF DFF_488(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g457),.DATA(g4642));
  MSFF DFF_489(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g468),.DATA(g6353));
  MSFF DFF_490(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g458),.DATA(g4643));
  MSFF DFF_491(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g471),.DATA(g6354));
  MSFF DFF_492(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g474),.DATA(g4644));
  MSFF DFF_493(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g480),.DATA(g6355));
  MSFF DFF_494(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g475),.DATA(g4645));
  MSFF DFF_495(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g483),.DATA(g6356));
  MSFF DFF_496(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g476),.DATA(g4646));
  MSFF DFF_497(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g486),.DATA(g6357));
  MSFF DFF_498(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g477),.DATA(g4647));
  MSFF DFF_499(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g489),.DATA(g6358));
  MSFF DFF_500(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g478),.DATA(g4648));
  MSFF DFF_501(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g492),.DATA(g6359));
  MSFF DFF_502(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g479),.DATA(g4649));
  MSFF DFF_503(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g495),.DATA(g6360));
  MSFF DFF_504(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g516),.DATA(g4650));
  MSFF DFF_505(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g518),.DATA(g6361));
  MSFF DFF_506(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g517),.DATA(g4651));
  MSFF DFF_507(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g521),.DATA(g6362));
  MSFF DFF_508(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g535),.DATA(g3844));
  MSFF DFF_509(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g536),.DATA(g6363));
  MSFF DFF_510(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g539),.DATA(g3845));
  MSFF DFF_511(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g540),.DATA(g6364));
  MSFF DFF_512(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g543),.DATA(g3846));
  MSFF DFF_513(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g544),.DATA(g6365));
  MSFF DFF_514(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g547),.DATA(g9026));
  MSFF DFF_515(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g550),.DATA(g9027));
  MSFF DFF_516(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g553),.DATA(g9028));
  MSFF DFF_517(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g556),.DATA(g3847));
  MSFF DFF_518(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g557),.DATA(g6366));
  MSFF DFF_519(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g566),.DATA(g3848));
  MSFF DFF_520(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g567),.DATA(g6367));
  MSFF DFF_521(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g579),.DATA(g3850));
  MSFF DFF_522(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g580),.DATA(g6368));
  MSFF DFF_523(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g583),.DATA(g3851));
  MSFF DFF_524(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g584),.DATA(g6369));
  MSFF DFF_525(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g587),.DATA(g3852));
  MSFF DFF_526(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g560),.DATA(g6370));
  MSFF DFF_527(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g563),.DATA(g9029));
  MSFF DFF_528(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g570),.DATA(g9030));
  MSFF DFF_529(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g588),.DATA(g9031));
  MSFF DFF_530(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g591),.DATA(g9032));
  MSFF DFF_531(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g573),.DATA(g9033));
  MSFF DFF_532(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g576),.DATA(g3849));
  MSFF DFF_533(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g595),.DATA(g576));
  MSFF DFF_534(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g596),.DATA(g6795));
  MSFF DFF_535(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g597),.DATA(g6796));
  MSFF DFF_536(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g598),.DATA(g6797));
  MSFF DFF_537(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g599),.DATA(g6798));
  MSFF DFF_538(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g600),.DATA(g6807));
  MSFF DFF_539(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g601),.DATA(g6799));
  MSFF DFF_540(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g602),.DATA(g6800));
  MSFF DFF_541(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g603),.DATA(g6801));
  MSFF DFF_542(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g604),.DATA(g6802));
  MSFF DFF_543(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g605),.DATA(g6803));
  MSFF DFF_544(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g606),.DATA(g6804));
  MSFF DFF_545(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g607),.DATA(g6805));
  MSFF DFF_546(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g608),.DATA(g6806));
  MSFF DFF_547(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g609),.DATA(g6808));
  MSFF DFF_548(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g610),.DATA(g6809));
  MSFF DFF_549(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g611),.DATA(g6810));
  MSFF DFF_550(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g612),.DATA(g6811));
  MSFF DFF_551(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g613),.DATA(g6820));
  MSFF DFF_552(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g614),.DATA(g6812));
  MSFF DFF_553(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g615),.DATA(g6813));
  MSFF DFF_554(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g616),.DATA(g6814));
  MSFF DFF_555(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g617),.DATA(g6815));
  MSFF DFF_556(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g618),.DATA(g6816));
  MSFF DFF_557(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g619),.DATA(g6817));
  MSFF DFF_558(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g620),.DATA(g6818));
  MSFF DFF_559(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g621),.DATA(g6819));
  MSFF DFF_560(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g622),.DATA(g6821));
  MSFF DFF_561(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g623),.DATA(g6822));
  MSFF DFF_562(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g624),.DATA(g6831));
  MSFF DFF_563(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g625),.DATA(g6823));
  MSFF DFF_564(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g626),.DATA(g6824));
  MSFF DFF_565(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g627),.DATA(g6825));
  MSFF DFF_566(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g628),.DATA(g6826));
  MSFF DFF_567(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g629),.DATA(g6827));
  MSFF DFF_568(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g630),.DATA(g6828));
  MSFF DFF_569(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g631),.DATA(g6829));
  MSFF DFF_570(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g632),.DATA(g6830));
  MSFF DFF_571(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g646),.DATA(g4652));
  MSFF DFF_572(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g652),.DATA(g646));
  MSFF DFF_573(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g661),.DATA(g7743));
  MSFF DFF_574(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g665),.DATA(g7744));
  MSFF DFF_575(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g669),.DATA(g7745));
  MSFF DFF_576(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g673),.DATA(g7746));
  MSFF DFF_577(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g677),.DATA(g7747));
  MSFF DFF_578(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g681),.DATA(g7748));
  MSFF DFF_579(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g685),.DATA(g7749));
  MSFF DFF_580(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g706),.DATA(g7750));
  MSFF DFF_581(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g710),.DATA(g7751));
  MSFF DFF_582(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g714),.DATA(g7752));
  MSFF DFF_583(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g718),.DATA(g7753));
  MSFF DFF_584(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g734),.DATA(g7755));
  MSFF DFF_585(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g730),.DATA(g7754));
  MSFF DFF_586(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g689),.DATA(g6371));
  MSFF DFF_587(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g758),.DATA(g6840));
  MSFF DFF_588(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g759),.DATA(g6832));
  MSFF DFF_589(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g760),.DATA(g6833));
  MSFF DFF_590(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g761),.DATA(g6834));
  MSFF DFF_591(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g762),.DATA(g6835));
  MSFF DFF_592(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g763),.DATA(g6836));
  MSFF DFF_593(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g764),.DATA(g6837));
  MSFF DFF_594(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g765),.DATA(g6838));
  MSFF DFF_595(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g766),.DATA(g6839));
  MSFF DFF_596(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g767),.DATA(g6841));
  MSFF DFF_597(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g768),.DATA(g6842));
  MSFF DFF_598(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g769),.DATA(g6843));
  MSFF DFF_599(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g770),.DATA(g6844));
  MSFF DFF_600(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g771),.DATA(g6845));
  MSFF DFF_601(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g772),.DATA(g6846));
  MSFF DFF_602(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g773),.DATA(g6847));
  MSFF DFF_603(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g774),.DATA(g6848));
  MSFF DFF_604(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g795),.DATA(g3854));
  MSFF DFF_605(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g792),.DATA(g5162));
  MSFF DFF_606(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g782),.DATA(g5734));
  MSFF DFF_607(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g799),.DATA(g7756));
  MSFF DFF_608(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g803),.DATA(g7757));
  MSFF DFF_609(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g806),.DATA(g7510));
  MSFF DFF_610(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g809),.DATA(g7511));
  MSFF DFF_611(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g812),.DATA(g7758));
  MSFF DFF_612(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g775),.DATA(g7759));
  MSFF DFF_613(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g778),.DATA(g7296));
  MSFF DFF_614(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g815),.DATA(g7760));
  MSFF DFF_615(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g819),.DATA(g7761));
  MSFF DFF_616(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g822),.DATA(g7512));
  MSFF DFF_617(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g825),.DATA(g7513));
  MSFF DFF_618(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g828),.DATA(g7762));
  MSFF DFF_619(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g786),.DATA(g7763));
  MSFF DFF_620(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g789),.DATA(g7297));
  MSFF DFF_621(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g955),.DATA(g3857));
  MSFF DFF_622(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g959),.DATA(g5169));
  MSFF DFF_623(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g945),.DATA(g5170));
  MSFF DFF_624(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g948),.DATA(g8664));
  MSFF DFF_625(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g949),.DATA(g8665));
  MSFF DFF_626(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g950),.DATA(g8666));
  MSFF DFF_627(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g951),.DATA(g8667));
  MSFF DFF_628(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g952),.DATA(g8668));
  MSFF DFF_629(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g953),.DATA(g8669));
  MSFF DFF_630(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g954),.DATA(g8670));
  MSFF DFF_631(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g943),.DATA(g8671));
  MSFF DFF_632(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g936),.DATA(g5168));
  MSFF DFF_633(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g940),.DATA(g5735));
  MSFF DFF_634(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g942),.DATA(g2652));
  MSFF DFF_635(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g944),.DATA(g6372));
  MSFF DFF_636(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g855),.DATA(g8220));
  MSFF DFF_637(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g859),.DATA(g8221));
  MSFF DFF_638(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g863),.DATA(g8222));
  MSFF DFF_639(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g831),.DATA(g2651));
  MSFF DFF_640(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g834),.DATA(g2650));
  MSFF DFF_641(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g837),.DATA(g2649));
  MSFF DFF_642(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g840),.DATA(g2648));
  MSFF DFF_643(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g843),.DATA(g2647));
  MSFF DFF_644(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g846),.DATA(g2646));
  MSFF DFF_645(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g849),.DATA(g2645));
  MSFF DFF_646(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g852),.DATA(g2644));
  MSFF DFF_647(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g890),.DATA(g7102));
  MSFF DFF_648(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g878),.DATA(g890));
  MSFF DFF_649(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g926),.DATA(g878));
  MSFF DFF_650(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g875),.DATA(g5165));
  MSFF DFF_651(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g866),.DATA(g5163));
  MSFF DFF_652(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g929),.DATA(g3856));
  MSFF DFF_653(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g933),.DATA(g5166));
  MSFF DFF_654(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g871),.DATA(g5167));
  MSFF DFF_655(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g874),.DATA(g4654));
  MSFF DFF_656(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g891),.DATA(g3855));
  MSFF DFF_657(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g896),.DATA(g891));
  MSFF DFF_658(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g901),.DATA(g896));
  MSFF DFF_659(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g906),.DATA(g901));
  MSFF DFF_660(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g911),.DATA(g906));
  MSFF DFF_661(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g916),.DATA(g911));
  MSFF DFF_662(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g921),.DATA(g916));
  MSFF DFF_663(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g883),.DATA(g921));
  MSFF DFF_664(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g887),.DATA(g7099));
  MSFF DFF_665(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g888),.DATA(g7100));
  MSFF DFF_666(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g889),.DATA(g7101));
  MSFF DFF_667(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g741),.DATA(g9386));
  MSFF DFF_668(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g746),.DATA(g8956));
//
  NOT NOT1_0(.VSS(VSS),.VDD(VDD),.Y(I5353),.A(g3833));
  NOT NOT1_1(.VSS(VSS),.VDD(VDD),.Y(g206),.A(I5353));
  NOT NOT1_2(.VSS(VSS),.VDD(VDD),.Y(I5356),.A(g3837));
  NOT NOT1_3(.VSS(VSS),.VDD(VDD),.Y(g291),.A(I5356));
  NOT NOT1_4(.VSS(VSS),.VDD(VDD),.Y(I5359),.A(g3839));
  NOT NOT1_5(.VSS(VSS),.VDD(VDD),.Y(g372),.A(I5359));
  NOT NOT1_6(.VSS(VSS),.VDD(VDD),.Y(I5362),.A(g3841));
  NOT NOT1_7(.VSS(VSS),.VDD(VDD),.Y(g453),.A(I5362));
  NOT NOT1_8(.VSS(VSS),.VDD(VDD),.Y(I5365),.A(g3843));
  NOT NOT1_9(.VSS(VSS),.VDD(VDD),.Y(g534),.A(I5365));
  NOT NOT1_10(.VSS(VSS),.VDD(VDD),.Y(I5368),.A(g3853));
  NOT NOT1_11(.VSS(VSS),.VDD(VDD),.Y(g594),.A(I5368));
  NOT NOT1_12(.VSS(VSS),.VDD(VDD),.Y(I5371),.A(g633));
  NOT NOT1_13(.VSS(VSS),.VDD(VDD),.Y(g636),.A(I5371));
  NOT NOT1_14(.VSS(VSS),.VDD(VDD),.Y(I5374),.A(g634));
  NOT NOT1_15(.VSS(VSS),.VDD(VDD),.Y(g639),.A(I5374));
  NOT NOT1_16(.VSS(VSS),.VDD(VDD),.Y(I5377),.A(g635));
  NOT NOT1_17(.VSS(VSS),.VDD(VDD),.Y(g642),.A(I5377));
  NOT NOT1_18(.VSS(VSS),.VDD(VDD),.Y(I5380),.A(g645));
  NOT NOT1_19(.VSS(VSS),.VDD(VDD),.Y(g649),.A(I5380));
  NOT NOT1_20(.VSS(VSS),.VDD(VDD),.Y(I5383),.A(g647));
  NOT NOT1_21(.VSS(VSS),.VDD(VDD),.Y(g655),.A(I5383));
  NOT NOT1_22(.VSS(VSS),.VDD(VDD),.Y(I5386),.A(g648));
  NOT NOT1_23(.VSS(VSS),.VDD(VDD),.Y(g658),.A(I5386));
  NOT NOT1_24(.VSS(VSS),.VDD(VDD),.Y(I5389),.A(g690));
  NOT NOT1_25(.VSS(VSS),.VDD(VDD),.Y(g691),.A(I5389));
  NOT NOT1_26(.VSS(VSS),.VDD(VDD),.Y(I5392),.A(g694));
  NOT NOT1_27(.VSS(VSS),.VDD(VDD),.Y(g695),.A(I5392));
  NOT NOT1_28(.VSS(VSS),.VDD(VDD),.Y(I5395),.A(g698));
  NOT NOT1_29(.VSS(VSS),.VDD(VDD),.Y(g699),.A(I5395));
  NOT NOT1_30(.VSS(VSS),.VDD(VDD),.Y(I5398),.A(g702));
  NOT NOT1_31(.VSS(VSS),.VDD(VDD),.Y(g703),.A(I5398));
  NOT NOT1_32(.VSS(VSS),.VDD(VDD),.Y(I5401),.A(g723));
  NOT NOT1_33(.VSS(VSS),.VDD(VDD),.Y(g724),.A(I5401));
  NOT NOT1_34(.VSS(VSS),.VDD(VDD),.Y(I5404),.A(g722));
  NOT NOT1_35(.VSS(VSS),.VDD(VDD),.Y(g738),.A(I5404));
  NOT NOT1_36(.VSS(VSS),.VDD(VDD),.Y(I5407),.A(g4653));
  NOT NOT1_37(.VSS(VSS),.VDD(VDD),.Y(g785),.A(I5407));
  NOT NOT1_38(.VSS(VSS),.VDD(VDD),.Y(I5410),.A(g8866));
  NOT NOT1_39(.VSS(VSS),.VDD(VDD),.Y(g1006),.A(I5410));
  NOT NOT1_40(.VSS(VSS),.VDD(VDD),.Y(I5413),.A(g1016));
  NOT NOT1_41(.VSS(VSS),.VDD(VDD),.Y(g1011),.A(I5413));
  NOT NOT1_42(.VSS(VSS),.VDD(VDD),.Y(I5416),.A(g8868));
  NOT NOT1_43(.VSS(VSS),.VDD(VDD),.Y(g1015),.A(I5416));
  NOT NOT1_44(.VSS(VSS),.VDD(VDD),.Y(I5419),.A(g1603));
  NOT NOT1_45(.VSS(VSS),.VDD(VDD),.Y(g1017),.A(I5419));
  NOT NOT1_46(.VSS(VSS),.VDD(VDD),.Y(I5422),.A(g1234));
  NOT NOT1_47(.VSS(VSS),.VDD(VDD),.Y(g1235),.A(I5422));
  NOT NOT1_48(.VSS(VSS),.VDD(VDD),.Y(I5425),.A(g1245));
  NOT NOT1_49(.VSS(VSS),.VDD(VDD),.Y(g1246),.A(I5425));
  NOT NOT1_50(.VSS(VSS),.VDD(VDD),.Y(I5428),.A(g49));
  NOT NOT1_51(.VSS(VSS),.VDD(VDD),.Y(g1555),.A(I5428));
  NOT NOT1_52(.VSS(VSS),.VDD(VDD),.Y(g1556),.A(g65));
  NOT NOT1_53(.VSS(VSS),.VDD(VDD),.Y(I5432),.A(g1176));
  NOT NOT1_54(.VSS(VSS),.VDD(VDD),.Y(g1557),.A(I5432));
  NOT NOT1_55(.VSS(VSS),.VDD(VDD),.Y(I5435),.A(g1461));
  NOT NOT1_56(.VSS(VSS),.VDD(VDD),.Y(g1558),.A(I5435));
  NOT NOT1_57(.VSS(VSS),.VDD(VDD),.Y(g1562),.A(g636));
  NOT NOT1_58(.VSS(VSS),.VDD(VDD),.Y(g1563),.A(g639));
  NOT NOT1_59(.VSS(VSS),.VDD(VDD),.Y(g1564),.A(g642));
  NOT NOT1_60(.VSS(VSS),.VDD(VDD),.Y(g1565),.A(g649));
  NOT NOT1_61(.VSS(VSS),.VDD(VDD),.Y(g1566),.A(g652));
  NOT NOT1_62(.VSS(VSS),.VDD(VDD),.Y(g1567),.A(g655));
  NOT NOT1_63(.VSS(VSS),.VDD(VDD),.Y(g1568),.A(g658));
  NOT NOT1_64(.VSS(VSS),.VDD(VDD),.Y(g1569),.A(g661));
  NOT NOT1_65(.VSS(VSS),.VDD(VDD),.Y(g1570),.A(g665));
  NOT NOT1_66(.VSS(VSS),.VDD(VDD),.Y(g1571),.A(g669));
  NOT NOT1_67(.VSS(VSS),.VDD(VDD),.Y(g1572),.A(g673));
  NOT NOT1_68(.VSS(VSS),.VDD(VDD),.Y(g1573),.A(g677));
  NOT NOT1_69(.VSS(VSS),.VDD(VDD),.Y(g1574),.A(g681));
  NOT NOT1_70(.VSS(VSS),.VDD(VDD),.Y(g1575),.A(g685));
  NOT NOT1_71(.VSS(VSS),.VDD(VDD),.Y(g1576),.A(g691));
  NOT NOT1_72(.VSS(VSS),.VDD(VDD),.Y(g1577),.A(g695));
  NOT NOT1_73(.VSS(VSS),.VDD(VDD),.Y(g1578),.A(g699));
  NOT NOT1_74(.VSS(VSS),.VDD(VDD),.Y(g1579),.A(g703));
  NOT NOT1_75(.VSS(VSS),.VDD(VDD),.Y(g1580),.A(g706));
  NOT NOT1_76(.VSS(VSS),.VDD(VDD),.Y(g1581),.A(g710));
  NOT NOT1_77(.VSS(VSS),.VDD(VDD),.Y(g1582),.A(g714));
  NOT NOT1_78(.VSS(VSS),.VDD(VDD),.Y(g1583),.A(g718));
  NOT NOT1_79(.VSS(VSS),.VDD(VDD),.Y(g1584),.A(g738));
  NOT NOT1_80(.VSS(VSS),.VDD(VDD),.Y(g1585),.A(g724));
  NOT NOT1_81(.VSS(VSS),.VDD(VDD),.Y(g1586),.A(g730));
  NOT NOT1_82(.VSS(VSS),.VDD(VDD),.Y(g1587),.A(g734));
  NOT NOT1_83(.VSS(VSS),.VDD(VDD),.Y(g1588),.A(g741));
  NOT NOT1_84(.VSS(VSS),.VDD(VDD),.Y(g1589),.A(g746));
  NOT NOT1_85(.VSS(VSS),.VDD(VDD),.Y(I5466),.A(g926));
  NOT NOT1_86(.VSS(VSS),.VDD(VDD),.Y(g1590),.A(I5466));
  NOT NOT1_87(.VSS(VSS),.VDD(VDD),.Y(g1597),.A(g973));
  NOT NOT1_88(.VSS(VSS),.VDD(VDD),.Y(g1600),.A(g976));
  NOT NOT1_89(.VSS(VSS),.VDD(VDD),.Y(I5471),.A(g1029));
  NOT NOT1_90(.VSS(VSS),.VDD(VDD),.Y(g1603),.A(I5471));
  NOT NOT1_91(.VSS(VSS),.VDD(VDD),.Y(g1611),.A(g1073));
  NOT NOT1_92(.VSS(VSS),.VDD(VDD),.Y(I5475),.A(g1084));
  NOT NOT1_93(.VSS(VSS),.VDD(VDD),.Y(g1612),.A(I5475));
  NOT NOT1_94(.VSS(VSS),.VDD(VDD),.Y(I5478),.A(g1148));
  NOT NOT1_95(.VSS(VSS),.VDD(VDD),.Y(g1616),.A(I5478));
  NOT NOT1_96(.VSS(VSS),.VDD(VDD),.Y(g1637),.A(g1087));
  NOT NOT1_97(.VSS(VSS),.VDD(VDD),.Y(g1638),.A(g1092));
  NOT NOT1_98(.VSS(VSS),.VDD(VDD),.Y(g1639),.A(g1207));
  NOT NOT1_99(.VSS(VSS),.VDD(VDD),.Y(g1643),.A(g1211));
  NOT NOT1_100(.VSS(VSS),.VDD(VDD),.Y(g1646),.A(g1214));
  NOT NOT1_101(.VSS(VSS),.VDD(VDD),.Y(g1649),.A(g1217));
  NOT NOT1_102(.VSS(VSS),.VDD(VDD),.Y(g1652),.A(g1220));
  NOT NOT1_103(.VSS(VSS),.VDD(VDD),.Y(g1655),.A(g1231));
  NOT NOT1_104(.VSS(VSS),.VDD(VDD),.Y(g1658),.A(g1313));
  NOT NOT1_105(.VSS(VSS),.VDD(VDD),.Y(g1661),.A(g1405));
  NOT NOT1_106(.VSS(VSS),.VDD(VDD),.Y(g1662),.A(g1412));
  NOT NOT1_107(.VSS(VSS),.VDD(VDD),.Y(g1663),.A(g1416));
  NOT NOT1_108(.VSS(VSS),.VDD(VDD),.Y(g1664),.A(g1462));
  NOT NOT1_109(.VSS(VSS),.VDD(VDD),.Y(g1665),.A(g1467));
  NOT NOT1_110(.VSS(VSS),.VDD(VDD),.Y(g1666),.A(g1472));
  NOT NOT1_111(.VSS(VSS),.VDD(VDD),.Y(g1667),.A(g1481));
  NOT NOT1_112(.VSS(VSS),.VDD(VDD),.Y(g1670),.A(g1489));
  NOT NOT1_113(.VSS(VSS),.VDD(VDD),.Y(g1671),.A(g1494));
  NOT NOT1_114(.VSS(VSS),.VDD(VDD),.Y(g1672),.A(g1499));
  NOT NOT1_115(.VSS(VSS),.VDD(VDD),.Y(g1673),.A(g1504));
  NOT NOT1_116(.VSS(VSS),.VDD(VDD),.Y(g1674),.A(g1514));
  NOT NOT1_117(.VSS(VSS),.VDD(VDD),.Y(g1675),.A(g1519));
  NOT NOT1_118(.VSS(VSS),.VDD(VDD),.Y(g1676),.A(g727));
  NOT NOT1_119(.VSS(VSS),.VDD(VDD),.Y(g1677),.A(g1532));
  NOT NOT1_120(.VSS(VSS),.VDD(VDD),.Y(I5512),.A(g557));
  NOT NOT1_121(.VSS(VSS),.VDD(VDD),.Y(g1679),.A(I5512));
  NOT NOT1_122(.VSS(VSS),.VDD(VDD),.Y(I5515),.A(g567));
  NOT NOT1_123(.VSS(VSS),.VDD(VDD),.Y(g1680),.A(I5515));
  NOT NOT1_124(.VSS(VSS),.VDD(VDD),.Y(g1681),.A(g929));
  NOT NOT1_125(.VSS(VSS),.VDD(VDD),.Y(g1683),.A(g795));
  NOT NOT1_126(.VSS(VSS),.VDD(VDD),.Y(g1684),.A(g1));
  NOT NOT1_127(.VSS(VSS),.VDD(VDD),.Y(I5528),.A(g43));
  NOT NOT1_128(.VSS(VSS),.VDD(VDD),.Y(g1685),.A(I5528));
  NOT NOT1_129(.VSS(VSS),.VDD(VDD),.Y(I5531),.A(g866));
  NOT NOT1_130(.VSS(VSS),.VDD(VDD),.Y(g1686),.A(I5531));
  NOT NOT1_131(.VSS(VSS),.VDD(VDD),.Y(g1687),.A(g10));
  NOT NOT1_132(.VSS(VSS),.VDD(VDD),.Y(I5535),.A(g48));
  NOT NOT1_133(.VSS(VSS),.VDD(VDD),.Y(g1688),.A(I5535));
  NOT NOT1_134(.VSS(VSS),.VDD(VDD),.Y(g1689),.A(g855));
  NOT NOT1_135(.VSS(VSS),.VDD(VDD),.Y(g1694),.A(g21));
  NOT NOT1_136(.VSS(VSS),.VDD(VDD),.Y(g1695),.A(g778));
  NOT NOT1_137(.VSS(VSS),.VDD(VDD),.Y(I5542),.A(g1272));
  NOT NOT1_138(.VSS(VSS),.VDD(VDD),.Y(g1698),.A(I5542));
  NOT NOT1_139(.VSS(VSS),.VDD(VDD),.Y(I5545),.A(g1276));
  NOT NOT1_140(.VSS(VSS),.VDD(VDD),.Y(g1701),.A(I5545));
  NOT NOT1_141(.VSS(VSS),.VDD(VDD),.Y(I5548),.A(g1280));
  NOT NOT1_142(.VSS(VSS),.VDD(VDD),.Y(g1704),.A(I5548));
  NOT NOT1_143(.VSS(VSS),.VDD(VDD),.Y(g1707),.A(g955));
  NOT NOT1_144(.VSS(VSS),.VDD(VDD),.Y(I5552),.A(g1284));
  NOT NOT1_145(.VSS(VSS),.VDD(VDD),.Y(g1708),.A(I5552));
  NOT NOT1_146(.VSS(VSS),.VDD(VDD),.Y(I5555),.A(g1288));
  NOT NOT1_147(.VSS(VSS),.VDD(VDD),.Y(g1711),.A(I5555));
  NOT NOT1_148(.VSS(VSS),.VDD(VDD),.Y(I5559),.A(g1292));
  NOT NOT1_149(.VSS(VSS),.VDD(VDD),.Y(g1715),.A(I5559));
  NOT NOT1_150(.VSS(VSS),.VDD(VDD),.Y(I5562),.A(g1300));
  NOT NOT1_151(.VSS(VSS),.VDD(VDD),.Y(g1718),.A(I5562));
  NOT NOT1_152(.VSS(VSS),.VDD(VDD),.Y(I5565),.A(g1296));
  NOT NOT1_153(.VSS(VSS),.VDD(VDD),.Y(g1721),.A(I5565));
  NOT NOT1_154(.VSS(VSS),.VDD(VDD),.Y(I5568),.A(g1409));
  NOT NOT1_155(.VSS(VSS),.VDD(VDD),.Y(g1724),.A(I5568));
  NOT NOT1_156(.VSS(VSS),.VDD(VDD),.Y(g1726),.A(g158));
  NOT NOT1_157(.VSS(VSS),.VDD(VDD),.Y(g1727),.A(g596));
  NOT NOT1_158(.VSS(VSS),.VDD(VDD),.Y(g1732),.A(g1439));
  NOT NOT1_159(.VSS(VSS),.VDD(VDD),.Y(I5577),.A(g172));
  NOT NOT1_160(.VSS(VSS),.VDD(VDD),.Y(g1736),.A(I5577));
  NOT NOT1_161(.VSS(VSS),.VDD(VDD),.Y(g1737),.A(g597));
  NOT NOT1_162(.VSS(VSS),.VDD(VDD),.Y(g1738),.A(g741));
  NOT NOT1_163(.VSS(VSS),.VDD(VDD),.Y(g1742),.A(g1486));
  NOT NOT1_164(.VSS(VSS),.VDD(VDD),.Y(g1743),.A(g598));
  NOT NOT1_165(.VSS(VSS),.VDD(VDD),.Y(g1744),.A(g600));
  NOT NOT1_166(.VSS(VSS),.VDD(VDD),.Y(g1745),.A(g746));
  NOT NOT1_167(.VSS(VSS),.VDD(VDD),.Y(g1746),.A(g290));
  NOT NOT1_168(.VSS(VSS),.VDD(VDD),.Y(g1747),.A(g599));
  NOT NOT1_169(.VSS(VSS),.VDD(VDD),.Y(g1748),.A(g601));
  NOT NOT1_170(.VSS(VSS),.VDD(VDD),.Y(g1749),.A(g371));
  NOT NOT1_171(.VSS(VSS),.VDD(VDD),.Y(g1750),.A(g602));
  NOT NOT1_172(.VSS(VSS),.VDD(VDD),.Y(g1751),.A(g452));
  NOT NOT1_173(.VSS(VSS),.VDD(VDD),.Y(g1752),.A(g603));
  NOT NOT1_174(.VSS(VSS),.VDD(VDD),.Y(g1756),.A(g533));
  NOT NOT1_175(.VSS(VSS),.VDD(VDD),.Y(g1757),.A(g604));
  NOT NOT1_176(.VSS(VSS),.VDD(VDD),.Y(g1758),.A(g1084));
  NOT NOT1_177(.VSS(VSS),.VDD(VDD),.Y(I5605),.A(g58));
  NOT NOT1_178(.VSS(VSS),.VDD(VDD),.Y(g1760),.A(I5605));
  NOT NOT1_179(.VSS(VSS),.VDD(VDD),.Y(g1768),.A(g605));
  NOT NOT1_180(.VSS(VSS),.VDD(VDD),.Y(I5609),.A(g16));
  NOT NOT1_181(.VSS(VSS),.VDD(VDD),.Y(g1769),.A(I5609));
  NOT NOT1_182(.VSS(VSS),.VDD(VDD),.Y(g1770),.A(g606));
  NOT NOT1_183(.VSS(VSS),.VDD(VDD),.Y(g1771),.A(g609));
  NOT NOT1_184(.VSS(VSS),.VDD(VDD),.Y(g1772),.A(g607));
  NOT NOT1_185(.VSS(VSS),.VDD(VDD),.Y(g1773),.A(g610));
  NOT NOT1_186(.VSS(VSS),.VDD(VDD),.Y(I5616),.A(g979));
  NOT NOT1_187(.VSS(VSS),.VDD(VDD),.Y(g1774),.A(I5616));
  NOT NOT1_188(.VSS(VSS),.VDD(VDD),.Y(g1776),.A(g608));
  NOT NOT1_189(.VSS(VSS),.VDD(VDD),.Y(g1777),.A(g611));
  NOT NOT1_190(.VSS(VSS),.VDD(VDD),.Y(g1778),.A(g613));
  NOT NOT1_191(.VSS(VSS),.VDD(VDD),.Y(g1779),.A(g612));
  NOT NOT1_192(.VSS(VSS),.VDD(VDD),.Y(g1780),.A(g614));
  NOT NOT1_193(.VSS(VSS),.VDD(VDD),.Y(g1781),.A(g622));
  NOT NOT1_194(.VSS(VSS),.VDD(VDD),.Y(g1782),.A(g624));
  NOT NOT1_195(.VSS(VSS),.VDD(VDD),.Y(I5633),.A(g891));
  NOT NOT1_196(.VSS(VSS),.VDD(VDD),.Y(g1783),.A(I5633));
  NOT NOT1_197(.VSS(VSS),.VDD(VDD),.Y(I5636),.A(g891));
  NOT NOT1_198(.VSS(VSS),.VDD(VDD),.Y(g1784),.A(I5636));
  NOT NOT1_199(.VSS(VSS),.VDD(VDD),.Y(g1785),.A(g615));
  NOT NOT1_200(.VSS(VSS),.VDD(VDD),.Y(g1786),.A(g623));
  NOT NOT1_201(.VSS(VSS),.VDD(VDD),.Y(g1787),.A(g625));
  NOT NOT1_202(.VSS(VSS),.VDD(VDD),.Y(g1788),.A(g984));
  NOT NOT1_203(.VSS(VSS),.VDD(VDD),.Y(g1789),.A(g1034));
  NOT NOT1_204(.VSS(VSS),.VDD(VDD),.Y(g1792),.A(g616));
  NOT NOT1_205(.VSS(VSS),.VDD(VDD),.Y(g1793),.A(g626));
  NOT NOT1_206(.VSS(VSS),.VDD(VDD),.Y(I5646),.A(g883));
  NOT NOT1_207(.VSS(VSS),.VDD(VDD),.Y(g1794),.A(I5646));
  NOT NOT1_208(.VSS(VSS),.VDD(VDD),.Y(I5649),.A(g1389));
  NOT NOT1_209(.VSS(VSS),.VDD(VDD),.Y(g1795),.A(I5649));
  NOT NOT1_210(.VSS(VSS),.VDD(VDD),.Y(g1796),.A(g617));
  NOT NOT1_211(.VSS(VSS),.VDD(VDD),.Y(g1797),.A(g627));
  NOT NOT1_212(.VSS(VSS),.VDD(VDD),.Y(I5654),.A(g921));
  NOT NOT1_213(.VSS(VSS),.VDD(VDD),.Y(g1798),.A(I5654));
  NOT NOT1_214(.VSS(VSS),.VDD(VDD),.Y(I5657),.A(g921));
  NOT NOT1_215(.VSS(VSS),.VDD(VDD),.Y(g1799),.A(I5657));
  NOT NOT1_216(.VSS(VSS),.VDD(VDD),.Y(g1800),.A(g1477));
  NOT NOT1_217(.VSS(VSS),.VDD(VDD),.Y(g1801),.A(g618));
  NOT NOT1_218(.VSS(VSS),.VDD(VDD),.Y(g1802),.A(g628));
  NOT NOT1_219(.VSS(VSS),.VDD(VDD),.Y(g1803),.A(g758));
  NOT NOT1_220(.VSS(VSS),.VDD(VDD),.Y(I5664),.A(g916));
  NOT NOT1_221(.VSS(VSS),.VDD(VDD),.Y(g1804),.A(I5664));
  NOT NOT1_222(.VSS(VSS),.VDD(VDD),.Y(I5667),.A(g916));
  NOT NOT1_223(.VSS(VSS),.VDD(VDD),.Y(g1805),.A(I5667));
  NOT NOT1_224(.VSS(VSS),.VDD(VDD),.Y(I5670),.A(g941));
  NOT NOT1_225(.VSS(VSS),.VDD(VDD),.Y(g1806),.A(I5670));
  NOT NOT1_226(.VSS(VSS),.VDD(VDD),.Y(g1807),.A(g619));
  NOT NOT1_227(.VSS(VSS),.VDD(VDD),.Y(g1808),.A(g629));
  NOT NOT1_228(.VSS(VSS),.VDD(VDD),.Y(g1809),.A(g759));
  NOT NOT1_229(.VSS(VSS),.VDD(VDD),.Y(I5676),.A(g911));
  NOT NOT1_230(.VSS(VSS),.VDD(VDD),.Y(g1810),.A(I5676));
  NOT NOT1_231(.VSS(VSS),.VDD(VDD),.Y(I5679),.A(g911));
  NOT NOT1_232(.VSS(VSS),.VDD(VDD),.Y(g1811),.A(I5679));
  NOT NOT1_233(.VSS(VSS),.VDD(VDD),.Y(I5682),.A(g168));
  NOT NOT1_234(.VSS(VSS),.VDD(VDD),.Y(g1812),.A(I5682));
  NOT NOT1_235(.VSS(VSS),.VDD(VDD),.Y(g1813),.A(g620));
  NOT NOT1_236(.VSS(VSS),.VDD(VDD),.Y(g1814),.A(g630));
  NOT NOT1_237(.VSS(VSS),.VDD(VDD),.Y(g1815),.A(g760));
  NOT NOT1_238(.VSS(VSS),.VDD(VDD),.Y(g1816),.A(g767));
  NOT NOT1_239(.VSS(VSS),.VDD(VDD),.Y(I5689),.A(g906));
  NOT NOT1_240(.VSS(VSS),.VDD(VDD),.Y(g1817),.A(I5689));
  NOT NOT1_241(.VSS(VSS),.VDD(VDD),.Y(I5692),.A(g906));
  NOT NOT1_242(.VSS(VSS),.VDD(VDD),.Y(g1818),.A(I5692));
  NOT NOT1_243(.VSS(VSS),.VDD(VDD),.Y(g1820),.A(g621));
  NOT NOT1_244(.VSS(VSS),.VDD(VDD),.Y(g1821),.A(g631));
  NOT NOT1_245(.VSS(VSS),.VDD(VDD),.Y(g1822),.A(g761));
  NOT NOT1_246(.VSS(VSS),.VDD(VDD),.Y(g1823),.A(g768));
  NOT NOT1_247(.VSS(VSS),.VDD(VDD),.Y(I5706),.A(g901));
  NOT NOT1_248(.VSS(VSS),.VDD(VDD),.Y(g1824),.A(I5706));
  NOT NOT1_249(.VSS(VSS),.VDD(VDD),.Y(I5709),.A(g901));
  NOT NOT1_250(.VSS(VSS),.VDD(VDD),.Y(g1825),.A(I5709));
  NOT NOT1_251(.VSS(VSS),.VDD(VDD),.Y(g1826),.A(g632));
  NOT NOT1_252(.VSS(VSS),.VDD(VDD),.Y(g1827),.A(g762));
  NOT NOT1_253(.VSS(VSS),.VDD(VDD),.Y(g1828),.A(g769));
  NOT NOT1_254(.VSS(VSS),.VDD(VDD),.Y(I5715),.A(g896));
  NOT NOT1_255(.VSS(VSS),.VDD(VDD),.Y(g1829),.A(I5715));
  NOT NOT1_256(.VSS(VSS),.VDD(VDD),.Y(I5718),.A(g896));
  NOT NOT1_257(.VSS(VSS),.VDD(VDD),.Y(g1830),.A(I5718));
  NOT NOT1_258(.VSS(VSS),.VDD(VDD),.Y(g1831),.A(g689));
  NOT NOT1_259(.VSS(VSS),.VDD(VDD),.Y(g1832),.A(g763));
  NOT NOT1_260(.VSS(VSS),.VDD(VDD),.Y(g1833),.A(g770));
  NOT NOT1_261(.VSS(VSS),.VDD(VDD),.Y(g1837),.A(g1007));
  NOT NOT1_262(.VSS(VSS),.VDD(VDD),.Y(g1838),.A(g1450));
  NOT NOT1_263(.VSS(VSS),.VDD(VDD),.Y(g1842),.A(g764));
  NOT NOT1_264(.VSS(VSS),.VDD(VDD),.Y(g1843),.A(g771));
  NOT NOT1_265(.VSS(VSS),.VDD(VDD),.Y(g1847),.A(g765));
  NOT NOT1_266(.VSS(VSS),.VDD(VDD),.Y(g1848),.A(g772));
  NOT NOT1_267(.VSS(VSS),.VDD(VDD),.Y(I5732),.A(g859));
  NOT NOT1_268(.VSS(VSS),.VDD(VDD),.Y(g1849),.A(I5732));
  NOT NOT1_269(.VSS(VSS),.VDD(VDD),.Y(g1852),.A(g887));
  NOT NOT1_270(.VSS(VSS),.VDD(VDD),.Y(g1853),.A(g766));
  NOT NOT1_271(.VSS(VSS),.VDD(VDD),.Y(g1854),.A(g773));
  NOT NOT1_272(.VSS(VSS),.VDD(VDD),.Y(g1855),.A(g866));
  NOT NOT1_273(.VSS(VSS),.VDD(VDD),.Y(g1856),.A(g774));
  NOT NOT1_274(.VSS(VSS),.VDD(VDD),.Y(g1857),.A(g889));
  NOT NOT1_275(.VSS(VSS),.VDD(VDD),.Y(g1860),.A(g162));
  NOT NOT1_276(.VSS(VSS),.VDD(VDD),.Y(g1863),.A(g68));
  NOT NOT1_277(.VSS(VSS),.VDD(VDD),.Y(g1864),.A(g162));
  NOT NOT1_278(.VSS(VSS),.VDD(VDD),.Y(g1865),.A(g1013));
  NOT NOT1_279(.VSS(VSS),.VDD(VDD),.Y(g1866),.A(g71));
  NOT NOT1_280(.VSS(VSS),.VDD(VDD),.Y(g1867),.A(g878));
  NOT NOT1_281(.VSS(VSS),.VDD(VDD),.Y(I5747),.A(g1260));
  NOT NOT1_282(.VSS(VSS),.VDD(VDD),.Y(g1868),.A(I5747));
  NOT NOT1_283(.VSS(VSS),.VDD(VDD),.Y(g1869),.A(g74));
  NOT NOT1_284(.VSS(VSS),.VDD(VDD),.Y(I5751),.A(g963));
  NOT NOT1_285(.VSS(VSS),.VDD(VDD),.Y(g1870),.A(I5751));
  NOT NOT1_286(.VSS(VSS),.VDD(VDD),.Y(I5754),.A(g966));
  NOT NOT1_287(.VSS(VSS),.VDD(VDD),.Y(g1871),.A(I5754));
  NOT NOT1_288(.VSS(VSS),.VDD(VDD),.Y(g1876),.A(g77));
  NOT NOT1_289(.VSS(VSS),.VDD(VDD),.Y(g1877),.A(g595));
  NOT NOT1_290(.VSS(VSS),.VDD(VDD),.Y(g1878),.A(g80));
  NOT NOT1_291(.VSS(VSS),.VDD(VDD),.Y(I5763),.A(g1207));
  NOT NOT1_292(.VSS(VSS),.VDD(VDD),.Y(g1879),.A(I5763));
  NOT NOT1_293(.VSS(VSS),.VDD(VDD),.Y(I5766),.A(g1254));
  NOT NOT1_294(.VSS(VSS),.VDD(VDD),.Y(g1886),.A(I5766));
  NOT NOT1_295(.VSS(VSS),.VDD(VDD),.Y(g1887),.A(g83));
  NOT NOT1_296(.VSS(VSS),.VDD(VDD),.Y(g1888),.A(g781));
  NOT NOT1_297(.VSS(VSS),.VDD(VDD),.Y(g1889),.A(g1018));
  NOT NOT1_298(.VSS(VSS),.VDD(VDD),.Y(I5772),.A(g1240));
  NOT NOT1_299(.VSS(VSS),.VDD(VDD),.Y(g1894),.A(I5772));
  NOT NOT1_300(.VSS(VSS),.VDD(VDD),.Y(I5775),.A(g1240));
  NOT NOT1_301(.VSS(VSS),.VDD(VDD),.Y(g1895),.A(I5775));
  NOT NOT1_302(.VSS(VSS),.VDD(VDD),.Y(g1896),.A(g86));
  NOT NOT1_303(.VSS(VSS),.VDD(VDD),.Y(g1897),.A(g789));
  NOT NOT1_304(.VSS(VSS),.VDD(VDD),.Y(I5781),.A(g979));
  NOT NOT1_305(.VSS(VSS),.VDD(VDD),.Y(g1901),.A(I5781));
  NOT NOT1_306(.VSS(VSS),.VDD(VDD),.Y(g1904),.A(g1021));
  NOT NOT1_307(.VSS(VSS),.VDD(VDD),.Y(g1907),.A(g52));
  NOT NOT1_308(.VSS(VSS),.VDD(VDD),.Y(g1908),.A(g812));
  NOT NOT1_309(.VSS(VSS),.VDD(VDD),.Y(g1909),.A(g998));
  NOT NOT1_310(.VSS(VSS),.VDD(VDD),.Y(I5789),.A(g1524));
  NOT NOT1_311(.VSS(VSS),.VDD(VDD),.Y(g1911),.A(I5789));
  NOT NOT1_312(.VSS(VSS),.VDD(VDD),.Y(g1912),.A(g1524));
  NOT NOT1_313(.VSS(VSS),.VDD(VDD),.Y(g1916),.A(g775));
  NOT NOT1_314(.VSS(VSS),.VDD(VDD),.Y(I5795),.A(g1236));
  NOT NOT1_315(.VSS(VSS),.VDD(VDD),.Y(g1917),.A(I5795));
  NOT NOT1_316(.VSS(VSS),.VDD(VDD),.Y(g1918),.A(g822));
  NOT NOT1_317(.VSS(VSS),.VDD(VDD),.Y(g1922),.A(g1251));
  NOT NOT1_318(.VSS(VSS),.VDD(VDD),.Y(I5801),.A(g1424));
  NOT NOT1_319(.VSS(VSS),.VDD(VDD),.Y(g1923),.A(I5801));
  NOT NOT1_320(.VSS(VSS),.VDD(VDD),.Y(g1924),.A(g174));
  NOT NOT1_321(.VSS(VSS),.VDD(VDD),.Y(g1925),.A(g825));
  NOT NOT1_322(.VSS(VSS),.VDD(VDD),.Y(g1926),.A(g874));
  NOT NOT1_323(.VSS(VSS),.VDD(VDD),.Y(g1929),.A(g1224));
  NOT NOT1_324(.VSS(VSS),.VDD(VDD),.Y(g1933),.A(g1247));
  NOT NOT1_325(.VSS(VSS),.VDD(VDD),.Y(g1934),.A(g154));
  NOT NOT1_326(.VSS(VSS),.VDD(VDD),.Y(g1935),.A(g1280));
  NOT NOT1_327(.VSS(VSS),.VDD(VDD),.Y(g1938),.A(g1288));
  NOT NOT1_328(.VSS(VSS),.VDD(VDD),.Y(I5812),.A(g1243));
  NOT NOT1_329(.VSS(VSS),.VDD(VDD),.Y(g1941),.A(I5812));
  NOT NOT1_330(.VSS(VSS),.VDD(VDD),.Y(g1942),.A(g828));
  NOT NOT1_331(.VSS(VSS),.VDD(VDD),.Y(g1943),.A(g1025));
  NOT NOT1_332(.VSS(VSS),.VDD(VDD),.Y(I5817),.A(g1081));
  NOT NOT1_333(.VSS(VSS),.VDD(VDD),.Y(g1944),.A(I5817));
  NOT NOT1_334(.VSS(VSS),.VDD(VDD),.Y(g1945),.A(g1081));
  NOT NOT1_335(.VSS(VSS),.VDD(VDD),.Y(g1948),.A(g1250));
  NOT NOT1_336(.VSS(VSS),.VDD(VDD),.Y(g1949),.A(g1292));
  NOT NOT1_337(.VSS(VSS),.VDD(VDD),.Y(g1952),.A(g1333));
  NOT NOT1_338(.VSS(VSS),.VDD(VDD),.Y(g1958),.A(g786));
  NOT NOT1_339(.VSS(VSS),.VDD(VDD),.Y(g1959),.A(g1252));
  NOT NOT1_340(.VSS(VSS),.VDD(VDD),.Y(g1960),.A(g1268));
  NOT NOT1_341(.VSS(VSS),.VDD(VDD),.Y(g1961),.A(g1345));
  NOT NOT1_342(.VSS(VSS),.VDD(VDD),.Y(g1967),.A(g1432));
  NOT NOT1_343(.VSS(VSS),.VDD(VDD),.Y(I5831),.A(g1194));
  NOT NOT1_344(.VSS(VSS),.VDD(VDD),.Y(g1970),.A(I5831));
  NOT NOT1_345(.VSS(VSS),.VDD(VDD),.Y(g1974),.A(g803));
  NOT NOT1_346(.VSS(VSS),.VDD(VDD),.Y(g1975),.A(g1253));
  NOT NOT1_347(.VSS(VSS),.VDD(VDD),.Y(g1976),.A(g1269));
  NOT NOT1_348(.VSS(VSS),.VDD(VDD),.Y(g1977),.A(g1357));
  NOT NOT1_349(.VSS(VSS),.VDD(VDD),.Y(I5839),.A(g1198));
  NOT NOT1_350(.VSS(VSS),.VDD(VDD),.Y(g1983),.A(I5839));
  NOT NOT1_351(.VSS(VSS),.VDD(VDD),.Y(I5842),.A(g68));
  NOT NOT1_352(.VSS(VSS),.VDD(VDD),.Y(g1987),.A(I5842));
  NOT NOT1_353(.VSS(VSS),.VDD(VDD),.Y(g2006),.A(g806));
  NOT NOT1_354(.VSS(VSS),.VDD(VDD),.Y(g2007),.A(g1223));
  NOT NOT1_355(.VSS(VSS),.VDD(VDD),.Y(I5847),.A(g1360));
  NOT NOT1_356(.VSS(VSS),.VDD(VDD),.Y(g2011),.A(I5847));
  NOT NOT1_357(.VSS(VSS),.VDD(VDD),.Y(g2015),.A(g33));
  NOT NOT1_358(.VSS(VSS),.VDD(VDD),.Y(I5852),.A(g1202));
  NOT NOT1_359(.VSS(VSS),.VDD(VDD),.Y(g2016),.A(I5852));
  NOT NOT1_360(.VSS(VSS),.VDD(VDD),.Y(I5855),.A(g71));
  NOT NOT1_361(.VSS(VSS),.VDD(VDD),.Y(g2020),.A(I5855));
  NOT NOT1_362(.VSS(VSS),.VDD(VDD),.Y(g2038),.A(g809));
  NOT NOT1_363(.VSS(VSS),.VDD(VDD),.Y(g2039),.A(g1228));
  NOT NOT1_364(.VSS(VSS),.VDD(VDD),.Y(I5861),.A(g1313));
  NOT NOT1_365(.VSS(VSS),.VDD(VDD),.Y(g2044),.A(I5861));
  NOT NOT1_366(.VSS(VSS),.VDD(VDD),.Y(I5865),.A(g1206));
  NOT NOT1_367(.VSS(VSS),.VDD(VDD),.Y(g2052),.A(I5865));
  NOT NOT1_368(.VSS(VSS),.VDD(VDD),.Y(I5868),.A(g74));
  NOT NOT1_369(.VSS(VSS),.VDD(VDD),.Y(g2057),.A(I5868));
  NOT NOT1_370(.VSS(VSS),.VDD(VDD),.Y(g2073),.A(g1254));
  NOT NOT1_371(.VSS(VSS),.VDD(VDD),.Y(I5872),.A(g77));
  NOT NOT1_372(.VSS(VSS),.VDD(VDD),.Y(g2074),.A(I5872));
  NOT NOT1_373(.VSS(VSS),.VDD(VDD),.Y(g2091),.A(g819));
  NOT NOT1_374(.VSS(VSS),.VDD(VDD),.Y(g2092),.A(g1225));
  NOT NOT1_375(.VSS(VSS),.VDD(VDD),.Y(g2096),.A(g1226));
  NOT NOT1_376(.VSS(VSS),.VDD(VDD),.Y(g2100),.A(g1227));
  NOT NOT1_377(.VSS(VSS),.VDD(VDD),.Y(I5879),.A(g1267));
  NOT NOT1_378(.VSS(VSS),.VDD(VDD),.Y(g2104),.A(I5879));
  NOT NOT1_379(.VSS(VSS),.VDD(VDD),.Y(g2105),.A(g1444));
  NOT NOT1_380(.VSS(VSS),.VDD(VDD),.Y(I5883),.A(g80));
  NOT NOT1_381(.VSS(VSS),.VDD(VDD),.Y(g2106),.A(I5883));
  NOT NOT1_382(.VSS(VSS),.VDD(VDD),.Y(g2128),.A(g1284));
  NOT NOT1_383(.VSS(VSS),.VDD(VDD),.Y(g2131),.A(g1300));
  NOT NOT1_384(.VSS(VSS),.VDD(VDD),.Y(g2134),.A(g1317));
  NOT NOT1_385(.VSS(VSS),.VDD(VDD),.Y(I5889),.A(g83));
  NOT NOT1_386(.VSS(VSS),.VDD(VDD),.Y(g2137),.A(I5889));
  NOT NOT1_387(.VSS(VSS),.VDD(VDD),.Y(g2145),.A(g1296));
  NOT NOT1_388(.VSS(VSS),.VDD(VDD),.Y(g2148),.A(g1304));
  NOT NOT1_389(.VSS(VSS),.VDD(VDD),.Y(I5894),.A(g86));
  NOT NOT1_390(.VSS(VSS),.VDD(VDD),.Y(g2149),.A(I5894));
  NOT NOT1_391(.VSS(VSS),.VDD(VDD),.Y(I5897),.A(g173));
  NOT NOT1_392(.VSS(VSS),.VDD(VDD),.Y(g2157),.A(I5897));
  NOT NOT1_393(.VSS(VSS),.VDD(VDD),.Y(g2161),.A(g1454));
  NOT NOT1_394(.VSS(VSS),.VDD(VDD),.Y(I5901),.A(g52));
  NOT NOT1_395(.VSS(VSS),.VDD(VDD),.Y(g2162),.A(I5901));
  NOT NOT1_396(.VSS(VSS),.VDD(VDD),.Y(g2170),.A(g1229));
  NOT NOT1_397(.VSS(VSS),.VDD(VDD),.Y(g2174),.A(g1319));
  NOT NOT1_398(.VSS(VSS),.VDD(VDD),.Y(g2177),.A(g1322));
  NOT NOT1_399(.VSS(VSS),.VDD(VDD),.Y(g2180),.A(g1318));
  NOT NOT1_400(.VSS(VSS),.VDD(VDD),.Y(I5908),.A(g196));
  NOT NOT1_401(.VSS(VSS),.VDD(VDD),.Y(g2183),.A(I5908));
  NOT NOT1_402(.VSS(VSS),.VDD(VDD),.Y(I5911),.A(g216));
  NOT NOT1_403(.VSS(VSS),.VDD(VDD),.Y(g2184),.A(I5911));
  NOT NOT1_404(.VSS(VSS),.VDD(VDD),.Y(I5914),.A(g1097));
  NOT NOT1_405(.VSS(VSS),.VDD(VDD),.Y(g2185),.A(I5914));
  NOT NOT1_406(.VSS(VSS),.VDD(VDD),.Y(g2202),.A(g1321));
  NOT NOT1_407(.VSS(VSS),.VDD(VDD),.Y(g2205),.A(g13));
  NOT NOT1_408(.VSS(VSS),.VDD(VDD),.Y(I5920),.A(g219));
  NOT NOT1_409(.VSS(VSS),.VDD(VDD),.Y(g2207),.A(I5920));
  NOT NOT1_410(.VSS(VSS),.VDD(VDD),.Y(I5923),.A(g252));
  NOT NOT1_411(.VSS(VSS),.VDD(VDD),.Y(g2208),.A(I5923));
  NOT NOT1_412(.VSS(VSS),.VDD(VDD),.Y(I5926),.A(g297));
  NOT NOT1_413(.VSS(VSS),.VDD(VDD),.Y(g2209),.A(I5926));
  NOT NOT1_414(.VSS(VSS),.VDD(VDD),.Y(g2210),.A(g1326));
  NOT NOT1_415(.VSS(VSS),.VDD(VDD),.Y(g2215),.A(g1416));
  NOT NOT1_416(.VSS(VSS),.VDD(VDD),.Y(I5933),.A(g1158));
  NOT NOT1_417(.VSS(VSS),.VDD(VDD),.Y(g2216),.A(I5933));
  NOT NOT1_418(.VSS(VSS),.VDD(VDD),.Y(I5936),.A(g222));
  NOT NOT1_419(.VSS(VSS),.VDD(VDD),.Y(g2221),.A(I5936));
  NOT NOT1_420(.VSS(VSS),.VDD(VDD),.Y(I5939),.A(g275));
  NOT NOT1_421(.VSS(VSS),.VDD(VDD),.Y(g2222),.A(I5939));
  NOT NOT1_422(.VSS(VSS),.VDD(VDD),.Y(I5942),.A(g300));
  NOT NOT1_423(.VSS(VSS),.VDD(VDD),.Y(g2223),.A(I5942));
  NOT NOT1_424(.VSS(VSS),.VDD(VDD),.Y(I5945),.A(g333));
  NOT NOT1_425(.VSS(VSS),.VDD(VDD),.Y(g2224),.A(I5945));
  NOT NOT1_426(.VSS(VSS),.VDD(VDD),.Y(I5948),.A(g378));
  NOT NOT1_427(.VSS(VSS),.VDD(VDD),.Y(g2225),.A(I5948));
  NOT NOT1_428(.VSS(VSS),.VDD(VDD),.Y(g2226),.A(g1320));
  NOT NOT1_429(.VSS(VSS),.VDD(VDD),.Y(I5954),.A(g89));
  NOT NOT1_430(.VSS(VSS),.VDD(VDD),.Y(g2231),.A(I5954));
  NOT NOT1_431(.VSS(VSS),.VDD(VDD),.Y(I5957),.A(g110));
  NOT NOT1_432(.VSS(VSS),.VDD(VDD),.Y(g2232),.A(I5957));
  NOT NOT1_433(.VSS(VSS),.VDD(VDD),.Y(I5960),.A(g187));
  NOT NOT1_434(.VSS(VSS),.VDD(VDD),.Y(g2233),.A(I5960));
  NOT NOT1_435(.VSS(VSS),.VDD(VDD),.Y(I5963),.A(g225));
  NOT NOT1_436(.VSS(VSS),.VDD(VDD),.Y(g2234),.A(I5963));
  NOT NOT1_437(.VSS(VSS),.VDD(VDD),.Y(I5966),.A(g278));
  NOT NOT1_438(.VSS(VSS),.VDD(VDD),.Y(g2235),.A(I5966));
  NOT NOT1_439(.VSS(VSS),.VDD(VDD),.Y(I5969),.A(g303));
  NOT NOT1_440(.VSS(VSS),.VDD(VDD),.Y(g2236),.A(I5969));
  NOT NOT1_441(.VSS(VSS),.VDD(VDD),.Y(I5972),.A(g356));
  NOT NOT1_442(.VSS(VSS),.VDD(VDD),.Y(g2237),.A(I5972));
  NOT NOT1_443(.VSS(VSS),.VDD(VDD),.Y(I5975),.A(g381));
  NOT NOT1_444(.VSS(VSS),.VDD(VDD),.Y(g2238),.A(I5975));
  NOT NOT1_445(.VSS(VSS),.VDD(VDD),.Y(I5978),.A(g414));
  NOT NOT1_446(.VSS(VSS),.VDD(VDD),.Y(g2239),.A(I5978));
  NOT NOT1_447(.VSS(VSS),.VDD(VDD),.Y(I5981),.A(g459));
  NOT NOT1_448(.VSS(VSS),.VDD(VDD),.Y(g2240),.A(I5981));
  NOT NOT1_449(.VSS(VSS),.VDD(VDD),.Y(I5984),.A(g540));
  NOT NOT1_450(.VSS(VSS),.VDD(VDD),.Y(g2241),.A(I5984));
  NOT NOT1_451(.VSS(VSS),.VDD(VDD),.Y(g2242),.A(g985));
  NOT NOT1_452(.VSS(VSS),.VDD(VDD),.Y(g2245),.A(g999));
  NOT NOT1_453(.VSS(VSS),.VDD(VDD),.Y(I5989),.A(g1460));
  NOT NOT1_454(.VSS(VSS),.VDD(VDD),.Y(g2246),.A(I5989));
  NOT NOT1_455(.VSS(VSS),.VDD(VDD),.Y(g2253),.A(g1323));
  NOT NOT1_456(.VSS(VSS),.VDD(VDD),.Y(g2256),.A(g1324));
  NOT NOT1_457(.VSS(VSS),.VDD(VDD),.Y(g2259),.A(g1325));
  NOT NOT1_458(.VSS(VSS),.VDD(VDD),.Y(g2263),.A(g1394));
  NOT NOT1_459(.VSS(VSS),.VDD(VDD),.Y(I5997),.A(g114));
  NOT NOT1_460(.VSS(VSS),.VDD(VDD),.Y(g2264),.A(I5997));
  NOT NOT1_461(.VSS(VSS),.VDD(VDD),.Y(I6000),.A(g202));
  NOT NOT1_462(.VSS(VSS),.VDD(VDD),.Y(g2265),.A(I6000));
  NOT NOT1_463(.VSS(VSS),.VDD(VDD),.Y(I6003),.A(g228));
  NOT NOT1_464(.VSS(VSS),.VDD(VDD),.Y(g2266),.A(I6003));
  NOT NOT1_465(.VSS(VSS),.VDD(VDD),.Y(I6006),.A(g306));
  NOT NOT1_466(.VSS(VSS),.VDD(VDD),.Y(g2267),.A(I6006));
  NOT NOT1_467(.VSS(VSS),.VDD(VDD),.Y(I6009),.A(g359));
  NOT NOT1_468(.VSS(VSS),.VDD(VDD),.Y(g2268),.A(I6009));
  NOT NOT1_469(.VSS(VSS),.VDD(VDD),.Y(I6012),.A(g384));
  NOT NOT1_470(.VSS(VSS),.VDD(VDD),.Y(g2269),.A(I6012));
  NOT NOT1_471(.VSS(VSS),.VDD(VDD),.Y(I6015),.A(g437));
  NOT NOT1_472(.VSS(VSS),.VDD(VDD),.Y(g2270),.A(I6015));
  NOT NOT1_473(.VSS(VSS),.VDD(VDD),.Y(I6018),.A(g462));
  NOT NOT1_474(.VSS(VSS),.VDD(VDD),.Y(g2271),.A(I6018));
  NOT NOT1_475(.VSS(VSS),.VDD(VDD),.Y(I6021),.A(g495));
  NOT NOT1_476(.VSS(VSS),.VDD(VDD),.Y(g2272),.A(I6021));
  NOT NOT1_477(.VSS(VSS),.VDD(VDD),.Y(I6024),.A(g544));
  NOT NOT1_478(.VSS(VSS),.VDD(VDD),.Y(g2273),.A(I6024));
  NOT NOT1_479(.VSS(VSS),.VDD(VDD),.Y(g2274),.A(g782));
  NOT NOT1_480(.VSS(VSS),.VDD(VDD),.Y(g2275),.A(g990));
  NOT NOT1_481(.VSS(VSS),.VDD(VDD),.Y(I6029),.A(g1207));
  NOT NOT1_482(.VSS(VSS),.VDD(VDD),.Y(g2276),.A(I6029));
  NOT NOT1_483(.VSS(VSS),.VDD(VDD),.Y(g2282),.A(g1400));
  NOT NOT1_484(.VSS(VSS),.VDD(VDD),.Y(I6033),.A(g3));
  NOT NOT1_485(.VSS(VSS),.VDD(VDD),.Y(g2283),.A(I6033));
  NOT NOT1_486(.VSS(VSS),.VDD(VDD),.Y(I6036),.A(g130));
  NOT NOT1_487(.VSS(VSS),.VDD(VDD),.Y(g2284),.A(I6036));
  NOT NOT1_488(.VSS(VSS),.VDD(VDD),.Y(I6039),.A(g207));
  NOT NOT1_489(.VSS(VSS),.VDD(VDD),.Y(g2285),.A(I6039));
  NOT NOT1_490(.VSS(VSS),.VDD(VDD),.Y(I6042),.A(g237));
  NOT NOT1_491(.VSS(VSS),.VDD(VDD),.Y(g2286),.A(I6042));
  NOT NOT1_492(.VSS(VSS),.VDD(VDD),.Y(I6045),.A(g309));
  NOT NOT1_493(.VSS(VSS),.VDD(VDD),.Y(g2287),.A(I6045));
  NOT NOT1_494(.VSS(VSS),.VDD(VDD),.Y(I6048),.A(g387));
  NOT NOT1_495(.VSS(VSS),.VDD(VDD),.Y(g2288),.A(I6048));
  NOT NOT1_496(.VSS(VSS),.VDD(VDD),.Y(I6051),.A(g440));
  NOT NOT1_497(.VSS(VSS),.VDD(VDD),.Y(g2289),.A(I6051));
  NOT NOT1_498(.VSS(VSS),.VDD(VDD),.Y(I6054),.A(g465));
  NOT NOT1_499(.VSS(VSS),.VDD(VDD),.Y(g2290),.A(I6054));
  NOT NOT1_500(.VSS(VSS),.VDD(VDD),.Y(I6057),.A(g518));
  NOT NOT1_501(.VSS(VSS),.VDD(VDD),.Y(g2291),.A(I6057));
  NOT NOT1_502(.VSS(VSS),.VDD(VDD),.Y(I6060),.A(g580));
  NOT NOT1_503(.VSS(VSS),.VDD(VDD),.Y(g2292),.A(I6060));
  NOT NOT1_504(.VSS(VSS),.VDD(VDD),.Y(g2293),.A(g888));
  NOT NOT1_505(.VSS(VSS),.VDD(VDD),.Y(g2295),.A(g995));
  NOT NOT1_506(.VSS(VSS),.VDD(VDD),.Y(I6072),.A(g1211));
  NOT NOT1_507(.VSS(VSS),.VDD(VDD),.Y(g2298),.A(I6072));
  NOT NOT1_508(.VSS(VSS),.VDD(VDD),.Y(I6075),.A(g2));
  NOT NOT1_509(.VSS(VSS),.VDD(VDD),.Y(g2306),.A(I6075));
  NOT NOT1_510(.VSS(VSS),.VDD(VDD),.Y(I6078),.A(g95));
  NOT NOT1_511(.VSS(VSS),.VDD(VDD),.Y(g2307),.A(I6078));
  NOT NOT1_512(.VSS(VSS),.VDD(VDD),.Y(I6081),.A(g118));
  NOT NOT1_513(.VSS(VSS),.VDD(VDD),.Y(g2308),.A(I6081));
  NOT NOT1_514(.VSS(VSS),.VDD(VDD),.Y(I6084),.A(g240));
  NOT NOT1_515(.VSS(VSS),.VDD(VDD),.Y(g2309),.A(I6084));
  NOT NOT1_516(.VSS(VSS),.VDD(VDD),.Y(I6087),.A(g318));
  NOT NOT1_517(.VSS(VSS),.VDD(VDD),.Y(g2310),.A(I6087));
  NOT NOT1_518(.VSS(VSS),.VDD(VDD),.Y(I6090),.A(g390));
  NOT NOT1_519(.VSS(VSS),.VDD(VDD),.Y(g2311),.A(I6090));
  NOT NOT1_520(.VSS(VSS),.VDD(VDD),.Y(I6093),.A(g468));
  NOT NOT1_521(.VSS(VSS),.VDD(VDD),.Y(g2312),.A(I6093));
  NOT NOT1_522(.VSS(VSS),.VDD(VDD),.Y(I6096),.A(g521));
  NOT NOT1_523(.VSS(VSS),.VDD(VDD),.Y(g2313),.A(I6096));
  NOT NOT1_524(.VSS(VSS),.VDD(VDD),.Y(I6099),.A(g584));
  NOT NOT1_525(.VSS(VSS),.VDD(VDD),.Y(g2314),.A(I6099));
  NOT NOT1_526(.VSS(VSS),.VDD(VDD),.Y(I6109),.A(g1214));
  NOT NOT1_527(.VSS(VSS),.VDD(VDD),.Y(g2316),.A(I6109));
  NOT NOT1_528(.VSS(VSS),.VDD(VDD),.Y(I6112),.A(g4));
  NOT NOT1_529(.VSS(VSS),.VDD(VDD),.Y(g2323),.A(I6112));
  NOT NOT1_530(.VSS(VSS),.VDD(VDD),.Y(I6115),.A(g134));
  NOT NOT1_531(.VSS(VSS),.VDD(VDD),.Y(g2324),.A(I6115));
  NOT NOT1_532(.VSS(VSS),.VDD(VDD),.Y(I6118),.A(g243));
  NOT NOT1_533(.VSS(VSS),.VDD(VDD),.Y(g2325),.A(I6118));
  NOT NOT1_534(.VSS(VSS),.VDD(VDD),.Y(I6121),.A(g321));
  NOT NOT1_535(.VSS(VSS),.VDD(VDD),.Y(g2326),.A(I6121));
  NOT NOT1_536(.VSS(VSS),.VDD(VDD),.Y(I6124),.A(g399));
  NOT NOT1_537(.VSS(VSS),.VDD(VDD),.Y(g2327),.A(I6124));
  NOT NOT1_538(.VSS(VSS),.VDD(VDD),.Y(I6127),.A(g471));
  NOT NOT1_539(.VSS(VSS),.VDD(VDD),.Y(g2328),.A(I6127));
  NOT NOT1_540(.VSS(VSS),.VDD(VDD),.Y(I6130),.A(g560));
  NOT NOT1_541(.VSS(VSS),.VDD(VDD),.Y(g2329),.A(I6130));
  NOT NOT1_542(.VSS(VSS),.VDD(VDD),.Y(g2331),.A(g933));
  NOT NOT1_543(.VSS(VSS),.VDD(VDD),.Y(g2332),.A(g926));
  NOT NOT1_544(.VSS(VSS),.VDD(VDD),.Y(I6143),.A(g1217));
  NOT NOT1_545(.VSS(VSS),.VDD(VDD),.Y(g2334),.A(I6143));
  NOT NOT1_546(.VSS(VSS),.VDD(VDD),.Y(g2340),.A(g1327));
  NOT NOT1_547(.VSS(VSS),.VDD(VDD),.Y(g2343),.A(g1392));
  NOT NOT1_548(.VSS(VSS),.VDD(VDD),.Y(I6148),.A(g5));
  NOT NOT1_549(.VSS(VSS),.VDD(VDD),.Y(g2344),.A(I6148));
  NOT NOT1_550(.VSS(VSS),.VDD(VDD),.Y(I6151),.A(g12));
  NOT NOT1_551(.VSS(VSS),.VDD(VDD),.Y(g2345),.A(I6151));
  NOT NOT1_552(.VSS(VSS),.VDD(VDD),.Y(I6154),.A(g122));
  NOT NOT1_553(.VSS(VSS),.VDD(VDD),.Y(g2346),.A(I6154));
  NOT NOT1_554(.VSS(VSS),.VDD(VDD),.Y(I6157),.A(g246));
  NOT NOT1_555(.VSS(VSS),.VDD(VDD),.Y(g2347),.A(I6157));
  NOT NOT1_556(.VSS(VSS),.VDD(VDD),.Y(I6160),.A(g324));
  NOT NOT1_557(.VSS(VSS),.VDD(VDD),.Y(g2348),.A(I6160));
  NOT NOT1_558(.VSS(VSS),.VDD(VDD),.Y(I6163),.A(g402));
  NOT NOT1_559(.VSS(VSS),.VDD(VDD),.Y(g2349),.A(I6163));
  NOT NOT1_560(.VSS(VSS),.VDD(VDD),.Y(I6166),.A(g480));
  NOT NOT1_561(.VSS(VSS),.VDD(VDD),.Y(g2350),.A(I6166));
  NOT NOT1_562(.VSS(VSS),.VDD(VDD),.Y(g2351),.A(g792));
  NOT NOT1_563(.VSS(VSS),.VDD(VDD),.Y(g2353),.A(g871));
  NOT NOT1_564(.VSS(VSS),.VDD(VDD),.Y(I6178),.A(g1220));
  NOT NOT1_565(.VSS(VSS),.VDD(VDD),.Y(g2354),.A(I6178));
  NOT NOT1_566(.VSS(VSS),.VDD(VDD),.Y(g2359),.A(g1397));
  NOT NOT1_567(.VSS(VSS),.VDD(VDD),.Y(g2360),.A(g1435));
  NOT NOT1_568(.VSS(VSS),.VDD(VDD),.Y(I6183),.A(g6));
  NOT NOT1_569(.VSS(VSS),.VDD(VDD),.Y(g2361),.A(I6183));
  NOT NOT1_570(.VSS(VSS),.VDD(VDD),.Y(I6186),.A(g138));
  NOT NOT1_571(.VSS(VSS),.VDD(VDD),.Y(g2362),.A(I6186));
  NOT NOT1_572(.VSS(VSS),.VDD(VDD),.Y(I6189),.A(g249));
  NOT NOT1_573(.VSS(VSS),.VDD(VDD),.Y(g2363),.A(I6189));
  NOT NOT1_574(.VSS(VSS),.VDD(VDD),.Y(I6192),.A(g327));
  NOT NOT1_575(.VSS(VSS),.VDD(VDD),.Y(g2364),.A(I6192));
  NOT NOT1_576(.VSS(VSS),.VDD(VDD),.Y(I6195),.A(g405));
  NOT NOT1_577(.VSS(VSS),.VDD(VDD),.Y(g2365),.A(I6195));
  NOT NOT1_578(.VSS(VSS),.VDD(VDD),.Y(I6198),.A(g483));
  NOT NOT1_579(.VSS(VSS),.VDD(VDD),.Y(g2366),.A(I6198));
  NOT NOT1_580(.VSS(VSS),.VDD(VDD),.Y(g2371),.A(g944));
  NOT NOT1_581(.VSS(VSS),.VDD(VDD),.Y(I6214),.A(g7));
  NOT NOT1_582(.VSS(VSS),.VDD(VDD),.Y(g2372),.A(I6214));
  NOT NOT1_583(.VSS(VSS),.VDD(VDD),.Y(I6217),.A(g105));
  NOT NOT1_584(.VSS(VSS),.VDD(VDD),.Y(g2373),.A(I6217));
  NOT NOT1_585(.VSS(VSS),.VDD(VDD),.Y(I6220),.A(g126));
  NOT NOT1_586(.VSS(VSS),.VDD(VDD),.Y(g2374),.A(I6220));
  NOT NOT1_587(.VSS(VSS),.VDD(VDD),.Y(I6223),.A(g330));
  NOT NOT1_588(.VSS(VSS),.VDD(VDD),.Y(g2375),.A(I6223));
  NOT NOT1_589(.VSS(VSS),.VDD(VDD),.Y(I6226),.A(g408));
  NOT NOT1_590(.VSS(VSS),.VDD(VDD),.Y(g2376),.A(I6226));
  NOT NOT1_591(.VSS(VSS),.VDD(VDD),.Y(I6229),.A(g486));
  NOT NOT1_592(.VSS(VSS),.VDD(VDD),.Y(g2377),.A(I6229));
  NOT NOT1_593(.VSS(VSS),.VDD(VDD),.Y(I6239),.A(g8));
  NOT NOT1_594(.VSS(VSS),.VDD(VDD),.Y(g2379),.A(I6239));
  NOT NOT1_595(.VSS(VSS),.VDD(VDD),.Y(I6242),.A(g1554));
  NOT NOT1_596(.VSS(VSS),.VDD(VDD),.Y(g2380),.A(I6242));
  NOT NOT1_597(.VSS(VSS),.VDD(VDD),.Y(I6245),.A(g142));
  NOT NOT1_598(.VSS(VSS),.VDD(VDD),.Y(g2381),.A(I6245));
  NOT NOT1_599(.VSS(VSS),.VDD(VDD),.Y(I6248),.A(g411));
  NOT NOT1_600(.VSS(VSS),.VDD(VDD),.Y(g2382),.A(I6248));
  NOT NOT1_601(.VSS(VSS),.VDD(VDD),.Y(I6251),.A(g489));
  NOT NOT1_602(.VSS(VSS),.VDD(VDD),.Y(g2383),.A(I6251));
  NOT NOT1_603(.VSS(VSS),.VDD(VDD),.Y(I6254),.A(g536));
  NOT NOT1_604(.VSS(VSS),.VDD(VDD),.Y(g2384),.A(I6254));
  NOT NOT1_605(.VSS(VSS),.VDD(VDD),.Y(g2389),.A(g1230));
  NOT NOT1_606(.VSS(VSS),.VDD(VDD),.Y(g2392),.A(g11));
  NOT NOT1_607(.VSS(VSS),.VDD(VDD),.Y(I6267),.A(g100));
  NOT NOT1_608(.VSS(VSS),.VDD(VDD),.Y(g2393),.A(I6267));
  NOT NOT1_609(.VSS(VSS),.VDD(VDD),.Y(I6270),.A(g492));
  NOT NOT1_610(.VSS(VSS),.VDD(VDD),.Y(g2394),.A(I6270));
  NOT NOT1_611(.VSS(VSS),.VDD(VDD),.Y(g2396),.A(g1033));
  NOT NOT1_612(.VSS(VSS),.VDD(VDD),.Y(g2397),.A(g1272));
  NOT NOT1_613(.VSS(VSS),.VDD(VDD),.Y(g2401),.A(g22));
  NOT NOT1_614(.VSS(VSS),.VDD(VDD),.Y(g2402),.A(g29));
  NOT NOT1_615(.VSS(VSS),.VDD(VDD),.Y(g2403),.A(g1176));
  NOT NOT1_616(.VSS(VSS),.VDD(VDD),.Y(g2404),.A(g1276));
  NOT NOT1_617(.VSS(VSS),.VDD(VDD),.Y(I6286),.A(g1307));
  NOT NOT1_618(.VSS(VSS),.VDD(VDD),.Y(g2407),.A(I6286));
  NOT NOT1_619(.VSS(VSS),.VDD(VDD),.Y(g2424),.A(g1329));
  NOT NOT1_620(.VSS(VSS),.VDD(VDD),.Y(g2452),.A(g23));
  NOT NOT1_621(.VSS(VSS),.VDD(VDD),.Y(I6291),.A(g46));
  NOT NOT1_622(.VSS(VSS),.VDD(VDD),.Y(g2453),.A(I6291));
  NOT NOT1_623(.VSS(VSS),.VDD(VDD),.Y(I6294),.A(g1330));
  NOT NOT1_624(.VSS(VSS),.VDD(VDD),.Y(g2454),.A(I6294));
  NOT NOT1_625(.VSS(VSS),.VDD(VDD),.Y(g2457),.A(g24));
  NOT NOT1_626(.VSS(VSS),.VDD(VDD),.Y(g2458),.A(g30));
  NOT NOT1_627(.VSS(VSS),.VDD(VDD),.Y(I6299),.A(g47));
  NOT NOT1_628(.VSS(VSS),.VDD(VDD),.Y(g2459),.A(I6299));
  NOT NOT1_629(.VSS(VSS),.VDD(VDD),.Y(I6302),.A(g1313));
  NOT NOT1_630(.VSS(VSS),.VDD(VDD),.Y(g2460),.A(I6302));
  NOT NOT1_631(.VSS(VSS),.VDD(VDD),.Y(I6305),.A(g1333));
  NOT NOT1_632(.VSS(VSS),.VDD(VDD),.Y(g2467),.A(I6305));
  NOT NOT1_633(.VSS(VSS),.VDD(VDD),.Y(g2470),.A(g42));
  NOT NOT1_634(.VSS(VSS),.VDD(VDD),.Y(I6309),.A(g1336));
  NOT NOT1_635(.VSS(VSS),.VDD(VDD),.Y(g2471),.A(I6309));
  NOT NOT1_636(.VSS(VSS),.VDD(VDD),.Y(g2477),.A(g25));
  NOT NOT1_637(.VSS(VSS),.VDD(VDD),.Y(g2478),.A(g31));
  NOT NOT1_638(.VSS(VSS),.VDD(VDD),.Y(g2479),.A(g32));
  NOT NOT1_639(.VSS(VSS),.VDD(VDD),.Y(g2480),.A(g44));
  NOT NOT1_640(.VSS(VSS),.VDD(VDD),.Y(I6317),.A(g1339));
  NOT NOT1_641(.VSS(VSS),.VDD(VDD),.Y(g2481),.A(I6317));
  NOT NOT1_642(.VSS(VSS),.VDD(VDD),.Y(g2484),.A(g45));
  NOT NOT1_643(.VSS(VSS),.VDD(VDD),.Y(g2485),.A(g62));
  NOT NOT1_644(.VSS(VSS),.VDD(VDD),.Y(g2486),.A(g959));
  NOT NOT1_645(.VSS(VSS),.VDD(VDD),.Y(I6323),.A(g1342));
  NOT NOT1_646(.VSS(VSS),.VDD(VDD),.Y(g2487),.A(I6323));
  NOT NOT1_647(.VSS(VSS),.VDD(VDD),.Y(I6326),.A(g1443));
  NOT NOT1_648(.VSS(VSS),.VDD(VDD),.Y(g2490),.A(I6326));
  NOT NOT1_649(.VSS(VSS),.VDD(VDD),.Y(g2494),.A(g9));
  NOT NOT1_650(.VSS(VSS),.VDD(VDD),.Y(g2495),.A(g26));
  NOT NOT1_651(.VSS(VSS),.VDD(VDD),.Y(g2496),.A(g942));
  NOT NOT1_652(.VSS(VSS),.VDD(VDD),.Y(g2497),.A(g945));
  NOT NOT1_653(.VSS(VSS),.VDD(VDD),.Y(I6333),.A(g1345));
  NOT NOT1_654(.VSS(VSS),.VDD(VDD),.Y(g2498),.A(I6333));
  NOT NOT1_655(.VSS(VSS),.VDD(VDD),.Y(g2501),.A(g27));
  NOT NOT1_656(.VSS(VSS),.VDD(VDD),.Y(I6337),.A(g1348));
  NOT NOT1_657(.VSS(VSS),.VDD(VDD),.Y(g2502),.A(I6337));
  NOT NOT1_658(.VSS(VSS),.VDD(VDD),.Y(g2505),.A(g28));
  NOT NOT1_659(.VSS(VSS),.VDD(VDD),.Y(I6341),.A(g1351));
  NOT NOT1_660(.VSS(VSS),.VDD(VDD),.Y(g2506),.A(I6341));
  NOT NOT1_661(.VSS(VSS),.VDD(VDD),.Y(g2509),.A(g37));
  NOT NOT1_662(.VSS(VSS),.VDD(VDD),.Y(g2510),.A(g58));
  NOT NOT1_663(.VSS(VSS),.VDD(VDD),.Y(g2511),.A(g1328));
  NOT NOT1_664(.VSS(VSS),.VDD(VDD),.Y(g2514),.A(g1330));
  NOT NOT1_665(.VSS(VSS),.VDD(VDD),.Y(I6348),.A(g1354));
  NOT NOT1_666(.VSS(VSS),.VDD(VDD),.Y(g2517),.A(I6348));
  NOT NOT1_667(.VSS(VSS),.VDD(VDD),.Y(g2520),.A(g41));
  NOT NOT1_668(.VSS(VSS),.VDD(VDD),.Y(g2522),.A(g1342));
  NOT NOT1_669(.VSS(VSS),.VDD(VDD),.Y(I6354),.A(g1357));
  NOT NOT1_670(.VSS(VSS),.VDD(VDD),.Y(g2525),.A(I6354));
  NOT NOT1_671(.VSS(VSS),.VDD(VDD),.Y(g2528),.A(g1260));
  NOT NOT1_672(.VSS(VSS),.VDD(VDD),.Y(I6358),.A(g13));
  NOT NOT1_673(.VSS(VSS),.VDD(VDD),.Y(g2532),.A(I6358));
  NOT NOT1_674(.VSS(VSS),.VDD(VDD),.Y(g2533),.A(g1336));
  NOT NOT1_675(.VSS(VSS),.VDD(VDD),.Y(g2536),.A(g1354));
  NOT NOT1_676(.VSS(VSS),.VDD(VDD),.Y(I6363),.A(g16));
  NOT NOT1_677(.VSS(VSS),.VDD(VDD),.Y(g2539),.A(I6363));
  NOT NOT1_678(.VSS(VSS),.VDD(VDD),.Y(g2540),.A(g1339));
  NOT NOT1_679(.VSS(VSS),.VDD(VDD),.Y(g2543),.A(g1348));
  NOT NOT1_680(.VSS(VSS),.VDD(VDD),.Y(I6368),.A(g20));
  NOT NOT1_681(.VSS(VSS),.VDD(VDD),.Y(g2546),.A(I6368));
  NOT NOT1_682(.VSS(VSS),.VDD(VDD),.Y(I6371),.A(g33));
  NOT NOT1_683(.VSS(VSS),.VDD(VDD),.Y(g2547),.A(I6371));
  NOT NOT1_684(.VSS(VSS),.VDD(VDD),.Y(g2548),.A(g1351));
  NOT NOT1_685(.VSS(VSS),.VDD(VDD),.Y(g2551),.A(g1360));
  NOT NOT1_686(.VSS(VSS),.VDD(VDD),.Y(I6376),.A(g38));
  NOT NOT1_687(.VSS(VSS),.VDD(VDD),.Y(g2554),.A(I6376));
  NOT NOT1_688(.VSS(VSS),.VDD(VDD),.Y(g2555),.A(g936));
  NOT NOT1_689(.VSS(VSS),.VDD(VDD),.Y(g2556),.A(g1190));
  NOT NOT1_690(.VSS(VSS),.VDD(VDD),.Y(g2557),.A(g940));
  NOT NOT1_691(.VSS(VSS),.VDD(VDD),.Y(g2561),.A(g1555));
  NOT NOT1_692(.VSS(VSS),.VDD(VDD),.Y(g2562),.A(g1652));
  NOT NOT1_693(.VSS(VSS),.VDD(VDD),.Y(g2573),.A(g1649));
  NOT NOT1_694(.VSS(VSS),.VDD(VDD),.Y(g2584),.A(g1646));
  NOT NOT1_695(.VSS(VSS),.VDD(VDD),.Y(g2595),.A(g1643));
  NOT NOT1_696(.VSS(VSS),.VDD(VDD),.Y(g2605),.A(g1639));
  NOT NOT1_697(.VSS(VSS),.VDD(VDD),.Y(g2614),.A(g1562));
  NOT NOT1_698(.VSS(VSS),.VDD(VDD),.Y(g2615),.A(g1563));
  NOT NOT1_699(.VSS(VSS),.VDD(VDD),.Y(g2616),.A(g1564));
  NOT NOT1_700(.VSS(VSS),.VDD(VDD),.Y(g2617),.A(g1565));
  NOT NOT1_701(.VSS(VSS),.VDD(VDD),.Y(g2618),.A(g1566));
  NOT NOT1_702(.VSS(VSS),.VDD(VDD),.Y(g2621),.A(g1567));
  NOT NOT1_703(.VSS(VSS),.VDD(VDD),.Y(g2622),.A(g1568));
  NOT NOT1_704(.VSS(VSS),.VDD(VDD),.Y(g2623),.A(g1585));
  NOT NOT1_705(.VSS(VSS),.VDD(VDD),.Y(g2624),.A(g1569));
  NOT NOT1_706(.VSS(VSS),.VDD(VDD),.Y(g2625),.A(g1570));
  NOT NOT1_707(.VSS(VSS),.VDD(VDD),.Y(g2626),.A(g1571));
  NOT NOT1_708(.VSS(VSS),.VDD(VDD),.Y(g2627),.A(g1572));
  NOT NOT1_709(.VSS(VSS),.VDD(VDD),.Y(g2628),.A(g1573));
  NOT NOT1_710(.VSS(VSS),.VDD(VDD),.Y(g2629),.A(g1574));
  NOT NOT1_711(.VSS(VSS),.VDD(VDD),.Y(g2630),.A(g1575));
  NOT NOT1_712(.VSS(VSS),.VDD(VDD),.Y(g2631),.A(g1586));
  NOT NOT1_713(.VSS(VSS),.VDD(VDD),.Y(g2632),.A(g1576));
  NOT NOT1_714(.VSS(VSS),.VDD(VDD),.Y(g2633),.A(g1577));
  NOT NOT1_715(.VSS(VSS),.VDD(VDD),.Y(g2634),.A(g1578));
  NOT NOT1_716(.VSS(VSS),.VDD(VDD),.Y(g2635),.A(g1579));
  NOT NOT1_717(.VSS(VSS),.VDD(VDD),.Y(g2636),.A(g1580));
  NOT NOT1_718(.VSS(VSS),.VDD(VDD),.Y(g2637),.A(g1581));
  NOT NOT1_719(.VSS(VSS),.VDD(VDD),.Y(g2638),.A(g1582));
  NOT NOT1_720(.VSS(VSS),.VDD(VDD),.Y(g2639),.A(g1583));
  NOT NOT1_721(.VSS(VSS),.VDD(VDD),.Y(g2640),.A(g1584));
  NOT NOT1_722(.VSS(VSS),.VDD(VDD),.Y(g2641),.A(g1587));
  NOT NOT1_723(.VSS(VSS),.VDD(VDD),.Y(g2642),.A(g1588));
  NOT NOT1_724(.VSS(VSS),.VDD(VDD),.Y(g2643),.A(g1589));
  NOT NOT1_725(.VSS(VSS),.VDD(VDD),.Y(I6416),.A(g1794));
  NOT NOT1_726(.VSS(VSS),.VDD(VDD),.Y(g2644),.A(I6416));
  NOT NOT1_727(.VSS(VSS),.VDD(VDD),.Y(I6419),.A(g1799));
  NOT NOT1_728(.VSS(VSS),.VDD(VDD),.Y(g2645),.A(I6419));
  NOT NOT1_729(.VSS(VSS),.VDD(VDD),.Y(I6422),.A(g1805));
  NOT NOT1_730(.VSS(VSS),.VDD(VDD),.Y(g2646),.A(I6422));
  NOT NOT1_731(.VSS(VSS),.VDD(VDD),.Y(I6425),.A(g1811));
  NOT NOT1_732(.VSS(VSS),.VDD(VDD),.Y(g2647),.A(I6425));
  NOT NOT1_733(.VSS(VSS),.VDD(VDD),.Y(I6428),.A(g1818));
  NOT NOT1_734(.VSS(VSS),.VDD(VDD),.Y(g2648),.A(I6428));
  NOT NOT1_735(.VSS(VSS),.VDD(VDD),.Y(I6431),.A(g1825));
  NOT NOT1_736(.VSS(VSS),.VDD(VDD),.Y(g2649),.A(I6431));
  NOT NOT1_737(.VSS(VSS),.VDD(VDD),.Y(I6434),.A(g1830));
  NOT NOT1_738(.VSS(VSS),.VDD(VDD),.Y(g2650),.A(I6434));
  NOT NOT1_739(.VSS(VSS),.VDD(VDD),.Y(I6437),.A(g1784));
  NOT NOT1_740(.VSS(VSS),.VDD(VDD),.Y(g2651),.A(I6437));
  NOT NOT1_741(.VSS(VSS),.VDD(VDD),.Y(I6440),.A(g1806));
  NOT NOT1_742(.VSS(VSS),.VDD(VDD),.Y(g2652),.A(I6440));
  NOT NOT1_743(.VSS(VSS),.VDD(VDD),.Y(I6443),.A(g1774));
  NOT NOT1_744(.VSS(VSS),.VDD(VDD),.Y(g2653),.A(I6443));
  NOT NOT1_745(.VSS(VSS),.VDD(VDD),.Y(I6446),.A(g1812));
  NOT NOT1_746(.VSS(VSS),.VDD(VDD),.Y(g2654),.A(I6446));
  NOT NOT1_747(.VSS(VSS),.VDD(VDD),.Y(g2655),.A(g1611));
  NOT NOT1_748(.VSS(VSS),.VDD(VDD),.Y(g2659),.A(g1655));
  NOT NOT1_749(.VSS(VSS),.VDD(VDD),.Y(I6451),.A(g1895));
  NOT NOT1_750(.VSS(VSS),.VDD(VDD),.Y(g2660),.A(I6451));
  NOT NOT1_751(.VSS(VSS),.VDD(VDD),.Y(I6454),.A(g1868));
  NOT NOT1_752(.VSS(VSS),.VDD(VDD),.Y(g2661),.A(I6454));
  NOT NOT1_753(.VSS(VSS),.VDD(VDD),.Y(I6457),.A(g1886));
  NOT NOT1_754(.VSS(VSS),.VDD(VDD),.Y(g2662),.A(I6457));
  NOT NOT1_755(.VSS(VSS),.VDD(VDD),.Y(I6460),.A(g2104));
  NOT NOT1_756(.VSS(VSS),.VDD(VDD),.Y(g2663),.A(I6460));
  NOT NOT1_757(.VSS(VSS),.VDD(VDD),.Y(I6463),.A(g1769));
  NOT NOT1_758(.VSS(VSS),.VDD(VDD),.Y(g2664),.A(I6463));
  NOT NOT1_759(.VSS(VSS),.VDD(VDD),.Y(g2665),.A(g1661));
  NOT NOT1_760(.VSS(VSS),.VDD(VDD),.Y(g2668),.A(g1662));
  NOT NOT1_761(.VSS(VSS),.VDD(VDD),.Y(I6468),.A(g1917));
  NOT NOT1_762(.VSS(VSS),.VDD(VDD),.Y(g2671),.A(I6468));
  NOT NOT1_763(.VSS(VSS),.VDD(VDD),.Y(I6471),.A(g1923));
  NOT NOT1_764(.VSS(VSS),.VDD(VDD),.Y(g2672),.A(I6471));
  NOT NOT1_765(.VSS(VSS),.VDD(VDD),.Y(I6474),.A(g1941));
  NOT NOT1_766(.VSS(VSS),.VDD(VDD),.Y(g2673),.A(I6474));
  NOT NOT1_767(.VSS(VSS),.VDD(VDD),.Y(g2674),.A(g1675));
  NOT NOT1_768(.VSS(VSS),.VDD(VDD),.Y(g2677),.A(g1664));
  NOT NOT1_769(.VSS(VSS),.VDD(VDD),.Y(g2680),.A(g1665));
  NOT NOT1_770(.VSS(VSS),.VDD(VDD),.Y(g2683),.A(g1666));
  NOT NOT1_771(.VSS(VSS),.VDD(VDD),.Y(g2686),.A(g1667));
  NOT NOT1_772(.VSS(VSS),.VDD(VDD),.Y(g2689),.A(g1670));
  NOT NOT1_773(.VSS(VSS),.VDD(VDD),.Y(g2692),.A(g1671));
  NOT NOT1_774(.VSS(VSS),.VDD(VDD),.Y(g2695),.A(g1672));
  NOT NOT1_775(.VSS(VSS),.VDD(VDD),.Y(g2698),.A(g1673));
  NOT NOT1_776(.VSS(VSS),.VDD(VDD),.Y(g2699),.A(g1674));
  NOT NOT1_777(.VSS(VSS),.VDD(VDD),.Y(g2700),.A(g1744));
  NOT NOT1_778(.VSS(VSS),.VDD(VDD),.Y(g2703),.A(g1809));
  NOT NOT1_779(.VSS(VSS),.VDD(VDD),.Y(g2706),.A(g1821));
  NOT NOT1_780(.VSS(VSS),.VDD(VDD),.Y(g2709),.A(g1747));
  NOT NOT1_781(.VSS(VSS),.VDD(VDD),.Y(g2712),.A(g2039));
  NOT NOT1_782(.VSS(VSS),.VDD(VDD),.Y(g2721),.A(g1803));
  NOT NOT1_783(.VSS(VSS),.VDD(VDD),.Y(g2724),.A(g1814));
  NOT NOT1_784(.VSS(VSS),.VDD(VDD),.Y(g2727),.A(g2424));
  NOT NOT1_785(.VSS(VSS),.VDD(VDD),.Y(g2728),.A(g2256));
  NOT NOT1_786(.VSS(VSS),.VDD(VDD),.Y(g2734),.A(g2170));
  NOT NOT1_787(.VSS(VSS),.VDD(VDD),.Y(g2743),.A(g1808));
  NOT NOT1_788(.VSS(VSS),.VDD(VDD),.Y(g2746),.A(g2259));
  NOT NOT1_789(.VSS(VSS),.VDD(VDD),.Y(g2752),.A(g2389));
  NOT NOT1_790(.VSS(VSS),.VDD(VDD),.Y(g2761),.A(g1820));
  NOT NOT1_791(.VSS(VSS),.VDD(VDD),.Y(g2764),.A(g1802));
  NOT NOT1_792(.VSS(VSS),.VDD(VDD),.Y(I6509),.A(g1684));
  NOT NOT1_793(.VSS(VSS),.VDD(VDD),.Y(g2767),.A(I6509));
  NOT NOT1_794(.VSS(VSS),.VDD(VDD),.Y(g2769),.A(g2424));
  NOT NOT1_795(.VSS(VSS),.VDD(VDD),.Y(g2770),.A(g2210));
  NOT NOT1_796(.VSS(VSS),.VDD(VDD),.Y(g2774),.A(g1813));
  NOT NOT1_797(.VSS(VSS),.VDD(VDD),.Y(g2777),.A(g1797));
  NOT NOT1_798(.VSS(VSS),.VDD(VDD),.Y(I6517),.A(g1687));
  NOT NOT1_799(.VSS(VSS),.VDD(VDD),.Y(g2780),.A(I6517));
  NOT NOT1_800(.VSS(VSS),.VDD(VDD),.Y(g2782),.A(g1616));
  NOT NOT1_801(.VSS(VSS),.VDD(VDD),.Y(g2784),.A(g2340));
  NOT NOT1_802(.VSS(VSS),.VDD(VDD),.Y(g2787),.A(g1807));
  NOT NOT1_803(.VSS(VSS),.VDD(VDD),.Y(g2790),.A(g1793));
  NOT NOT1_804(.VSS(VSS),.VDD(VDD),.Y(I6532),.A(g1694));
  NOT NOT1_805(.VSS(VSS),.VDD(VDD),.Y(g2793),.A(I6532));
  NOT NOT1_806(.VSS(VSS),.VDD(VDD),.Y(g2794),.A(g2185));
  NOT NOT1_807(.VSS(VSS),.VDD(VDD),.Y(g2795),.A(g1801));
  NOT NOT1_808(.VSS(VSS),.VDD(VDD),.Y(g2798),.A(g1787));
  NOT NOT1_809(.VSS(VSS),.VDD(VDD),.Y(g2804),.A(g1796));
  NOT NOT1_810(.VSS(VSS),.VDD(VDD),.Y(g2807),.A(g1782));
  NOT NOT1_811(.VSS(VSS),.VDD(VDD),.Y(g2810),.A(g1922));
  NOT NOT1_812(.VSS(VSS),.VDD(VDD),.Y(g2816),.A(g1685));
  NOT NOT1_813(.VSS(VSS),.VDD(VDD),.Y(g2817),.A(g1849));
  NOT NOT1_814(.VSS(VSS),.VDD(VDD),.Y(g2818),.A(g1792));
  NOT NOT1_815(.VSS(VSS),.VDD(VDD),.Y(g2821),.A(g1786));
  NOT NOT1_816(.VSS(VSS),.VDD(VDD),.Y(g2824),.A(g1688));
  NOT NOT1_817(.VSS(VSS),.VDD(VDD),.Y(I6553),.A(g2246));
  NOT NOT1_818(.VSS(VSS),.VDD(VDD),.Y(g2825),.A(I6553));
  NOT NOT1_819(.VSS(VSS),.VDD(VDD),.Y(g2826),.A(g2183));
  NOT NOT1_820(.VSS(VSS),.VDD(VDD),.Y(g2828),.A(g1980));
  NOT NOT1_821(.VSS(VSS),.VDD(VDD),.Y(g2829),.A(g1785));
  NOT NOT1_822(.VSS(VSS),.VDD(VDD),.Y(g2832),.A(g2184));
  NOT NOT1_823(.VSS(VSS),.VDD(VDD),.Y(I6561),.A(g1715));
  NOT NOT1_824(.VSS(VSS),.VDD(VDD),.Y(g2833),.A(I6561));
  NOT NOT1_825(.VSS(VSS),.VDD(VDD),.Y(I6564),.A(g2073));
  NOT NOT1_826(.VSS(VSS),.VDD(VDD),.Y(g2834),.A(I6564));
  NOT NOT1_827(.VSS(VSS),.VDD(VDD),.Y(g2837),.A(g1780));
  NOT NOT1_828(.VSS(VSS),.VDD(VDD),.Y(g2840),.A(g2207));
  NOT NOT1_829(.VSS(VSS),.VDD(VDD),.Y(g2841),.A(g2208));
  NOT NOT1_830(.VSS(VSS),.VDD(VDD),.Y(g2842),.A(g2209));
  NOT NOT1_831(.VSS(VSS),.VDD(VDD),.Y(I6571),.A(g1711));
  NOT NOT1_832(.VSS(VSS),.VDD(VDD),.Y(g2843),.A(I6571));
  NOT NOT1_833(.VSS(VSS),.VDD(VDD),.Y(I6574),.A(g576));
  NOT NOT1_834(.VSS(VSS),.VDD(VDD),.Y(g2844),.A(I6574));
  NOT NOT1_835(.VSS(VSS),.VDD(VDD),.Y(I6578),.A(g1603));
  NOT NOT1_836(.VSS(VSS),.VDD(VDD),.Y(g2862),.A(I6578));
  NOT NOT1_837(.VSS(VSS),.VDD(VDD),.Y(g2863),.A(g1778));
  NOT NOT1_838(.VSS(VSS),.VDD(VDD),.Y(g2866),.A(g2221));
  NOT NOT1_839(.VSS(VSS),.VDD(VDD),.Y(g2867),.A(g2222));
  NOT NOT1_840(.VSS(VSS),.VDD(VDD),.Y(g2868),.A(g2223));
  NOT NOT1_841(.VSS(VSS),.VDD(VDD),.Y(g2869),.A(g2224));
  NOT NOT1_842(.VSS(VSS),.VDD(VDD),.Y(g2870),.A(g2225));
  NOT NOT1_843(.VSS(VSS),.VDD(VDD),.Y(I6587),.A(g1708));
  NOT NOT1_844(.VSS(VSS),.VDD(VDD),.Y(g2871),.A(I6587));
  NOT NOT1_845(.VSS(VSS),.VDD(VDD),.Y(I6590),.A(g2467));
  NOT NOT1_846(.VSS(VSS),.VDD(VDD),.Y(g2872),.A(I6590));
  NOT NOT1_847(.VSS(VSS),.VDD(VDD),.Y(g2873),.A(g1779));
  NOT NOT1_848(.VSS(VSS),.VDD(VDD),.Y(g2876),.A(g2231));
  NOT NOT1_849(.VSS(VSS),.VDD(VDD),.Y(g2877),.A(g2232));
  NOT NOT1_850(.VSS(VSS),.VDD(VDD),.Y(g2878),.A(g2233));
  NOT NOT1_851(.VSS(VSS),.VDD(VDD),.Y(I6597),.A(g1970));
  NOT NOT1_852(.VSS(VSS),.VDD(VDD),.Y(g2879),.A(I6597));
  NOT NOT1_853(.VSS(VSS),.VDD(VDD),.Y(g2880),.A(g2234));
  NOT NOT1_854(.VSS(VSS),.VDD(VDD),.Y(g2881),.A(g2235));
  NOT NOT1_855(.VSS(VSS),.VDD(VDD),.Y(g2882),.A(g2236));
  NOT NOT1_856(.VSS(VSS),.VDD(VDD),.Y(g2883),.A(g2237));
  NOT NOT1_857(.VSS(VSS),.VDD(VDD),.Y(g2884),.A(g2238));
  NOT NOT1_858(.VSS(VSS),.VDD(VDD),.Y(g2885),.A(g2239));
  NOT NOT1_859(.VSS(VSS),.VDD(VDD),.Y(g2886),.A(g2240));
  NOT NOT1_860(.VSS(VSS),.VDD(VDD),.Y(g2887),.A(g2241));
  NOT NOT1_861(.VSS(VSS),.VDD(VDD),.Y(I6608),.A(g1612));
  NOT NOT1_862(.VSS(VSS),.VDD(VDD),.Y(g2888),.A(I6608));
  NOT NOT1_863(.VSS(VSS),.VDD(VDD),.Y(g2890),.A(g2264));
  NOT NOT1_864(.VSS(VSS),.VDD(VDD),.Y(g2891),.A(g2265));
  NOT NOT1_865(.VSS(VSS),.VDD(VDD),.Y(g2892),.A(g2266));
  NOT NOT1_866(.VSS(VSS),.VDD(VDD),.Y(I6615),.A(g1983));
  NOT NOT1_867(.VSS(VSS),.VDD(VDD),.Y(g2893),.A(I6615));
  NOT NOT1_868(.VSS(VSS),.VDD(VDD),.Y(g2894),.A(g2267));
  NOT NOT1_869(.VSS(VSS),.VDD(VDD),.Y(g2895),.A(g2268));
  NOT NOT1_870(.VSS(VSS),.VDD(VDD),.Y(g2896),.A(g2269));
  NOT NOT1_871(.VSS(VSS),.VDD(VDD),.Y(g2897),.A(g2270));
  NOT NOT1_872(.VSS(VSS),.VDD(VDD),.Y(g2898),.A(g2271));
  NOT NOT1_873(.VSS(VSS),.VDD(VDD),.Y(g2899),.A(g2272));
  NOT NOT1_874(.VSS(VSS),.VDD(VDD),.Y(g2900),.A(g2273));
  NOT NOT1_875(.VSS(VSS),.VDD(VDD),.Y(g2901),.A(g2284));
  NOT NOT1_876(.VSS(VSS),.VDD(VDD),.Y(g2902),.A(g2285));
  NOT NOT1_877(.VSS(VSS),.VDD(VDD),.Y(g2903),.A(g2286));
  NOT NOT1_878(.VSS(VSS),.VDD(VDD),.Y(g2904),.A(g2287));
  NOT NOT1_879(.VSS(VSS),.VDD(VDD),.Y(I6629),.A(g2052));
  NOT NOT1_880(.VSS(VSS),.VDD(VDD),.Y(g2905),.A(I6629));
  NOT NOT1_881(.VSS(VSS),.VDD(VDD),.Y(g2906),.A(g2288));
  NOT NOT1_882(.VSS(VSS),.VDD(VDD),.Y(g2907),.A(g2289));
  NOT NOT1_883(.VSS(VSS),.VDD(VDD),.Y(g2908),.A(g2290));
  NOT NOT1_884(.VSS(VSS),.VDD(VDD),.Y(g2909),.A(g2291));
  NOT NOT1_885(.VSS(VSS),.VDD(VDD),.Y(I6636),.A(g1704));
  NOT NOT1_886(.VSS(VSS),.VDD(VDD),.Y(g2910),.A(I6636));
  NOT NOT1_887(.VSS(VSS),.VDD(VDD),.Y(g2911),.A(g2292));
  NOT NOT1_888(.VSS(VSS),.VDD(VDD),.Y(g2913),.A(g2307));
  NOT NOT1_889(.VSS(VSS),.VDD(VDD),.Y(g2914),.A(g2308));
  NOT NOT1_890(.VSS(VSS),.VDD(VDD),.Y(I6643),.A(g1970));
  NOT NOT1_891(.VSS(VSS),.VDD(VDD),.Y(g2915),.A(I6643));
  NOT NOT1_892(.VSS(VSS),.VDD(VDD),.Y(I6646),.A(g2246));
  NOT NOT1_893(.VSS(VSS),.VDD(VDD),.Y(g2916),.A(I6646));
  NOT NOT1_894(.VSS(VSS),.VDD(VDD),.Y(g2917),.A(g2309));
  NOT NOT1_895(.VSS(VSS),.VDD(VDD),.Y(g2918),.A(g2310));
  NOT NOT1_896(.VSS(VSS),.VDD(VDD),.Y(g2919),.A(g2311));
  NOT NOT1_897(.VSS(VSS),.VDD(VDD),.Y(I6652),.A(g2016));
  NOT NOT1_898(.VSS(VSS),.VDD(VDD),.Y(g2920),.A(I6652));
  NOT NOT1_899(.VSS(VSS),.VDD(VDD),.Y(g2921),.A(g2312));
  NOT NOT1_900(.VSS(VSS),.VDD(VDD),.Y(g2922),.A(g2313));
  NOT NOT1_901(.VSS(VSS),.VDD(VDD),.Y(I6657),.A(g1701));
  NOT NOT1_902(.VSS(VSS),.VDD(VDD),.Y(g2923),.A(I6657));
  NOT NOT1_903(.VSS(VSS),.VDD(VDD),.Y(g2924),.A(g2314));
  NOT NOT1_904(.VSS(VSS),.VDD(VDD),.Y(g2925),.A(g2324));
  NOT NOT1_905(.VSS(VSS),.VDD(VDD),.Y(g2926),.A(g2325));
  NOT NOT1_906(.VSS(VSS),.VDD(VDD),.Y(I6663),.A(g2246));
  NOT NOT1_907(.VSS(VSS),.VDD(VDD),.Y(g2927),.A(I6663));
  NOT NOT1_908(.VSS(VSS),.VDD(VDD),.Y(g2928),.A(g2326));
  NOT NOT1_909(.VSS(VSS),.VDD(VDD),.Y(g2929),.A(g2327));
  NOT NOT1_910(.VSS(VSS),.VDD(VDD),.Y(g2930),.A(g2328));
  NOT NOT1_911(.VSS(VSS),.VDD(VDD),.Y(I6669),.A(g1698));
  NOT NOT1_912(.VSS(VSS),.VDD(VDD),.Y(g2931),.A(I6669));
  NOT NOT1_913(.VSS(VSS),.VDD(VDD),.Y(g2932),.A(g2329));
  NOT NOT1_914(.VSS(VSS),.VDD(VDD),.Y(I6673),.A(g2246));
  NOT NOT1_915(.VSS(VSS),.VDD(VDD),.Y(g2933),.A(I6673));
  NOT NOT1_916(.VSS(VSS),.VDD(VDD),.Y(I6676),.A(g1603));
  NOT NOT1_917(.VSS(VSS),.VDD(VDD),.Y(g2934),.A(I6676));
  NOT NOT1_918(.VSS(VSS),.VDD(VDD),.Y(I6680),.A(g1558));
  NOT NOT1_919(.VSS(VSS),.VDD(VDD),.Y(g2936),.A(I6680));
  NOT NOT1_920(.VSS(VSS),.VDD(VDD),.Y(g2937),.A(g2346));
  NOT NOT1_921(.VSS(VSS),.VDD(VDD),.Y(g2938),.A(g2347));
  NOT NOT1_922(.VSS(VSS),.VDD(VDD),.Y(g2939),.A(g2348));
  NOT NOT1_923(.VSS(VSS),.VDD(VDD),.Y(I6686),.A(g2246));
  NOT NOT1_924(.VSS(VSS),.VDD(VDD),.Y(g2940),.A(I6686));
  NOT NOT1_925(.VSS(VSS),.VDD(VDD),.Y(g2941),.A(g2349));
  NOT NOT1_926(.VSS(VSS),.VDD(VDD),.Y(g2942),.A(g2350));
  NOT NOT1_927(.VSS(VSS),.VDD(VDD),.Y(g2943),.A(g2362));
  NOT NOT1_928(.VSS(VSS),.VDD(VDD),.Y(g2944),.A(g2363));
  NOT NOT1_929(.VSS(VSS),.VDD(VDD),.Y(g2945),.A(g2364));
  NOT NOT1_930(.VSS(VSS),.VDD(VDD),.Y(g2946),.A(g2365));
  NOT NOT1_931(.VSS(VSS),.VDD(VDD),.Y(I6695),.A(g2246));
  NOT NOT1_932(.VSS(VSS),.VDD(VDD),.Y(g2947),.A(I6695));
  NOT NOT1_933(.VSS(VSS),.VDD(VDD),.Y(g2948),.A(g2366));
  NOT NOT1_934(.VSS(VSS),.VDD(VDD),.Y(g2953),.A(g2373));
  NOT NOT1_935(.VSS(VSS),.VDD(VDD),.Y(g2954),.A(g2374));
  NOT NOT1_936(.VSS(VSS),.VDD(VDD),.Y(I6703),.A(g1983));
  NOT NOT1_937(.VSS(VSS),.VDD(VDD),.Y(g2955),.A(I6703));
  NOT NOT1_938(.VSS(VSS),.VDD(VDD),.Y(g2956),.A(g2375));
  NOT NOT1_939(.VSS(VSS),.VDD(VDD),.Y(g2957),.A(g2376));
  NOT NOT1_940(.VSS(VSS),.VDD(VDD),.Y(g2958),.A(g2377));
  NOT NOT1_941(.VSS(VSS),.VDD(VDD),.Y(g2959),.A(g1926));
  NOT NOT1_942(.VSS(VSS),.VDD(VDD),.Y(g2960),.A(g2381));
  NOT NOT1_943(.VSS(VSS),.VDD(VDD),.Y(I6711),.A(g1726));
  NOT NOT1_944(.VSS(VSS),.VDD(VDD),.Y(g2961),.A(I6711));
  NOT NOT1_945(.VSS(VSS),.VDD(VDD),.Y(g2962),.A(g2382));
  NOT NOT1_946(.VSS(VSS),.VDD(VDD),.Y(g2963),.A(g2383));
  NOT NOT1_947(.VSS(VSS),.VDD(VDD),.Y(I6716),.A(g1721));
  NOT NOT1_948(.VSS(VSS),.VDD(VDD),.Y(g2964),.A(I6716));
  NOT NOT1_949(.VSS(VSS),.VDD(VDD),.Y(g2965),.A(g2384));
  NOT NOT1_950(.VSS(VSS),.VDD(VDD),.Y(g2966),.A(g1856));
  NOT NOT1_951(.VSS(VSS),.VDD(VDD),.Y(g2969),.A(g2393));
  NOT NOT1_952(.VSS(VSS),.VDD(VDD),.Y(g2970),.A(g2394));
  NOT NOT1_953(.VSS(VSS),.VDD(VDD),.Y(I6723),.A(g2052));
  NOT NOT1_954(.VSS(VSS),.VDD(VDD),.Y(g2971),.A(I6723));
  NOT NOT1_955(.VSS(VSS),.VDD(VDD),.Y(g2973),.A(g1854));
  NOT NOT1_956(.VSS(VSS),.VDD(VDD),.Y(I6728),.A(g1959));
  NOT NOT1_957(.VSS(VSS),.VDD(VDD),.Y(g2976),.A(I6728));
  NOT NOT1_958(.VSS(VSS),.VDD(VDD),.Y(g2982),.A(g1848));
  NOT NOT1_959(.VSS(VSS),.VDD(VDD),.Y(I6733),.A(g1718));
  NOT NOT1_960(.VSS(VSS),.VDD(VDD),.Y(g2985),.A(I6733));
  NOT NOT1_961(.VSS(VSS),.VDD(VDD),.Y(g2989),.A(g1843));
  NOT NOT1_962(.VSS(VSS),.VDD(VDD),.Y(g2992),.A(g1833));
  NOT NOT1_963(.VSS(VSS),.VDD(VDD),.Y(g2996),.A(g1828));
  NOT NOT1_964(.VSS(VSS),.VDD(VDD),.Y(g2999),.A(g1823));
  NOT NOT1_965(.VSS(VSS),.VDD(VDD),.Y(g3008),.A(g1816));
  NOT NOT1_966(.VSS(VSS),.VDD(VDD),.Y(I6764),.A(g1955));
  NOT NOT1_967(.VSS(VSS),.VDD(VDD),.Y(g3013),.A(I6764));
  NOT NOT1_968(.VSS(VSS),.VDD(VDD),.Y(I6767),.A(g1933));
  NOT NOT1_969(.VSS(VSS),.VDD(VDD),.Y(g3014),.A(I6767));
  NOT NOT1_970(.VSS(VSS),.VDD(VDD),.Y(I6770),.A(g1590));
  NOT NOT1_971(.VSS(VSS),.VDD(VDD),.Y(g3018),.A(I6770));
  NOT NOT1_972(.VSS(VSS),.VDD(VDD),.Y(g3019),.A(g2007));
  NOT NOT1_973(.VSS(VSS),.VDD(VDD),.Y(g3029),.A(g1929));
  NOT NOT1_974(.VSS(VSS),.VDD(VDD),.Y(g3038),.A(g2092));
  NOT NOT1_975(.VSS(VSS),.VDD(VDD),.Y(g3047),.A(g1736));
  NOT NOT1_976(.VSS(VSS),.VDD(VDD),.Y(I6784),.A(g2052));
  NOT NOT1_977(.VSS(VSS),.VDD(VDD),.Y(g3048),.A(I6784));
  NOT NOT1_978(.VSS(VSS),.VDD(VDD),.Y(I6788),.A(g1681));
  NOT NOT1_979(.VSS(VSS),.VDD(VDD),.Y(g3050),.A(I6788));
  NOT NOT1_980(.VSS(VSS),.VDD(VDD),.Y(I6791),.A(g1967));
  NOT NOT1_981(.VSS(VSS),.VDD(VDD),.Y(g3051),.A(I6791));
  NOT NOT1_982(.VSS(VSS),.VDD(VDD),.Y(g3052),.A(g2096));
  NOT NOT1_983(.VSS(VSS),.VDD(VDD),.Y(I6795),.A(g1683));
  NOT NOT1_984(.VSS(VSS),.VDD(VDD),.Y(g3061),.A(I6795));
  NOT NOT1_985(.VSS(VSS),.VDD(VDD),.Y(g3062),.A(g2100));
  NOT NOT1_986(.VSS(VSS),.VDD(VDD),.Y(g3071),.A(g1948));
  NOT NOT1_987(.VSS(VSS),.VDD(VDD),.Y(I6800),.A(g2016));
  NOT NOT1_988(.VSS(VSS),.VDD(VDD),.Y(g3074),.A(I6800));
  NOT NOT1_989(.VSS(VSS),.VDD(VDD),.Y(g3075),.A(g2216));
  NOT NOT1_990(.VSS(VSS),.VDD(VDD),.Y(g3076),.A(g1831));
  NOT NOT1_991(.VSS(VSS),.VDD(VDD),.Y(I6805),.A(g1603));
  NOT NOT1_992(.VSS(VSS),.VDD(VDD),.Y(g3077),.A(I6805));
  NOT NOT1_993(.VSS(VSS),.VDD(VDD),.Y(g3078),.A(g1603));
  NOT NOT1_994(.VSS(VSS),.VDD(VDD),.Y(g3079),.A(g1603));
  NOT NOT1_995(.VSS(VSS),.VDD(VDD),.Y(g3080),.A(g1679));
  NOT NOT1_996(.VSS(VSS),.VDD(VDD),.Y(g3082),.A(g1680));
  NOT NOT1_997(.VSS(VSS),.VDD(VDD),.Y(I6820),.A(g1707));
  NOT NOT1_998(.VSS(VSS),.VDD(VDD),.Y(g3084),.A(I6820));
  NOT NOT1_999(.VSS(VSS),.VDD(VDD),.Y(g3085),.A(g1945));
  NOT NOT1_1000(.VSS(VSS),.VDD(VDD),.Y(g3086),.A(g1852));
  NOT NOT1_1001(.VSS(VSS),.VDD(VDD),.Y(g3091),.A(g1603));
  NOT NOT1_1002(.VSS(VSS),.VDD(VDD),.Y(I6826),.A(g2185));
  NOT NOT1_1003(.VSS(VSS),.VDD(VDD),.Y(g3092),.A(I6826));
  NOT NOT1_1004(.VSS(VSS),.VDD(VDD),.Y(g3093),.A(g1686));
  NOT NOT1_1005(.VSS(VSS),.VDD(VDD),.Y(I6831),.A(g2185));
  NOT NOT1_1006(.VSS(VSS),.VDD(VDD),.Y(g3095),.A(I6831));
  NOT NOT1_1007(.VSS(VSS),.VDD(VDD),.Y(I6834),.A(g287));
  NOT NOT1_1008(.VSS(VSS),.VDD(VDD),.Y(g3096),.A(I6834));
  NOT NOT1_1009(.VSS(VSS),.VDD(VDD),.Y(g3124),.A(g1857));
  NOT NOT1_1010(.VSS(VSS),.VDD(VDD),.Y(I6839),.A(g2185));
  NOT NOT1_1011(.VSS(VSS),.VDD(VDD),.Y(g3128),.A(I6839));
  NOT NOT1_1012(.VSS(VSS),.VDD(VDD),.Y(I6849),.A(g368));
  NOT NOT1_1013(.VSS(VSS),.VDD(VDD),.Y(g3130),.A(I6849));
  NOT NOT1_1014(.VSS(VSS),.VDD(VDD),.Y(I6853),.A(g2185));
  NOT NOT1_1015(.VSS(VSS),.VDD(VDD),.Y(g3158),.A(I6853));
  NOT NOT1_1016(.VSS(VSS),.VDD(VDD),.Y(I6856),.A(g449));
  NOT NOT1_1017(.VSS(VSS),.VDD(VDD),.Y(g3159),.A(I6856));
  NOT NOT1_1018(.VSS(VSS),.VDD(VDD),.Y(I6860),.A(g2185));
  NOT NOT1_1019(.VSS(VSS),.VDD(VDD),.Y(g3187),.A(I6860));
  NOT NOT1_1020(.VSS(VSS),.VDD(VDD),.Y(I6864),.A(g2528));
  NOT NOT1_1021(.VSS(VSS),.VDD(VDD),.Y(g3189),.A(I6864));
  NOT NOT1_1022(.VSS(VSS),.VDD(VDD),.Y(I6868),.A(g530));
  NOT NOT1_1023(.VSS(VSS),.VDD(VDD),.Y(g3191),.A(I6868));
  NOT NOT1_1024(.VSS(VSS),.VDD(VDD),.Y(I6872),.A(g2185));
  NOT NOT1_1025(.VSS(VSS),.VDD(VDD),.Y(g3219),.A(I6872));
  NOT NOT1_1026(.VSS(VSS),.VDD(VDD),.Y(g3220),.A(g1889));
  NOT NOT1_1027(.VSS(VSS),.VDD(VDD),.Y(I6887),.A(g2528));
  NOT NOT1_1028(.VSS(VSS),.VDD(VDD),.Y(g3230),.A(I6887));
  NOT NOT1_1029(.VSS(VSS),.VDD(VDD),.Y(I6894),.A(g1863));
  NOT NOT1_1030(.VSS(VSS),.VDD(VDD),.Y(g3238),.A(I6894));
  NOT NOT1_1031(.VSS(VSS),.VDD(VDD),.Y(I6900),.A(g1866));
  NOT NOT1_1032(.VSS(VSS),.VDD(VDD),.Y(g3264),.A(I6900));
  NOT NOT1_1033(.VSS(VSS),.VDD(VDD),.Y(g3285),.A(g1689));
  NOT NOT1_1034(.VSS(VSS),.VDD(VDD),.Y(I6911),.A(g1869));
  NOT NOT1_1035(.VSS(VSS),.VDD(VDD),.Y(g3287),.A(I6911));
  NOT NOT1_1036(.VSS(VSS),.VDD(VDD),.Y(I6930),.A(g1876));
  NOT NOT1_1037(.VSS(VSS),.VDD(VDD),.Y(g3316),.A(I6930));
  NOT NOT1_1038(.VSS(VSS),.VDD(VDD),.Y(g3338),.A(g1901));
  NOT NOT1_1039(.VSS(VSS),.VDD(VDD),.Y(g3340),.A(g2474));
  NOT NOT1_1040(.VSS(VSS),.VDD(VDD),.Y(I6936),.A(g1878));
  NOT NOT1_1041(.VSS(VSS),.VDD(VDD),.Y(g3341),.A(I6936));
  NOT NOT1_1042(.VSS(VSS),.VDD(VDD),.Y(I6946),.A(g1887));
  NOT NOT1_1043(.VSS(VSS),.VDD(VDD),.Y(g3359),.A(I6946));
  NOT NOT1_1044(.VSS(VSS),.VDD(VDD),.Y(I6949),.A(g2148));
  NOT NOT1_1045(.VSS(VSS),.VDD(VDD),.Y(g3390),.A(I6949));
  NOT NOT1_1046(.VSS(VSS),.VDD(VDD),.Y(I6952),.A(g1896));
  NOT NOT1_1047(.VSS(VSS),.VDD(VDD),.Y(g3398),.A(I6952));
  NOT NOT1_1048(.VSS(VSS),.VDD(VDD),.Y(I6956),.A(g1907));
  NOT NOT1_1049(.VSS(VSS),.VDD(VDD),.Y(g3430),.A(I6956));
  NOT NOT1_1050(.VSS(VSS),.VDD(VDD),.Y(I6959),.A(g1558));
  NOT NOT1_1051(.VSS(VSS),.VDD(VDD),.Y(g3461),.A(I6959));
  NOT NOT1_1052(.VSS(VSS),.VDD(VDD),.Y(g3462),.A(g1743));
  NOT NOT1_1053(.VSS(VSS),.VDD(VDD),.Y(I6963),.A(g1558));
  NOT NOT1_1054(.VSS(VSS),.VDD(VDD),.Y(g3465),.A(I6963));
  NOT NOT1_1055(.VSS(VSS),.VDD(VDD),.Y(g3485),.A(g1737));
  NOT NOT1_1056(.VSS(VSS),.VDD(VDD),.Y(g3488),.A(g1727));
  NOT NOT1_1057(.VSS(VSS),.VDD(VDD),.Y(g3491),.A(g1800));
  NOT NOT1_1058(.VSS(VSS),.VDD(VDD),.Y(I6970),.A(g1872));
  NOT NOT1_1059(.VSS(VSS),.VDD(VDD),.Y(g3492),.A(I6970));
  NOT NOT1_1060(.VSS(VSS),.VDD(VDD),.Y(g3495),.A(g1616));
  NOT NOT1_1061(.VSS(VSS),.VDD(VDD),.Y(I6974),.A(g2528));
  NOT NOT1_1062(.VSS(VSS),.VDD(VDD),.Y(g3496),.A(I6974));
  NOT NOT1_1063(.VSS(VSS),.VDD(VDD),.Y(g3497),.A(g2185));
  NOT NOT1_1064(.VSS(VSS),.VDD(VDD),.Y(g3498),.A(g1616));
  NOT NOT1_1065(.VSS(VSS),.VDD(VDD),.Y(g3499),.A(g2185));
  NOT NOT1_1066(.VSS(VSS),.VDD(VDD),.Y(g3500),.A(g1616));
  NOT NOT1_1067(.VSS(VSS),.VDD(VDD),.Y(g3501),.A(g2185));
  NOT NOT1_1068(.VSS(VSS),.VDD(VDD),.Y(g3502),.A(g1616));
  NOT NOT1_1069(.VSS(VSS),.VDD(VDD),.Y(g3503),.A(g2407));
  NOT NOT1_1070(.VSS(VSS),.VDD(VDD),.Y(g3506),.A(g1781));
  NOT NOT1_1071(.VSS(VSS),.VDD(VDD),.Y(g3510),.A(g2185));
  NOT NOT1_1072(.VSS(VSS),.VDD(VDD),.Y(g3511),.A(g1616));
  NOT NOT1_1073(.VSS(VSS),.VDD(VDD),.Y(g3512),.A(g1616));
  NOT NOT1_1074(.VSS(VSS),.VDD(VDD),.Y(g3513),.A(g2407));
  NOT NOT1_1075(.VSS(VSS),.VDD(VDD),.Y(g3514),.A(g2424));
  NOT NOT1_1076(.VSS(VSS),.VDD(VDD),.Y(g3517),.A(g2283));
  NOT NOT1_1077(.VSS(VSS),.VDD(VDD),.Y(g3519),.A(g2185));
  NOT NOT1_1078(.VSS(VSS),.VDD(VDD),.Y(g3520),.A(g1616));
  NOT NOT1_1079(.VSS(VSS),.VDD(VDD),.Y(g3521),.A(g2185));
  NOT NOT1_1080(.VSS(VSS),.VDD(VDD),.Y(g3522),.A(g2407));
  NOT NOT1_1081(.VSS(VSS),.VDD(VDD),.Y(g3523),.A(g2407));
  NOT NOT1_1082(.VSS(VSS),.VDD(VDD),.Y(g3524),.A(g2306));
  NOT NOT1_1083(.VSS(VSS),.VDD(VDD),.Y(g3526),.A(g2185));
  NOT NOT1_1084(.VSS(VSS),.VDD(VDD),.Y(g3527),.A(g1616));
  NOT NOT1_1085(.VSS(VSS),.VDD(VDD),.Y(g3529),.A(g2323));
  NOT NOT1_1086(.VSS(VSS),.VDD(VDD),.Y(g3530),.A(g2185));
  NOT NOT1_1087(.VSS(VSS),.VDD(VDD),.Y(g3531),.A(g1616));
  NOT NOT1_1088(.VSS(VSS),.VDD(VDD),.Y(g3532),.A(g2407));
  NOT NOT1_1089(.VSS(VSS),.VDD(VDD),.Y(g3533),.A(g2397));
  NOT NOT1_1090(.VSS(VSS),.VDD(VDD),.Y(g3539),.A(g2424));
  NOT NOT1_1091(.VSS(VSS),.VDD(VDD),.Y(g3540),.A(g2424));
  NOT NOT1_1092(.VSS(VSS),.VDD(VDD),.Y(g3542),.A(g1777));
  NOT NOT1_1093(.VSS(VSS),.VDD(VDD),.Y(g3545),.A(g2344));
  NOT NOT1_1094(.VSS(VSS),.VDD(VDD),.Y(I7029),.A(g2392));
  NOT NOT1_1095(.VSS(VSS),.VDD(VDD),.Y(g3546),.A(I7029));
  NOT NOT1_1096(.VSS(VSS),.VDD(VDD),.Y(g3547),.A(g2345));
  NOT NOT1_1097(.VSS(VSS),.VDD(VDD),.Y(g3548),.A(g2185));
  NOT NOT1_1098(.VSS(VSS),.VDD(VDD),.Y(g3549),.A(g2404));
  NOT NOT1_1099(.VSS(VSS),.VDD(VDD),.Y(I7036),.A(g2454));
  NOT NOT1_1100(.VSS(VSS),.VDD(VDD),.Y(g3556),.A(I7036));
  NOT NOT1_1101(.VSS(VSS),.VDD(VDD),.Y(g3557),.A(g1773));
  NOT NOT1_1102(.VSS(VSS),.VDD(VDD),.Y(g3560),.A(g2361));
  NOT NOT1_1103(.VSS(VSS),.VDD(VDD),.Y(I7041),.A(g2401));
  NOT NOT1_1104(.VSS(VSS),.VDD(VDD),.Y(g3561),.A(I7041));
  NOT NOT1_1105(.VSS(VSS),.VDD(VDD),.Y(I7044),.A(g2402));
  NOT NOT1_1106(.VSS(VSS),.VDD(VDD),.Y(g3562),.A(I7044));
  NOT NOT1_1107(.VSS(VSS),.VDD(VDD),.Y(g3563),.A(g2007));
  NOT NOT1_1108(.VSS(VSS),.VDD(VDD),.Y(g3567),.A(g2407));
  NOT NOT1_1109(.VSS(VSS),.VDD(VDD),.Y(g3568),.A(g1935));
  NOT NOT1_1110(.VSS(VSS),.VDD(VDD),.Y(g3573),.A(g2424));
  NOT NOT1_1111(.VSS(VSS),.VDD(VDD),.Y(g3574),.A(g1771));
  NOT NOT1_1112(.VSS(VSS),.VDD(VDD),.Y(g3577),.A(g2372));
  NOT NOT1_1113(.VSS(VSS),.VDD(VDD),.Y(I7053),.A(g2452));
  NOT NOT1_1114(.VSS(VSS),.VDD(VDD),.Y(g3578),.A(I7053));
  NOT NOT1_1115(.VSS(VSS),.VDD(VDD),.Y(g3579),.A(g1929));
  NOT NOT1_1116(.VSS(VSS),.VDD(VDD),.Y(g3582),.A(g2407));
  NOT NOT1_1117(.VSS(VSS),.VDD(VDD),.Y(g3583),.A(g2128));
  NOT NOT1_1118(.VSS(VSS),.VDD(VDD),.Y(g3587),.A(g1964));
  NOT NOT1_1119(.VSS(VSS),.VDD(VDD),.Y(g3588),.A(g2379));
  NOT NOT1_1120(.VSS(VSS),.VDD(VDD),.Y(I7061),.A(g2457));
  NOT NOT1_1121(.VSS(VSS),.VDD(VDD),.Y(g3589),.A(I7061));
  NOT NOT1_1122(.VSS(VSS),.VDD(VDD),.Y(I7064),.A(g2458));
  NOT NOT1_1123(.VSS(VSS),.VDD(VDD),.Y(g3590),.A(I7064));
  NOT NOT1_1124(.VSS(VSS),.VDD(VDD),.Y(g3591),.A(g1789));
  NOT NOT1_1125(.VSS(VSS),.VDD(VDD),.Y(g3603),.A(g2092));
  NOT NOT1_1126(.VSS(VSS),.VDD(VDD),.Y(g3604),.A(g2407));
  NOT NOT1_1127(.VSS(VSS),.VDD(VDD),.Y(g3605),.A(g1938));
  NOT NOT1_1128(.VSS(VSS),.VDD(VDD),.Y(g3610),.A(g2424));
  NOT NOT1_1129(.VSS(VSS),.VDD(VDD),.Y(I7079),.A(g2532));
  NOT NOT1_1130(.VSS(VSS),.VDD(VDD),.Y(g3611),.A(I7079));
  NOT NOT1_1131(.VSS(VSS),.VDD(VDD),.Y(I7082),.A(g2470));
  NOT NOT1_1132(.VSS(VSS),.VDD(VDD),.Y(g3612),.A(I7082));
  NOT NOT1_1133(.VSS(VSS),.VDD(VDD),.Y(g3617),.A(g1655));
  NOT NOT1_1134(.VSS(VSS),.VDD(VDD),.Y(g3629),.A(g2424));
  NOT NOT1_1135(.VSS(VSS),.VDD(VDD),.Y(I7095),.A(g2539));
  NOT NOT1_1136(.VSS(VSS),.VDD(VDD),.Y(g3630),.A(I7095));
  NOT NOT1_1137(.VSS(VSS),.VDD(VDD),.Y(I7098),.A(g2477));
  NOT NOT1_1138(.VSS(VSS),.VDD(VDD),.Y(g3631),.A(I7098));
  NOT NOT1_1139(.VSS(VSS),.VDD(VDD),.Y(I7101),.A(g2478));
  NOT NOT1_1140(.VSS(VSS),.VDD(VDD),.Y(g3632),.A(I7101));
  NOT NOT1_1141(.VSS(VSS),.VDD(VDD),.Y(I7104),.A(g2479));
  NOT NOT1_1142(.VSS(VSS),.VDD(VDD),.Y(g3633),.A(I7104));
  NOT NOT1_1143(.VSS(VSS),.VDD(VDD),.Y(I7107),.A(g2480));
  NOT NOT1_1144(.VSS(VSS),.VDD(VDD),.Y(g3634),.A(I7107));
  NOT NOT1_1145(.VSS(VSS),.VDD(VDD),.Y(g3635),.A(g1949));
  NOT NOT1_1146(.VSS(VSS),.VDD(VDD),.Y(g3639),.A(g2424));
  NOT NOT1_1147(.VSS(VSS),.VDD(VDD),.Y(I7112),.A(g2546));
  NOT NOT1_1148(.VSS(VSS),.VDD(VDD),.Y(g3640),.A(I7112));
  NOT NOT1_1149(.VSS(VSS),.VDD(VDD),.Y(I7115),.A(g2547));
  NOT NOT1_1150(.VSS(VSS),.VDD(VDD),.Y(g3641),.A(I7115));
  NOT NOT1_1151(.VSS(VSS),.VDD(VDD),.Y(I7118),.A(g2484));
  NOT NOT1_1152(.VSS(VSS),.VDD(VDD),.Y(g3642),.A(I7118));
  NOT NOT1_1153(.VSS(VSS),.VDD(VDD),.Y(g3643),.A(g2453));
  NOT NOT1_1154(.VSS(VSS),.VDD(VDD),.Y(g3644),.A(g2131));
  NOT NOT1_1155(.VSS(VSS),.VDD(VDD),.Y(g3647),.A(g2424));
  NOT NOT1_1156(.VSS(VSS),.VDD(VDD),.Y(g3648),.A(g2424));
  NOT NOT1_1157(.VSS(VSS),.VDD(VDD),.Y(g3649),.A(g2424));
  NOT NOT1_1158(.VSS(VSS),.VDD(VDD),.Y(I7126),.A(g2494));
  NOT NOT1_1159(.VSS(VSS),.VDD(VDD),.Y(g3650),.A(I7126));
  NOT NOT1_1160(.VSS(VSS),.VDD(VDD),.Y(I7129),.A(g2495));
  NOT NOT1_1161(.VSS(VSS),.VDD(VDD),.Y(g3651),.A(I7129));
  NOT NOT1_1162(.VSS(VSS),.VDD(VDD),.Y(I7132),.A(g2554));
  NOT NOT1_1163(.VSS(VSS),.VDD(VDD),.Y(g3652),.A(I7132));
  NOT NOT1_1164(.VSS(VSS),.VDD(VDD),.Y(g3653),.A(g2459));
  NOT NOT1_1165(.VSS(VSS),.VDD(VDD),.Y(g3654),.A(g2521));
  NOT NOT1_1166(.VSS(VSS),.VDD(VDD),.Y(g3655),.A(g1844));
  NOT NOT1_1167(.VSS(VSS),.VDD(VDD),.Y(I7145),.A(g2501));
  NOT NOT1_1168(.VSS(VSS),.VDD(VDD),.Y(g3657),.A(I7145));
  NOT NOT1_1169(.VSS(VSS),.VDD(VDD),.Y(g3659),.A(g2293));
  NOT NOT1_1170(.VSS(VSS),.VDD(VDD),.Y(g3666),.A(g2134));
  NOT NOT1_1171(.VSS(VSS),.VDD(VDD),.Y(I7164),.A(g2157));
  NOT NOT1_1172(.VSS(VSS),.VDD(VDD),.Y(g3674),.A(I7164));
  NOT NOT1_1173(.VSS(VSS),.VDD(VDD),.Y(I7167),.A(g2505));
  NOT NOT1_1174(.VSS(VSS),.VDD(VDD),.Y(g3675),.A(I7167));
  NOT NOT1_1175(.VSS(VSS),.VDD(VDD),.Y(g3676),.A(g2380));
  NOT NOT1_1176(.VSS(VSS),.VDD(VDD),.Y(g3677),.A(g2485));
  NOT NOT1_1177(.VSS(VSS),.VDD(VDD),.Y(g3684),.A(g2180));
  NOT NOT1_1178(.VSS(VSS),.VDD(VDD),.Y(I7195),.A(g1795));
  NOT NOT1_1179(.VSS(VSS),.VDD(VDD),.Y(g3691),.A(I7195));
  NOT NOT1_1180(.VSS(VSS),.VDD(VDD),.Y(I7198),.A(g2509));
  NOT NOT1_1181(.VSS(VSS),.VDD(VDD),.Y(g3692),.A(I7198));
  NOT NOT1_1182(.VSS(VSS),.VDD(VDD),.Y(g3693),.A(g2424));
  NOT NOT1_1183(.VSS(VSS),.VDD(VDD),.Y(g3694),.A(g2174));
  NOT NOT1_1184(.VSS(VSS),.VDD(VDD),.Y(g3700),.A(g2514));
  NOT NOT1_1185(.VSS(VSS),.VDD(VDD),.Y(I7204),.A(g2520));
  NOT NOT1_1186(.VSS(VSS),.VDD(VDD),.Y(g3705),.A(I7204));
  NOT NOT1_1187(.VSS(VSS),.VDD(VDD),.Y(g3707),.A(g2226));
  NOT NOT1_1188(.VSS(VSS),.VDD(VDD),.Y(g3712),.A(g1952));
  NOT NOT1_1189(.VSS(VSS),.VDD(VDD),.Y(g3716),.A(g2522));
  NOT NOT1_1190(.VSS(VSS),.VDD(VDD),.Y(I7211),.A(g1742));
  NOT NOT1_1191(.VSS(VSS),.VDD(VDD),.Y(g3721),.A(I7211));
  NOT NOT1_1192(.VSS(VSS),.VDD(VDD),.Y(g3723),.A(g2096));
  NOT NOT1_1193(.VSS(VSS),.VDD(VDD),.Y(g3728),.A(g2202));
  NOT NOT1_1194(.VSS(VSS),.VDD(VDD),.Y(g3732),.A(g2533));
  NOT NOT1_1195(.VSS(VSS),.VDD(VDD),.Y(g3735),.A(g1961));
  NOT NOT1_1196(.VSS(VSS),.VDD(VDD),.Y(g3739),.A(g2536));
  NOT NOT1_1197(.VSS(VSS),.VDD(VDD),.Y(g3743),.A(g1776));
  NOT NOT1_1198(.VSS(VSS),.VDD(VDD),.Y(g3746),.A(g2100));
  NOT NOT1_1199(.VSS(VSS),.VDD(VDD),.Y(g3750),.A(g2177));
  NOT NOT1_1200(.VSS(VSS),.VDD(VDD),.Y(g3753),.A(g2540));
  NOT NOT1_1201(.VSS(VSS),.VDD(VDD),.Y(g3754),.A(g2543));
  NOT NOT1_1202(.VSS(VSS),.VDD(VDD),.Y(g3757),.A(g1977));
  NOT NOT1_1203(.VSS(VSS),.VDD(VDD),.Y(g3761),.A(g1772));
  NOT NOT1_1204(.VSS(VSS),.VDD(VDD),.Y(g3764),.A(g2039));
  NOT NOT1_1205(.VSS(VSS),.VDD(VDD),.Y(g3768),.A(g2253));
  NOT NOT1_1206(.VSS(VSS),.VDD(VDD),.Y(g3769),.A(g2548));
  NOT NOT1_1207(.VSS(VSS),.VDD(VDD),.Y(g3770),.A(g2551));
  NOT NOT1_1208(.VSS(VSS),.VDD(VDD),.Y(g3771),.A(g1853));
  NOT NOT1_1209(.VSS(VSS),.VDD(VDD),.Y(g3774),.A(g1770));
  NOT NOT1_1210(.VSS(VSS),.VDD(VDD),.Y(g3777),.A(g2170));
  NOT NOT1_1211(.VSS(VSS),.VDD(VDD),.Y(g3778),.A(g2145));
  NOT NOT1_1212(.VSS(VSS),.VDD(VDD),.Y(g3779),.A(g2511));
  NOT NOT1_1213(.VSS(VSS),.VDD(VDD),.Y(g3780),.A(g1847));
  NOT NOT1_1214(.VSS(VSS),.VDD(VDD),.Y(I7255),.A(g1955));
  NOT NOT1_1215(.VSS(VSS),.VDD(VDD),.Y(g3783),.A(I7255));
  NOT NOT1_1216(.VSS(VSS),.VDD(VDD),.Y(g3784),.A(g1768));
  NOT NOT1_1217(.VSS(VSS),.VDD(VDD),.Y(g3787),.A(g1842));
  NOT NOT1_1218(.VSS(VSS),.VDD(VDD),.Y(g3798),.A(g1757));
  NOT NOT1_1219(.VSS(VSS),.VDD(VDD),.Y(I7262),.A(g2514));
  NOT NOT1_1220(.VSS(VSS),.VDD(VDD),.Y(g3801),.A(I7262));
  NOT NOT1_1221(.VSS(VSS),.VDD(VDD),.Y(g3802),.A(g1832));
  NOT NOT1_1222(.VSS(VSS),.VDD(VDD),.Y(g3805),.A(g1752));
  NOT NOT1_1223(.VSS(VSS),.VDD(VDD),.Y(g3808),.A(g1827));
  NOT NOT1_1224(.VSS(VSS),.VDD(VDD),.Y(g3812),.A(g1750));
  NOT NOT1_1225(.VSS(VSS),.VDD(VDD),.Y(g3815),.A(g1822));
  NOT NOT1_1226(.VSS(VSS),.VDD(VDD),.Y(g3819),.A(g1748));
  NOT NOT1_1227(.VSS(VSS),.VDD(VDD),.Y(g3822),.A(g1815));
  NOT NOT1_1228(.VSS(VSS),.VDD(VDD),.Y(g3825),.A(g1826));
  NOT NOT1_1229(.VSS(VSS),.VDD(VDD),.Y(I7287),.A(g2561));
  NOT NOT1_1230(.VSS(VSS),.VDD(VDD),.Y(g3828),.A(I7287));
  NOT NOT1_1231(.VSS(VSS),.VDD(VDD),.Y(I7290),.A(g2936));
  NOT NOT1_1232(.VSS(VSS),.VDD(VDD),.Y(g3829),.A(I7290));
  NOT NOT1_1233(.VSS(VSS),.VDD(VDD),.Y(I7293),.A(g2955));
  NOT NOT1_1234(.VSS(VSS),.VDD(VDD),.Y(g3830),.A(I7293));
  NOT NOT1_1235(.VSS(VSS),.VDD(VDD),.Y(I7296),.A(g2915));
  NOT NOT1_1236(.VSS(VSS),.VDD(VDD),.Y(g3831),.A(I7296));
  NOT NOT1_1237(.VSS(VSS),.VDD(VDD),.Y(I7299),.A(g2961));
  NOT NOT1_1238(.VSS(VSS),.VDD(VDD),.Y(g3832),.A(I7299));
  NOT NOT1_1239(.VSS(VSS),.VDD(VDD),.Y(I7302),.A(g2825));
  NOT NOT1_1240(.VSS(VSS),.VDD(VDD),.Y(g3833),.A(I7302));
  NOT NOT1_1241(.VSS(VSS),.VDD(VDD),.Y(I7305),.A(g3048));
  NOT NOT1_1242(.VSS(VSS),.VDD(VDD),.Y(g3834),.A(I7305));
  NOT NOT1_1243(.VSS(VSS),.VDD(VDD),.Y(I7308),.A(g3074));
  NOT NOT1_1244(.VSS(VSS),.VDD(VDD),.Y(g3835),.A(I7308));
  NOT NOT1_1245(.VSS(VSS),.VDD(VDD),.Y(I7311),.A(g2879));
  NOT NOT1_1246(.VSS(VSS),.VDD(VDD),.Y(g3836),.A(I7311));
  NOT NOT1_1247(.VSS(VSS),.VDD(VDD),.Y(I7314),.A(g2916));
  NOT NOT1_1248(.VSS(VSS),.VDD(VDD),.Y(g3837),.A(I7314));
  NOT NOT1_1249(.VSS(VSS),.VDD(VDD),.Y(I7317),.A(g2893));
  NOT NOT1_1250(.VSS(VSS),.VDD(VDD),.Y(g3838),.A(I7317));
  NOT NOT1_1251(.VSS(VSS),.VDD(VDD),.Y(I7320),.A(g2927));
  NOT NOT1_1252(.VSS(VSS),.VDD(VDD),.Y(g3839),.A(I7320));
  NOT NOT1_1253(.VSS(VSS),.VDD(VDD),.Y(I7323),.A(g2905));
  NOT NOT1_1254(.VSS(VSS),.VDD(VDD),.Y(g3840),.A(I7323));
  NOT NOT1_1255(.VSS(VSS),.VDD(VDD),.Y(I7326),.A(g2940));
  NOT NOT1_1256(.VSS(VSS),.VDD(VDD),.Y(g3841),.A(I7326));
  NOT NOT1_1257(.VSS(VSS),.VDD(VDD),.Y(I7329),.A(g2920));
  NOT NOT1_1258(.VSS(VSS),.VDD(VDD),.Y(g3842),.A(I7329));
  NOT NOT1_1259(.VSS(VSS),.VDD(VDD),.Y(I7332),.A(g2947));
  NOT NOT1_1260(.VSS(VSS),.VDD(VDD),.Y(g3843),.A(I7332));
  NOT NOT1_1261(.VSS(VSS),.VDD(VDD),.Y(I7335),.A(g2910));
  NOT NOT1_1262(.VSS(VSS),.VDD(VDD),.Y(g3844),.A(I7335));
  NOT NOT1_1263(.VSS(VSS),.VDD(VDD),.Y(I7338),.A(g2923));
  NOT NOT1_1264(.VSS(VSS),.VDD(VDD),.Y(g3845),.A(I7338));
  NOT NOT1_1265(.VSS(VSS),.VDD(VDD),.Y(I7341),.A(g2931));
  NOT NOT1_1266(.VSS(VSS),.VDD(VDD),.Y(g3846),.A(I7341));
  NOT NOT1_1267(.VSS(VSS),.VDD(VDD),.Y(I7344),.A(g2964));
  NOT NOT1_1268(.VSS(VSS),.VDD(VDD),.Y(g3847),.A(I7344));
  NOT NOT1_1269(.VSS(VSS),.VDD(VDD),.Y(I7347),.A(g2985));
  NOT NOT1_1270(.VSS(VSS),.VDD(VDD),.Y(g3848),.A(I7347));
  NOT NOT1_1271(.VSS(VSS),.VDD(VDD),.Y(I7350),.A(g2971));
  NOT NOT1_1272(.VSS(VSS),.VDD(VDD),.Y(g3849),.A(I7350));
  NOT NOT1_1273(.VSS(VSS),.VDD(VDD),.Y(I7353),.A(g2833));
  NOT NOT1_1274(.VSS(VSS),.VDD(VDD),.Y(g3850),.A(I7353));
  NOT NOT1_1275(.VSS(VSS),.VDD(VDD),.Y(I7356),.A(g2843));
  NOT NOT1_1276(.VSS(VSS),.VDD(VDD),.Y(g3851),.A(I7356));
  NOT NOT1_1277(.VSS(VSS),.VDD(VDD),.Y(I7359),.A(g2871));
  NOT NOT1_1278(.VSS(VSS),.VDD(VDD),.Y(g3852),.A(I7359));
  NOT NOT1_1279(.VSS(VSS),.VDD(VDD),.Y(I7362),.A(g2933));
  NOT NOT1_1280(.VSS(VSS),.VDD(VDD),.Y(g3853),.A(I7362));
  NOT NOT1_1281(.VSS(VSS),.VDD(VDD),.Y(I7365),.A(g3061));
  NOT NOT1_1282(.VSS(VSS),.VDD(VDD),.Y(g3854),.A(I7365));
  NOT NOT1_1283(.VSS(VSS),.VDD(VDD),.Y(I7368),.A(g3018));
  NOT NOT1_1284(.VSS(VSS),.VDD(VDD),.Y(g3855),.A(I7368));
  NOT NOT1_1285(.VSS(VSS),.VDD(VDD),.Y(I7371),.A(g3050));
  NOT NOT1_1286(.VSS(VSS),.VDD(VDD),.Y(g3856),.A(I7371));
  NOT NOT1_1287(.VSS(VSS),.VDD(VDD),.Y(I7374),.A(g3084));
  NOT NOT1_1288(.VSS(VSS),.VDD(VDD),.Y(g3857),.A(I7374));
  NOT NOT1_1289(.VSS(VSS),.VDD(VDD),.Y(I7377),.A(g3189));
  NOT NOT1_1290(.VSS(VSS),.VDD(VDD),.Y(g3858),.A(I7377));
  NOT NOT1_1291(.VSS(VSS),.VDD(VDD),.Y(I7380),.A(g3461));
  NOT NOT1_1292(.VSS(VSS),.VDD(VDD),.Y(g3859),.A(I7380));
  NOT NOT1_1293(.VSS(VSS),.VDD(VDD),.Y(I7383),.A(g3465));
  NOT NOT1_1294(.VSS(VSS),.VDD(VDD),.Y(g3860),.A(I7383));
  NOT NOT1_1295(.VSS(VSS),.VDD(VDD),.Y(I7386),.A(g3013));
  NOT NOT1_1296(.VSS(VSS),.VDD(VDD),.Y(g3861),.A(I7386));
  NOT NOT1_1297(.VSS(VSS),.VDD(VDD),.Y(I7389),.A(g3496));
  NOT NOT1_1298(.VSS(VSS),.VDD(VDD),.Y(g3862),.A(I7389));
  NOT NOT1_1299(.VSS(VSS),.VDD(VDD),.Y(I7392),.A(g3230));
  NOT NOT1_1300(.VSS(VSS),.VDD(VDD),.Y(g3863),.A(I7392));
  NOT NOT1_1301(.VSS(VSS),.VDD(VDD),.Y(g3864),.A(g2943));
  NOT NOT1_1302(.VSS(VSS),.VDD(VDD),.Y(g3865),.A(g2944));
  NOT NOT1_1303(.VSS(VSS),.VDD(VDD),.Y(g3866),.A(g2945));
  NOT NOT1_1304(.VSS(VSS),.VDD(VDD),.Y(g3867),.A(g2946));
  NOT NOT1_1305(.VSS(VSS),.VDD(VDD),.Y(g3868),.A(g2948));
  NOT NOT1_1306(.VSS(VSS),.VDD(VDD),.Y(I7400),.A(g3075));
  NOT NOT1_1307(.VSS(VSS),.VDD(VDD),.Y(g3869),.A(I7400));
  NOT NOT1_1308(.VSS(VSS),.VDD(VDD),.Y(g3870),.A(g3466));
  NOT NOT1_1309(.VSS(VSS),.VDD(VDD),.Y(g3871),.A(g2953));
  NOT NOT1_1310(.VSS(VSS),.VDD(VDD),.Y(g3872),.A(g2954));
  NOT NOT1_1311(.VSS(VSS),.VDD(VDD),.Y(g3873),.A(g2956));
  NOT NOT1_1312(.VSS(VSS),.VDD(VDD),.Y(g3874),.A(g2957));
  NOT NOT1_1313(.VSS(VSS),.VDD(VDD),.Y(g3875),.A(g2958));
  NOT NOT1_1314(.VSS(VSS),.VDD(VDD),.Y(g3876),.A(g3466));
  NOT NOT1_1315(.VSS(VSS),.VDD(VDD),.Y(g3877),.A(g2960));
  NOT NOT1_1316(.VSS(VSS),.VDD(VDD),.Y(g3878),.A(g2962));
  NOT NOT1_1317(.VSS(VSS),.VDD(VDD),.Y(g3879),.A(g2963));
  NOT NOT1_1318(.VSS(VSS),.VDD(VDD),.Y(g3880),.A(g2965));
  NOT NOT1_1319(.VSS(VSS),.VDD(VDD),.Y(g3881),.A(g2969));
  NOT NOT1_1320(.VSS(VSS),.VDD(VDD),.Y(g3882),.A(g2970));
  NOT NOT1_1321(.VSS(VSS),.VDD(VDD),.Y(I7417),.A(g3659));
  NOT NOT1_1322(.VSS(VSS),.VDD(VDD),.Y(g3884),.A(I7417));
  NOT NOT1_1323(.VSS(VSS),.VDD(VDD),.Y(g3888),.A(g3097));
  NOT NOT1_1324(.VSS(VSS),.VDD(VDD),.Y(g3891),.A(g3097));
  NOT NOT1_1325(.VSS(VSS),.VDD(VDD),.Y(g3892),.A(g3131));
  NOT NOT1_1326(.VSS(VSS),.VDD(VDD),.Y(I7473),.A(g3546));
  NOT NOT1_1327(.VSS(VSS),.VDD(VDD),.Y(g3896),.A(I7473));
  NOT NOT1_1328(.VSS(VSS),.VDD(VDD),.Y(g3897),.A(g3131));
  NOT NOT1_1329(.VSS(VSS),.VDD(VDD),.Y(g3898),.A(g3160));
  NOT NOT1_1330(.VSS(VSS),.VDD(VDD),.Y(I7492),.A(g3561));
  NOT NOT1_1331(.VSS(VSS),.VDD(VDD),.Y(g3901),.A(I7492));
  NOT NOT1_1332(.VSS(VSS),.VDD(VDD),.Y(I7495),.A(g3562));
  NOT NOT1_1333(.VSS(VSS),.VDD(VDD),.Y(g3902),.A(I7495));
  NOT NOT1_1334(.VSS(VSS),.VDD(VDD),.Y(I7498),.A(g2752));
  NOT NOT1_1335(.VSS(VSS),.VDD(VDD),.Y(g3903),.A(I7498));
  NOT NOT1_1336(.VSS(VSS),.VDD(VDD),.Y(g3904),.A(g3160));
  NOT NOT1_1337(.VSS(VSS),.VDD(VDD),.Y(g3905),.A(g3192));
  NOT NOT1_1338(.VSS(VSS),.VDD(VDD),.Y(I7517),.A(g3578));
  NOT NOT1_1339(.VSS(VSS),.VDD(VDD),.Y(g3908),.A(I7517));
  NOT NOT1_1340(.VSS(VSS),.VDD(VDD),.Y(I7520),.A(g2734));
  NOT NOT1_1341(.VSS(VSS),.VDD(VDD),.Y(g3909),.A(I7520));
  NOT NOT1_1342(.VSS(VSS),.VDD(VDD),.Y(I7523),.A(g2562));
  NOT NOT1_1343(.VSS(VSS),.VDD(VDD),.Y(g3910),.A(I7523));
  NOT NOT1_1344(.VSS(VSS),.VDD(VDD),.Y(I7526),.A(g2752));
  NOT NOT1_1345(.VSS(VSS),.VDD(VDD),.Y(g3911),.A(I7526));
  NOT NOT1_1346(.VSS(VSS),.VDD(VDD),.Y(g3912),.A(g3192));
  NOT NOT1_1347(.VSS(VSS),.VDD(VDD),.Y(g3913),.A(g2834));
  NOT NOT1_1348(.VSS(VSS),.VDD(VDD),.Y(I7545),.A(g3589));
  NOT NOT1_1349(.VSS(VSS),.VDD(VDD),.Y(g3916),.A(I7545));
  NOT NOT1_1350(.VSS(VSS),.VDD(VDD),.Y(I7548),.A(g3590));
  NOT NOT1_1351(.VSS(VSS),.VDD(VDD),.Y(g3917),.A(I7548));
  NOT NOT1_1352(.VSS(VSS),.VDD(VDD),.Y(I7551),.A(g2712));
  NOT NOT1_1353(.VSS(VSS),.VDD(VDD),.Y(g3918),.A(I7551));
  NOT NOT1_1354(.VSS(VSS),.VDD(VDD),.Y(I7554),.A(g2573));
  NOT NOT1_1355(.VSS(VSS),.VDD(VDD),.Y(g3919),.A(I7554));
  NOT NOT1_1356(.VSS(VSS),.VDD(VDD),.Y(g3920),.A(g3097));
  NOT NOT1_1357(.VSS(VSS),.VDD(VDD),.Y(I7558),.A(g2734));
  NOT NOT1_1358(.VSS(VSS),.VDD(VDD),.Y(g3921),.A(I7558));
  NOT NOT1_1359(.VSS(VSS),.VDD(VDD),.Y(I7561),.A(g2562));
  NOT NOT1_1360(.VSS(VSS),.VDD(VDD),.Y(g3922),.A(I7561));
  NOT NOT1_1361(.VSS(VSS),.VDD(VDD),.Y(I7564),.A(g2752));
  NOT NOT1_1362(.VSS(VSS),.VDD(VDD),.Y(g3923),.A(I7564));
  NOT NOT1_1363(.VSS(VSS),.VDD(VDD),.Y(I7581),.A(g3612));
  NOT NOT1_1364(.VSS(VSS),.VDD(VDD),.Y(g3926),.A(I7581));
  NOT NOT1_1365(.VSS(VSS),.VDD(VDD),.Y(I7584),.A(g3062));
  NOT NOT1_1366(.VSS(VSS),.VDD(VDD),.Y(g3927),.A(I7584));
  NOT NOT1_1367(.VSS(VSS),.VDD(VDD),.Y(g3928),.A(g3097));
  NOT NOT1_1368(.VSS(VSS),.VDD(VDD),.Y(I7588),.A(g2584));
  NOT NOT1_1369(.VSS(VSS),.VDD(VDD),.Y(g3929),.A(I7588));
  NOT NOT1_1370(.VSS(VSS),.VDD(VDD),.Y(g3930),.A(g3097));
  NOT NOT1_1371(.VSS(VSS),.VDD(VDD),.Y(I7592),.A(g2712));
  NOT NOT1_1372(.VSS(VSS),.VDD(VDD),.Y(g3931),.A(I7592));
  NOT NOT1_1373(.VSS(VSS),.VDD(VDD),.Y(I7595),.A(g2573));
  NOT NOT1_1374(.VSS(VSS),.VDD(VDD),.Y(g3932),.A(I7595));
  NOT NOT1_1375(.VSS(VSS),.VDD(VDD),.Y(g3933),.A(g3131));
  NOT NOT1_1376(.VSS(VSS),.VDD(VDD),.Y(I7599),.A(g2734));
  NOT NOT1_1377(.VSS(VSS),.VDD(VDD),.Y(g3934),.A(I7599));
  NOT NOT1_1378(.VSS(VSS),.VDD(VDD),.Y(I7602),.A(g2562));
  NOT NOT1_1379(.VSS(VSS),.VDD(VDD),.Y(g3935),.A(I7602));
  NOT NOT1_1380(.VSS(VSS),.VDD(VDD),.Y(I7605),.A(g2752));
  NOT NOT1_1381(.VSS(VSS),.VDD(VDD),.Y(g3936),.A(I7605));
  NOT NOT1_1382(.VSS(VSS),.VDD(VDD),.Y(g3937),.A(g2845));
  NOT NOT1_1383(.VSS(VSS),.VDD(VDD),.Y(I7623),.A(g3631));
  NOT NOT1_1384(.VSS(VSS),.VDD(VDD),.Y(g3940),.A(I7623));
  NOT NOT1_1385(.VSS(VSS),.VDD(VDD),.Y(I7626),.A(g3632));
  NOT NOT1_1386(.VSS(VSS),.VDD(VDD),.Y(g3941),.A(I7626));
  NOT NOT1_1387(.VSS(VSS),.VDD(VDD),.Y(I7629),.A(g3633));
  NOT NOT1_1388(.VSS(VSS),.VDD(VDD),.Y(g3942),.A(I7629));
  NOT NOT1_1389(.VSS(VSS),.VDD(VDD),.Y(I7632),.A(g3634));
  NOT NOT1_1390(.VSS(VSS),.VDD(VDD),.Y(g3943),.A(I7632));
  NOT NOT1_1391(.VSS(VSS),.VDD(VDD),.Y(I7635),.A(g3052));
  NOT NOT1_1392(.VSS(VSS),.VDD(VDD),.Y(g3944),.A(I7635));
  NOT NOT1_1393(.VSS(VSS),.VDD(VDD),.Y(g3945),.A(g3097));
  NOT NOT1_1394(.VSS(VSS),.VDD(VDD),.Y(g3946),.A(g3097));
  NOT NOT1_1395(.VSS(VSS),.VDD(VDD),.Y(I7640),.A(g3062));
  NOT NOT1_1396(.VSS(VSS),.VDD(VDD),.Y(g3947),.A(I7640));
  NOT NOT1_1397(.VSS(VSS),.VDD(VDD),.Y(g3948),.A(g3131));
  NOT NOT1_1398(.VSS(VSS),.VDD(VDD),.Y(I7644),.A(g2584));
  NOT NOT1_1399(.VSS(VSS),.VDD(VDD),.Y(g3949),.A(I7644));
  NOT NOT1_1400(.VSS(VSS),.VDD(VDD),.Y(g3950),.A(g3131));
  NOT NOT1_1401(.VSS(VSS),.VDD(VDD),.Y(I7648),.A(g2712));
  NOT NOT1_1402(.VSS(VSS),.VDD(VDD),.Y(g3951),.A(I7648));
  NOT NOT1_1403(.VSS(VSS),.VDD(VDD),.Y(I7651),.A(g2573));
  NOT NOT1_1404(.VSS(VSS),.VDD(VDD),.Y(g3952),.A(I7651));
  NOT NOT1_1405(.VSS(VSS),.VDD(VDD),.Y(g3953),.A(g3160));
  NOT NOT1_1406(.VSS(VSS),.VDD(VDD),.Y(I7655),.A(g2734));
  NOT NOT1_1407(.VSS(VSS),.VDD(VDD),.Y(g3954),.A(I7655));
  NOT NOT1_1408(.VSS(VSS),.VDD(VDD),.Y(I7658),.A(g2562));
  NOT NOT1_1409(.VSS(VSS),.VDD(VDD),.Y(g3955),.A(I7658));
  NOT NOT1_1410(.VSS(VSS),.VDD(VDD),.Y(g3956),.A(g2845));
  NOT NOT1_1411(.VSS(VSS),.VDD(VDD),.Y(I7662),.A(g3642));
  NOT NOT1_1412(.VSS(VSS),.VDD(VDD),.Y(g3957),.A(I7662));
  NOT NOT1_1413(.VSS(VSS),.VDD(VDD),.Y(g3958),.A(g3097));
  NOT NOT1_1414(.VSS(VSS),.VDD(VDD),.Y(g3959),.A(g3097));
  NOT NOT1_1415(.VSS(VSS),.VDD(VDD),.Y(I7667),.A(g3052));
  NOT NOT1_1416(.VSS(VSS),.VDD(VDD),.Y(g3960),.A(I7667));
  NOT NOT1_1417(.VSS(VSS),.VDD(VDD),.Y(g3961),.A(g3131));
  NOT NOT1_1418(.VSS(VSS),.VDD(VDD),.Y(g3962),.A(g3131));
  NOT NOT1_1419(.VSS(VSS),.VDD(VDD),.Y(I7672),.A(g3062));
  NOT NOT1_1420(.VSS(VSS),.VDD(VDD),.Y(g3963),.A(I7672));
  NOT NOT1_1421(.VSS(VSS),.VDD(VDD),.Y(g3964),.A(g3160));
  NOT NOT1_1422(.VSS(VSS),.VDD(VDD),.Y(I7676),.A(g2584));
  NOT NOT1_1423(.VSS(VSS),.VDD(VDD),.Y(g3965),.A(I7676));
  NOT NOT1_1424(.VSS(VSS),.VDD(VDD),.Y(g3966),.A(g3160));
  NOT NOT1_1425(.VSS(VSS),.VDD(VDD),.Y(I7680),.A(g2712));
  NOT NOT1_1426(.VSS(VSS),.VDD(VDD),.Y(g3967),.A(I7680));
  NOT NOT1_1427(.VSS(VSS),.VDD(VDD),.Y(I7683),.A(g2573));
  NOT NOT1_1428(.VSS(VSS),.VDD(VDD),.Y(g3968),.A(I7683));
  NOT NOT1_1429(.VSS(VSS),.VDD(VDD),.Y(g3969),.A(g3192));
  NOT NOT1_1430(.VSS(VSS),.VDD(VDD),.Y(g3970),.A(g2845));
  NOT NOT1_1431(.VSS(VSS),.VDD(VDD),.Y(I7688),.A(g3650));
  NOT NOT1_1432(.VSS(VSS),.VDD(VDD),.Y(g3971),.A(I7688));
  NOT NOT1_1433(.VSS(VSS),.VDD(VDD),.Y(I7691),.A(g3651));
  NOT NOT1_1434(.VSS(VSS),.VDD(VDD),.Y(g3972),.A(I7691));
  NOT NOT1_1435(.VSS(VSS),.VDD(VDD),.Y(g3973),.A(g3097));
  NOT NOT1_1436(.VSS(VSS),.VDD(VDD),.Y(g3974),.A(g3131));
  NOT NOT1_1437(.VSS(VSS),.VDD(VDD),.Y(g3975),.A(g3131));
  NOT NOT1_1438(.VSS(VSS),.VDD(VDD),.Y(I7697),.A(g3052));
  NOT NOT1_1439(.VSS(VSS),.VDD(VDD),.Y(g3976),.A(I7697));
  NOT NOT1_1440(.VSS(VSS),.VDD(VDD),.Y(g3977),.A(g3160));
  NOT NOT1_1441(.VSS(VSS),.VDD(VDD),.Y(g3978),.A(g3160));
  NOT NOT1_1442(.VSS(VSS),.VDD(VDD),.Y(I7702),.A(g3062));
  NOT NOT1_1443(.VSS(VSS),.VDD(VDD),.Y(g3979),.A(I7702));
  NOT NOT1_1444(.VSS(VSS),.VDD(VDD),.Y(g3980),.A(g3192));
  NOT NOT1_1445(.VSS(VSS),.VDD(VDD),.Y(I7706),.A(g2584));
  NOT NOT1_1446(.VSS(VSS),.VDD(VDD),.Y(g3981),.A(I7706));
  NOT NOT1_1447(.VSS(VSS),.VDD(VDD),.Y(g3982),.A(g3192));
  NOT NOT1_1448(.VSS(VSS),.VDD(VDD),.Y(g3983),.A(g2845));
  NOT NOT1_1449(.VSS(VSS),.VDD(VDD),.Y(I7712),.A(g3657));
  NOT NOT1_1450(.VSS(VSS),.VDD(VDD),.Y(g3985),.A(I7712));
  NOT NOT1_1451(.VSS(VSS),.VDD(VDD),.Y(I7716),.A(g3038));
  NOT NOT1_1452(.VSS(VSS),.VDD(VDD),.Y(g3987),.A(I7716));
  NOT NOT1_1453(.VSS(VSS),.VDD(VDD),.Y(g3988),.A(g3097));
  NOT NOT1_1454(.VSS(VSS),.VDD(VDD),.Y(g3989),.A(g3131));
  NOT NOT1_1455(.VSS(VSS),.VDD(VDD),.Y(g3990),.A(g3160));
  NOT NOT1_1456(.VSS(VSS),.VDD(VDD),.Y(g3991),.A(g3160));
  NOT NOT1_1457(.VSS(VSS),.VDD(VDD),.Y(I7723),.A(g3052));
  NOT NOT1_1458(.VSS(VSS),.VDD(VDD),.Y(g3992),.A(I7723));
  NOT NOT1_1459(.VSS(VSS),.VDD(VDD),.Y(g3993),.A(g3192));
  NOT NOT1_1460(.VSS(VSS),.VDD(VDD),.Y(g3994),.A(g3192));
  NOT NOT1_1461(.VSS(VSS),.VDD(VDD),.Y(I7728),.A(g3675));
  NOT NOT1_1462(.VSS(VSS),.VDD(VDD),.Y(g3995),.A(I7728));
  NOT NOT1_1463(.VSS(VSS),.VDD(VDD),.Y(I7731),.A(g3029));
  NOT NOT1_1464(.VSS(VSS),.VDD(VDD),.Y(g3996),.A(I7731));
  NOT NOT1_1465(.VSS(VSS),.VDD(VDD),.Y(I7734),.A(g2595));
  NOT NOT1_1466(.VSS(VSS),.VDD(VDD),.Y(g3997),.A(I7734));
  NOT NOT1_1467(.VSS(VSS),.VDD(VDD),.Y(g3998),.A(g3097));
  NOT NOT1_1468(.VSS(VSS),.VDD(VDD),.Y(I7738),.A(g3038));
  NOT NOT1_1469(.VSS(VSS),.VDD(VDD),.Y(g3999),.A(I7738));
  NOT NOT1_1470(.VSS(VSS),.VDD(VDD),.Y(g4000),.A(g3131));
  NOT NOT1_1471(.VSS(VSS),.VDD(VDD),.Y(g4001),.A(g3160));
  NOT NOT1_1472(.VSS(VSS),.VDD(VDD),.Y(g4002),.A(g3192));
  NOT NOT1_1473(.VSS(VSS),.VDD(VDD),.Y(g4003),.A(g3192));
  NOT NOT1_1474(.VSS(VSS),.VDD(VDD),.Y(g4004),.A(g2845));
  NOT NOT1_1475(.VSS(VSS),.VDD(VDD),.Y(I7746),.A(g3591));
  NOT NOT1_1476(.VSS(VSS),.VDD(VDD),.Y(g4005),.A(I7746));
  NOT NOT1_1477(.VSS(VSS),.VDD(VDD),.Y(I7749),.A(g3692));
  NOT NOT1_1478(.VSS(VSS),.VDD(VDD),.Y(g4006),.A(I7749));
  NOT NOT1_1479(.VSS(VSS),.VDD(VDD),.Y(I7752),.A(g3591));
  NOT NOT1_1480(.VSS(VSS),.VDD(VDD),.Y(g4007),.A(I7752));
  NOT NOT1_1481(.VSS(VSS),.VDD(VDD),.Y(I7755),.A(g3019));
  NOT NOT1_1482(.VSS(VSS),.VDD(VDD),.Y(g4008),.A(I7755));
  NOT NOT1_1483(.VSS(VSS),.VDD(VDD),.Y(I7758),.A(g2605));
  NOT NOT1_1484(.VSS(VSS),.VDD(VDD),.Y(g4009),.A(I7758));
  NOT NOT1_1485(.VSS(VSS),.VDD(VDD),.Y(g4010),.A(g3097));
  NOT NOT1_1486(.VSS(VSS),.VDD(VDD),.Y(I7762),.A(g3029));
  NOT NOT1_1487(.VSS(VSS),.VDD(VDD),.Y(g4011),.A(I7762));
  NOT NOT1_1488(.VSS(VSS),.VDD(VDD),.Y(I7765),.A(g2595));
  NOT NOT1_1489(.VSS(VSS),.VDD(VDD),.Y(g4012),.A(I7765));
  NOT NOT1_1490(.VSS(VSS),.VDD(VDD),.Y(g4013),.A(g3131));
  NOT NOT1_1491(.VSS(VSS),.VDD(VDD),.Y(I7769),.A(g3038));
  NOT NOT1_1492(.VSS(VSS),.VDD(VDD),.Y(g4014),.A(I7769));
  NOT NOT1_1493(.VSS(VSS),.VDD(VDD),.Y(g4015),.A(g3160));
  NOT NOT1_1494(.VSS(VSS),.VDD(VDD),.Y(g4016),.A(g3192));
  NOT NOT1_1495(.VSS(VSS),.VDD(VDD),.Y(g4017),.A(g2845));
  NOT NOT1_1496(.VSS(VSS),.VDD(VDD),.Y(I7775),.A(g3705));
  NOT NOT1_1497(.VSS(VSS),.VDD(VDD),.Y(g4018),.A(I7775));
  NOT NOT1_1498(.VSS(VSS),.VDD(VDD),.Y(I7778),.A(g3019));
  NOT NOT1_1499(.VSS(VSS),.VDD(VDD),.Y(g4019),.A(I7778));
  NOT NOT1_1500(.VSS(VSS),.VDD(VDD),.Y(I7781),.A(g2605));
  NOT NOT1_1501(.VSS(VSS),.VDD(VDD),.Y(g4020),.A(I7781));
  NOT NOT1_1502(.VSS(VSS),.VDD(VDD),.Y(g4021),.A(g3131));
  NOT NOT1_1503(.VSS(VSS),.VDD(VDD),.Y(I7785),.A(g3029));
  NOT NOT1_1504(.VSS(VSS),.VDD(VDD),.Y(g4022),.A(I7785));
  NOT NOT1_1505(.VSS(VSS),.VDD(VDD),.Y(I7788),.A(g2595));
  NOT NOT1_1506(.VSS(VSS),.VDD(VDD),.Y(g4023),.A(I7788));
  NOT NOT1_1507(.VSS(VSS),.VDD(VDD),.Y(g4024),.A(g3160));
  NOT NOT1_1508(.VSS(VSS),.VDD(VDD),.Y(I7792),.A(g3038));
  NOT NOT1_1509(.VSS(VSS),.VDD(VDD),.Y(g4025),.A(I7792));
  NOT NOT1_1510(.VSS(VSS),.VDD(VDD),.Y(g4026),.A(g3192));
  NOT NOT1_1511(.VSS(VSS),.VDD(VDD),.Y(g4027),.A(g2845));
  NOT NOT1_1512(.VSS(VSS),.VDD(VDD),.Y(I7797),.A(g3019));
  NOT NOT1_1513(.VSS(VSS),.VDD(VDD),.Y(g4028),.A(I7797));
  NOT NOT1_1514(.VSS(VSS),.VDD(VDD),.Y(I7800),.A(g2605));
  NOT NOT1_1515(.VSS(VSS),.VDD(VDD),.Y(g4029),.A(I7800));
  NOT NOT1_1516(.VSS(VSS),.VDD(VDD),.Y(g4030),.A(g3160));
  NOT NOT1_1517(.VSS(VSS),.VDD(VDD),.Y(I7804),.A(g3029));
  NOT NOT1_1518(.VSS(VSS),.VDD(VDD),.Y(g4031),.A(I7804));
  NOT NOT1_1519(.VSS(VSS),.VDD(VDD),.Y(I7807),.A(g2595));
  NOT NOT1_1520(.VSS(VSS),.VDD(VDD),.Y(g4032),.A(I7807));
  NOT NOT1_1521(.VSS(VSS),.VDD(VDD),.Y(g4033),.A(g3192));
  NOT NOT1_1522(.VSS(VSS),.VDD(VDD),.Y(I7811),.A(g3019));
  NOT NOT1_1523(.VSS(VSS),.VDD(VDD),.Y(g4034),.A(I7811));
  NOT NOT1_1524(.VSS(VSS),.VDD(VDD),.Y(I7814),.A(g2605));
  NOT NOT1_1525(.VSS(VSS),.VDD(VDD),.Y(g4035),.A(I7814));
  NOT NOT1_1526(.VSS(VSS),.VDD(VDD),.Y(g4036),.A(g3192));
  NOT NOT1_1527(.VSS(VSS),.VDD(VDD),.Y(g4037),.A(g2845));
  NOT NOT1_1528(.VSS(VSS),.VDD(VDD),.Y(g4041),.A(g2605));
  NOT NOT1_1529(.VSS(VSS),.VDD(VDD),.Y(g4044),.A(g2595));
  NOT NOT1_1530(.VSS(VSS),.VDD(VDD),.Y(g4050),.A(g3080));
  NOT NOT1_1531(.VSS(VSS),.VDD(VDD),.Y(g4051),.A(g3093));
  NOT NOT1_1532(.VSS(VSS),.VDD(VDD),.Y(g4056),.A(g3082));
  NOT NOT1_1533(.VSS(VSS),.VDD(VDD),.Y(I7832),.A(g2768));
  NOT NOT1_1534(.VSS(VSS),.VDD(VDD),.Y(g4057),.A(I7832));
  NOT NOT1_1535(.VSS(VSS),.VDD(VDD),.Y(I7838),.A(g2781));
  NOT NOT1_1536(.VSS(VSS),.VDD(VDD),.Y(g4065),.A(I7838));
  NOT NOT1_1537(.VSS(VSS),.VDD(VDD),.Y(I7844),.A(g3784));
  NOT NOT1_1538(.VSS(VSS),.VDD(VDD),.Y(g4069),.A(I7844));
  NOT NOT1_1539(.VSS(VSS),.VDD(VDD),.Y(I7847),.A(g3798));
  NOT NOT1_1540(.VSS(VSS),.VDD(VDD),.Y(g4070),.A(I7847));
  NOT NOT1_1541(.VSS(VSS),.VDD(VDD),.Y(I7850),.A(g2795));
  NOT NOT1_1542(.VSS(VSS),.VDD(VDD),.Y(g4071),.A(I7850));
  NOT NOT1_1543(.VSS(VSS),.VDD(VDD),.Y(I7856),.A(g3805));
  NOT NOT1_1544(.VSS(VSS),.VDD(VDD),.Y(g4075),.A(I7856));
  NOT NOT1_1545(.VSS(VSS),.VDD(VDD),.Y(I7859),.A(g2804));
  NOT NOT1_1546(.VSS(VSS),.VDD(VDD),.Y(g4076),.A(I7859));
  NOT NOT1_1547(.VSS(VSS),.VDD(VDD),.Y(I7864),.A(g3812));
  NOT NOT1_1548(.VSS(VSS),.VDD(VDD),.Y(g4079),.A(I7864));
  NOT NOT1_1549(.VSS(VSS),.VDD(VDD),.Y(I7867),.A(g2818));
  NOT NOT1_1550(.VSS(VSS),.VDD(VDD),.Y(g4080),.A(I7867));
  NOT NOT1_1551(.VSS(VSS),.VDD(VDD),.Y(I7870),.A(g2827));
  NOT NOT1_1552(.VSS(VSS),.VDD(VDD),.Y(g4081),.A(I7870));
  NOT NOT1_1553(.VSS(VSS),.VDD(VDD),.Y(I7875),.A(g3819));
  NOT NOT1_1554(.VSS(VSS),.VDD(VDD),.Y(g4084),.A(I7875));
  NOT NOT1_1555(.VSS(VSS),.VDD(VDD),.Y(I7878),.A(g2829));
  NOT NOT1_1556(.VSS(VSS),.VDD(VDD),.Y(g4085),.A(I7878));
  NOT NOT1_1557(.VSS(VSS),.VDD(VDD),.Y(I7882),.A(g2700));
  NOT NOT1_1558(.VSS(VSS),.VDD(VDD),.Y(g4087),.A(I7882));
  NOT NOT1_1559(.VSS(VSS),.VDD(VDD),.Y(I7885),.A(g2837));
  NOT NOT1_1560(.VSS(VSS),.VDD(VDD),.Y(g4088),.A(I7885));
  NOT NOT1_1561(.VSS(VSS),.VDD(VDD),.Y(I7888),.A(g3505));
  NOT NOT1_1562(.VSS(VSS),.VDD(VDD),.Y(g4089),.A(I7888));
  NOT NOT1_1563(.VSS(VSS),.VDD(VDD),.Y(I7899),.A(g3743));
  NOT NOT1_1564(.VSS(VSS),.VDD(VDD),.Y(g4092),.A(I7899));
  NOT NOT1_1565(.VSS(VSS),.VDD(VDD),.Y(I7902),.A(g2709));
  NOT NOT1_1566(.VSS(VSS),.VDD(VDD),.Y(g4093),.A(I7902));
  NOT NOT1_1567(.VSS(VSS),.VDD(VDD),.Y(I7905),.A(g2863));
  NOT NOT1_1568(.VSS(VSS),.VDD(VDD),.Y(g4094),.A(I7905));
  NOT NOT1_1569(.VSS(VSS),.VDD(VDD),.Y(I7908),.A(g3516));
  NOT NOT1_1570(.VSS(VSS),.VDD(VDD),.Y(g4095),.A(I7908));
  NOT NOT1_1571(.VSS(VSS),.VDD(VDD),.Y(I7911),.A(g2767));
  NOT NOT1_1572(.VSS(VSS),.VDD(VDD),.Y(g4096),.A(I7911));
  NOT NOT1_1573(.VSS(VSS),.VDD(VDD),.Y(I7919),.A(g3761));
  NOT NOT1_1574(.VSS(VSS),.VDD(VDD),.Y(g4102),.A(I7919));
  NOT NOT1_1575(.VSS(VSS),.VDD(VDD),.Y(I7922),.A(g3462));
  NOT NOT1_1576(.VSS(VSS),.VDD(VDD),.Y(g4103),.A(I7922));
  NOT NOT1_1577(.VSS(VSS),.VDD(VDD),.Y(I7925),.A(g2761));
  NOT NOT1_1578(.VSS(VSS),.VDD(VDD),.Y(g4104),.A(I7925));
  NOT NOT1_1579(.VSS(VSS),.VDD(VDD),.Y(I7928),.A(g2873));
  NOT NOT1_1580(.VSS(VSS),.VDD(VDD),.Y(g4105),.A(I7928));
  NOT NOT1_1581(.VSS(VSS),.VDD(VDD),.Y(I7931),.A(g2780));
  NOT NOT1_1582(.VSS(VSS),.VDD(VDD),.Y(g4106),.A(I7931));
  NOT NOT1_1583(.VSS(VSS),.VDD(VDD),.Y(I7944),.A(g3774));
  NOT NOT1_1584(.VSS(VSS),.VDD(VDD),.Y(g4111),.A(I7944));
  NOT NOT1_1585(.VSS(VSS),.VDD(VDD),.Y(I7947),.A(g3485));
  NOT NOT1_1586(.VSS(VSS),.VDD(VDD),.Y(g4112),.A(I7947));
  NOT NOT1_1587(.VSS(VSS),.VDD(VDD),.Y(I7950),.A(g2774));
  NOT NOT1_1588(.VSS(VSS),.VDD(VDD),.Y(g4113),.A(I7950));
  NOT NOT1_1589(.VSS(VSS),.VDD(VDD),.Y(I7953),.A(g3542));
  NOT NOT1_1590(.VSS(VSS),.VDD(VDD),.Y(g4114),.A(I7953));
  NOT NOT1_1591(.VSS(VSS),.VDD(VDD),.Y(I7956),.A(g2810));
  NOT NOT1_1592(.VSS(VSS),.VDD(VDD),.Y(g4115),.A(I7956));
  NOT NOT1_1593(.VSS(VSS),.VDD(VDD),.Y(I7959),.A(g2793));
  NOT NOT1_1594(.VSS(VSS),.VDD(VDD),.Y(g4116),.A(I7959));
  NOT NOT1_1595(.VSS(VSS),.VDD(VDD),.Y(I7964),.A(g3488));
  NOT NOT1_1596(.VSS(VSS),.VDD(VDD),.Y(g4119),.A(I7964));
  NOT NOT1_1597(.VSS(VSS),.VDD(VDD),.Y(I7967),.A(g2787));
  NOT NOT1_1598(.VSS(VSS),.VDD(VDD),.Y(g4120),.A(I7967));
  NOT NOT1_1599(.VSS(VSS),.VDD(VDD),.Y(I7970),.A(g3557));
  NOT NOT1_1600(.VSS(VSS),.VDD(VDD),.Y(g4121),.A(I7970));
  NOT NOT1_1601(.VSS(VSS),.VDD(VDD),.Y(I7973),.A(g3071));
  NOT NOT1_1602(.VSS(VSS),.VDD(VDD),.Y(g4122),.A(I7973));
  NOT NOT1_1603(.VSS(VSS),.VDD(VDD),.Y(I7978),.A(g3574));
  NOT NOT1_1604(.VSS(VSS),.VDD(VDD),.Y(g4125),.A(I7978));
  NOT NOT1_1605(.VSS(VSS),.VDD(VDD),.Y(I7981),.A(g3555));
  NOT NOT1_1606(.VSS(VSS),.VDD(VDD),.Y(g4126),.A(I7981));
  NOT NOT1_1607(.VSS(VSS),.VDD(VDD),.Y(I7987),.A(g3528));
  NOT NOT1_1608(.VSS(VSS),.VDD(VDD),.Y(g4130),.A(I7987));
  NOT NOT1_1609(.VSS(VSS),.VDD(VDD),.Y(g4134),.A(g3676));
  NOT NOT1_1610(.VSS(VSS),.VDD(VDD),.Y(I8011),.A(g3225));
  NOT NOT1_1611(.VSS(VSS),.VDD(VDD),.Y(g4146),.A(I8011));
  NOT NOT1_1612(.VSS(VSS),.VDD(VDD),.Y(I8024),.A(g3076));
  NOT NOT1_1613(.VSS(VSS),.VDD(VDD),.Y(g4153),.A(I8024));
  NOT NOT1_1614(.VSS(VSS),.VDD(VDD),.Y(I8084),.A(g3706));
  NOT NOT1_1615(.VSS(VSS),.VDD(VDD),.Y(g4191),.A(I8084));
  NOT NOT1_1616(.VSS(VSS),.VDD(VDD),.Y(I8094),.A(g2976));
  NOT NOT1_1617(.VSS(VSS),.VDD(VDD),.Y(g4195),.A(I8094));
  NOT NOT1_1618(.VSS(VSS),.VDD(VDD),.Y(I8097),.A(g3237));
  NOT NOT1_1619(.VSS(VSS),.VDD(VDD),.Y(g4196),.A(I8097));
  NOT NOT1_1620(.VSS(VSS),.VDD(VDD),.Y(g4197),.A(g3591));
  NOT NOT1_1621(.VSS(VSS),.VDD(VDD),.Y(I8101),.A(g3259));
  NOT NOT1_1622(.VSS(VSS),.VDD(VDD),.Y(g4198),.A(I8101));
  NOT NOT1_1623(.VSS(VSS),.VDD(VDD),.Y(I8105),.A(g3339));
  NOT NOT1_1624(.VSS(VSS),.VDD(VDD),.Y(g4200),.A(I8105));
  NOT NOT1_1625(.VSS(VSS),.VDD(VDD),.Y(g4202),.A(g2810));
  NOT NOT1_1626(.VSS(VSS),.VDD(VDD),.Y(g4226),.A(g3591));
  NOT NOT1_1627(.VSS(VSS),.VDD(VDD),.Y(I8140),.A(g3429));
  NOT NOT1_1628(.VSS(VSS),.VDD(VDD),.Y(g4229),.A(I8140));
  NOT NOT1_1629(.VSS(VSS),.VDD(VDD),.Y(I8161),.A(g3517));
  NOT NOT1_1630(.VSS(VSS),.VDD(VDD),.Y(g4242),.A(I8161));
  NOT NOT1_1631(.VSS(VSS),.VDD(VDD),.Y(I8172),.A(g3524));
  NOT NOT1_1632(.VSS(VSS),.VDD(VDD),.Y(g4245),.A(I8172));
  NOT NOT1_1633(.VSS(VSS),.VDD(VDD),.Y(I8177),.A(g2810));
  NOT NOT1_1634(.VSS(VSS),.VDD(VDD),.Y(g4250),.A(I8177));
  NOT NOT1_1635(.VSS(VSS),.VDD(VDD),.Y(I8180),.A(g3529));
  NOT NOT1_1636(.VSS(VSS),.VDD(VDD),.Y(g4251),.A(I8180));
  NOT NOT1_1637(.VSS(VSS),.VDD(VDD),.Y(g4253),.A(g2734));
  NOT NOT1_1638(.VSS(VSS),.VDD(VDD),.Y(I8190),.A(g3545));
  NOT NOT1_1639(.VSS(VSS),.VDD(VDD),.Y(g4257),.A(I8190));
  NOT NOT1_1640(.VSS(VSS),.VDD(VDD),.Y(I8193),.A(g3547));
  NOT NOT1_1641(.VSS(VSS),.VDD(VDD),.Y(g4258),.A(I8193));
  NOT NOT1_1642(.VSS(VSS),.VDD(VDD),.Y(I8196),.A(g3654));
  NOT NOT1_1643(.VSS(VSS),.VDD(VDD),.Y(g4259),.A(I8196));
  NOT NOT1_1644(.VSS(VSS),.VDD(VDD),.Y(g4265),.A(g3591));
  NOT NOT1_1645(.VSS(VSS),.VDD(VDD),.Y(I8202),.A(g3560));
  NOT NOT1_1646(.VSS(VSS),.VDD(VDD),.Y(g4266),.A(I8202));
  NOT NOT1_1647(.VSS(VSS),.VDD(VDD),.Y(I8205),.A(g2655));
  NOT NOT1_1648(.VSS(VSS),.VDD(VDD),.Y(g4267),.A(I8205));
  NOT NOT1_1649(.VSS(VSS),.VDD(VDD),.Y(g4270),.A(g2573));
  NOT NOT1_1650(.VSS(VSS),.VDD(VDD),.Y(I8215),.A(g3577));
  NOT NOT1_1651(.VSS(VSS),.VDD(VDD),.Y(g4273),.A(I8215));
  NOT NOT1_1652(.VSS(VSS),.VDD(VDD),.Y(I8218),.A(g3002));
  NOT NOT1_1653(.VSS(VSS),.VDD(VDD),.Y(g4274),.A(I8218));
  NOT NOT1_1654(.VSS(VSS),.VDD(VDD),.Y(g4275),.A(g3790));
  NOT NOT1_1655(.VSS(VSS),.VDD(VDD),.Y(g4279),.A(g3340));
  NOT NOT1_1656(.VSS(VSS),.VDD(VDD),.Y(g4281),.A(g2562));
  NOT NOT1_1657(.VSS(VSS),.VDD(VDD),.Y(I8233),.A(g3588));
  NOT NOT1_1658(.VSS(VSS),.VDD(VDD),.Y(g4285),.A(I8233));
  NOT NOT1_1659(.VSS(VSS),.VDD(VDD),.Y(g4286),.A(g3790));
  NOT NOT1_1660(.VSS(VSS),.VDD(VDD),.Y(g4296),.A(g3790));
  NOT NOT1_1661(.VSS(VSS),.VDD(VDD),.Y(I8261),.A(g3643));
  NOT NOT1_1662(.VSS(VSS),.VDD(VDD),.Y(g4300),.A(I8261));
  NOT NOT1_1663(.VSS(VSS),.VDD(VDD),.Y(I8264),.A(g3653));
  NOT NOT1_1664(.VSS(VSS),.VDD(VDD),.Y(g4301),.A(I8264));
  NOT NOT1_1665(.VSS(VSS),.VDD(VDD),.Y(I8268),.A(g2801));
  NOT NOT1_1666(.VSS(VSS),.VDD(VDD),.Y(g4303),.A(I8268));
  NOT NOT1_1667(.VSS(VSS),.VDD(VDD),.Y(I8273),.A(g2976));
  NOT NOT1_1668(.VSS(VSS),.VDD(VDD),.Y(g4306),.A(I8273));
  NOT NOT1_1669(.VSS(VSS),.VDD(VDD),.Y(g4307),.A(g3700));
  NOT NOT1_1670(.VSS(VSS),.VDD(VDD),.Y(I8277),.A(g3504));
  NOT NOT1_1671(.VSS(VSS),.VDD(VDD),.Y(g4308),.A(I8277));
  NOT NOT1_1672(.VSS(VSS),.VDD(VDD),.Y(I8282),.A(g3515));
  NOT NOT1_1673(.VSS(VSS),.VDD(VDD),.Y(g4311),.A(I8282));
  NOT NOT1_1674(.VSS(VSS),.VDD(VDD),.Y(I8291),.A(g878));
  NOT NOT1_1675(.VSS(VSS),.VDD(VDD),.Y(g4316),.A(I8291));
  NOT NOT1_1676(.VSS(VSS),.VDD(VDD),.Y(g4328),.A(g3086));
  NOT NOT1_1677(.VSS(VSS),.VDD(VDD),.Y(g4335),.A(g3659));
  NOT NOT1_1678(.VSS(VSS),.VDD(VDD),.Y(I8308),.A(g3674));
  NOT NOT1_1679(.VSS(VSS),.VDD(VDD),.Y(g4341),.A(I8308));
  NOT NOT1_1680(.VSS(VSS),.VDD(VDD),.Y(g4344),.A(g3124));
  NOT NOT1_1681(.VSS(VSS),.VDD(VDD),.Y(I8315),.A(g3691));
  NOT NOT1_1682(.VSS(VSS),.VDD(VDD),.Y(g4350),.A(I8315));
  NOT NOT1_1683(.VSS(VSS),.VDD(VDD),.Y(g4353),.A(g3665));
  NOT NOT1_1684(.VSS(VSS),.VDD(VDD),.Y(g4357),.A(g3679));
  NOT NOT1_1685(.VSS(VSS),.VDD(VDD),.Y(g4358),.A(g3680));
  NOT NOT1_1686(.VSS(VSS),.VDD(VDD),.Y(I8333),.A(g3721));
  NOT NOT1_1687(.VSS(VSS),.VDD(VDD),.Y(g4360),.A(I8333));
  NOT NOT1_1688(.VSS(VSS),.VDD(VDD),.Y(g4362),.A(g2810));
  NOT NOT1_1689(.VSS(VSS),.VDD(VDD),.Y(I8351),.A(g1160));
  NOT NOT1_1690(.VSS(VSS),.VDD(VDD),.Y(g4370),.A(I8351));
  NOT NOT1_1691(.VSS(VSS),.VDD(VDD),.Y(I8354),.A(g1163));
  NOT NOT1_1692(.VSS(VSS),.VDD(VDD),.Y(g4371),.A(I8354));
  NOT NOT1_1693(.VSS(VSS),.VDD(VDD),.Y(I8357),.A(g1182));
  NOT NOT1_1694(.VSS(VSS),.VDD(VDD),.Y(g4372),.A(I8357));
  NOT NOT1_1695(.VSS(VSS),.VDD(VDD),.Y(I8360),.A(g1186));
  NOT NOT1_1696(.VSS(VSS),.VDD(VDD),.Y(g4373),.A(I8360));
  NOT NOT1_1697(.VSS(VSS),.VDD(VDD),.Y(g4381),.A(g3466));
  NOT NOT1_1698(.VSS(VSS),.VDD(VDD),.Y(I8373),.A(g3783));
  NOT NOT1_1699(.VSS(VSS),.VDD(VDD),.Y(g4382),.A(I8373));
  NOT NOT1_1700(.VSS(VSS),.VDD(VDD),.Y(I8428),.A(g3611));
  NOT NOT1_1701(.VSS(VSS),.VDD(VDD),.Y(g4426),.A(I8428));
  NOT NOT1_1702(.VSS(VSS),.VDD(VDD),.Y(I8446),.A(g3014));
  NOT NOT1_1703(.VSS(VSS),.VDD(VDD),.Y(g4438),.A(I8446));
  NOT NOT1_1704(.VSS(VSS),.VDD(VDD),.Y(I8449),.A(g3630));
  NOT NOT1_1705(.VSS(VSS),.VDD(VDD),.Y(g4443),.A(I8449));
  NOT NOT1_1706(.VSS(VSS),.VDD(VDD),.Y(I8452),.A(g2816));
  NOT NOT1_1707(.VSS(VSS),.VDD(VDD),.Y(g4444),.A(I8452));
  NOT NOT1_1708(.VSS(VSS),.VDD(VDD),.Y(g4455),.A(g3811));
  NOT NOT1_1709(.VSS(VSS),.VDD(VDD),.Y(I8477),.A(g3014));
  NOT NOT1_1710(.VSS(VSS),.VDD(VDD),.Y(g4457),.A(I8477));
  NOT NOT1_1711(.VSS(VSS),.VDD(VDD),.Y(I8480),.A(g3640));
  NOT NOT1_1712(.VSS(VSS),.VDD(VDD),.Y(g4462),.A(I8480));
  NOT NOT1_1713(.VSS(VSS),.VDD(VDD),.Y(I8483),.A(g3641));
  NOT NOT1_1714(.VSS(VSS),.VDD(VDD),.Y(g4463),.A(I8483));
  NOT NOT1_1715(.VSS(VSS),.VDD(VDD),.Y(I8486),.A(g2824));
  NOT NOT1_1716(.VSS(VSS),.VDD(VDD),.Y(g4464),.A(I8486));
  NOT NOT1_1717(.VSS(VSS),.VDD(VDD),.Y(g4465),.A(g3677));
  NOT NOT1_1718(.VSS(VSS),.VDD(VDD),.Y(g4475),.A(g3818));
  NOT NOT1_1719(.VSS(VSS),.VDD(VDD),.Y(I8517),.A(g3014));
  NOT NOT1_1720(.VSS(VSS),.VDD(VDD),.Y(g4477),.A(I8517));
  NOT NOT1_1721(.VSS(VSS),.VDD(VDD),.Y(I8520),.A(g3652));
  NOT NOT1_1722(.VSS(VSS),.VDD(VDD),.Y(g4482),.A(I8520));
  NOT NOT1_1723(.VSS(VSS),.VDD(VDD),.Y(g4489),.A(g2826));
  NOT NOT1_1724(.VSS(VSS),.VDD(VDD),.Y(I8543),.A(g2810));
  NOT NOT1_1725(.VSS(VSS),.VDD(VDD),.Y(g4493),.A(I8543));
  NOT NOT1_1726(.VSS(VSS),.VDD(VDD),.Y(g4500),.A(g2832));
  NOT NOT1_1727(.VSS(VSS),.VDD(VDD),.Y(g4501),.A(g2801));
  NOT NOT1_1728(.VSS(VSS),.VDD(VDD),.Y(I8565),.A(g3071));
  NOT NOT1_1729(.VSS(VSS),.VDD(VDD),.Y(g4503),.A(I8565));
  NOT NOT1_1730(.VSS(VSS),.VDD(VDD),.Y(g4510),.A(g2840));
  NOT NOT1_1731(.VSS(VSS),.VDD(VDD),.Y(g4511),.A(g2841));
  NOT NOT1_1732(.VSS(VSS),.VDD(VDD),.Y(g4512),.A(g2842));
  NOT NOT1_1733(.VSS(VSS),.VDD(VDD),.Y(g4521),.A(g2866));
  NOT NOT1_1734(.VSS(VSS),.VDD(VDD),.Y(g4522),.A(g2867));
  NOT NOT1_1735(.VSS(VSS),.VDD(VDD),.Y(g4523),.A(g2868));
  NOT NOT1_1736(.VSS(VSS),.VDD(VDD),.Y(g4524),.A(g2869));
  NOT NOT1_1737(.VSS(VSS),.VDD(VDD),.Y(g4525),.A(g2870));
  NOT NOT1_1738(.VSS(VSS),.VDD(VDD),.Y(g4527),.A(g3466));
  NOT NOT1_1739(.VSS(VSS),.VDD(VDD),.Y(g4535),.A(g2876));
  NOT NOT1_1740(.VSS(VSS),.VDD(VDD),.Y(g4536),.A(g2877));
  NOT NOT1_1741(.VSS(VSS),.VDD(VDD),.Y(g4537),.A(g2878));
  NOT NOT1_1742(.VSS(VSS),.VDD(VDD),.Y(g4538),.A(g2880));
  NOT NOT1_1743(.VSS(VSS),.VDD(VDD),.Y(g4539),.A(g2881));
  NOT NOT1_1744(.VSS(VSS),.VDD(VDD),.Y(g4540),.A(g2882));
  NOT NOT1_1745(.VSS(VSS),.VDD(VDD),.Y(g4541),.A(g2883));
  NOT NOT1_1746(.VSS(VSS),.VDD(VDD),.Y(g4542),.A(g2884));
  NOT NOT1_1747(.VSS(VSS),.VDD(VDD),.Y(g4543),.A(g2885));
  NOT NOT1_1748(.VSS(VSS),.VDD(VDD),.Y(g4544),.A(g2886));
  NOT NOT1_1749(.VSS(VSS),.VDD(VDD),.Y(g4545),.A(g2887));
  NOT NOT1_1750(.VSS(VSS),.VDD(VDD),.Y(g4547),.A(g3466));
  NOT NOT1_1751(.VSS(VSS),.VDD(VDD),.Y(g4552),.A(g2890));
  NOT NOT1_1752(.VSS(VSS),.VDD(VDD),.Y(g4553),.A(g2891));
  NOT NOT1_1753(.VSS(VSS),.VDD(VDD),.Y(g4554),.A(g2892));
  NOT NOT1_1754(.VSS(VSS),.VDD(VDD),.Y(g4555),.A(g2894));
  NOT NOT1_1755(.VSS(VSS),.VDD(VDD),.Y(g4556),.A(g2895));
  NOT NOT1_1756(.VSS(VSS),.VDD(VDD),.Y(g4557),.A(g2896));
  NOT NOT1_1757(.VSS(VSS),.VDD(VDD),.Y(g4558),.A(g2897));
  NOT NOT1_1758(.VSS(VSS),.VDD(VDD),.Y(g4559),.A(g2898));
  NOT NOT1_1759(.VSS(VSS),.VDD(VDD),.Y(g4560),.A(g2899));
  NOT NOT1_1760(.VSS(VSS),.VDD(VDD),.Y(g4561),.A(g2900));
  NOT NOT1_1761(.VSS(VSS),.VDD(VDD),.Y(g4562),.A(g3466));
  NOT NOT1_1762(.VSS(VSS),.VDD(VDD),.Y(I8665),.A(g3051));
  NOT NOT1_1763(.VSS(VSS),.VDD(VDD),.Y(g4564),.A(I8665));
  NOT NOT1_1764(.VSS(VSS),.VDD(VDD),.Y(g4565),.A(g2901));
  NOT NOT1_1765(.VSS(VSS),.VDD(VDD),.Y(g4566),.A(g2902));
  NOT NOT1_1766(.VSS(VSS),.VDD(VDD),.Y(g4567),.A(g2903));
  NOT NOT1_1767(.VSS(VSS),.VDD(VDD),.Y(g4568),.A(g2904));
  NOT NOT1_1768(.VSS(VSS),.VDD(VDD),.Y(g4569),.A(g2906));
  NOT NOT1_1769(.VSS(VSS),.VDD(VDD),.Y(g4570),.A(g2907));
  NOT NOT1_1770(.VSS(VSS),.VDD(VDD),.Y(g4571),.A(g2908));
  NOT NOT1_1771(.VSS(VSS),.VDD(VDD),.Y(g4572),.A(g2909));
  NOT NOT1_1772(.VSS(VSS),.VDD(VDD),.Y(g4573),.A(g2911));
  NOT NOT1_1773(.VSS(VSS),.VDD(VDD),.Y(g4574),.A(g3466));
  NOT NOT1_1774(.VSS(VSS),.VDD(VDD),.Y(g4576),.A(g2913));
  NOT NOT1_1775(.VSS(VSS),.VDD(VDD),.Y(g4577),.A(g2914));
  NOT NOT1_1776(.VSS(VSS),.VDD(VDD),.Y(g4578),.A(g2917));
  NOT NOT1_1777(.VSS(VSS),.VDD(VDD),.Y(g4579),.A(g2918));
  NOT NOT1_1778(.VSS(VSS),.VDD(VDD),.Y(g4580),.A(g2919));
  NOT NOT1_1779(.VSS(VSS),.VDD(VDD),.Y(g4581),.A(g2921));
  NOT NOT1_1780(.VSS(VSS),.VDD(VDD),.Y(g4582),.A(g2922));
  NOT NOT1_1781(.VSS(VSS),.VDD(VDD),.Y(g4583),.A(g2924));
  NOT NOT1_1782(.VSS(VSS),.VDD(VDD),.Y(g4584),.A(g3466));
  NOT NOT1_1783(.VSS(VSS),.VDD(VDD),.Y(g4585),.A(g2925));
  NOT NOT1_1784(.VSS(VSS),.VDD(VDD),.Y(g4586),.A(g2926));
  NOT NOT1_1785(.VSS(VSS),.VDD(VDD),.Y(g4587),.A(g2928));
  NOT NOT1_1786(.VSS(VSS),.VDD(VDD),.Y(g4588),.A(g2929));
  NOT NOT1_1787(.VSS(VSS),.VDD(VDD),.Y(g4589),.A(g2930));
  NOT NOT1_1788(.VSS(VSS),.VDD(VDD),.Y(g4590),.A(g2932));
  NOT NOT1_1789(.VSS(VSS),.VDD(VDD),.Y(g4591),.A(g2937));
  NOT NOT1_1790(.VSS(VSS),.VDD(VDD),.Y(g4592),.A(g2938));
  NOT NOT1_1791(.VSS(VSS),.VDD(VDD),.Y(g4593),.A(g2939));
  NOT NOT1_1792(.VSS(VSS),.VDD(VDD),.Y(g4594),.A(g2941));
  NOT NOT1_1793(.VSS(VSS),.VDD(VDD),.Y(g4595),.A(g2942));
  NOT NOT1_1794(.VSS(VSS),.VDD(VDD),.Y(g4596),.A(g3466));
  NOT NOT1_1795(.VSS(VSS),.VDD(VDD),.Y(I8706),.A(g3828));
  NOT NOT1_1796(.VSS(VSS),.VDD(VDD),.Y(g4597),.A(I8706));
  NOT NOT1_1797(.VSS(VSS),.VDD(VDD),.Y(I8709),.A(g4191));
  NOT NOT1_1798(.VSS(VSS),.VDD(VDD),.Y(g4598),.A(I8709));
  NOT NOT1_1799(.VSS(VSS),.VDD(VDD),.Y(I8712),.A(g4007));
  NOT NOT1_1800(.VSS(VSS),.VDD(VDD),.Y(g4599),.A(I8712));
  NOT NOT1_1801(.VSS(VSS),.VDD(VDD),.Y(I8715),.A(g3903));
  NOT NOT1_1802(.VSS(VSS),.VDD(VDD),.Y(g4600),.A(I8715));
  NOT NOT1_1803(.VSS(VSS),.VDD(VDD),.Y(I8718),.A(g3909));
  NOT NOT1_1804(.VSS(VSS),.VDD(VDD),.Y(g4601),.A(I8718));
  NOT NOT1_1805(.VSS(VSS),.VDD(VDD),.Y(I8721),.A(g3918));
  NOT NOT1_1806(.VSS(VSS),.VDD(VDD),.Y(g4602),.A(I8721));
  NOT NOT1_1807(.VSS(VSS),.VDD(VDD),.Y(I8724),.A(g3927));
  NOT NOT1_1808(.VSS(VSS),.VDD(VDD),.Y(g4603),.A(I8724));
  NOT NOT1_1809(.VSS(VSS),.VDD(VDD),.Y(I8727),.A(g3944));
  NOT NOT1_1810(.VSS(VSS),.VDD(VDD),.Y(g4604),.A(I8727));
  NOT NOT1_1811(.VSS(VSS),.VDD(VDD),.Y(I8730),.A(g3987));
  NOT NOT1_1812(.VSS(VSS),.VDD(VDD),.Y(g4605),.A(I8730));
  NOT NOT1_1813(.VSS(VSS),.VDD(VDD),.Y(I8733),.A(g3996));
  NOT NOT1_1814(.VSS(VSS),.VDD(VDD),.Y(g4606),.A(I8733));
  NOT NOT1_1815(.VSS(VSS),.VDD(VDD),.Y(I8736),.A(g4008));
  NOT NOT1_1816(.VSS(VSS),.VDD(VDD),.Y(g4607),.A(I8736));
  NOT NOT1_1817(.VSS(VSS),.VDD(VDD),.Y(I8739),.A(g3910));
  NOT NOT1_1818(.VSS(VSS),.VDD(VDD),.Y(g4608),.A(I8739));
  NOT NOT1_1819(.VSS(VSS),.VDD(VDD),.Y(I8742),.A(g3919));
  NOT NOT1_1820(.VSS(VSS),.VDD(VDD),.Y(g4609),.A(I8742));
  NOT NOT1_1821(.VSS(VSS),.VDD(VDD),.Y(I8745),.A(g3929));
  NOT NOT1_1822(.VSS(VSS),.VDD(VDD),.Y(g4610),.A(I8745));
  NOT NOT1_1823(.VSS(VSS),.VDD(VDD),.Y(I8748),.A(g3997));
  NOT NOT1_1824(.VSS(VSS),.VDD(VDD),.Y(g4611),.A(I8748));
  NOT NOT1_1825(.VSS(VSS),.VDD(VDD),.Y(I8751),.A(g4009));
  NOT NOT1_1826(.VSS(VSS),.VDD(VDD),.Y(g4612),.A(I8751));
  NOT NOT1_1827(.VSS(VSS),.VDD(VDD),.Y(I8754),.A(g3911));
  NOT NOT1_1828(.VSS(VSS),.VDD(VDD),.Y(g4613),.A(I8754));
  NOT NOT1_1829(.VSS(VSS),.VDD(VDD),.Y(I8757),.A(g3921));
  NOT NOT1_1830(.VSS(VSS),.VDD(VDD),.Y(g4614),.A(I8757));
  NOT NOT1_1831(.VSS(VSS),.VDD(VDD),.Y(I8760),.A(g3931));
  NOT NOT1_1832(.VSS(VSS),.VDD(VDD),.Y(g4615),.A(I8760));
  NOT NOT1_1833(.VSS(VSS),.VDD(VDD),.Y(I8763),.A(g3947));
  NOT NOT1_1834(.VSS(VSS),.VDD(VDD),.Y(g4616),.A(I8763));
  NOT NOT1_1835(.VSS(VSS),.VDD(VDD),.Y(I8766),.A(g3960));
  NOT NOT1_1836(.VSS(VSS),.VDD(VDD),.Y(g4617),.A(I8766));
  NOT NOT1_1837(.VSS(VSS),.VDD(VDD),.Y(I8769),.A(g3999));
  NOT NOT1_1838(.VSS(VSS),.VDD(VDD),.Y(g4618),.A(I8769));
  NOT NOT1_1839(.VSS(VSS),.VDD(VDD),.Y(I8772),.A(g4011));
  NOT NOT1_1840(.VSS(VSS),.VDD(VDD),.Y(g4619),.A(I8772));
  NOT NOT1_1841(.VSS(VSS),.VDD(VDD),.Y(I8775),.A(g4019));
  NOT NOT1_1842(.VSS(VSS),.VDD(VDD),.Y(g4620),.A(I8775));
  NOT NOT1_1843(.VSS(VSS),.VDD(VDD),.Y(I8778),.A(g3922));
  NOT NOT1_1844(.VSS(VSS),.VDD(VDD),.Y(g4621),.A(I8778));
  NOT NOT1_1845(.VSS(VSS),.VDD(VDD),.Y(I8781),.A(g3932));
  NOT NOT1_1846(.VSS(VSS),.VDD(VDD),.Y(g4622),.A(I8781));
  NOT NOT1_1847(.VSS(VSS),.VDD(VDD),.Y(I8784),.A(g3949));
  NOT NOT1_1848(.VSS(VSS),.VDD(VDD),.Y(g4623),.A(I8784));
  NOT NOT1_1849(.VSS(VSS),.VDD(VDD),.Y(I8787),.A(g4012));
  NOT NOT1_1850(.VSS(VSS),.VDD(VDD),.Y(g4624),.A(I8787));
  NOT NOT1_1851(.VSS(VSS),.VDD(VDD),.Y(I8790),.A(g4020));
  NOT NOT1_1852(.VSS(VSS),.VDD(VDD),.Y(g4625),.A(I8790));
  NOT NOT1_1853(.VSS(VSS),.VDD(VDD),.Y(I8793),.A(g3923));
  NOT NOT1_1854(.VSS(VSS),.VDD(VDD),.Y(g4626),.A(I8793));
  NOT NOT1_1855(.VSS(VSS),.VDD(VDD),.Y(I8796),.A(g3934));
  NOT NOT1_1856(.VSS(VSS),.VDD(VDD),.Y(g4627),.A(I8796));
  NOT NOT1_1857(.VSS(VSS),.VDD(VDD),.Y(I8799),.A(g3951));
  NOT NOT1_1858(.VSS(VSS),.VDD(VDD),.Y(g4628),.A(I8799));
  NOT NOT1_1859(.VSS(VSS),.VDD(VDD),.Y(I8802),.A(g3963));
  NOT NOT1_1860(.VSS(VSS),.VDD(VDD),.Y(g4629),.A(I8802));
  NOT NOT1_1861(.VSS(VSS),.VDD(VDD),.Y(I8805),.A(g3976));
  NOT NOT1_1862(.VSS(VSS),.VDD(VDD),.Y(g4630),.A(I8805));
  NOT NOT1_1863(.VSS(VSS),.VDD(VDD),.Y(I8808),.A(g4014));
  NOT NOT1_1864(.VSS(VSS),.VDD(VDD),.Y(g4631),.A(I8808));
  NOT NOT1_1865(.VSS(VSS),.VDD(VDD),.Y(I8811),.A(g4022));
  NOT NOT1_1866(.VSS(VSS),.VDD(VDD),.Y(g4632),.A(I8811));
  NOT NOT1_1867(.VSS(VSS),.VDD(VDD),.Y(I8814),.A(g4028));
  NOT NOT1_1868(.VSS(VSS),.VDD(VDD),.Y(g4633),.A(I8814));
  NOT NOT1_1869(.VSS(VSS),.VDD(VDD),.Y(I8817),.A(g3935));
  NOT NOT1_1870(.VSS(VSS),.VDD(VDD),.Y(g4634),.A(I8817));
  NOT NOT1_1871(.VSS(VSS),.VDD(VDD),.Y(I8820),.A(g3952));
  NOT NOT1_1872(.VSS(VSS),.VDD(VDD),.Y(g4635),.A(I8820));
  NOT NOT1_1873(.VSS(VSS),.VDD(VDD),.Y(I8823),.A(g3965));
  NOT NOT1_1874(.VSS(VSS),.VDD(VDD),.Y(g4636),.A(I8823));
  NOT NOT1_1875(.VSS(VSS),.VDD(VDD),.Y(I8826),.A(g4023));
  NOT NOT1_1876(.VSS(VSS),.VDD(VDD),.Y(g4637),.A(I8826));
  NOT NOT1_1877(.VSS(VSS),.VDD(VDD),.Y(I8829),.A(g4029));
  NOT NOT1_1878(.VSS(VSS),.VDD(VDD),.Y(g4638),.A(I8829));
  NOT NOT1_1879(.VSS(VSS),.VDD(VDD),.Y(I8832),.A(g3936));
  NOT NOT1_1880(.VSS(VSS),.VDD(VDD),.Y(g4639),.A(I8832));
  NOT NOT1_1881(.VSS(VSS),.VDD(VDD),.Y(I8835),.A(g3954));
  NOT NOT1_1882(.VSS(VSS),.VDD(VDD),.Y(g4640),.A(I8835));
  NOT NOT1_1883(.VSS(VSS),.VDD(VDD),.Y(I8838),.A(g3967));
  NOT NOT1_1884(.VSS(VSS),.VDD(VDD),.Y(g4641),.A(I8838));
  NOT NOT1_1885(.VSS(VSS),.VDD(VDD),.Y(I8841),.A(g3979));
  NOT NOT1_1886(.VSS(VSS),.VDD(VDD),.Y(g4642),.A(I8841));
  NOT NOT1_1887(.VSS(VSS),.VDD(VDD),.Y(I8844),.A(g3992));
  NOT NOT1_1888(.VSS(VSS),.VDD(VDD),.Y(g4643),.A(I8844));
  NOT NOT1_1889(.VSS(VSS),.VDD(VDD),.Y(I8847),.A(g4025));
  NOT NOT1_1890(.VSS(VSS),.VDD(VDD),.Y(g4644),.A(I8847));
  NOT NOT1_1891(.VSS(VSS),.VDD(VDD),.Y(I8850),.A(g4031));
  NOT NOT1_1892(.VSS(VSS),.VDD(VDD),.Y(g4645),.A(I8850));
  NOT NOT1_1893(.VSS(VSS),.VDD(VDD),.Y(I8853),.A(g4034));
  NOT NOT1_1894(.VSS(VSS),.VDD(VDD),.Y(g4646),.A(I8853));
  NOT NOT1_1895(.VSS(VSS),.VDD(VDD),.Y(I8856),.A(g3955));
  NOT NOT1_1896(.VSS(VSS),.VDD(VDD),.Y(g4647),.A(I8856));
  NOT NOT1_1897(.VSS(VSS),.VDD(VDD),.Y(I8859),.A(g3968));
  NOT NOT1_1898(.VSS(VSS),.VDD(VDD),.Y(g4648),.A(I8859));
  NOT NOT1_1899(.VSS(VSS),.VDD(VDD),.Y(I8862),.A(g3981));
  NOT NOT1_1900(.VSS(VSS),.VDD(VDD),.Y(g4649),.A(I8862));
  NOT NOT1_1901(.VSS(VSS),.VDD(VDD),.Y(I8865),.A(g4032));
  NOT NOT1_1902(.VSS(VSS),.VDD(VDD),.Y(g4650),.A(I8865));
  NOT NOT1_1903(.VSS(VSS),.VDD(VDD),.Y(I8868),.A(g4035));
  NOT NOT1_1904(.VSS(VSS),.VDD(VDD),.Y(g4651),.A(I8868));
  NOT NOT1_1905(.VSS(VSS),.VDD(VDD),.Y(I8871),.A(g3869));
  NOT NOT1_1906(.VSS(VSS),.VDD(VDD),.Y(g4652),.A(I8871));
  NOT NOT1_1907(.VSS(VSS),.VDD(VDD),.Y(I8874),.A(g3884));
  NOT NOT1_1908(.VSS(VSS),.VDD(VDD),.Y(g4653),.A(I8874));
  NOT NOT1_1909(.VSS(VSS),.VDD(VDD),.Y(I8877),.A(g4274));
  NOT NOT1_1910(.VSS(VSS),.VDD(VDD),.Y(g4654),.A(I8877));
  NOT NOT1_1911(.VSS(VSS),.VDD(VDD),.Y(I8880),.A(g4303));
  NOT NOT1_1912(.VSS(VSS),.VDD(VDD),.Y(g4655),.A(I8880));
  NOT NOT1_1913(.VSS(VSS),.VDD(VDD),.Y(I8883),.A(g4198));
  NOT NOT1_1914(.VSS(VSS),.VDD(VDD),.Y(g4656),.A(I8883));
  NOT NOT1_1915(.VSS(VSS),.VDD(VDD),.Y(I8886),.A(g4308));
  NOT NOT1_1916(.VSS(VSS),.VDD(VDD),.Y(g4657),.A(I8886));
  NOT NOT1_1917(.VSS(VSS),.VDD(VDD),.Y(I8889),.A(g4311));
  NOT NOT1_1918(.VSS(VSS),.VDD(VDD),.Y(g4658),.A(I8889));
  NOT NOT1_1919(.VSS(VSS),.VDD(VDD),.Y(I8892),.A(g4115));
  NOT NOT1_1920(.VSS(VSS),.VDD(VDD),.Y(g4659),.A(I8892));
  NOT NOT1_1921(.VSS(VSS),.VDD(VDD),.Y(I8895),.A(g4130));
  NOT NOT1_1922(.VSS(VSS),.VDD(VDD),.Y(g4660),.A(I8895));
  NOT NOT1_1923(.VSS(VSS),.VDD(VDD),.Y(I8898),.A(g4089));
  NOT NOT1_1924(.VSS(VSS),.VDD(VDD),.Y(g4661),.A(I8898));
  NOT NOT1_1925(.VSS(VSS),.VDD(VDD),.Y(I8901),.A(g4122));
  NOT NOT1_1926(.VSS(VSS),.VDD(VDD),.Y(g4662),.A(I8901));
  NOT NOT1_1927(.VSS(VSS),.VDD(VDD),.Y(I8904),.A(g4126));
  NOT NOT1_1928(.VSS(VSS),.VDD(VDD),.Y(g4663),.A(I8904));
  NOT NOT1_1929(.VSS(VSS),.VDD(VDD),.Y(I8907),.A(g4095));
  NOT NOT1_1930(.VSS(VSS),.VDD(VDD),.Y(g4664),.A(I8907));
  NOT NOT1_1931(.VSS(VSS),.VDD(VDD),.Y(I8910),.A(g4200));
  NOT NOT1_1932(.VSS(VSS),.VDD(VDD),.Y(g4665),.A(I8910));
  NOT NOT1_1933(.VSS(VSS),.VDD(VDD),.Y(I8913),.A(g4306));
  NOT NOT1_1934(.VSS(VSS),.VDD(VDD),.Y(g4666),.A(I8913));
  NOT NOT1_1935(.VSS(VSS),.VDD(VDD),.Y(I8916),.A(g4195));
  NOT NOT1_1936(.VSS(VSS),.VDD(VDD),.Y(g4667),.A(I8916));
  NOT NOT1_1937(.VSS(VSS),.VDD(VDD),.Y(I8919),.A(g4196));
  NOT NOT1_1938(.VSS(VSS),.VDD(VDD),.Y(g4668),.A(I8919));
  NOT NOT1_1939(.VSS(VSS),.VDD(VDD),.Y(I8922),.A(g4229));
  NOT NOT1_1940(.VSS(VSS),.VDD(VDD),.Y(g4669),.A(I8922));
  NOT NOT1_1941(.VSS(VSS),.VDD(VDD),.Y(I8925),.A(g4482));
  NOT NOT1_1942(.VSS(VSS),.VDD(VDD),.Y(g4670),.A(I8925));
  NOT NOT1_1943(.VSS(VSS),.VDD(VDD),.Y(I8928),.A(g4153));
  NOT NOT1_1944(.VSS(VSS),.VDD(VDD),.Y(g4673),.A(I8928));
  NOT NOT1_1945(.VSS(VSS),.VDD(VDD),.Y(I8932),.A(g4096));
  NOT NOT1_1946(.VSS(VSS),.VDD(VDD),.Y(g4677),.A(I8932));
  NOT NOT1_1947(.VSS(VSS),.VDD(VDD),.Y(I8935),.A(g4005));
  NOT NOT1_1948(.VSS(VSS),.VDD(VDD),.Y(g4678),.A(I8935));
  NOT NOT1_1949(.VSS(VSS),.VDD(VDD),.Y(I8945),.A(g4106));
  NOT NOT1_1950(.VSS(VSS),.VDD(VDD),.Y(g4680),.A(I8945));
  NOT NOT1_1951(.VSS(VSS),.VDD(VDD),.Y(I8949),.A(g4116));
  NOT NOT1_1952(.VSS(VSS),.VDD(VDD),.Y(g4684),.A(I8949));
  NOT NOT1_1953(.VSS(VSS),.VDD(VDD),.Y(I8952),.A(g4197));
  NOT NOT1_1954(.VSS(VSS),.VDD(VDD),.Y(g4685),.A(I8952));
  NOT NOT1_1955(.VSS(VSS),.VDD(VDD),.Y(I8962),.A(g4553));
  NOT NOT1_1956(.VSS(VSS),.VDD(VDD),.Y(g4687),.A(I8962));
  NOT NOT1_1957(.VSS(VSS),.VDD(VDD),.Y(I8966),.A(g4444));
  NOT NOT1_1958(.VSS(VSS),.VDD(VDD),.Y(g4689),.A(I8966));
  NOT NOT1_1959(.VSS(VSS),.VDD(VDD),.Y(I8971),.A(g4464));
  NOT NOT1_1960(.VSS(VSS),.VDD(VDD),.Y(g4692),.A(I8971));
  NOT NOT1_1961(.VSS(VSS),.VDD(VDD),.Y(I8974),.A(g3871));
  NOT NOT1_1962(.VSS(VSS),.VDD(VDD),.Y(g4693),.A(I8974));
  NOT NOT1_1963(.VSS(VSS),.VDD(VDD),.Y(I8977),.A(g3877));
  NOT NOT1_1964(.VSS(VSS),.VDD(VDD),.Y(g4694),.A(I8977));
  NOT NOT1_1965(.VSS(VSS),.VDD(VDD),.Y(I8980),.A(g4535));
  NOT NOT1_1966(.VSS(VSS),.VDD(VDD),.Y(g4695),.A(I8980));
  NOT NOT1_1967(.VSS(VSS),.VDD(VDD),.Y(I8983),.A(g4536));
  NOT NOT1_1968(.VSS(VSS),.VDD(VDD),.Y(g4696),.A(I8983));
  NOT NOT1_1969(.VSS(VSS),.VDD(VDD),.Y(I8986),.A(g4552));
  NOT NOT1_1970(.VSS(VSS),.VDD(VDD),.Y(g4697),.A(I8986));
  NOT NOT1_1971(.VSS(VSS),.VDD(VDD),.Y(I8989),.A(g4537));
  NOT NOT1_1972(.VSS(VSS),.VDD(VDD),.Y(g4698),.A(I8989));
  NOT NOT1_1973(.VSS(VSS),.VDD(VDD),.Y(I8994),.A(g4565));
  NOT NOT1_1974(.VSS(VSS),.VDD(VDD),.Y(g4701),.A(I8994));
  NOT NOT1_1975(.VSS(VSS),.VDD(VDD),.Y(I8998),.A(g4576));
  NOT NOT1_1976(.VSS(VSS),.VDD(VDD),.Y(g4703),.A(I8998));
  NOT NOT1_1977(.VSS(VSS),.VDD(VDD),.Y(I9001),.A(g4577));
  NOT NOT1_1978(.VSS(VSS),.VDD(VDD),.Y(g4704),.A(I9001));
  NOT NOT1_1979(.VSS(VSS),.VDD(VDD),.Y(I9005),.A(g4585));
  NOT NOT1_1980(.VSS(VSS),.VDD(VDD),.Y(g4706),.A(I9005));
  NOT NOT1_1981(.VSS(VSS),.VDD(VDD),.Y(I9009),.A(g4591));
  NOT NOT1_1982(.VSS(VSS),.VDD(VDD),.Y(g4710),.A(I9009));
  NOT NOT1_1983(.VSS(VSS),.VDD(VDD),.Y(I9014),.A(g3864));
  NOT NOT1_1984(.VSS(VSS),.VDD(VDD),.Y(g4713),.A(I9014));
  NOT NOT1_1985(.VSS(VSS),.VDD(VDD),.Y(I9018),.A(g3872));
  NOT NOT1_1986(.VSS(VSS),.VDD(VDD),.Y(g4718),.A(I9018));
  NOT NOT1_1987(.VSS(VSS),.VDD(VDD),.Y(I9021),.A(g4489));
  NOT NOT1_1988(.VSS(VSS),.VDD(VDD),.Y(g4719),.A(I9021));
  NOT NOT1_1989(.VSS(VSS),.VDD(VDD),.Y(I9025),.A(g4462));
  NOT NOT1_1990(.VSS(VSS),.VDD(VDD),.Y(g4721),.A(I9025));
  NOT NOT1_1991(.VSS(VSS),.VDD(VDD),.Y(I9034),.A(g4317));
  NOT NOT1_1992(.VSS(VSS),.VDD(VDD),.Y(g4732),.A(I9034));
  NOT NOT1_1993(.VSS(VSS),.VDD(VDD),.Y(g4733),.A(g4202));
  NOT NOT1_1994(.VSS(VSS),.VDD(VDD),.Y(I9050),.A(g3881));
  NOT NOT1_1995(.VSS(VSS),.VDD(VDD),.Y(g4738),.A(I9050));
  NOT NOT1_1996(.VSS(VSS),.VDD(VDD),.Y(I9053),.A(g4327));
  NOT NOT1_1997(.VSS(VSS),.VDD(VDD),.Y(g4739),.A(I9053));
  NOT NOT1_1998(.VSS(VSS),.VDD(VDD),.Y(I9064),.A(g4302));
  NOT NOT1_1999(.VSS(VSS),.VDD(VDD),.Y(g4742),.A(I9064));
  NOT NOT1_2000(.VSS(VSS),.VDD(VDD),.Y(I9076),.A(g4353));
  NOT NOT1_2001(.VSS(VSS),.VDD(VDD),.Y(g4746),.A(I9076));
  NOT NOT1_2002(.VSS(VSS),.VDD(VDD),.Y(g4748),.A(g4465));
  NOT NOT1_2003(.VSS(VSS),.VDD(VDD),.Y(I9081),.A(g4357));
  NOT NOT1_2004(.VSS(VSS),.VDD(VDD),.Y(g4776),.A(I9081));
  NOT NOT1_2005(.VSS(VSS),.VDD(VDD),.Y(I9084),.A(g4358));
  NOT NOT1_2006(.VSS(VSS),.VDD(VDD),.Y(g4777),.A(I9084));
  NOT NOT1_2007(.VSS(VSS),.VDD(VDD),.Y(I9089),.A(g4566));
  NOT NOT1_2008(.VSS(VSS),.VDD(VDD),.Y(g4780),.A(I9089));
  NOT NOT1_2009(.VSS(VSS),.VDD(VDD),.Y(I9095),.A(g4283));
  NOT NOT1_2010(.VSS(VSS),.VDD(VDD),.Y(g4784),.A(I9095));
  NOT NOT1_2011(.VSS(VSS),.VDD(VDD),.Y(I9103),.A(g4374));
  NOT NOT1_2012(.VSS(VSS),.VDD(VDD),.Y(g4788),.A(I9103));
  NOT NOT1_2013(.VSS(VSS),.VDD(VDD),.Y(I9111),.A(g4232));
  NOT NOT1_2014(.VSS(VSS),.VDD(VDD),.Y(g4792),.A(I9111));
  NOT NOT1_2015(.VSS(VSS),.VDD(VDD),.Y(I9116),.A(g4297));
  NOT NOT1_2016(.VSS(VSS),.VDD(VDD),.Y(g4795),.A(I9116));
  NOT NOT1_2017(.VSS(VSS),.VDD(VDD),.Y(I9123),.A(g4455));
  NOT NOT1_2018(.VSS(VSS),.VDD(VDD),.Y(g4800),.A(I9123));
  NOT NOT1_2019(.VSS(VSS),.VDD(VDD),.Y(I9126),.A(g3870));
  NOT NOT1_2020(.VSS(VSS),.VDD(VDD),.Y(g4801),.A(I9126));
  NOT NOT1_2021(.VSS(VSS),.VDD(VDD),.Y(I9129),.A(g4475));
  NOT NOT1_2022(.VSS(VSS),.VDD(VDD),.Y(g4802),.A(I9129));
  NOT NOT1_2023(.VSS(VSS),.VDD(VDD),.Y(I9132),.A(g4284));
  NOT NOT1_2024(.VSS(VSS),.VDD(VDD),.Y(g4803),.A(I9132));
  NOT NOT1_2025(.VSS(VSS),.VDD(VDD),.Y(I9136),.A(g4280));
  NOT NOT1_2026(.VSS(VSS),.VDD(VDD),.Y(g4805),.A(I9136));
  NOT NOT1_2027(.VSS(VSS),.VDD(VDD),.Y(I9139),.A(g4364));
  NOT NOT1_2028(.VSS(VSS),.VDD(VDD),.Y(g4806),.A(I9139));
  NOT NOT1_2029(.VSS(VSS),.VDD(VDD),.Y(I9142),.A(g4236));
  NOT NOT1_2030(.VSS(VSS),.VDD(VDD),.Y(g4807),.A(I9142));
  NOT NOT1_2031(.VSS(VSS),.VDD(VDD),.Y(I9145),.A(g4264));
  NOT NOT1_2032(.VSS(VSS),.VDD(VDD),.Y(g4808),.A(I9145));
  NOT NOT1_2033(.VSS(VSS),.VDD(VDD),.Y(I9148),.A(g4354));
  NOT NOT1_2034(.VSS(VSS),.VDD(VDD),.Y(g4809),.A(I9148));
  NOT NOT1_2035(.VSS(VSS),.VDD(VDD),.Y(I9158),.A(g4256));
  NOT NOT1_2036(.VSS(VSS),.VDD(VDD),.Y(g4811),.A(I9158));
  NOT NOT1_2037(.VSS(VSS),.VDD(VDD),.Y(I9162),.A(g4272));
  NOT NOT1_2038(.VSS(VSS),.VDD(VDD),.Y(g4813),.A(I9162));
  NOT NOT1_2039(.VSS(VSS),.VDD(VDD),.Y(I9177),.A(g4299));
  NOT NOT1_2040(.VSS(VSS),.VDD(VDD),.Y(g4822),.A(I9177));
  NOT NOT1_2041(.VSS(VSS),.VDD(VDD),.Y(g4841),.A(g4250));
  NOT NOT1_2042(.VSS(VSS),.VDD(VDD),.Y(I9209),.A(g4349));
  NOT NOT1_2043(.VSS(VSS),.VDD(VDD),.Y(g4867),.A(I9209));
  NOT NOT1_2044(.VSS(VSS),.VDD(VDD),.Y(I9217),.A(g4443));
  NOT NOT1_2045(.VSS(VSS),.VDD(VDD),.Y(g4873),.A(I9217));
  NOT NOT1_2046(.VSS(VSS),.VDD(VDD),.Y(g4882),.A(g4069));
  NOT NOT1_2047(.VSS(VSS),.VDD(VDD),.Y(g4885),.A(g4070));
  NOT NOT1_2048(.VSS(VSS),.VDD(VDD),.Y(g4886),.A(g4071));
  NOT NOT1_2049(.VSS(VSS),.VDD(VDD),.Y(g4890),.A(g4075));
  NOT NOT1_2050(.VSS(VSS),.VDD(VDD),.Y(g4891),.A(g4076));
  NOT NOT1_2051(.VSS(VSS),.VDD(VDD),.Y(I9250),.A(g4134));
  NOT NOT1_2052(.VSS(VSS),.VDD(VDD),.Y(g4892),.A(I9250));
  NOT NOT1_2053(.VSS(VSS),.VDD(VDD),.Y(g4895),.A(g4078));
  NOT NOT1_2054(.VSS(VSS),.VDD(VDD),.Y(g4898),.A(g4079));
  NOT NOT1_2055(.VSS(VSS),.VDD(VDD),.Y(g4899),.A(g4080));
  NOT NOT1_2056(.VSS(VSS),.VDD(VDD),.Y(I9258),.A(g4249));
  NOT NOT1_2057(.VSS(VSS),.VDD(VDD),.Y(g4900),.A(I9258));
  NOT NOT1_2058(.VSS(VSS),.VDD(VDD),.Y(g4903),.A(g4084));
  NOT NOT1_2059(.VSS(VSS),.VDD(VDD),.Y(g4904),.A(g4085));
  NOT NOT1_2060(.VSS(VSS),.VDD(VDD),.Y(g4907),.A(g4087));
  NOT NOT1_2061(.VSS(VSS),.VDD(VDD),.Y(g4908),.A(g4088));
  NOT NOT1_2062(.VSS(VSS),.VDD(VDD),.Y(I9271),.A(g4263));
  NOT NOT1_2063(.VSS(VSS),.VDD(VDD),.Y(g4909),.A(I9271));
  NOT NOT1_2064(.VSS(VSS),.VDD(VDD),.Y(g4913),.A(g4092));
  NOT NOT1_2065(.VSS(VSS),.VDD(VDD),.Y(g4914),.A(g4093));
  NOT NOT1_2066(.VSS(VSS),.VDD(VDD),.Y(g4915),.A(g4094));
  NOT NOT1_2067(.VSS(VSS),.VDD(VDD),.Y(g4916),.A(g4202));
  NOT NOT1_2068(.VSS(VSS),.VDD(VDD),.Y(g4917),.A(g4102));
  NOT NOT1_2069(.VSS(VSS),.VDD(VDD),.Y(g4918),.A(g4103));
  NOT NOT1_2070(.VSS(VSS),.VDD(VDD),.Y(g4919),.A(g4104));
  NOT NOT1_2071(.VSS(VSS),.VDD(VDD),.Y(g4920),.A(g4105));
  NOT NOT1_2072(.VSS(VSS),.VDD(VDD),.Y(g4921),.A(g4202));
  NOT NOT1_2073(.VSS(VSS),.VDD(VDD),.Y(g4922),.A(g4111));
  NOT NOT1_2074(.VSS(VSS),.VDD(VDD),.Y(g4923),.A(g4112));
  NOT NOT1_2075(.VSS(VSS),.VDD(VDD),.Y(g4924),.A(g4113));
  NOT NOT1_2076(.VSS(VSS),.VDD(VDD),.Y(g4925),.A(g4114));
  NOT NOT1_2077(.VSS(VSS),.VDD(VDD),.Y(g4926),.A(g4202));
  NOT NOT1_2078(.VSS(VSS),.VDD(VDD),.Y(g4928),.A(g4119));
  NOT NOT1_2079(.VSS(VSS),.VDD(VDD),.Y(g4929),.A(g4120));
  NOT NOT1_2080(.VSS(VSS),.VDD(VDD),.Y(g4930),.A(g4121));
  NOT NOT1_2081(.VSS(VSS),.VDD(VDD),.Y(I9301),.A(g4295));
  NOT NOT1_2082(.VSS(VSS),.VDD(VDD),.Y(g4931),.A(I9301));
  NOT NOT1_2083(.VSS(VSS),.VDD(VDD),.Y(g4932),.A(g4202));
  NOT NOT1_2084(.VSS(VSS),.VDD(VDD),.Y(g4934),.A(g4125));
  NOT NOT1_2085(.VSS(VSS),.VDD(VDD),.Y(g4935),.A(g4202));
  NOT NOT1_2086(.VSS(VSS),.VDD(VDD),.Y(I9310),.A(g4268));
  NOT NOT1_2087(.VSS(VSS),.VDD(VDD),.Y(g4938),.A(I9310));
  NOT NOT1_2088(.VSS(VSS),.VDD(VDD),.Y(g4960),.A(g4259));
  NOT NOT1_2089(.VSS(VSS),.VDD(VDD),.Y(g4963),.A(g4328));
  NOT NOT1_2090(.VSS(VSS),.VDD(VDD),.Y(I9325),.A(g4242));
  NOT NOT1_2091(.VSS(VSS),.VDD(VDD),.Y(g5000),.A(I9325));
  NOT NOT1_2092(.VSS(VSS),.VDD(VDD),.Y(g5002),.A(g4335));
  NOT NOT1_2093(.VSS(VSS),.VDD(VDD),.Y(I9333),.A(g4245));
  NOT NOT1_2094(.VSS(VSS),.VDD(VDD),.Y(g5006),.A(I9333));
  NOT NOT1_2095(.VSS(VSS),.VDD(VDD),.Y(I9336),.A(g4493));
  NOT NOT1_2096(.VSS(VSS),.VDD(VDD),.Y(g5007),.A(I9336));
  NOT NOT1_2097(.VSS(VSS),.VDD(VDD),.Y(g5009),.A(g4344));
  NOT NOT1_2098(.VSS(VSS),.VDD(VDD),.Y(I9341),.A(g4251));
  NOT NOT1_2099(.VSS(VSS),.VDD(VDD),.Y(g5013),.A(I9341));
  NOT NOT1_2100(.VSS(VSS),.VDD(VDD),.Y(I9344),.A(g4341));
  NOT NOT1_2101(.VSS(VSS),.VDD(VDD),.Y(g5014),.A(I9344));
  NOT NOT1_2102(.VSS(VSS),.VDD(VDD),.Y(I9347),.A(g3896));
  NOT NOT1_2103(.VSS(VSS),.VDD(VDD),.Y(g5015),.A(I9347));
  NOT NOT1_2104(.VSS(VSS),.VDD(VDD),.Y(I9350),.A(g4503));
  NOT NOT1_2105(.VSS(VSS),.VDD(VDD),.Y(g5016),.A(I9350));
  NOT NOT1_2106(.VSS(VSS),.VDD(VDD),.Y(g5022),.A(g4438));
  NOT NOT1_2107(.VSS(VSS),.VDD(VDD),.Y(I9360),.A(g4257));
  NOT NOT1_2108(.VSS(VSS),.VDD(VDD),.Y(g5024),.A(I9360));
  NOT NOT1_2109(.VSS(VSS),.VDD(VDD),.Y(I9363),.A(g4258));
  NOT NOT1_2110(.VSS(VSS),.VDD(VDD),.Y(g5025),.A(I9363));
  NOT NOT1_2111(.VSS(VSS),.VDD(VDD),.Y(I9366),.A(g4350));
  NOT NOT1_2112(.VSS(VSS),.VDD(VDD),.Y(g5026),.A(I9366));
  NOT NOT1_2113(.VSS(VSS),.VDD(VDD),.Y(I9369),.A(g3901));
  NOT NOT1_2114(.VSS(VSS),.VDD(VDD),.Y(g5027),.A(I9369));
  NOT NOT1_2115(.VSS(VSS),.VDD(VDD),.Y(I9372),.A(g3902));
  NOT NOT1_2116(.VSS(VSS),.VDD(VDD),.Y(g5028),.A(I9372));
  NOT NOT1_2117(.VSS(VSS),.VDD(VDD),.Y(g5037),.A(g4438));
  NOT NOT1_2118(.VSS(VSS),.VDD(VDD),.Y(g5038),.A(g4457));
  NOT NOT1_2119(.VSS(VSS),.VDD(VDD),.Y(I9393),.A(g4266));
  NOT NOT1_2120(.VSS(VSS),.VDD(VDD),.Y(g5041),.A(I9393));
  NOT NOT1_2121(.VSS(VSS),.VDD(VDD),.Y(I9396),.A(g3908));
  NOT NOT1_2122(.VSS(VSS),.VDD(VDD),.Y(g5042),.A(I9396));
  NOT NOT1_2123(.VSS(VSS),.VDD(VDD),.Y(I9407),.A(g4232));
  NOT NOT1_2124(.VSS(VSS),.VDD(VDD),.Y(g5051),.A(I9407));
  NOT NOT1_2125(.VSS(VSS),.VDD(VDD),.Y(g5053),.A(g4438));
  NOT NOT1_2126(.VSS(VSS),.VDD(VDD),.Y(g5054),.A(g4457));
  NOT NOT1_2127(.VSS(VSS),.VDD(VDD),.Y(g5055),.A(g4477));
  NOT NOT1_2128(.VSS(VSS),.VDD(VDD),.Y(I9416),.A(g4273));
  NOT NOT1_2129(.VSS(VSS),.VDD(VDD),.Y(g5058),.A(I9416));
  NOT NOT1_2130(.VSS(VSS),.VDD(VDD),.Y(I9419),.A(g3916));
  NOT NOT1_2131(.VSS(VSS),.VDD(VDD),.Y(g5059),.A(I9419));
  NOT NOT1_2132(.VSS(VSS),.VDD(VDD),.Y(I9422),.A(g4360));
  NOT NOT1_2133(.VSS(VSS),.VDD(VDD),.Y(g5060),.A(I9422));
  NOT NOT1_2134(.VSS(VSS),.VDD(VDD),.Y(I9425),.A(g3917));
  NOT NOT1_2135(.VSS(VSS),.VDD(VDD),.Y(g5061),.A(I9425));
  NOT NOT1_2136(.VSS(VSS),.VDD(VDD),.Y(g5071),.A(g4438));
  NOT NOT1_2137(.VSS(VSS),.VDD(VDD),.Y(g5072),.A(g4457));
  NOT NOT1_2138(.VSS(VSS),.VDD(VDD),.Y(g5073),.A(g4477));
  NOT NOT1_2139(.VSS(VSS),.VDD(VDD),.Y(I9440),.A(g4285));
  NOT NOT1_2140(.VSS(VSS),.VDD(VDD),.Y(g5074),.A(I9440));
  NOT NOT1_2141(.VSS(VSS),.VDD(VDD),.Y(I9443),.A(g4564));
  NOT NOT1_2142(.VSS(VSS),.VDD(VDD),.Y(g5075),.A(I9443));
  NOT NOT1_2143(.VSS(VSS),.VDD(VDD),.Y(I9446),.A(g3926));
  NOT NOT1_2144(.VSS(VSS),.VDD(VDD),.Y(g5076),.A(I9446));
  NOT NOT1_2145(.VSS(VSS),.VDD(VDD),.Y(g5083),.A(g4457));
  NOT NOT1_2146(.VSS(VSS),.VDD(VDD),.Y(g5084),.A(g4477));
  NOT NOT1_2147(.VSS(VSS),.VDD(VDD),.Y(I9457),.A(g3940));
  NOT NOT1_2148(.VSS(VSS),.VDD(VDD),.Y(g5085),.A(I9457));
  NOT NOT1_2149(.VSS(VSS),.VDD(VDD),.Y(I9460),.A(g3941));
  NOT NOT1_2150(.VSS(VSS),.VDD(VDD),.Y(g5086),.A(I9460));
  NOT NOT1_2151(.VSS(VSS),.VDD(VDD),.Y(I9463),.A(g3942));
  NOT NOT1_2152(.VSS(VSS),.VDD(VDD),.Y(g5087),.A(I9463));
  NOT NOT1_2153(.VSS(VSS),.VDD(VDD),.Y(I9466),.A(g3943));
  NOT NOT1_2154(.VSS(VSS),.VDD(VDD),.Y(g5088),.A(I9466));
  NOT NOT1_2155(.VSS(VSS),.VDD(VDD),.Y(g5099),.A(g4477));
  NOT NOT1_2156(.VSS(VSS),.VDD(VDD),.Y(I9484),.A(g3957));
  NOT NOT1_2157(.VSS(VSS),.VDD(VDD),.Y(g5100),.A(I9484));
  NOT NOT1_2158(.VSS(VSS),.VDD(VDD),.Y(g5101),.A(g4259));
  NOT NOT1_2159(.VSS(VSS),.VDD(VDD),.Y(I9493),.A(g4426));
  NOT NOT1_2160(.VSS(VSS),.VDD(VDD),.Y(g5109),.A(I9493));
  NOT NOT1_2161(.VSS(VSS),.VDD(VDD),.Y(I9496),.A(g3971));
  NOT NOT1_2162(.VSS(VSS),.VDD(VDD),.Y(g5112),.A(I9496));
  NOT NOT1_2163(.VSS(VSS),.VDD(VDD),.Y(I9499),.A(g4382));
  NOT NOT1_2164(.VSS(VSS),.VDD(VDD),.Y(g5113),.A(I9499));
  NOT NOT1_2165(.VSS(VSS),.VDD(VDD),.Y(I9502),.A(g3972));
  NOT NOT1_2166(.VSS(VSS),.VDD(VDD),.Y(g5114),.A(I9502));
  NOT NOT1_2167(.VSS(VSS),.VDD(VDD),.Y(I9505),.A(g4300));
  NOT NOT1_2168(.VSS(VSS),.VDD(VDD),.Y(g5115),.A(I9505));
  NOT NOT1_2169(.VSS(VSS),.VDD(VDD),.Y(I9512),.A(g3985));
  NOT NOT1_2170(.VSS(VSS),.VDD(VDD),.Y(g5120),.A(I9512));
  NOT NOT1_2171(.VSS(VSS),.VDD(VDD),.Y(I9515),.A(g4301));
  NOT NOT1_2172(.VSS(VSS),.VDD(VDD),.Y(g5121),.A(I9515));
  NOT NOT1_2173(.VSS(VSS),.VDD(VDD),.Y(I9520),.A(g3995));
  NOT NOT1_2174(.VSS(VSS),.VDD(VDD),.Y(g5124),.A(I9520));
  NOT NOT1_2175(.VSS(VSS),.VDD(VDD),.Y(I9525),.A(g4413));
  NOT NOT1_2176(.VSS(VSS),.VDD(VDD),.Y(g5127),.A(I9525));
  NOT NOT1_2177(.VSS(VSS),.VDD(VDD),.Y(I9528),.A(g4006));
  NOT NOT1_2178(.VSS(VSS),.VDD(VDD),.Y(g5128),.A(I9528));
  NOT NOT1_2179(.VSS(VSS),.VDD(VDD),.Y(I9531),.A(g4463));
  NOT NOT1_2180(.VSS(VSS),.VDD(VDD),.Y(g5129),.A(I9531));
  NOT NOT1_2181(.VSS(VSS),.VDD(VDD),.Y(I9539),.A(g4018));
  NOT NOT1_2182(.VSS(VSS),.VDD(VDD),.Y(g5137),.A(I9539));
  NOT NOT1_2183(.VSS(VSS),.VDD(VDD),.Y(I9543),.A(g4279));
  NOT NOT1_2184(.VSS(VSS),.VDD(VDD),.Y(g5139),.A(I9543));
  NOT NOT1_2185(.VSS(VSS),.VDD(VDD),.Y(I9555),.A(g4892));
  NOT NOT1_2186(.VSS(VSS),.VDD(VDD),.Y(g5143),.A(I9555));
  NOT NOT1_2187(.VSS(VSS),.VDD(VDD),.Y(I9558),.A(g4597));
  NOT NOT1_2188(.VSS(VSS),.VDD(VDD),.Y(g5144),.A(I9558));
  NOT NOT1_2189(.VSS(VSS),.VDD(VDD),.Y(I9561),.A(g4695));
  NOT NOT1_2190(.VSS(VSS),.VDD(VDD),.Y(g5145),.A(I9561));
  NOT NOT1_2191(.VSS(VSS),.VDD(VDD),.Y(I9564),.A(g4703));
  NOT NOT1_2192(.VSS(VSS),.VDD(VDD),.Y(g5146),.A(I9564));
  NOT NOT1_2193(.VSS(VSS),.VDD(VDD),.Y(I9567),.A(g4693));
  NOT NOT1_2194(.VSS(VSS),.VDD(VDD),.Y(g5147),.A(I9567));
  NOT NOT1_2195(.VSS(VSS),.VDD(VDD),.Y(I9570),.A(g4696));
  NOT NOT1_2196(.VSS(VSS),.VDD(VDD),.Y(g5148),.A(I9570));
  NOT NOT1_2197(.VSS(VSS),.VDD(VDD),.Y(I9573),.A(g4701));
  NOT NOT1_2198(.VSS(VSS),.VDD(VDD),.Y(g5149),.A(I9573));
  NOT NOT1_2199(.VSS(VSS),.VDD(VDD),.Y(I9576),.A(g4706));
  NOT NOT1_2200(.VSS(VSS),.VDD(VDD),.Y(g5150),.A(I9576));
  NOT NOT1_2201(.VSS(VSS),.VDD(VDD),.Y(I9579),.A(g4713));
  NOT NOT1_2202(.VSS(VSS),.VDD(VDD),.Y(g5151),.A(I9579));
  NOT NOT1_2203(.VSS(VSS),.VDD(VDD),.Y(I9582),.A(g4694));
  NOT NOT1_2204(.VSS(VSS),.VDD(VDD),.Y(g5152),.A(I9582));
  NOT NOT1_2205(.VSS(VSS),.VDD(VDD),.Y(I9585),.A(g4697));
  NOT NOT1_2206(.VSS(VSS),.VDD(VDD),.Y(g5153),.A(I9585));
  NOT NOT1_2207(.VSS(VSS),.VDD(VDD),.Y(I9588),.A(g4704));
  NOT NOT1_2208(.VSS(VSS),.VDD(VDD),.Y(g5154),.A(I9588));
  NOT NOT1_2209(.VSS(VSS),.VDD(VDD),.Y(I9591),.A(g4710));
  NOT NOT1_2210(.VSS(VSS),.VDD(VDD),.Y(g5155),.A(I9591));
  NOT NOT1_2211(.VSS(VSS),.VDD(VDD),.Y(I9594),.A(g4718));
  NOT NOT1_2212(.VSS(VSS),.VDD(VDD),.Y(g5156),.A(I9594));
  NOT NOT1_2213(.VSS(VSS),.VDD(VDD),.Y(I9597),.A(g4738));
  NOT NOT1_2214(.VSS(VSS),.VDD(VDD),.Y(g5157),.A(I9597));
  NOT NOT1_2215(.VSS(VSS),.VDD(VDD),.Y(I9600),.A(g4698));
  NOT NOT1_2216(.VSS(VSS),.VDD(VDD),.Y(g5158),.A(I9600));
  NOT NOT1_2217(.VSS(VSS),.VDD(VDD),.Y(I9603),.A(g4719));
  NOT NOT1_2218(.VSS(VSS),.VDD(VDD),.Y(g5159),.A(I9603));
  NOT NOT1_2219(.VSS(VSS),.VDD(VDD),.Y(I9606),.A(g4687));
  NOT NOT1_2220(.VSS(VSS),.VDD(VDD),.Y(g5160),.A(I9606));
  NOT NOT1_2221(.VSS(VSS),.VDD(VDD),.Y(I9609),.A(g4780));
  NOT NOT1_2222(.VSS(VSS),.VDD(VDD),.Y(g5161),.A(I9609));
  NOT NOT1_2223(.VSS(VSS),.VDD(VDD),.Y(I9612),.A(g4776));
  NOT NOT1_2224(.VSS(VSS),.VDD(VDD),.Y(g5162),.A(I9612));
  NOT NOT1_2225(.VSS(VSS),.VDD(VDD),.Y(I9615),.A(g4739));
  NOT NOT1_2226(.VSS(VSS),.VDD(VDD),.Y(g5163),.A(I9615));
  NOT NOT1_2227(.VSS(VSS),.VDD(VDD),.Y(I9618),.A(g4742));
  NOT NOT1_2228(.VSS(VSS),.VDD(VDD),.Y(g5164),.A(I9618));
  NOT NOT1_2229(.VSS(VSS),.VDD(VDD),.Y(I9621),.A(g4732));
  NOT NOT1_2230(.VSS(VSS),.VDD(VDD),.Y(g5165),.A(I9621));
  NOT NOT1_2231(.VSS(VSS),.VDD(VDD),.Y(I9624),.A(g4746));
  NOT NOT1_2232(.VSS(VSS),.VDD(VDD),.Y(g5166),.A(I9624));
  NOT NOT1_2233(.VSS(VSS),.VDD(VDD),.Y(I9627),.A(g4777));
  NOT NOT1_2234(.VSS(VSS),.VDD(VDD),.Y(g5167),.A(I9627));
  NOT NOT1_2235(.VSS(VSS),.VDD(VDD),.Y(I9630),.A(g4867));
  NOT NOT1_2236(.VSS(VSS),.VDD(VDD),.Y(g5168),.A(I9630));
  NOT NOT1_2237(.VSS(VSS),.VDD(VDD),.Y(I9633),.A(g4800));
  NOT NOT1_2238(.VSS(VSS),.VDD(VDD),.Y(g5169),.A(I9633));
  NOT NOT1_2239(.VSS(VSS),.VDD(VDD),.Y(I9636),.A(g4802));
  NOT NOT1_2240(.VSS(VSS),.VDD(VDD),.Y(g5170),.A(I9636));
  NOT NOT1_2241(.VSS(VSS),.VDD(VDD),.Y(I9639),.A(g4685));
  NOT NOT1_2242(.VSS(VSS),.VDD(VDD),.Y(g5171),.A(I9639));
  NOT NOT1_2243(.VSS(VSS),.VDD(VDD),.Y(I9642),.A(g4788));
  NOT NOT1_2244(.VSS(VSS),.VDD(VDD),.Y(g5172),.A(I9642));
  NOT NOT1_2245(.VSS(VSS),.VDD(VDD),.Y(I9645),.A(g4900));
  NOT NOT1_2246(.VSS(VSS),.VDD(VDD),.Y(g5173),.A(I9645));
  NOT NOT1_2247(.VSS(VSS),.VDD(VDD),.Y(I9648),.A(g4795));
  NOT NOT1_2248(.VSS(VSS),.VDD(VDD),.Y(g5174),.A(I9648));
  NOT NOT1_2249(.VSS(VSS),.VDD(VDD),.Y(I9651),.A(g4805));
  NOT NOT1_2250(.VSS(VSS),.VDD(VDD),.Y(g5175),.A(I9651));
  NOT NOT1_2251(.VSS(VSS),.VDD(VDD),.Y(I9654),.A(g4792));
  NOT NOT1_2252(.VSS(VSS),.VDD(VDD),.Y(g5176),.A(I9654));
  NOT NOT1_2253(.VSS(VSS),.VDD(VDD),.Y(I9657),.A(g4784));
  NOT NOT1_2254(.VSS(VSS),.VDD(VDD),.Y(g5177),.A(I9657));
  NOT NOT1_2255(.VSS(VSS),.VDD(VDD),.Y(I9660),.A(g4806));
  NOT NOT1_2256(.VSS(VSS),.VDD(VDD),.Y(g5178),.A(I9660));
  NOT NOT1_2257(.VSS(VSS),.VDD(VDD),.Y(I9663),.A(g4809));
  NOT NOT1_2258(.VSS(VSS),.VDD(VDD),.Y(g5179),.A(I9663));
  NOT NOT1_2259(.VSS(VSS),.VDD(VDD),.Y(I9666),.A(g4931));
  NOT NOT1_2260(.VSS(VSS),.VDD(VDD),.Y(g5180),.A(I9666));
  NOT NOT1_2261(.VSS(VSS),.VDD(VDD),.Y(I9669),.A(g4909));
  NOT NOT1_2262(.VSS(VSS),.VDD(VDD),.Y(g5181),.A(I9669));
  NOT NOT1_2263(.VSS(VSS),.VDD(VDD),.Y(I9672),.A(g4803));
  NOT NOT1_2264(.VSS(VSS),.VDD(VDD),.Y(g5182),.A(I9672));
  NOT NOT1_2265(.VSS(VSS),.VDD(VDD),.Y(I9675),.A(g4807));
  NOT NOT1_2266(.VSS(VSS),.VDD(VDD),.Y(g5183),.A(I9675));
  NOT NOT1_2267(.VSS(VSS),.VDD(VDD),.Y(I9678),.A(g4808));
  NOT NOT1_2268(.VSS(VSS),.VDD(VDD),.Y(g5184),.A(I9678));
  NOT NOT1_2269(.VSS(VSS),.VDD(VDD),.Y(I9681),.A(g4811));
  NOT NOT1_2270(.VSS(VSS),.VDD(VDD),.Y(g5185),.A(I9681));
  NOT NOT1_2271(.VSS(VSS),.VDD(VDD),.Y(I9684),.A(g4813));
  NOT NOT1_2272(.VSS(VSS),.VDD(VDD),.Y(g5186),.A(I9684));
  NOT NOT1_2273(.VSS(VSS),.VDD(VDD),.Y(I9687),.A(g4822));
  NOT NOT1_2274(.VSS(VSS),.VDD(VDD),.Y(g5187),.A(I9687));
  NOT NOT1_2275(.VSS(VSS),.VDD(VDD),.Y(g5190),.A(g4938));
  NOT NOT1_2276(.VSS(VSS),.VDD(VDD),.Y(g5191),.A(g4969));
  NOT NOT1_2277(.VSS(VSS),.VDD(VDD),.Y(g5192),.A(g4841));
  NOT NOT1_2278(.VSS(VSS),.VDD(VDD),.Y(g5197),.A(g4938));
  NOT NOT1_2279(.VSS(VSS),.VDD(VDD),.Y(g5198),.A(g4969));
  NOT NOT1_2280(.VSS(VSS),.VDD(VDD),.Y(g5199),.A(g4841));
  NOT NOT1_2281(.VSS(VSS),.VDD(VDD),.Y(g5206),.A(g4938));
  NOT NOT1_2282(.VSS(VSS),.VDD(VDD),.Y(g5207),.A(g4673));
  NOT NOT1_2283(.VSS(VSS),.VDD(VDD),.Y(g5224),.A(g5114));
  NOT NOT1_2284(.VSS(VSS),.VDD(VDD),.Y(I9752),.A(g4705));
  NOT NOT1_2285(.VSS(VSS),.VDD(VDD),.Y(g5240),.A(I9752));
  NOT NOT1_2286(.VSS(VSS),.VDD(VDD),.Y(I9760),.A(g4838));
  NOT NOT1_2287(.VSS(VSS),.VDD(VDD),.Y(g5246),.A(I9760));
  NOT NOT1_2288(.VSS(VSS),.VDD(VDD),.Y(I9774),.A(g4678));
  NOT NOT1_2289(.VSS(VSS),.VDD(VDD),.Y(g5258),.A(I9774));
  NOT NOT1_2290(.VSS(VSS),.VDD(VDD),.Y(g5261),.A(g4748));
  NOT NOT1_2291(.VSS(VSS),.VDD(VDD),.Y(I9782),.A(g4720));
  NOT NOT1_2292(.VSS(VSS),.VDD(VDD),.Y(g5266),.A(I9782));
  NOT NOT1_2293(.VSS(VSS),.VDD(VDD),.Y(I9785),.A(g4747));
  NOT NOT1_2294(.VSS(VSS),.VDD(VDD),.Y(g5267),.A(I9785));
  NOT NOT1_2295(.VSS(VSS),.VDD(VDD),.Y(I9788),.A(g4711));
  NOT NOT1_2296(.VSS(VSS),.VDD(VDD),.Y(g5268),.A(I9788));
  NOT NOT1_2297(.VSS(VSS),.VDD(VDD),.Y(I9791),.A(g4779));
  NOT NOT1_2298(.VSS(VSS),.VDD(VDD),.Y(g5269),.A(I9791));
  NOT NOT1_2299(.VSS(VSS),.VDD(VDD),.Y(I9794),.A(g4778));
  NOT NOT1_2300(.VSS(VSS),.VDD(VDD),.Y(g5278),.A(I9794));
  NOT NOT1_2301(.VSS(VSS),.VDD(VDD),.Y(g5285),.A(g4841));
  NOT NOT1_2302(.VSS(VSS),.VDD(VDD),.Y(g5286),.A(g4714));
  NOT NOT1_2303(.VSS(VSS),.VDD(VDD),.Y(g5294),.A(g5087));
  NOT NOT1_2304(.VSS(VSS),.VDD(VDD),.Y(I9804),.A(g5113));
  NOT NOT1_2305(.VSS(VSS),.VDD(VDD),.Y(g5299),.A(I9804));
  NOT NOT1_2306(.VSS(VSS),.VDD(VDD),.Y(g5302),.A(g5028));
  NOT NOT1_2307(.VSS(VSS),.VDD(VDD),.Y(g5309),.A(g4969));
  NOT NOT1_2308(.VSS(VSS),.VDD(VDD),.Y(g5311),.A(g4938));
  NOT NOT1_2309(.VSS(VSS),.VDD(VDD),.Y(g5335),.A(g4677));
  NOT NOT1_2310(.VSS(VSS),.VDD(VDD),.Y(I9819),.A(g4691));
  NOT NOT1_2311(.VSS(VSS),.VDD(VDD),.Y(g5344),.A(I9819));
  NOT NOT1_2312(.VSS(VSS),.VDD(VDD),.Y(I9823),.A(g5138));
  NOT NOT1_2313(.VSS(VSS),.VDD(VDD),.Y(g5362),.A(I9823));
  NOT NOT1_2314(.VSS(VSS),.VDD(VDD),.Y(g5364),.A(g5124));
  NOT NOT1_2315(.VSS(VSS),.VDD(VDD),.Y(I9834),.A(g4782));
  NOT NOT1_2316(.VSS(VSS),.VDD(VDD),.Y(g5367),.A(I9834));
  NOT NOT1_2317(.VSS(VSS),.VDD(VDD),.Y(I9837),.A(g4781));
  NOT NOT1_2318(.VSS(VSS),.VDD(VDD),.Y(g5384),.A(I9837));
  NOT NOT1_2319(.VSS(VSS),.VDD(VDD),.Y(I9840),.A(g4702));
  NOT NOT1_2320(.VSS(VSS),.VDD(VDD),.Y(g5395),.A(I9840));
  NOT NOT1_2321(.VSS(VSS),.VDD(VDD),.Y(g5396),.A(g4692));
  NOT NOT1_2322(.VSS(VSS),.VDD(VDD),.Y(g5397),.A(g5076));
  NOT NOT1_2323(.VSS(VSS),.VDD(VDD),.Y(I9845),.A(g4728));
  NOT NOT1_2324(.VSS(VSS),.VDD(VDD),.Y(g5401),.A(I9845));
  NOT NOT1_2325(.VSS(VSS),.VDD(VDD),.Y(g5402),.A(g5000));
  NOT NOT1_2326(.VSS(VSS),.VDD(VDD),.Y(g5403),.A(g5088));
  NOT NOT1_2327(.VSS(VSS),.VDD(VDD),.Y(I9850),.A(g4798));
  NOT NOT1_2328(.VSS(VSS),.VDD(VDD),.Y(g5412),.A(I9850));
  NOT NOT1_2329(.VSS(VSS),.VDD(VDD),.Y(g5417),.A(g5006));
  NOT NOT1_2330(.VSS(VSS),.VDD(VDD),.Y(g5418),.A(g5100));
  NOT NOT1_2331(.VSS(VSS),.VDD(VDD),.Y(g5426),.A(g5013));
  NOT NOT1_2332(.VSS(VSS),.VDD(VDD),.Y(g5427),.A(g5115));
  NOT NOT1_2333(.VSS(VSS),.VDD(VDD),.Y(g5433),.A(g5024));
  NOT NOT1_2334(.VSS(VSS),.VDD(VDD),.Y(g5434),.A(g5112));
  NOT NOT1_2335(.VSS(VSS),.VDD(VDD),.Y(g5435),.A(g5121));
  NOT NOT1_2336(.VSS(VSS),.VDD(VDD),.Y(g5437),.A(g5041));
  NOT NOT1_2337(.VSS(VSS),.VDD(VDD),.Y(g5439),.A(g5058));
  NOT NOT1_2338(.VSS(VSS),.VDD(VDD),.Y(g5444),.A(g5074));
  NOT NOT1_2339(.VSS(VSS),.VDD(VDD),.Y(g5445),.A(g5059));
  NOT NOT1_2340(.VSS(VSS),.VDD(VDD),.Y(g5448),.A(g5137));
  NOT NOT1_2341(.VSS(VSS),.VDD(VDD),.Y(g5453),.A(g4680));
  NOT NOT1_2342(.VSS(VSS),.VDD(VDD),.Y(g5459),.A(g4882));
  NOT NOT1_2343(.VSS(VSS),.VDD(VDD),.Y(g5460),.A(g4684));
  NOT NOT1_2344(.VSS(VSS),.VDD(VDD),.Y(g5461),.A(g4885));
  NOT NOT1_2345(.VSS(VSS),.VDD(VDD),.Y(g5462),.A(g4886));
  NOT NOT1_2346(.VSS(VSS),.VDD(VDD),.Y(g5463),.A(g5085));
  NOT NOT1_2347(.VSS(VSS),.VDD(VDD),.Y(g5466),.A(g4890));
  NOT NOT1_2348(.VSS(VSS),.VDD(VDD),.Y(g5467),.A(g4891));
  NOT NOT1_2349(.VSS(VSS),.VDD(VDD),.Y(I9884),.A(g4868));
  NOT NOT1_2350(.VSS(VSS),.VDD(VDD),.Y(g5468),.A(I9884));
  NOT NOT1_2351(.VSS(VSS),.VDD(VDD),.Y(g5469),.A(g4898));
  NOT NOT1_2352(.VSS(VSS),.VDD(VDD),.Y(g5470),.A(g4899));
  NOT NOT1_2353(.VSS(VSS),.VDD(VDD),.Y(I9889),.A(g4819));
  NOT NOT1_2354(.VSS(VSS),.VDD(VDD),.Y(g5471),.A(I9889));
  NOT NOT1_2355(.VSS(VSS),.VDD(VDD),.Y(I9892),.A(g4879));
  NOT NOT1_2356(.VSS(VSS),.VDD(VDD),.Y(g5472),.A(I9892));
  NOT NOT1_2357(.VSS(VSS),.VDD(VDD),.Y(g5473),.A(g4903));
  NOT NOT1_2358(.VSS(VSS),.VDD(VDD),.Y(g5474),.A(g4904));
  NOT NOT1_2359(.VSS(VSS),.VDD(VDD),.Y(g5476),.A(g4907));
  NOT NOT1_2360(.VSS(VSS),.VDD(VDD),.Y(g5477),.A(g4908));
  NOT NOT1_2361(.VSS(VSS),.VDD(VDD),.Y(g5478),.A(g5025));
  NOT NOT1_2362(.VSS(VSS),.VDD(VDD),.Y(g5480),.A(g4913));
  NOT NOT1_2363(.VSS(VSS),.VDD(VDD),.Y(g5481),.A(g4914));
  NOT NOT1_2364(.VSS(VSS),.VDD(VDD),.Y(g5482),.A(g4915));
  NOT NOT1_2365(.VSS(VSS),.VDD(VDD),.Y(I9907),.A(g4837));
  NOT NOT1_2366(.VSS(VSS),.VDD(VDD),.Y(g5487),.A(I9907));
  NOT NOT1_2367(.VSS(VSS),.VDD(VDD),.Y(I9910),.A(g4681));
  NOT NOT1_2368(.VSS(VSS),.VDD(VDD),.Y(g5488),.A(I9910));
  NOT NOT1_2369(.VSS(VSS),.VDD(VDD),.Y(g5490),.A(g4917));
  NOT NOT1_2370(.VSS(VSS),.VDD(VDD),.Y(g5491),.A(g4918));
  NOT NOT1_2371(.VSS(VSS),.VDD(VDD),.Y(g5492),.A(g4919));
  NOT NOT1_2372(.VSS(VSS),.VDD(VDD),.Y(g5493),.A(g4920));
  NOT NOT1_2373(.VSS(VSS),.VDD(VDD),.Y(I9918),.A(g4968));
  NOT NOT1_2374(.VSS(VSS),.VDD(VDD),.Y(g5494),.A(I9918));
  NOT NOT1_2375(.VSS(VSS),.VDD(VDD),.Y(g5514),.A(g4922));
  NOT NOT1_2376(.VSS(VSS),.VDD(VDD),.Y(g5515),.A(g4923));
  NOT NOT1_2377(.VSS(VSS),.VDD(VDD),.Y(g5516),.A(g4924));
  NOT NOT1_2378(.VSS(VSS),.VDD(VDD),.Y(g5517),.A(g4925));
  NOT NOT1_2379(.VSS(VSS),.VDD(VDD),.Y(I9929),.A(g5052));
  NOT NOT1_2380(.VSS(VSS),.VDD(VDD),.Y(g5519),.A(I9929));
  NOT NOT1_2381(.VSS(VSS),.VDD(VDD),.Y(g5520),.A(g4928));
  NOT NOT1_2382(.VSS(VSS),.VDD(VDD),.Y(g5521),.A(g4929));
  NOT NOT1_2383(.VSS(VSS),.VDD(VDD),.Y(g5522),.A(g4930));
  NOT NOT1_2384(.VSS(VSS),.VDD(VDD),.Y(I9935),.A(g4812));
  NOT NOT1_2385(.VSS(VSS),.VDD(VDD),.Y(g5523),.A(I9935));
  NOT NOT1_2386(.VSS(VSS),.VDD(VDD),.Y(I9938),.A(g4878));
  NOT NOT1_2387(.VSS(VSS),.VDD(VDD),.Y(g5524),.A(I9938));
  NOT NOT1_2388(.VSS(VSS),.VDD(VDD),.Y(g5525),.A(g4934));
  NOT NOT1_2389(.VSS(VSS),.VDD(VDD),.Y(g5526),.A(g5086));
  NOT NOT1_2390(.VSS(VSS),.VDD(VDD),.Y(g5529),.A(g4689));
  NOT NOT1_2391(.VSS(VSS),.VDD(VDD),.Y(g5541),.A(g4814));
  NOT NOT1_2392(.VSS(VSS),.VDD(VDD),.Y(g5542),.A(g5061));
  NOT NOT1_2393(.VSS(VSS),.VDD(VDD),.Y(I9974),.A(g4676));
  NOT NOT1_2394(.VSS(VSS),.VDD(VDD),.Y(g5551),.A(I9974));
  NOT NOT1_2395(.VSS(VSS),.VDD(VDD),.Y(I10028),.A(g4825));
  NOT NOT1_2396(.VSS(VSS),.VDD(VDD),.Y(g5569),.A(I10028));
  NOT NOT1_2397(.VSS(VSS),.VDD(VDD),.Y(I10032),.A(g1236));
  NOT NOT1_2398(.VSS(VSS),.VDD(VDD),.Y(g5571),.A(I10032));
  NOT NOT1_2399(.VSS(VSS),.VDD(VDD),.Y(g5574),.A(g4969));
  NOT NOT1_2400(.VSS(VSS),.VDD(VDD),.Y(I10046),.A(g4840));
  NOT NOT1_2401(.VSS(VSS),.VDD(VDD),.Y(g5577),.A(I10046));
  NOT NOT1_2402(.VSS(VSS),.VDD(VDD),.Y(g5578),.A(g4841));
  NOT NOT1_2403(.VSS(VSS),.VDD(VDD),.Y(g5580),.A(g4938));
  NOT NOT1_2404(.VSS(VSS),.VDD(VDD),.Y(g5581),.A(g4969));
  NOT NOT1_2405(.VSS(VSS),.VDD(VDD),.Y(g5582),.A(g4969));
  NOT NOT1_2406(.VSS(VSS),.VDD(VDD),.Y(g5584),.A(g4841));
  NOT NOT1_2407(.VSS(VSS),.VDD(VDD),.Y(g5586),.A(g4938));
  NOT NOT1_2408(.VSS(VSS),.VDD(VDD),.Y(g5587),.A(g4938));
  NOT NOT1_2409(.VSS(VSS),.VDD(VDD),.Y(g5591),.A(g4841));
  NOT NOT1_2410(.VSS(VSS),.VDD(VDD),.Y(g5592),.A(g4969));
  NOT NOT1_2411(.VSS(VSS),.VDD(VDD),.Y(g5596),.A(g4841));
  NOT NOT1_2412(.VSS(VSS),.VDD(VDD),.Y(g5597),.A(g4969));
  NOT NOT1_2413(.VSS(VSS),.VDD(VDD),.Y(g5598),.A(g4938));
  NOT NOT1_2414(.VSS(VSS),.VDD(VDD),.Y(g5600),.A(g5128));
  NOT NOT1_2415(.VSS(VSS),.VDD(VDD),.Y(g5603),.A(g4938));
  NOT NOT1_2416(.VSS(VSS),.VDD(VDD),.Y(g5604),.A(g4969));
  NOT NOT1_2417(.VSS(VSS),.VDD(VDD),.Y(g5606),.A(g4748));
  NOT NOT1_2418(.VSS(VSS),.VDD(VDD),.Y(g5607),.A(g4938));
  NOT NOT1_2419(.VSS(VSS),.VDD(VDD),.Y(g5608),.A(g4969));
  NOT NOT1_2420(.VSS(VSS),.VDD(VDD),.Y(g5609),.A(g4748));
  NOT NOT1_2421(.VSS(VSS),.VDD(VDD),.Y(g5610),.A(g4938));
  NOT NOT1_2422(.VSS(VSS),.VDD(VDD),.Y(g5611),.A(g4969));
  NOT NOT1_2423(.VSS(VSS),.VDD(VDD),.Y(g5612),.A(g4814));
  NOT NOT1_2424(.VSS(VSS),.VDD(VDD),.Y(g5613),.A(g4748));
  NOT NOT1_2425(.VSS(VSS),.VDD(VDD),.Y(g5616),.A(g4938));
  NOT NOT1_2426(.VSS(VSS),.VDD(VDD),.Y(g5617),.A(g4969));
  NOT NOT1_2427(.VSS(VSS),.VDD(VDD),.Y(g5618),.A(g5015));
  NOT NOT1_2428(.VSS(VSS),.VDD(VDD),.Y(g5621),.A(g4748));
  NOT NOT1_2429(.VSS(VSS),.VDD(VDD),.Y(g5622),.A(g4938));
  NOT NOT1_2430(.VSS(VSS),.VDD(VDD),.Y(g5623),.A(g4969));
  NOT NOT1_2431(.VSS(VSS),.VDD(VDD),.Y(g5626),.A(g4748));
  NOT NOT1_2432(.VSS(VSS),.VDD(VDD),.Y(g5627),.A(g4673));
  NOT NOT1_2433(.VSS(VSS),.VDD(VDD),.Y(g5628),.A(g4748));
  NOT NOT1_2434(.VSS(VSS),.VDD(VDD),.Y(g5631),.A(g4938));
  NOT NOT1_2435(.VSS(VSS),.VDD(VDD),.Y(g5633),.A(g4895));
  NOT NOT1_2436(.VSS(VSS),.VDD(VDD),.Y(g5638),.A(g4748));
  NOT NOT1_2437(.VSS(VSS),.VDD(VDD),.Y(g5639),.A(g4748));
  NOT NOT1_2438(.VSS(VSS),.VDD(VDD),.Y(I10125),.A(g5127));
  NOT NOT1_2439(.VSS(VSS),.VDD(VDD),.Y(g5642),.A(I10125));
  NOT NOT1_2440(.VSS(VSS),.VDD(VDD),.Y(I10128),.A(g4688));
  NOT NOT1_2441(.VSS(VSS),.VDD(VDD),.Y(g5643),.A(I10128));
  NOT NOT1_2442(.VSS(VSS),.VDD(VDD),.Y(g5644),.A(g4748));
  NOT NOT1_2443(.VSS(VSS),.VDD(VDD),.Y(g5645),.A(g4748));
  NOT NOT1_2444(.VSS(VSS),.VDD(VDD),.Y(g5648),.A(g4748));
  NOT NOT1_2445(.VSS(VSS),.VDD(VDD),.Y(g5649),.A(g4748));
  NOT NOT1_2446(.VSS(VSS),.VDD(VDD),.Y(I10135),.A(g4960));
  NOT NOT1_2447(.VSS(VSS),.VDD(VDD),.Y(g5652),.A(I10135));
  NOT NOT1_2448(.VSS(VSS),.VDD(VDD),.Y(g5653),.A(g4748));
  NOT NOT1_2449(.VSS(VSS),.VDD(VDD),.Y(g5654),.A(g4748));
  NOT NOT1_2450(.VSS(VSS),.VDD(VDD),.Y(g5658),.A(g4748));
  NOT NOT1_2451(.VSS(VSS),.VDD(VDD),.Y(g5662),.A(g5027));
  NOT NOT1_2452(.VSS(VSS),.VDD(VDD),.Y(g5665),.A(g4748));
  NOT NOT1_2453(.VSS(VSS),.VDD(VDD),.Y(I10151),.A(g5007));
  NOT NOT1_2454(.VSS(VSS),.VDD(VDD),.Y(g5668),.A(I10151));
  NOT NOT1_2455(.VSS(VSS),.VDD(VDD),.Y(I10154),.A(g5109));
  NOT NOT1_2456(.VSS(VSS),.VDD(VDD),.Y(g5669),.A(I10154));
  NOT NOT1_2457(.VSS(VSS),.VDD(VDD),.Y(I10157),.A(g5109));
  NOT NOT1_2458(.VSS(VSS),.VDD(VDD),.Y(g5670),.A(I10157));
  NOT NOT1_2459(.VSS(VSS),.VDD(VDD),.Y(I10160),.A(g5139));
  NOT NOT1_2460(.VSS(VSS),.VDD(VDD),.Y(g5671),.A(I10160));
  NOT NOT1_2461(.VSS(VSS),.VDD(VDD),.Y(g5674),.A(g5042));
  NOT NOT1_2462(.VSS(VSS),.VDD(VDD),.Y(I10166),.A(g5016));
  NOT NOT1_2463(.VSS(VSS),.VDD(VDD),.Y(g5677),.A(I10166));
  NOT NOT1_2464(.VSS(VSS),.VDD(VDD),.Y(I10169),.A(g4873));
  NOT NOT1_2465(.VSS(VSS),.VDD(VDD),.Y(g5678),.A(I10169));
  NOT NOT1_2466(.VSS(VSS),.VDD(VDD),.Y(I10172),.A(g4873));
  NOT NOT1_2467(.VSS(VSS),.VDD(VDD),.Y(g5679),.A(I10172));
  NOT NOT1_2468(.VSS(VSS),.VDD(VDD),.Y(g5680),.A(g5101));
  NOT NOT1_2469(.VSS(VSS),.VDD(VDD),.Y(I10177),.A(g4721));
  NOT NOT1_2470(.VSS(VSS),.VDD(VDD),.Y(g5682),.A(I10177));
  NOT NOT1_2471(.VSS(VSS),.VDD(VDD),.Y(I10180),.A(g4721));
  NOT NOT1_2472(.VSS(VSS),.VDD(VDD),.Y(g5683),.A(I10180));
  NOT NOT1_2473(.VSS(VSS),.VDD(VDD),.Y(I10183),.A(g5129));
  NOT NOT1_2474(.VSS(VSS),.VDD(VDD),.Y(g5684),.A(I10183));
  NOT NOT1_2475(.VSS(VSS),.VDD(VDD),.Y(I10186),.A(g5129));
  NOT NOT1_2476(.VSS(VSS),.VDD(VDD),.Y(g5685),.A(I10186));
  NOT NOT1_2477(.VSS(VSS),.VDD(VDD),.Y(I10190),.A(g4670));
  NOT NOT1_2478(.VSS(VSS),.VDD(VDD),.Y(g5687),.A(I10190));
  NOT NOT1_2479(.VSS(VSS),.VDD(VDD),.Y(I10193),.A(g4670));
  NOT NOT1_2480(.VSS(VSS),.VDD(VDD),.Y(g5688),.A(I10193));
  NOT NOT1_2481(.VSS(VSS),.VDD(VDD),.Y(g5690),.A(g4748));
  NOT NOT1_2482(.VSS(VSS),.VDD(VDD),.Y(I10204),.A(g5060));
  NOT NOT1_2483(.VSS(VSS),.VDD(VDD),.Y(g5693),.A(I10204));
  NOT NOT1_2484(.VSS(VSS),.VDD(VDD),.Y(I10207),.A(g5075));
  NOT NOT1_2485(.VSS(VSS),.VDD(VDD),.Y(g5696),.A(I10207));
  NOT NOT1_2486(.VSS(VSS),.VDD(VDD),.Y(g5701),.A(g5120));
  NOT NOT1_2487(.VSS(VSS),.VDD(VDD),.Y(g5705),.A(g4841));
  NOT NOT1_2488(.VSS(VSS),.VDD(VDD),.Y(g5709),.A(g4841));
  NOT NOT1_2489(.VSS(VSS),.VDD(VDD),.Y(g5713),.A(g4841));
  NOT NOT1_2490(.VSS(VSS),.VDD(VDD),.Y(g5717),.A(g4969));
  NOT NOT1_2491(.VSS(VSS),.VDD(VDD),.Y(g5718),.A(g4841));
  NOT NOT1_2492(.VSS(VSS),.VDD(VDD),.Y(I10236),.A(g5014));
  NOT NOT1_2493(.VSS(VSS),.VDD(VDD),.Y(g5719),.A(I10236));
  NOT NOT1_2494(.VSS(VSS),.VDD(VDD),.Y(g5723),.A(g4938));
  NOT NOT1_2495(.VSS(VSS),.VDD(VDD),.Y(g5724),.A(g4969));
  NOT NOT1_2496(.VSS(VSS),.VDD(VDD),.Y(g5725),.A(g4841));
  NOT NOT1_2497(.VSS(VSS),.VDD(VDD),.Y(I10243),.A(g5026));
  NOT NOT1_2498(.VSS(VSS),.VDD(VDD),.Y(g5726),.A(I10243));
  NOT NOT1_2499(.VSS(VSS),.VDD(VDD),.Y(g5729),.A(g5144));
  NOT NOT1_2500(.VSS(VSS),.VDD(VDD),.Y(I10247),.A(g5266));
  NOT NOT1_2501(.VSS(VSS),.VDD(VDD),.Y(g5730),.A(I10247));
  NOT NOT1_2502(.VSS(VSS),.VDD(VDD),.Y(I10250),.A(g5268));
  NOT NOT1_2503(.VSS(VSS),.VDD(VDD),.Y(g5731),.A(I10250));
  NOT NOT1_2504(.VSS(VSS),.VDD(VDD),.Y(I10253),.A(g5240));
  NOT NOT1_2505(.VSS(VSS),.VDD(VDD),.Y(g5732),.A(I10253));
  NOT NOT1_2506(.VSS(VSS),.VDD(VDD),.Y(I10256),.A(g5401));
  NOT NOT1_2507(.VSS(VSS),.VDD(VDD),.Y(g5733),.A(I10256));
  NOT NOT1_2508(.VSS(VSS),.VDD(VDD),.Y(I10259),.A(g5362));
  NOT NOT1_2509(.VSS(VSS),.VDD(VDD),.Y(g5734),.A(I10259));
  NOT NOT1_2510(.VSS(VSS),.VDD(VDD),.Y(I10262),.A(g5551));
  NOT NOT1_2511(.VSS(VSS),.VDD(VDD),.Y(g5735),.A(I10262));
  NOT NOT1_2512(.VSS(VSS),.VDD(VDD),.Y(I10265),.A(g5468));
  NOT NOT1_2513(.VSS(VSS),.VDD(VDD),.Y(g5736),.A(I10265));
  NOT NOT1_2514(.VSS(VSS),.VDD(VDD),.Y(I10268),.A(g5471));
  NOT NOT1_2515(.VSS(VSS),.VDD(VDD),.Y(g5737),.A(I10268));
  NOT NOT1_2516(.VSS(VSS),.VDD(VDD),.Y(I10271),.A(g5487));
  NOT NOT1_2517(.VSS(VSS),.VDD(VDD),.Y(g5738),.A(I10271));
  NOT NOT1_2518(.VSS(VSS),.VDD(VDD),.Y(I10274),.A(g5524));
  NOT NOT1_2519(.VSS(VSS),.VDD(VDD),.Y(g5739),.A(I10274));
  NOT NOT1_2520(.VSS(VSS),.VDD(VDD),.Y(I10277),.A(g5472));
  NOT NOT1_2521(.VSS(VSS),.VDD(VDD),.Y(g5740),.A(I10277));
  NOT NOT1_2522(.VSS(VSS),.VDD(VDD),.Y(I10280),.A(g5488));
  NOT NOT1_2523(.VSS(VSS),.VDD(VDD),.Y(g5741),.A(I10280));
  NOT NOT1_2524(.VSS(VSS),.VDD(VDD),.Y(I10283),.A(g5643));
  NOT NOT1_2525(.VSS(VSS),.VDD(VDD),.Y(g5742),.A(I10283));
  NOT NOT1_2526(.VSS(VSS),.VDD(VDD),.Y(I10286),.A(g5519));
  NOT NOT1_2527(.VSS(VSS),.VDD(VDD),.Y(g5743),.A(I10286));
  NOT NOT1_2528(.VSS(VSS),.VDD(VDD),.Y(I10289),.A(g5569));
  NOT NOT1_2529(.VSS(VSS),.VDD(VDD),.Y(g5744),.A(I10289));
  NOT NOT1_2530(.VSS(VSS),.VDD(VDD),.Y(I10292),.A(g5577));
  NOT NOT1_2531(.VSS(VSS),.VDD(VDD),.Y(g5745),.A(I10292));
  NOT NOT1_2532(.VSS(VSS),.VDD(VDD),.Y(I10295),.A(g5523));
  NOT NOT1_2533(.VSS(VSS),.VDD(VDD),.Y(g5746),.A(I10295));
  NOT NOT1_2534(.VSS(VSS),.VDD(VDD),.Y(g5749),.A(g5207));
  NOT NOT1_2535(.VSS(VSS),.VDD(VDD),.Y(g5754),.A(g5403));
  NOT NOT1_2536(.VSS(VSS),.VDD(VDD),.Y(g5755),.A(g5494));
  NOT NOT1_2537(.VSS(VSS),.VDD(VDD),.Y(I10343),.A(g5704));
  NOT NOT1_2538(.VSS(VSS),.VDD(VDD),.Y(g5756),.A(I10343));
  NOT NOT1_2539(.VSS(VSS),.VDD(VDD),.Y(g5757),.A(g5261));
  NOT NOT1_2540(.VSS(VSS),.VDD(VDD),.Y(I10347),.A(g5706));
  NOT NOT1_2541(.VSS(VSS),.VDD(VDD),.Y(g5758),.A(I10347));
  NOT NOT1_2542(.VSS(VSS),.VDD(VDD),.Y(I10350),.A(g5707));
  NOT NOT1_2543(.VSS(VSS),.VDD(VDD),.Y(g5759),.A(I10350));
  NOT NOT1_2544(.VSS(VSS),.VDD(VDD),.Y(I10353),.A(g5710));
  NOT NOT1_2545(.VSS(VSS),.VDD(VDD),.Y(g5760),.A(I10353));
  NOT NOT1_2546(.VSS(VSS),.VDD(VDD),.Y(I10356),.A(g5711));
  NOT NOT1_2547(.VSS(VSS),.VDD(VDD),.Y(g5761),.A(I10356));
  NOT NOT1_2548(.VSS(VSS),.VDD(VDD),.Y(I10366),.A(g5715));
  NOT NOT1_2549(.VSS(VSS),.VDD(VDD),.Y(g5763),.A(I10366));
  NOT NOT1_2550(.VSS(VSS),.VDD(VDD),.Y(I10369),.A(g5716));
  NOT NOT1_2551(.VSS(VSS),.VDD(VDD),.Y(g5764),.A(I10369));
  NOT NOT1_2552(.VSS(VSS),.VDD(VDD),.Y(I10373),.A(g5722));
  NOT NOT1_2553(.VSS(VSS),.VDD(VDD),.Y(g5766),.A(I10373));
  NOT NOT1_2554(.VSS(VSS),.VDD(VDD),.Y(I10377),.A(g5188));
  NOT NOT1_2555(.VSS(VSS),.VDD(VDD),.Y(g5768),.A(I10377));
  NOT NOT1_2556(.VSS(VSS),.VDD(VDD),.Y(I10380),.A(g5448));
  NOT NOT1_2557(.VSS(VSS),.VDD(VDD),.Y(g5769),.A(I10380));
  NOT NOT1_2558(.VSS(VSS),.VDD(VDD),.Y(I10384),.A(g5193));
  NOT NOT1_2559(.VSS(VSS),.VDD(VDD),.Y(g5779),.A(I10384));
  NOT NOT1_2560(.VSS(VSS),.VDD(VDD),.Y(I10387),.A(g5194));
  NOT NOT1_2561(.VSS(VSS),.VDD(VDD),.Y(g5780),.A(I10387));
  NOT NOT1_2562(.VSS(VSS),.VDD(VDD),.Y(I10390),.A(g5195));
  NOT NOT1_2563(.VSS(VSS),.VDD(VDD),.Y(g5781),.A(I10390));
  NOT NOT1_2564(.VSS(VSS),.VDD(VDD),.Y(I10393),.A(g5196));
  NOT NOT1_2565(.VSS(VSS),.VDD(VDD),.Y(g5782),.A(I10393));
  NOT NOT1_2566(.VSS(VSS),.VDD(VDD),.Y(I10397),.A(g5200));
  NOT NOT1_2567(.VSS(VSS),.VDD(VDD),.Y(g5784),.A(I10397));
  NOT NOT1_2568(.VSS(VSS),.VDD(VDD),.Y(I10400),.A(g5201));
  NOT NOT1_2569(.VSS(VSS),.VDD(VDD),.Y(g5785),.A(I10400));
  NOT NOT1_2570(.VSS(VSS),.VDD(VDD),.Y(I10403),.A(g5202));
  NOT NOT1_2571(.VSS(VSS),.VDD(VDD),.Y(g5786),.A(I10403));
  NOT NOT1_2572(.VSS(VSS),.VDD(VDD),.Y(I10406),.A(g5203));
  NOT NOT1_2573(.VSS(VSS),.VDD(VDD),.Y(g5787),.A(I10406));
  NOT NOT1_2574(.VSS(VSS),.VDD(VDD),.Y(I10409),.A(g5204));
  NOT NOT1_2575(.VSS(VSS),.VDD(VDD),.Y(g5788),.A(I10409));
  NOT NOT1_2576(.VSS(VSS),.VDD(VDD),.Y(I10412),.A(g5205));
  NOT NOT1_2577(.VSS(VSS),.VDD(VDD),.Y(g5789),.A(I10412));
  NOT NOT1_2578(.VSS(VSS),.VDD(VDD),.Y(I10415),.A(g5397));
  NOT NOT1_2579(.VSS(VSS),.VDD(VDD),.Y(g5790),.A(I10415));
  NOT NOT1_2580(.VSS(VSS),.VDD(VDD),.Y(I10418),.A(g5453));
  NOT NOT1_2581(.VSS(VSS),.VDD(VDD),.Y(g5793),.A(I10418));
  NOT NOT1_2582(.VSS(VSS),.VDD(VDD),.Y(I10421),.A(g5208));
  NOT NOT1_2583(.VSS(VSS),.VDD(VDD),.Y(g5794),.A(I10421));
  NOT NOT1_2584(.VSS(VSS),.VDD(VDD),.Y(I10424),.A(g5209));
  NOT NOT1_2585(.VSS(VSS),.VDD(VDD),.Y(g5795),.A(I10424));
  NOT NOT1_2586(.VSS(VSS),.VDD(VDD),.Y(I10427),.A(g5210));
  NOT NOT1_2587(.VSS(VSS),.VDD(VDD),.Y(g5796),.A(I10427));
  NOT NOT1_2588(.VSS(VSS),.VDD(VDD),.Y(I10430),.A(g5211));
  NOT NOT1_2589(.VSS(VSS),.VDD(VDD),.Y(g5797),.A(I10430));
  NOT NOT1_2590(.VSS(VSS),.VDD(VDD),.Y(I10433),.A(g5212));
  NOT NOT1_2591(.VSS(VSS),.VDD(VDD),.Y(g5798),.A(I10433));
  NOT NOT1_2592(.VSS(VSS),.VDD(VDD),.Y(I10436),.A(g5213));
  NOT NOT1_2593(.VSS(VSS),.VDD(VDD),.Y(g5799),.A(I10436));
  NOT NOT1_2594(.VSS(VSS),.VDD(VDD),.Y(I10439),.A(g5214));
  NOT NOT1_2595(.VSS(VSS),.VDD(VDD),.Y(g5800),.A(I10439));
  NOT NOT1_2596(.VSS(VSS),.VDD(VDD),.Y(I10442),.A(g5215));
  NOT NOT1_2597(.VSS(VSS),.VDD(VDD),.Y(g5801),.A(I10442));
  NOT NOT1_2598(.VSS(VSS),.VDD(VDD),.Y(I10445),.A(g5418));
  NOT NOT1_2599(.VSS(VSS),.VDD(VDD),.Y(g5802),.A(I10445));
  NOT NOT1_2600(.VSS(VSS),.VDD(VDD),.Y(I10448),.A(g5335));
  NOT NOT1_2601(.VSS(VSS),.VDD(VDD),.Y(g5805),.A(I10448));
  NOT NOT1_2602(.VSS(VSS),.VDD(VDD),.Y(I10451),.A(g5216));
  NOT NOT1_2603(.VSS(VSS),.VDD(VDD),.Y(g5806),.A(I10451));
  NOT NOT1_2604(.VSS(VSS),.VDD(VDD),.Y(I10454),.A(g5217));
  NOT NOT1_2605(.VSS(VSS),.VDD(VDD),.Y(g5807),.A(I10454));
  NOT NOT1_2606(.VSS(VSS),.VDD(VDD),.Y(I10457),.A(g5218));
  NOT NOT1_2607(.VSS(VSS),.VDD(VDD),.Y(g5808),.A(I10457));
  NOT NOT1_2608(.VSS(VSS),.VDD(VDD),.Y(I10460),.A(g5219));
  NOT NOT1_2609(.VSS(VSS),.VDD(VDD),.Y(g5809),.A(I10460));
  NOT NOT1_2610(.VSS(VSS),.VDD(VDD),.Y(I10463),.A(g5220));
  NOT NOT1_2611(.VSS(VSS),.VDD(VDD),.Y(g5810),.A(I10463));
  NOT NOT1_2612(.VSS(VSS),.VDD(VDD),.Y(I10466),.A(g5221));
  NOT NOT1_2613(.VSS(VSS),.VDD(VDD),.Y(g5811),.A(I10466));
  NOT NOT1_2614(.VSS(VSS),.VDD(VDD),.Y(I10469),.A(g5222));
  NOT NOT1_2615(.VSS(VSS),.VDD(VDD),.Y(g5812),.A(I10469));
  NOT NOT1_2616(.VSS(VSS),.VDD(VDD),.Y(I10472),.A(g5223));
  NOT NOT1_2617(.VSS(VSS),.VDD(VDD),.Y(g5813),.A(I10472));
  NOT NOT1_2618(.VSS(VSS),.VDD(VDD),.Y(I10475),.A(g5529));
  NOT NOT1_2619(.VSS(VSS),.VDD(VDD),.Y(g5814),.A(I10475));
  NOT NOT1_2620(.VSS(VSS),.VDD(VDD),.Y(I10479),.A(g5227));
  NOT NOT1_2621(.VSS(VSS),.VDD(VDD),.Y(g5818),.A(I10479));
  NOT NOT1_2622(.VSS(VSS),.VDD(VDD),.Y(I10482),.A(g5228));
  NOT NOT1_2623(.VSS(VSS),.VDD(VDD),.Y(g5819),.A(I10482));
  NOT NOT1_2624(.VSS(VSS),.VDD(VDD),.Y(I10485),.A(g5229));
  NOT NOT1_2625(.VSS(VSS),.VDD(VDD),.Y(g5820),.A(I10485));
  NOT NOT1_2626(.VSS(VSS),.VDD(VDD),.Y(I10488),.A(g5230));
  NOT NOT1_2627(.VSS(VSS),.VDD(VDD),.Y(g5821),.A(I10488));
  NOT NOT1_2628(.VSS(VSS),.VDD(VDD),.Y(I10491),.A(g5231));
  NOT NOT1_2629(.VSS(VSS),.VDD(VDD),.Y(g5822),.A(I10491));
  NOT NOT1_2630(.VSS(VSS),.VDD(VDD),.Y(I10494),.A(g5232));
  NOT NOT1_2631(.VSS(VSS),.VDD(VDD),.Y(g5823),.A(I10494));
  NOT NOT1_2632(.VSS(VSS),.VDD(VDD),.Y(I10497),.A(g5233));
  NOT NOT1_2633(.VSS(VSS),.VDD(VDD),.Y(g5824),.A(I10497));
  NOT NOT1_2634(.VSS(VSS),.VDD(VDD),.Y(I10500),.A(g5234));
  NOT NOT1_2635(.VSS(VSS),.VDD(VDD),.Y(g5825),.A(I10500));
  NOT NOT1_2636(.VSS(VSS),.VDD(VDD),.Y(I10503),.A(g5235));
  NOT NOT1_2637(.VSS(VSS),.VDD(VDD),.Y(g5826),.A(I10503));
  NOT NOT1_2638(.VSS(VSS),.VDD(VDD),.Y(I10506),.A(g5236));
  NOT NOT1_2639(.VSS(VSS),.VDD(VDD),.Y(g5827),.A(I10506));
  NOT NOT1_2640(.VSS(VSS),.VDD(VDD),.Y(I10509),.A(g5237));
  NOT NOT1_2641(.VSS(VSS),.VDD(VDD),.Y(g5828),.A(I10509));
  NOT NOT1_2642(.VSS(VSS),.VDD(VDD),.Y(I10512),.A(g5238));
  NOT NOT1_2643(.VSS(VSS),.VDD(VDD),.Y(g5829),.A(I10512));
  NOT NOT1_2644(.VSS(VSS),.VDD(VDD),.Y(I10516),.A(g5241));
  NOT NOT1_2645(.VSS(VSS),.VDD(VDD),.Y(g5831),.A(I10516));
  NOT NOT1_2646(.VSS(VSS),.VDD(VDD),.Y(I10519),.A(g5242));
  NOT NOT1_2647(.VSS(VSS),.VDD(VDD),.Y(g5832),.A(I10519));
  NOT NOT1_2648(.VSS(VSS),.VDD(VDD),.Y(I10522),.A(g5243));
  NOT NOT1_2649(.VSS(VSS),.VDD(VDD),.Y(g5833),.A(I10522));
  NOT NOT1_2650(.VSS(VSS),.VDD(VDD),.Y(I10525),.A(g5244));
  NOT NOT1_2651(.VSS(VSS),.VDD(VDD),.Y(g5834),.A(I10525));
  NOT NOT1_2652(.VSS(VSS),.VDD(VDD),.Y(I10528),.A(g5245));
  NOT NOT1_2653(.VSS(VSS),.VDD(VDD),.Y(g5835),.A(I10528));
  NOT NOT1_2654(.VSS(VSS),.VDD(VDD),.Y(g5836),.A(g5529));
  NOT NOT1_2655(.VSS(VSS),.VDD(VDD),.Y(I10532),.A(g5253));
  NOT NOT1_2656(.VSS(VSS),.VDD(VDD),.Y(g5839),.A(I10532));
  NOT NOT1_2657(.VSS(VSS),.VDD(VDD),.Y(I10535),.A(g5254));
  NOT NOT1_2658(.VSS(VSS),.VDD(VDD),.Y(g5840),.A(I10535));
  NOT NOT1_2659(.VSS(VSS),.VDD(VDD),.Y(I10538),.A(g5255));
  NOT NOT1_2660(.VSS(VSS),.VDD(VDD),.Y(g5841),.A(I10538));
  NOT NOT1_2661(.VSS(VSS),.VDD(VDD),.Y(I10541),.A(g5256));
  NOT NOT1_2662(.VSS(VSS),.VDD(VDD),.Y(g5842),.A(I10541));
  NOT NOT1_2663(.VSS(VSS),.VDD(VDD),.Y(g5843),.A(g5367));
  NOT NOT1_2664(.VSS(VSS),.VDD(VDD),.Y(I10545),.A(g5259));
  NOT NOT1_2665(.VSS(VSS),.VDD(VDD),.Y(g5844),.A(I10545));
  NOT NOT1_2666(.VSS(VSS),.VDD(VDD),.Y(I10548),.A(g5260));
  NOT NOT1_2667(.VSS(VSS),.VDD(VDD),.Y(g5845),.A(I10548));
  NOT NOT1_2668(.VSS(VSS),.VDD(VDD),.Y(g5846),.A(g5367));
  NOT NOT1_2669(.VSS(VSS),.VDD(VDD),.Y(I10552),.A(g5396));
  NOT NOT1_2670(.VSS(VSS),.VDD(VDD),.Y(g5847),.A(I10552));
  NOT NOT1_2671(.VSS(VSS),.VDD(VDD),.Y(I10555),.A(g5529));
  NOT NOT1_2672(.VSS(VSS),.VDD(VDD),.Y(g5868),.A(I10555));
  NOT NOT1_2673(.VSS(VSS),.VDD(VDD),.Y(I10558),.A(g5264));
  NOT NOT1_2674(.VSS(VSS),.VDD(VDD),.Y(g5871),.A(I10558));
  NOT NOT1_2675(.VSS(VSS),.VDD(VDD),.Y(I10561),.A(g5265));
  NOT NOT1_2676(.VSS(VSS),.VDD(VDD),.Y(g5872),.A(I10561));
  NOT NOT1_2677(.VSS(VSS),.VDD(VDD),.Y(g5873),.A(g5367));
  NOT NOT1_2678(.VSS(VSS),.VDD(VDD),.Y(I10565),.A(g5402));
  NOT NOT1_2679(.VSS(VSS),.VDD(VDD),.Y(g5874),.A(I10565));
  NOT NOT1_2680(.VSS(VSS),.VDD(VDD),.Y(I10569),.A(g5417));
  NOT NOT1_2681(.VSS(VSS),.VDD(VDD),.Y(g5897),.A(I10569));
  NOT NOT1_2682(.VSS(VSS),.VDD(VDD),.Y(g5916),.A(g5384));
  NOT NOT1_2683(.VSS(VSS),.VDD(VDD),.Y(g5917),.A(g5412));
  NOT NOT1_2684(.VSS(VSS),.VDD(VDD),.Y(I10574),.A(g5426));
  NOT NOT1_2685(.VSS(VSS),.VDD(VDD),.Y(g5918),.A(I10574));
  NOT NOT1_2686(.VSS(VSS),.VDD(VDD),.Y(g5938),.A(g5412));
  NOT NOT1_2687(.VSS(VSS),.VDD(VDD),.Y(I10579),.A(g5433));
  NOT NOT1_2688(.VSS(VSS),.VDD(VDD),.Y(g5939),.A(I10579));
  NOT NOT1_2689(.VSS(VSS),.VDD(VDD),.Y(I10582),.A(g5437));
  NOT NOT1_2690(.VSS(VSS),.VDD(VDD),.Y(g5956),.A(I10582));
  NOT NOT1_2691(.VSS(VSS),.VDD(VDD),.Y(I10587),.A(g5439));
  NOT NOT1_2692(.VSS(VSS),.VDD(VDD),.Y(g5971),.A(I10587));
  NOT NOT1_2693(.VSS(VSS),.VDD(VDD),.Y(g5987),.A(g5294));
  NOT NOT1_2694(.VSS(VSS),.VDD(VDD),.Y(I10592),.A(g5444));
  NOT NOT1_2695(.VSS(VSS),.VDD(VDD),.Y(g5988),.A(I10592));
  NOT NOT1_2696(.VSS(VSS),.VDD(VDD),.Y(g6004),.A(g5494));
  NOT NOT1_2697(.VSS(VSS),.VDD(VDD),.Y(g6007),.A(g5494));
  NOT NOT1_2698(.VSS(VSS),.VDD(VDD),.Y(g6008),.A(g5367));
  NOT NOT1_2699(.VSS(VSS),.VDD(VDD),.Y(I10605),.A(g5440));
  NOT NOT1_2700(.VSS(VSS),.VDD(VDD),.Y(g6009),.A(I10605));
  NOT NOT1_2701(.VSS(VSS),.VDD(VDD),.Y(I10608),.A(g5701));
  NOT NOT1_2702(.VSS(VSS),.VDD(VDD),.Y(g6010),.A(I10608));
  NOT NOT1_2703(.VSS(VSS),.VDD(VDD),.Y(g6011),.A(g5494));
  NOT NOT1_2704(.VSS(VSS),.VDD(VDD),.Y(g6012),.A(g5367));
  NOT NOT1_2705(.VSS(VSS),.VDD(VDD),.Y(I10614),.A(g5302));
  NOT NOT1_2706(.VSS(VSS),.VDD(VDD),.Y(g6014),.A(I10614));
  NOT NOT1_2707(.VSS(VSS),.VDD(VDD),.Y(I10617),.A(g5677));
  NOT NOT1_2708(.VSS(VSS),.VDD(VDD),.Y(g6015),.A(I10617));
  NOT NOT1_2709(.VSS(VSS),.VDD(VDD),.Y(g6018),.A(g5494));
  NOT NOT1_2710(.VSS(VSS),.VDD(VDD),.Y(g6019),.A(g5367));
  NOT NOT1_2711(.VSS(VSS),.VDD(VDD),.Y(g6020),.A(g5367));
  NOT NOT1_2712(.VSS(VSS),.VDD(VDD),.Y(g6024),.A(g5494));
  NOT NOT1_2713(.VSS(VSS),.VDD(VDD),.Y(g6025),.A(g5367));
  NOT NOT1_2714(.VSS(VSS),.VDD(VDD),.Y(g6026),.A(g5384));
  NOT NOT1_2715(.VSS(VSS),.VDD(VDD),.Y(g6027),.A(g5384));
  NOT NOT1_2716(.VSS(VSS),.VDD(VDD),.Y(g6028),.A(g5529));
  NOT NOT1_2717(.VSS(VSS),.VDD(VDD),.Y(g6032),.A(g5494));
  NOT NOT1_2718(.VSS(VSS),.VDD(VDD),.Y(g6033),.A(g5384));
  NOT NOT1_2719(.VSS(VSS),.VDD(VDD),.Y(I10639),.A(g5224));
  NOT NOT1_2720(.VSS(VSS),.VDD(VDD),.Y(g6034),.A(I10639));
  NOT NOT1_2721(.VSS(VSS),.VDD(VDD),.Y(g6035),.A(g5494));
  NOT NOT1_2722(.VSS(VSS),.VDD(VDD),.Y(I10643),.A(g5267));
  NOT NOT1_2723(.VSS(VSS),.VDD(VDD),.Y(g6036),.A(I10643));
  NOT NOT1_2724(.VSS(VSS),.VDD(VDD),.Y(I10646),.A(g5364));
  NOT NOT1_2725(.VSS(VSS),.VDD(VDD),.Y(g6037),.A(I10646));
  NOT NOT1_2726(.VSS(VSS),.VDD(VDD),.Y(I10649),.A(g5657));
  NOT NOT1_2727(.VSS(VSS),.VDD(VDD),.Y(g6038),.A(I10649));
  NOT NOT1_2728(.VSS(VSS),.VDD(VDD),.Y(g6048),.A(g5246));
  NOT NOT1_2729(.VSS(VSS),.VDD(VDD),.Y(g6050),.A(g5246));
  NOT NOT1_2730(.VSS(VSS),.VDD(VDD),.Y(g6051),.A(g5246));
  NOT NOT1_2731(.VSS(VSS),.VDD(VDD),.Y(g6059),.A(g5317));
  NOT NOT1_2732(.VSS(VSS),.VDD(VDD),.Y(I10675),.A(g5662));
  NOT NOT1_2733(.VSS(VSS),.VDD(VDD),.Y(g6062),.A(I10675));
  NOT NOT1_2734(.VSS(VSS),.VDD(VDD),.Y(I10678),.A(g5566));
  NOT NOT1_2735(.VSS(VSS),.VDD(VDD),.Y(g6063),.A(I10678));
  NOT NOT1_2736(.VSS(VSS),.VDD(VDD),.Y(I10681),.A(g5686));
  NOT NOT1_2737(.VSS(VSS),.VDD(VDD),.Y(g6064),.A(I10681));
  NOT NOT1_2738(.VSS(VSS),.VDD(VDD),.Y(I10684),.A(g5258));
  NOT NOT1_2739(.VSS(VSS),.VDD(VDD),.Y(g6065),.A(I10684));
  NOT NOT1_2740(.VSS(VSS),.VDD(VDD),.Y(I10687),.A(g5674));
  NOT NOT1_2741(.VSS(VSS),.VDD(VDD),.Y(g6068),.A(I10687));
  NOT NOT1_2742(.VSS(VSS),.VDD(VDD),.Y(I10690),.A(g5538));
  NOT NOT1_2743(.VSS(VSS),.VDD(VDD),.Y(g6069),.A(I10690));
  NOT NOT1_2744(.VSS(VSS),.VDD(VDD),.Y(g6070),.A(g5317));
  NOT NOT1_2745(.VSS(VSS),.VDD(VDD),.Y(I10694),.A(g5445));
  NOT NOT1_2746(.VSS(VSS),.VDD(VDD),.Y(g6071),.A(I10694));
  NOT NOT1_2747(.VSS(VSS),.VDD(VDD),.Y(g6072),.A(g5345));
  NOT NOT1_2748(.VSS(VSS),.VDD(VDD),.Y(g6073),.A(g5384));
  NOT NOT1_2749(.VSS(VSS),.VDD(VDD),.Y(g6074),.A(g5317));
  NOT NOT1_2750(.VSS(VSS),.VDD(VDD),.Y(g6075),.A(g5345));
  NOT NOT1_2751(.VSS(VSS),.VDD(VDD),.Y(g6076),.A(g5287));
  NOT NOT1_2752(.VSS(VSS),.VDD(VDD),.Y(I10702),.A(g5529));
  NOT NOT1_2753(.VSS(VSS),.VDD(VDD),.Y(g6083),.A(I10702));
  NOT NOT1_2754(.VSS(VSS),.VDD(VDD),.Y(I10705),.A(g5463));
  NOT NOT1_2755(.VSS(VSS),.VDD(VDD),.Y(g6087),.A(I10705));
  NOT NOT1_2756(.VSS(VSS),.VDD(VDD),.Y(I10708),.A(g5545));
  NOT NOT1_2757(.VSS(VSS),.VDD(VDD),.Y(g6088),.A(I10708));
  NOT NOT1_2758(.VSS(VSS),.VDD(VDD),.Y(g6089),.A(g5317));
  NOT NOT1_2759(.VSS(VSS),.VDD(VDD),.Y(g6090),.A(g5529));
  NOT NOT1_2760(.VSS(VSS),.VDD(VDD),.Y(g6092),.A(g5317));
  NOT NOT1_2761(.VSS(VSS),.VDD(VDD),.Y(g6093),.A(g5345));
  NOT NOT1_2762(.VSS(VSS),.VDD(VDD),.Y(I10716),.A(g5537));
  NOT NOT1_2763(.VSS(VSS),.VDD(VDD),.Y(g6094),.A(I10716));
  NOT NOT1_2764(.VSS(VSS),.VDD(VDD),.Y(I10719),.A(g5559));
  NOT NOT1_2765(.VSS(VSS),.VDD(VDD),.Y(g6095),.A(I10719));
  NOT NOT1_2766(.VSS(VSS),.VDD(VDD),.Y(g6096),.A(g5317));
  NOT NOT1_2767(.VSS(VSS),.VDD(VDD),.Y(g6097),.A(g5345));
  NOT NOT1_2768(.VSS(VSS),.VDD(VDD),.Y(g6101),.A(g5317));
  NOT NOT1_2769(.VSS(VSS),.VDD(VDD),.Y(g6102),.A(g5345));
  NOT NOT1_2770(.VSS(VSS),.VDD(VDD),.Y(g6103),.A(g5317));
  NOT NOT1_2771(.VSS(VSS),.VDD(VDD),.Y(g6104),.A(g5345));
  NOT NOT1_2772(.VSS(VSS),.VDD(VDD),.Y(g6106),.A(g5345));
  NOT NOT1_2773(.VSS(VSS),.VDD(VDD),.Y(g6108),.A(g5345));
  NOT NOT1_2774(.VSS(VSS),.VDD(VDD),.Y(g6110),.A(g5335));
  NOT NOT1_2775(.VSS(VSS),.VDD(VDD),.Y(g6111),.A(g5453));
  NOT NOT1_2776(.VSS(VSS),.VDD(VDD),.Y(I10739),.A(g5572));
  NOT NOT1_2777(.VSS(VSS),.VDD(VDD),.Y(g6117),.A(I10739));
  NOT NOT1_2778(.VSS(VSS),.VDD(VDD),.Y(g6118),.A(g5549));
  NOT NOT1_2779(.VSS(VSS),.VDD(VDD),.Y(I10752),.A(g5618));
  NOT NOT1_2780(.VSS(VSS),.VDD(VDD),.Y(g6122),.A(I10752));
  NOT NOT1_2781(.VSS(VSS),.VDD(VDD),.Y(I10758),.A(g5662));
  NOT NOT1_2782(.VSS(VSS),.VDD(VDD),.Y(g6129),.A(I10758));
  NOT NOT1_2783(.VSS(VSS),.VDD(VDD),.Y(I10761),.A(g5302));
  NOT NOT1_2784(.VSS(VSS),.VDD(VDD),.Y(g6130),.A(I10761));
  NOT NOT1_2785(.VSS(VSS),.VDD(VDD),.Y(g6131),.A(g5529));
  NOT NOT1_2786(.VSS(VSS),.VDD(VDD),.Y(I10766),.A(g5674));
  NOT NOT1_2787(.VSS(VSS),.VDD(VDD),.Y(g6133),.A(I10766));
  NOT NOT1_2788(.VSS(VSS),.VDD(VDD),.Y(g6134),.A(g5428));
  NOT NOT1_2789(.VSS(VSS),.VDD(VDD),.Y(I10770),.A(g5441));
  NOT NOT1_2790(.VSS(VSS),.VDD(VDD),.Y(g6135),.A(I10770));
  NOT NOT1_2791(.VSS(VSS),.VDD(VDD),.Y(I10773),.A(g5708));
  NOT NOT1_2792(.VSS(VSS),.VDD(VDD),.Y(g6136),.A(I10773));
  NOT NOT1_2793(.VSS(VSS),.VDD(VDD),.Y(I10776),.A(g5576));
  NOT NOT1_2794(.VSS(VSS),.VDD(VDD),.Y(g6137),.A(I10776));
  NOT NOT1_2795(.VSS(VSS),.VDD(VDD),.Y(I10780),.A(g5445));
  NOT NOT1_2796(.VSS(VSS),.VDD(VDD),.Y(g6139),.A(I10780));
  NOT NOT1_2797(.VSS(VSS),.VDD(VDD),.Y(I10783),.A(g5542));
  NOT NOT1_2798(.VSS(VSS),.VDD(VDD),.Y(g6140),.A(I10783));
  NOT NOT1_2799(.VSS(VSS),.VDD(VDD),.Y(I10786),.A(g5452));
  NOT NOT1_2800(.VSS(VSS),.VDD(VDD),.Y(g6141),.A(I10786));
  NOT NOT1_2801(.VSS(VSS),.VDD(VDD),.Y(I10796),.A(g5397));
  NOT NOT1_2802(.VSS(VSS),.VDD(VDD),.Y(g6143),.A(I10796));
  NOT NOT1_2803(.VSS(VSS),.VDD(VDD),.Y(I10801),.A(g5463));
  NOT NOT1_2804(.VSS(VSS),.VDD(VDD),.Y(g6146),.A(I10801));
  NOT NOT1_2805(.VSS(VSS),.VDD(VDD),.Y(I10804),.A(g5526));
  NOT NOT1_2806(.VSS(VSS),.VDD(VDD),.Y(g6147),.A(I10804));
  NOT NOT1_2807(.VSS(VSS),.VDD(VDD),.Y(I10807),.A(g5294));
  NOT NOT1_2808(.VSS(VSS),.VDD(VDD),.Y(g6148),.A(I10807));
  NOT NOT1_2809(.VSS(VSS),.VDD(VDD),.Y(I10810),.A(g5403));
  NOT NOT1_2810(.VSS(VSS),.VDD(VDD),.Y(g6149),.A(I10810));
  NOT NOT1_2811(.VSS(VSS),.VDD(VDD),.Y(g6150),.A(g5287));
  NOT NOT1_2812(.VSS(VSS),.VDD(VDD),.Y(I10815),.A(g5418));
  NOT NOT1_2813(.VSS(VSS),.VDD(VDD),.Y(g6152),.A(I10815));
  NOT NOT1_2814(.VSS(VSS),.VDD(VDD),.Y(I10826),.A(g5434));
  NOT NOT1_2815(.VSS(VSS),.VDD(VDD),.Y(g6155),.A(I10826));
  NOT NOT1_2816(.VSS(VSS),.VDD(VDD),.Y(I10829),.A(g5224));
  NOT NOT1_2817(.VSS(VSS),.VDD(VDD),.Y(g6156),.A(I10829));
  NOT NOT1_2818(.VSS(VSS),.VDD(VDD),.Y(I10842),.A(g5701));
  NOT NOT1_2819(.VSS(VSS),.VDD(VDD),.Y(g6161),.A(I10842));
  NOT NOT1_2820(.VSS(VSS),.VDD(VDD),.Y(I10862),.A(g5364));
  NOT NOT1_2821(.VSS(VSS),.VDD(VDD),.Y(g6167),.A(I10862));
  NOT NOT1_2822(.VSS(VSS),.VDD(VDD),.Y(I10882),.A(g5600));
  NOT NOT1_2823(.VSS(VSS),.VDD(VDD),.Y(g6173),.A(I10882));
  NOT NOT1_2824(.VSS(VSS),.VDD(VDD),.Y(I10896),.A(g5475));
  NOT NOT1_2825(.VSS(VSS),.VDD(VDD),.Y(g6179),.A(I10896));
  NOT NOT1_2826(.VSS(VSS),.VDD(VDD),.Y(I10914),.A(g5448));
  NOT NOT1_2827(.VSS(VSS),.VDD(VDD),.Y(g6183),.A(I10914));
  NOT NOT1_2828(.VSS(VSS),.VDD(VDD),.Y(I10919),.A(g5479));
  NOT NOT1_2829(.VSS(VSS),.VDD(VDD),.Y(g6186),.A(I10919));
  NOT NOT1_2830(.VSS(VSS),.VDD(VDD),.Y(I10930),.A(g5600));
  NOT NOT1_2831(.VSS(VSS),.VDD(VDD),.Y(g6189),.A(I10930));
  NOT NOT1_2832(.VSS(VSS),.VDD(VDD),.Y(I10933),.A(g5668));
  NOT NOT1_2833(.VSS(VSS),.VDD(VDD),.Y(g6190),.A(I10933));
  NOT NOT1_2834(.VSS(VSS),.VDD(VDD),.Y(I10937),.A(g5560));
  NOT NOT1_2835(.VSS(VSS),.VDD(VDD),.Y(g6194),.A(I10937));
  NOT NOT1_2836(.VSS(VSS),.VDD(VDD),.Y(I10940),.A(g5489));
  NOT NOT1_2837(.VSS(VSS),.VDD(VDD),.Y(g6195),.A(I10940));
  NOT NOT1_2838(.VSS(VSS),.VDD(VDD),.Y(g6198),.A(g5335));
  NOT NOT1_2839(.VSS(VSS),.VDD(VDD),.Y(I10946),.A(g5563));
  NOT NOT1_2840(.VSS(VSS),.VDD(VDD),.Y(g6201),.A(I10946));
  NOT NOT1_2841(.VSS(VSS),.VDD(VDD),.Y(I10949),.A(g5513));
  NOT NOT1_2842(.VSS(VSS),.VDD(VDD),.Y(g6202),.A(I10949));
  NOT NOT1_2843(.VSS(VSS),.VDD(VDD),.Y(g6205),.A(g5628));
  NOT NOT1_2844(.VSS(VSS),.VDD(VDD),.Y(g6206),.A(g5639));
  NOT NOT1_2845(.VSS(VSS),.VDD(VDD),.Y(I10962),.A(g5719));
  NOT NOT1_2846(.VSS(VSS),.VDD(VDD),.Y(g6207),.A(I10962));
  NOT NOT1_2847(.VSS(VSS),.VDD(VDD),.Y(I10965),.A(g5719));
  NOT NOT1_2848(.VSS(VSS),.VDD(VDD),.Y(g6208),.A(I10965));
  NOT NOT1_2849(.VSS(VSS),.VDD(VDD),.Y(I10969),.A(g5606));
  NOT NOT1_2850(.VSS(VSS),.VDD(VDD),.Y(g6210),.A(I10969));
  NOT NOT1_2851(.VSS(VSS),.VDD(VDD),.Y(g6211),.A(g5645));
  NOT NOT1_2852(.VSS(VSS),.VDD(VDD),.Y(I10973),.A(g5726));
  NOT NOT1_2853(.VSS(VSS),.VDD(VDD),.Y(g6212),.A(I10973));
  NOT NOT1_2854(.VSS(VSS),.VDD(VDD),.Y(I10976),.A(g5726));
  NOT NOT1_2855(.VSS(VSS),.VDD(VDD),.Y(g6213),.A(I10976));
  NOT NOT1_2856(.VSS(VSS),.VDD(VDD),.Y(I10987),.A(g5609));
  NOT NOT1_2857(.VSS(VSS),.VDD(VDD),.Y(g6216),.A(I10987));
  NOT NOT1_2858(.VSS(VSS),.VDD(VDD),.Y(g6217),.A(g5649));
  NOT NOT1_2859(.VSS(VSS),.VDD(VDD),.Y(I10998),.A(g5672));
  NOT NOT1_2860(.VSS(VSS),.VDD(VDD),.Y(g6219),.A(I10998));
  NOT NOT1_2861(.VSS(VSS),.VDD(VDD),.Y(I11001),.A(g5698));
  NOT NOT1_2862(.VSS(VSS),.VDD(VDD),.Y(g6220),.A(I11001));
  NOT NOT1_2863(.VSS(VSS),.VDD(VDD),.Y(I11004),.A(g5613));
  NOT NOT1_2864(.VSS(VSS),.VDD(VDD),.Y(g6221),.A(I11004));
  NOT NOT1_2865(.VSS(VSS),.VDD(VDD),.Y(g6222),.A(g5654));
  NOT NOT1_2866(.VSS(VSS),.VDD(VDD),.Y(I11008),.A(g5693));
  NOT NOT1_2867(.VSS(VSS),.VDD(VDD),.Y(g6223),.A(I11008));
  NOT NOT1_2868(.VSS(VSS),.VDD(VDD),.Y(I11011),.A(g5693));
  NOT NOT1_2869(.VSS(VSS),.VDD(VDD),.Y(g6224),.A(I11011));
  NOT NOT1_2870(.VSS(VSS),.VDD(VDD),.Y(I11014),.A(g5621));
  NOT NOT1_2871(.VSS(VSS),.VDD(VDD),.Y(g6225),.A(I11014));
  NOT NOT1_2872(.VSS(VSS),.VDD(VDD),.Y(g6226),.A(g5658));
  NOT NOT1_2873(.VSS(VSS),.VDD(VDD),.Y(I11018),.A(g5626));
  NOT NOT1_2874(.VSS(VSS),.VDD(VDD),.Y(g6227),.A(I11018));
  NOT NOT1_2875(.VSS(VSS),.VDD(VDD),.Y(I11021),.A(g5627));
  NOT NOT1_2876(.VSS(VSS),.VDD(VDD),.Y(g6228),.A(I11021));
  NOT NOT1_2877(.VSS(VSS),.VDD(VDD),.Y(g6229),.A(g5665));
  NOT NOT1_2878(.VSS(VSS),.VDD(VDD),.Y(I11025),.A(g5638));
  NOT NOT1_2879(.VSS(VSS),.VDD(VDD),.Y(g6230),.A(I11025));
  NOT NOT1_2880(.VSS(VSS),.VDD(VDD),.Y(I11028),.A(g5642));
  NOT NOT1_2881(.VSS(VSS),.VDD(VDD),.Y(g6231),.A(I11028));
  NOT NOT1_2882(.VSS(VSS),.VDD(VDD),.Y(I11031),.A(g5335));
  NOT NOT1_2883(.VSS(VSS),.VDD(VDD),.Y(g6232),.A(I11031));
  NOT NOT1_2884(.VSS(VSS),.VDD(VDD),.Y(I11034),.A(g5644));
  NOT NOT1_2885(.VSS(VSS),.VDD(VDD),.Y(g6235),.A(I11034));
  NOT NOT1_2886(.VSS(VSS),.VDD(VDD),.Y(I11037),.A(g5299));
  NOT NOT1_2887(.VSS(VSS),.VDD(VDD),.Y(g6236),.A(I11037));
  NOT NOT1_2888(.VSS(VSS),.VDD(VDD),.Y(I11040),.A(g5299));
  NOT NOT1_2889(.VSS(VSS),.VDD(VDD),.Y(g6237),.A(I11040));
  NOT NOT1_2890(.VSS(VSS),.VDD(VDD),.Y(I11043),.A(g5648));
  NOT NOT1_2891(.VSS(VSS),.VDD(VDD),.Y(g6238),.A(I11043));
  NOT NOT1_2892(.VSS(VSS),.VDD(VDD),.Y(I11047),.A(g5653));
  NOT NOT1_2893(.VSS(VSS),.VDD(VDD),.Y(g6242),.A(I11047));
  NOT NOT1_2894(.VSS(VSS),.VDD(VDD),.Y(I11050),.A(g5335));
  NOT NOT1_2895(.VSS(VSS),.VDD(VDD),.Y(g6243),.A(I11050));
  NOT NOT1_2896(.VSS(VSS),.VDD(VDD),.Y(g6244),.A(g5670));
  NOT NOT1_2897(.VSS(VSS),.VDD(VDD),.Y(g6245),.A(g5690));
  NOT NOT1_2898(.VSS(VSS),.VDD(VDD),.Y(I11055),.A(g5696));
  NOT NOT1_2899(.VSS(VSS),.VDD(VDD),.Y(g6246),.A(I11055));
  NOT NOT1_2900(.VSS(VSS),.VDD(VDD),.Y(g6250),.A(g5679));
  NOT NOT1_2901(.VSS(VSS),.VDD(VDD),.Y(I11060),.A(g5453));
  NOT NOT1_2902(.VSS(VSS),.VDD(VDD),.Y(g6251),.A(I11060));
  NOT NOT1_2903(.VSS(VSS),.VDD(VDD),.Y(g6252),.A(g5418));
  NOT NOT1_2904(.VSS(VSS),.VDD(VDD),.Y(g6253),.A(g5403));
  NOT NOT1_2905(.VSS(VSS),.VDD(VDD),.Y(g6254),.A(g5683));
  NOT NOT1_2906(.VSS(VSS),.VDD(VDD),.Y(I11066),.A(g5460));
  NOT NOT1_2907(.VSS(VSS),.VDD(VDD),.Y(g6255),.A(I11066));
  NOT NOT1_2908(.VSS(VSS),.VDD(VDD),.Y(I11069),.A(g5671));
  NOT NOT1_2909(.VSS(VSS),.VDD(VDD),.Y(g6256),.A(I11069));
  NOT NOT1_2910(.VSS(VSS),.VDD(VDD),.Y(g6257),.A(g5685));
  NOT NOT1_2911(.VSS(VSS),.VDD(VDD),.Y(g6258),.A(g5427));
  NOT NOT1_2912(.VSS(VSS),.VDD(VDD),.Y(g6263),.A(g5688));
  NOT NOT1_2913(.VSS(VSS),.VDD(VDD),.Y(g6264),.A(g5403));
  NOT NOT1_2914(.VSS(VSS),.VDD(VDD),.Y(I11086),.A(g5397));
  NOT NOT1_2915(.VSS(VSS),.VDD(VDD),.Y(g6267),.A(I11086));
  NOT NOT1_2916(.VSS(VSS),.VDD(VDD),.Y(I11090),.A(g1000));
  NOT NOT1_2917(.VSS(VSS),.VDD(VDD),.Y(g6269),.A(I11090));
  NOT NOT1_2918(.VSS(VSS),.VDD(VDD),.Y(I11129),.A(g5418));
  NOT NOT1_2919(.VSS(VSS),.VDD(VDD),.Y(g6278),.A(I11129));
  NOT NOT1_2920(.VSS(VSS),.VDD(VDD),.Y(I11132),.A(g5624));
  NOT NOT1_2921(.VSS(VSS),.VDD(VDD),.Y(g6279),.A(I11132));
  NOT NOT1_2922(.VSS(VSS),.VDD(VDD),.Y(I11191),.A(g6155));
  NOT NOT1_2923(.VSS(VSS),.VDD(VDD),.Y(g6288),.A(I11191));
  NOT NOT1_2924(.VSS(VSS),.VDD(VDD),.Y(I11194),.A(g6243));
  NOT NOT1_2925(.VSS(VSS),.VDD(VDD),.Y(g6289),.A(I11194));
  NOT NOT1_2926(.VSS(VSS),.VDD(VDD),.Y(I11197),.A(g6122));
  NOT NOT1_2927(.VSS(VSS),.VDD(VDD),.Y(g6290),.A(I11197));
  NOT NOT1_2928(.VSS(VSS),.VDD(VDD),.Y(I11200),.A(g6251));
  NOT NOT1_2929(.VSS(VSS),.VDD(VDD),.Y(g6291),.A(I11200));
  NOT NOT1_2930(.VSS(VSS),.VDD(VDD),.Y(I11203),.A(g6129));
  NOT NOT1_2931(.VSS(VSS),.VDD(VDD),.Y(g6292),.A(I11203));
  NOT NOT1_2932(.VSS(VSS),.VDD(VDD),.Y(I11206),.A(g6133));
  NOT NOT1_2933(.VSS(VSS),.VDD(VDD),.Y(g6293),.A(I11206));
  NOT NOT1_2934(.VSS(VSS),.VDD(VDD),.Y(I11209),.A(g6139));
  NOT NOT1_2935(.VSS(VSS),.VDD(VDD),.Y(g6294),.A(I11209));
  NOT NOT1_2936(.VSS(VSS),.VDD(VDD),.Y(I11212),.A(g6146));
  NOT NOT1_2937(.VSS(VSS),.VDD(VDD),.Y(g6295),.A(I11212));
  NOT NOT1_2938(.VSS(VSS),.VDD(VDD),.Y(I11215),.A(g6156));
  NOT NOT1_2939(.VSS(VSS),.VDD(VDD),.Y(g6296),.A(I11215));
  NOT NOT1_2940(.VSS(VSS),.VDD(VDD),.Y(I11218),.A(g6161));
  NOT NOT1_2941(.VSS(VSS),.VDD(VDD),.Y(g6297),.A(I11218));
  NOT NOT1_2942(.VSS(VSS),.VDD(VDD),.Y(I11221),.A(g6167));
  NOT NOT1_2943(.VSS(VSS),.VDD(VDD),.Y(g6298),.A(I11221));
  NOT NOT1_2944(.VSS(VSS),.VDD(VDD),.Y(I11224),.A(g6255));
  NOT NOT1_2945(.VSS(VSS),.VDD(VDD),.Y(g6299),.A(I11224));
  NOT NOT1_2946(.VSS(VSS),.VDD(VDD),.Y(I11227),.A(g6130));
  NOT NOT1_2947(.VSS(VSS),.VDD(VDD),.Y(g6300),.A(I11227));
  NOT NOT1_2948(.VSS(VSS),.VDD(VDD),.Y(I11230),.A(g6140));
  NOT NOT1_2949(.VSS(VSS),.VDD(VDD),.Y(g6301),.A(I11230));
  NOT NOT1_2950(.VSS(VSS),.VDD(VDD),.Y(I11233),.A(g6147));
  NOT NOT1_2951(.VSS(VSS),.VDD(VDD),.Y(g6302),.A(I11233));
  NOT NOT1_2952(.VSS(VSS),.VDD(VDD),.Y(I11236),.A(g6148));
  NOT NOT1_2953(.VSS(VSS),.VDD(VDD),.Y(g6303),.A(I11236));
  NOT NOT1_2954(.VSS(VSS),.VDD(VDD),.Y(I11239),.A(g6173));
  NOT NOT1_2955(.VSS(VSS),.VDD(VDD),.Y(g6304),.A(I11239));
  NOT NOT1_2956(.VSS(VSS),.VDD(VDD),.Y(I11242),.A(g6183));
  NOT NOT1_2957(.VSS(VSS),.VDD(VDD),.Y(g6305),.A(I11242));
  NOT NOT1_2958(.VSS(VSS),.VDD(VDD),.Y(I11245),.A(g6143));
  NOT NOT1_2959(.VSS(VSS),.VDD(VDD),.Y(g6306),.A(I11245));
  NOT NOT1_2960(.VSS(VSS),.VDD(VDD),.Y(I11248),.A(g6149));
  NOT NOT1_2961(.VSS(VSS),.VDD(VDD),.Y(g6307),.A(I11248));
  NOT NOT1_2962(.VSS(VSS),.VDD(VDD),.Y(I11251),.A(g6152));
  NOT NOT1_2963(.VSS(VSS),.VDD(VDD),.Y(g6308),.A(I11251));
  NOT NOT1_2964(.VSS(VSS),.VDD(VDD),.Y(I11254),.A(g5793));
  NOT NOT1_2965(.VSS(VSS),.VDD(VDD),.Y(g6309),.A(I11254));
  NOT NOT1_2966(.VSS(VSS),.VDD(VDD),.Y(I11257),.A(g5805));
  NOT NOT1_2967(.VSS(VSS),.VDD(VDD),.Y(g6310),.A(I11257));
  NOT NOT1_2968(.VSS(VSS),.VDD(VDD),.Y(I11260),.A(g5779));
  NOT NOT1_2969(.VSS(VSS),.VDD(VDD),.Y(g6311),.A(I11260));
  NOT NOT1_2970(.VSS(VSS),.VDD(VDD),.Y(I11263),.A(g5784));
  NOT NOT1_2971(.VSS(VSS),.VDD(VDD),.Y(g6312),.A(I11263));
  NOT NOT1_2972(.VSS(VSS),.VDD(VDD),.Y(I11266),.A(g5794));
  NOT NOT1_2973(.VSS(VSS),.VDD(VDD),.Y(g6313),.A(I11266));
  NOT NOT1_2974(.VSS(VSS),.VDD(VDD),.Y(I11269),.A(g5756));
  NOT NOT1_2975(.VSS(VSS),.VDD(VDD),.Y(g6314),.A(I11269));
  NOT NOT1_2976(.VSS(VSS),.VDD(VDD),.Y(I11272),.A(g5758));
  NOT NOT1_2977(.VSS(VSS),.VDD(VDD),.Y(g6315),.A(I11272));
  NOT NOT1_2978(.VSS(VSS),.VDD(VDD),.Y(I11275),.A(g5768));
  NOT NOT1_2979(.VSS(VSS),.VDD(VDD),.Y(g6316),.A(I11275));
  NOT NOT1_2980(.VSS(VSS),.VDD(VDD),.Y(I11278),.A(g5780));
  NOT NOT1_2981(.VSS(VSS),.VDD(VDD),.Y(g6317),.A(I11278));
  NOT NOT1_2982(.VSS(VSS),.VDD(VDD),.Y(I11281),.A(g5785));
  NOT NOT1_2983(.VSS(VSS),.VDD(VDD),.Y(g6318),.A(I11281));
  NOT NOT1_2984(.VSS(VSS),.VDD(VDD),.Y(I11284),.A(g5795));
  NOT NOT1_2985(.VSS(VSS),.VDD(VDD),.Y(g6319),.A(I11284));
  NOT NOT1_2986(.VSS(VSS),.VDD(VDD),.Y(I11287),.A(g5806));
  NOT NOT1_2987(.VSS(VSS),.VDD(VDD),.Y(g6320),.A(I11287));
  NOT NOT1_2988(.VSS(VSS),.VDD(VDD),.Y(I11290),.A(g5818));
  NOT NOT1_2989(.VSS(VSS),.VDD(VDD),.Y(g6321),.A(I11290));
  NOT NOT1_2990(.VSS(VSS),.VDD(VDD),.Y(I11293),.A(g5824));
  NOT NOT1_2991(.VSS(VSS),.VDD(VDD),.Y(g6322),.A(I11293));
  NOT NOT1_2992(.VSS(VSS),.VDD(VDD),.Y(I11296),.A(g5831));
  NOT NOT1_2993(.VSS(VSS),.VDD(VDD),.Y(g6323),.A(I11296));
  NOT NOT1_2994(.VSS(VSS),.VDD(VDD),.Y(I11299),.A(g5786));
  NOT NOT1_2995(.VSS(VSS),.VDD(VDD),.Y(g6324),.A(I11299));
  NOT NOT1_2996(.VSS(VSS),.VDD(VDD),.Y(I11302),.A(g5796));
  NOT NOT1_2997(.VSS(VSS),.VDD(VDD),.Y(g6325),.A(I11302));
  NOT NOT1_2998(.VSS(VSS),.VDD(VDD),.Y(I11305),.A(g5807));
  NOT NOT1_2999(.VSS(VSS),.VDD(VDD),.Y(g6326),.A(I11305));
  NOT NOT1_3000(.VSS(VSS),.VDD(VDD),.Y(I11308),.A(g5759));
  NOT NOT1_3001(.VSS(VSS),.VDD(VDD),.Y(g6327),.A(I11308));
  NOT NOT1_3002(.VSS(VSS),.VDD(VDD),.Y(I11311),.A(g5760));
  NOT NOT1_3003(.VSS(VSS),.VDD(VDD),.Y(g6328),.A(I11311));
  NOT NOT1_3004(.VSS(VSS),.VDD(VDD),.Y(I11314),.A(g5781));
  NOT NOT1_3005(.VSS(VSS),.VDD(VDD),.Y(g6329),.A(I11314));
  NOT NOT1_3006(.VSS(VSS),.VDD(VDD),.Y(I11317),.A(g5787));
  NOT NOT1_3007(.VSS(VSS),.VDD(VDD),.Y(g6330),.A(I11317));
  NOT NOT1_3008(.VSS(VSS),.VDD(VDD),.Y(I11320),.A(g5797));
  NOT NOT1_3009(.VSS(VSS),.VDD(VDD),.Y(g6331),.A(I11320));
  NOT NOT1_3010(.VSS(VSS),.VDD(VDD),.Y(I11323),.A(g5808));
  NOT NOT1_3011(.VSS(VSS),.VDD(VDD),.Y(g6332),.A(I11323));
  NOT NOT1_3012(.VSS(VSS),.VDD(VDD),.Y(I11326),.A(g5819));
  NOT NOT1_3013(.VSS(VSS),.VDD(VDD),.Y(g6333),.A(I11326));
  NOT NOT1_3014(.VSS(VSS),.VDD(VDD),.Y(I11329),.A(g5825));
  NOT NOT1_3015(.VSS(VSS),.VDD(VDD),.Y(g6334),.A(I11329));
  NOT NOT1_3016(.VSS(VSS),.VDD(VDD),.Y(I11332),.A(g5832));
  NOT NOT1_3017(.VSS(VSS),.VDD(VDD),.Y(g6335),.A(I11332));
  NOT NOT1_3018(.VSS(VSS),.VDD(VDD),.Y(I11335),.A(g5839));
  NOT NOT1_3019(.VSS(VSS),.VDD(VDD),.Y(g6336),.A(I11335));
  NOT NOT1_3020(.VSS(VSS),.VDD(VDD),.Y(I11338),.A(g5798));
  NOT NOT1_3021(.VSS(VSS),.VDD(VDD),.Y(g6337),.A(I11338));
  NOT NOT1_3022(.VSS(VSS),.VDD(VDD),.Y(I11341),.A(g5809));
  NOT NOT1_3023(.VSS(VSS),.VDD(VDD),.Y(g6338),.A(I11341));
  NOT NOT1_3024(.VSS(VSS),.VDD(VDD),.Y(I11344),.A(g5820));
  NOT NOT1_3025(.VSS(VSS),.VDD(VDD),.Y(g6339),.A(I11344));
  NOT NOT1_3026(.VSS(VSS),.VDD(VDD),.Y(I11347),.A(g5761));
  NOT NOT1_3027(.VSS(VSS),.VDD(VDD),.Y(g6340),.A(I11347));
  NOT NOT1_3028(.VSS(VSS),.VDD(VDD),.Y(I11350),.A(g5763));
  NOT NOT1_3029(.VSS(VSS),.VDD(VDD),.Y(g6341),.A(I11350));
  NOT NOT1_3030(.VSS(VSS),.VDD(VDD),.Y(I11353),.A(g5788));
  NOT NOT1_3031(.VSS(VSS),.VDD(VDD),.Y(g6342),.A(I11353));
  NOT NOT1_3032(.VSS(VSS),.VDD(VDD),.Y(I11356),.A(g5799));
  NOT NOT1_3033(.VSS(VSS),.VDD(VDD),.Y(g6343),.A(I11356));
  NOT NOT1_3034(.VSS(VSS),.VDD(VDD),.Y(I11359),.A(g5810));
  NOT NOT1_3035(.VSS(VSS),.VDD(VDD),.Y(g6344),.A(I11359));
  NOT NOT1_3036(.VSS(VSS),.VDD(VDD),.Y(I11362),.A(g5821));
  NOT NOT1_3037(.VSS(VSS),.VDD(VDD),.Y(g6345),.A(I11362));
  NOT NOT1_3038(.VSS(VSS),.VDD(VDD),.Y(I11365),.A(g5826));
  NOT NOT1_3039(.VSS(VSS),.VDD(VDD),.Y(g6346),.A(I11365));
  NOT NOT1_3040(.VSS(VSS),.VDD(VDD),.Y(I11368),.A(g5833));
  NOT NOT1_3041(.VSS(VSS),.VDD(VDD),.Y(g6347),.A(I11368));
  NOT NOT1_3042(.VSS(VSS),.VDD(VDD),.Y(I11371),.A(g5840));
  NOT NOT1_3043(.VSS(VSS),.VDD(VDD),.Y(g6348),.A(I11371));
  NOT NOT1_3044(.VSS(VSS),.VDD(VDD),.Y(I11374),.A(g5844));
  NOT NOT1_3045(.VSS(VSS),.VDD(VDD),.Y(g6349),.A(I11374));
  NOT NOT1_3046(.VSS(VSS),.VDD(VDD),.Y(I11377),.A(g5811));
  NOT NOT1_3047(.VSS(VSS),.VDD(VDD),.Y(g6350),.A(I11377));
  NOT NOT1_3048(.VSS(VSS),.VDD(VDD),.Y(I11380),.A(g5822));
  NOT NOT1_3049(.VSS(VSS),.VDD(VDD),.Y(g6351),.A(I11380));
  NOT NOT1_3050(.VSS(VSS),.VDD(VDD),.Y(I11383),.A(g5827));
  NOT NOT1_3051(.VSS(VSS),.VDD(VDD),.Y(g6352),.A(I11383));
  NOT NOT1_3052(.VSS(VSS),.VDD(VDD),.Y(I11386),.A(g5764));
  NOT NOT1_3053(.VSS(VSS),.VDD(VDD),.Y(g6353),.A(I11386));
  NOT NOT1_3054(.VSS(VSS),.VDD(VDD),.Y(I11389),.A(g5766));
  NOT NOT1_3055(.VSS(VSS),.VDD(VDD),.Y(g6354),.A(I11389));
  NOT NOT1_3056(.VSS(VSS),.VDD(VDD),.Y(I11392),.A(g5800));
  NOT NOT1_3057(.VSS(VSS),.VDD(VDD),.Y(g6355),.A(I11392));
  NOT NOT1_3058(.VSS(VSS),.VDD(VDD),.Y(I11395),.A(g5812));
  NOT NOT1_3059(.VSS(VSS),.VDD(VDD),.Y(g6356),.A(I11395));
  NOT NOT1_3060(.VSS(VSS),.VDD(VDD),.Y(I11398),.A(g5823));
  NOT NOT1_3061(.VSS(VSS),.VDD(VDD),.Y(g6357),.A(I11398));
  NOT NOT1_3062(.VSS(VSS),.VDD(VDD),.Y(I11401),.A(g5828));
  NOT NOT1_3063(.VSS(VSS),.VDD(VDD),.Y(g6358),.A(I11401));
  NOT NOT1_3064(.VSS(VSS),.VDD(VDD),.Y(I11404),.A(g5834));
  NOT NOT1_3065(.VSS(VSS),.VDD(VDD),.Y(g6359),.A(I11404));
  NOT NOT1_3066(.VSS(VSS),.VDD(VDD),.Y(I11407),.A(g5841));
  NOT NOT1_3067(.VSS(VSS),.VDD(VDD),.Y(g6360),.A(I11407));
  NOT NOT1_3068(.VSS(VSS),.VDD(VDD),.Y(I11410),.A(g5845));
  NOT NOT1_3069(.VSS(VSS),.VDD(VDD),.Y(g6361),.A(I11410));
  NOT NOT1_3070(.VSS(VSS),.VDD(VDD),.Y(I11413),.A(g5871));
  NOT NOT1_3071(.VSS(VSS),.VDD(VDD),.Y(g6362),.A(I11413));
  NOT NOT1_3072(.VSS(VSS),.VDD(VDD),.Y(I11416),.A(g5829));
  NOT NOT1_3073(.VSS(VSS),.VDD(VDD),.Y(g6363),.A(I11416));
  NOT NOT1_3074(.VSS(VSS),.VDD(VDD),.Y(I11419),.A(g5835));
  NOT NOT1_3075(.VSS(VSS),.VDD(VDD),.Y(g6364),.A(I11419));
  NOT NOT1_3076(.VSS(VSS),.VDD(VDD),.Y(I11422),.A(g5842));
  NOT NOT1_3077(.VSS(VSS),.VDD(VDD),.Y(g6365),.A(I11422));
  NOT NOT1_3078(.VSS(VSS),.VDD(VDD),.Y(I11425),.A(g5872));
  NOT NOT1_3079(.VSS(VSS),.VDD(VDD),.Y(g6366),.A(I11425));
  NOT NOT1_3080(.VSS(VSS),.VDD(VDD),.Y(I11428),.A(g5813));
  NOT NOT1_3081(.VSS(VSS),.VDD(VDD),.Y(g6367),.A(I11428));
  NOT NOT1_3082(.VSS(VSS),.VDD(VDD),.Y(I11431),.A(g5782));
  NOT NOT1_3083(.VSS(VSS),.VDD(VDD),.Y(g6368),.A(I11431));
  NOT NOT1_3084(.VSS(VSS),.VDD(VDD),.Y(I11434),.A(g5789));
  NOT NOT1_3085(.VSS(VSS),.VDD(VDD),.Y(g6369),.A(I11434));
  NOT NOT1_3086(.VSS(VSS),.VDD(VDD),.Y(I11437),.A(g5801));
  NOT NOT1_3087(.VSS(VSS),.VDD(VDD),.Y(g6370),.A(I11437));
  NOT NOT1_3088(.VSS(VSS),.VDD(VDD),.Y(I11440),.A(g6009));
  NOT NOT1_3089(.VSS(VSS),.VDD(VDD),.Y(g6371),.A(I11440));
  NOT NOT1_3090(.VSS(VSS),.VDD(VDD),.Y(I11443),.A(g6038));
  NOT NOT1_3091(.VSS(VSS),.VDD(VDD),.Y(g6372),.A(I11443));
  NOT NOT1_3092(.VSS(VSS),.VDD(VDD),.Y(I11446),.A(g6062));
  NOT NOT1_3093(.VSS(VSS),.VDD(VDD),.Y(g6373),.A(I11446));
  NOT NOT1_3094(.VSS(VSS),.VDD(VDD),.Y(I11449),.A(g6068));
  NOT NOT1_3095(.VSS(VSS),.VDD(VDD),.Y(g6374),.A(I11449));
  NOT NOT1_3096(.VSS(VSS),.VDD(VDD),.Y(I11452),.A(g6071));
  NOT NOT1_3097(.VSS(VSS),.VDD(VDD),.Y(g6375),.A(I11452));
  NOT NOT1_3098(.VSS(VSS),.VDD(VDD),.Y(I11455),.A(g6087));
  NOT NOT1_3099(.VSS(VSS),.VDD(VDD),.Y(g6376),.A(I11455));
  NOT NOT1_3100(.VSS(VSS),.VDD(VDD),.Y(I11458),.A(g6063));
  NOT NOT1_3101(.VSS(VSS),.VDD(VDD),.Y(g6377),.A(I11458));
  NOT NOT1_3102(.VSS(VSS),.VDD(VDD),.Y(I11461),.A(g6094));
  NOT NOT1_3103(.VSS(VSS),.VDD(VDD),.Y(g6378),.A(I11461));
  NOT NOT1_3104(.VSS(VSS),.VDD(VDD),.Y(I11464),.A(g6088));
  NOT NOT1_3105(.VSS(VSS),.VDD(VDD),.Y(g6379),.A(I11464));
  NOT NOT1_3106(.VSS(VSS),.VDD(VDD),.Y(I11467),.A(g6064));
  NOT NOT1_3107(.VSS(VSS),.VDD(VDD),.Y(g6380),.A(I11467));
  NOT NOT1_3108(.VSS(VSS),.VDD(VDD),.Y(I11470),.A(g6095));
  NOT NOT1_3109(.VSS(VSS),.VDD(VDD),.Y(g6381),.A(I11470));
  NOT NOT1_3110(.VSS(VSS),.VDD(VDD),.Y(I11473),.A(g6069));
  NOT NOT1_3111(.VSS(VSS),.VDD(VDD),.Y(g6382),.A(I11473));
  NOT NOT1_3112(.VSS(VSS),.VDD(VDD),.Y(I11476),.A(g6194));
  NOT NOT1_3113(.VSS(VSS),.VDD(VDD),.Y(g6383),.A(I11476));
  NOT NOT1_3114(.VSS(VSS),.VDD(VDD),.Y(I11479),.A(g6201));
  NOT NOT1_3115(.VSS(VSS),.VDD(VDD),.Y(g6384),.A(I11479));
  NOT NOT1_3116(.VSS(VSS),.VDD(VDD),.Y(I11482),.A(g6117));
  NOT NOT1_3117(.VSS(VSS),.VDD(VDD),.Y(g6385),.A(I11482));
  NOT NOT1_3118(.VSS(VSS),.VDD(VDD),.Y(I11485),.A(g6137));
  NOT NOT1_3119(.VSS(VSS),.VDD(VDD),.Y(g6386),.A(I11485));
  NOT NOT1_3120(.VSS(VSS),.VDD(VDD),.Y(I11488),.A(g6034));
  NOT NOT1_3121(.VSS(VSS),.VDD(VDD),.Y(g6387),.A(I11488));
  NOT NOT1_3122(.VSS(VSS),.VDD(VDD),.Y(I11491),.A(g6010));
  NOT NOT1_3123(.VSS(VSS),.VDD(VDD),.Y(g6388),.A(I11491));
  NOT NOT1_3124(.VSS(VSS),.VDD(VDD),.Y(I11494),.A(g6037));
  NOT NOT1_3125(.VSS(VSS),.VDD(VDD),.Y(g6389),.A(I11494));
  NOT NOT1_3126(.VSS(VSS),.VDD(VDD),.Y(I11497),.A(g6014));
  NOT NOT1_3127(.VSS(VSS),.VDD(VDD),.Y(g6390),.A(I11497));
  NOT NOT1_3128(.VSS(VSS),.VDD(VDD),.Y(I11500),.A(g6219));
  NOT NOT1_3129(.VSS(VSS),.VDD(VDD),.Y(g6391),.A(I11500));
  NOT NOT1_3130(.VSS(VSS),.VDD(VDD),.Y(I11503),.A(g6220));
  NOT NOT1_3131(.VSS(VSS),.VDD(VDD),.Y(g6392),.A(I11503));
  NOT NOT1_3132(.VSS(VSS),.VDD(VDD),.Y(I11506),.A(g6189));
  NOT NOT1_3133(.VSS(VSS),.VDD(VDD),.Y(g6393),.A(I11506));
  NOT NOT1_3134(.VSS(VSS),.VDD(VDD),.Y(I11512),.A(g5874));
  NOT NOT1_3135(.VSS(VSS),.VDD(VDD),.Y(g6397),.A(I11512));
  NOT NOT1_3136(.VSS(VSS),.VDD(VDD),.Y(I11515),.A(g5897));
  NOT NOT1_3137(.VSS(VSS),.VDD(VDD),.Y(g6398),.A(I11515));
  NOT NOT1_3138(.VSS(VSS),.VDD(VDD),.Y(I11522),.A(g5847));
  NOT NOT1_3139(.VSS(VSS),.VDD(VDD),.Y(g6403),.A(I11522));
  NOT NOT1_3140(.VSS(VSS),.VDD(VDD),.Y(I11525),.A(g5874));
  NOT NOT1_3141(.VSS(VSS),.VDD(VDD),.Y(g6404),.A(I11525));
  NOT NOT1_3142(.VSS(VSS),.VDD(VDD),.Y(I11533),.A(g5847));
  NOT NOT1_3143(.VSS(VSS),.VDD(VDD),.Y(g6410),.A(I11533));
  NOT NOT1_3144(.VSS(VSS),.VDD(VDD),.Y(I11556),.A(g6065));
  NOT NOT1_3145(.VSS(VSS),.VDD(VDD),.Y(g6425),.A(I11556));
  NOT NOT1_3146(.VSS(VSS),.VDD(VDD),.Y(I11559),.A(g6065));
  NOT NOT1_3147(.VSS(VSS),.VDD(VDD),.Y(g6426),.A(I11559));
  NOT NOT1_3148(.VSS(VSS),.VDD(VDD),.Y(I11562),.A(g5939));
  NOT NOT1_3149(.VSS(VSS),.VDD(VDD),.Y(g6427),.A(I11562));
  NOT NOT1_3150(.VSS(VSS),.VDD(VDD),.Y(I11569),.A(g6279));
  NOT NOT1_3151(.VSS(VSS),.VDD(VDD),.Y(g6432),.A(I11569));
  NOT NOT1_3152(.VSS(VSS),.VDD(VDD),.Y(I11586),.A(g6256));
  NOT NOT1_3153(.VSS(VSS),.VDD(VDD),.Y(g6441),.A(I11586));
  NOT NOT1_3154(.VSS(VSS),.VDD(VDD),.Y(I11591),.A(g5814));
  NOT NOT1_3155(.VSS(VSS),.VDD(VDD),.Y(g6446),.A(I11591));
  NOT NOT1_3156(.VSS(VSS),.VDD(VDD),.Y(I11596),.A(g6228));
  NOT NOT1_3157(.VSS(VSS),.VDD(VDD),.Y(g6449),.A(I11596));
  NOT NOT1_3158(.VSS(VSS),.VDD(VDD),.Y(I11607),.A(g5767));
  NOT NOT1_3159(.VSS(VSS),.VDD(VDD),.Y(g6461),.A(I11607));
  NOT NOT1_3160(.VSS(VSS),.VDD(VDD),.Y(I11622),.A(g5847));
  NOT NOT1_3161(.VSS(VSS),.VDD(VDD),.Y(g6468),.A(I11622));
  NOT NOT1_3162(.VSS(VSS),.VDD(VDD),.Y(I11627),.A(g5874));
  NOT NOT1_3163(.VSS(VSS),.VDD(VDD),.Y(g6471),.A(I11627));
  NOT NOT1_3164(.VSS(VSS),.VDD(VDD),.Y(I11633),.A(g5897));
  NOT NOT1_3165(.VSS(VSS),.VDD(VDD),.Y(g6475),.A(I11633));
  NOT NOT1_3166(.VSS(VSS),.VDD(VDD),.Y(I11638),.A(g5847));
  NOT NOT1_3167(.VSS(VSS),.VDD(VDD),.Y(g6478),.A(I11638));
  NOT NOT1_3168(.VSS(VSS),.VDD(VDD),.Y(I11641),.A(g5918));
  NOT NOT1_3169(.VSS(VSS),.VDD(VDD),.Y(g6481),.A(I11641));
  NOT NOT1_3170(.VSS(VSS),.VDD(VDD),.Y(I11645),.A(g5874));
  NOT NOT1_3171(.VSS(VSS),.VDD(VDD),.Y(g6483),.A(I11645));
  NOT NOT1_3172(.VSS(VSS),.VDD(VDD),.Y(I11648),.A(g6028));
  NOT NOT1_3173(.VSS(VSS),.VDD(VDD),.Y(g6486),.A(I11648));
  NOT NOT1_3174(.VSS(VSS),.VDD(VDD),.Y(I11652),.A(g5939));
  NOT NOT1_3175(.VSS(VSS),.VDD(VDD),.Y(g6488),.A(I11652));
  NOT NOT1_3176(.VSS(VSS),.VDD(VDD),.Y(I11656),.A(g5772));
  NOT NOT1_3177(.VSS(VSS),.VDD(VDD),.Y(g6490),.A(I11656));
  NOT NOT1_3178(.VSS(VSS),.VDD(VDD),.Y(I11659),.A(g5897));
  NOT NOT1_3179(.VSS(VSS),.VDD(VDD),.Y(g6493),.A(I11659));
  NOT NOT1_3180(.VSS(VSS),.VDD(VDD),.Y(I11662),.A(g5956));
  NOT NOT1_3181(.VSS(VSS),.VDD(VDD),.Y(g6496),.A(I11662));
  NOT NOT1_3182(.VSS(VSS),.VDD(VDD),.Y(I11666),.A(g5772));
  NOT NOT1_3183(.VSS(VSS),.VDD(VDD),.Y(g6498),.A(I11666));
  NOT NOT1_3184(.VSS(VSS),.VDD(VDD),.Y(I11669),.A(g5918));
  NOT NOT1_3185(.VSS(VSS),.VDD(VDD),.Y(g6501),.A(I11669));
  NOT NOT1_3186(.VSS(VSS),.VDD(VDD),.Y(I11672),.A(g5971));
  NOT NOT1_3187(.VSS(VSS),.VDD(VDD),.Y(g6502),.A(I11672));
  NOT NOT1_3188(.VSS(VSS),.VDD(VDD),.Y(I11677),.A(g6076));
  NOT NOT1_3189(.VSS(VSS),.VDD(VDD),.Y(g6505),.A(I11677));
  NOT NOT1_3190(.VSS(VSS),.VDD(VDD),.Y(I11680),.A(g5939));
  NOT NOT1_3191(.VSS(VSS),.VDD(VDD),.Y(g6506),.A(I11680));
  NOT NOT1_3192(.VSS(VSS),.VDD(VDD),.Y(I11683),.A(g5988));
  NOT NOT1_3193(.VSS(VSS),.VDD(VDD),.Y(g6507),.A(I11683));
  NOT NOT1_3194(.VSS(VSS),.VDD(VDD),.Y(I11686),.A(g6076));
  NOT NOT1_3195(.VSS(VSS),.VDD(VDD),.Y(g6508),.A(I11686));
  NOT NOT1_3196(.VSS(VSS),.VDD(VDD),.Y(I11689),.A(g5956));
  NOT NOT1_3197(.VSS(VSS),.VDD(VDD),.Y(g6509),.A(I11689));
  NOT NOT1_3198(.VSS(VSS),.VDD(VDD),.Y(I11693),.A(g6076));
  NOT NOT1_3199(.VSS(VSS),.VDD(VDD),.Y(g6511),.A(I11693));
  NOT NOT1_3200(.VSS(VSS),.VDD(VDD),.Y(I11696),.A(g5971));
  NOT NOT1_3201(.VSS(VSS),.VDD(VDD),.Y(g6514),.A(I11696));
  NOT NOT1_3202(.VSS(VSS),.VDD(VDD),.Y(g6515),.A(g6125));
  NOT NOT1_3203(.VSS(VSS),.VDD(VDD),.Y(I11701),.A(g5772));
  NOT NOT1_3204(.VSS(VSS),.VDD(VDD),.Y(g6517),.A(I11701));
  NOT NOT1_3205(.VSS(VSS),.VDD(VDD),.Y(I11704),.A(g6076));
  NOT NOT1_3206(.VSS(VSS),.VDD(VDD),.Y(g6520),.A(I11704));
  NOT NOT1_3207(.VSS(VSS),.VDD(VDD),.Y(I11707),.A(g5988));
  NOT NOT1_3208(.VSS(VSS),.VDD(VDD),.Y(g6523),.A(I11707));
  NOT NOT1_3209(.VSS(VSS),.VDD(VDD),.Y(I11710),.A(g6098));
  NOT NOT1_3210(.VSS(VSS),.VDD(VDD),.Y(g6524),.A(I11710));
  NOT NOT1_3211(.VSS(VSS),.VDD(VDD),.Y(I11714),.A(g5772));
  NOT NOT1_3212(.VSS(VSS),.VDD(VDD),.Y(g6538),.A(I11714));
  NOT NOT1_3213(.VSS(VSS),.VDD(VDD),.Y(I11718),.A(g6115));
  NOT NOT1_3214(.VSS(VSS),.VDD(VDD),.Y(g6542),.A(I11718));
  NOT NOT1_3215(.VSS(VSS),.VDD(VDD),.Y(I11722),.A(g5772));
  NOT NOT1_3216(.VSS(VSS),.VDD(VDD),.Y(g6552),.A(I11722));
  NOT NOT1_3217(.VSS(VSS),.VDD(VDD),.Y(I11725),.A(g6036));
  NOT NOT1_3218(.VSS(VSS),.VDD(VDD),.Y(g6553),.A(I11725));
  NOT NOT1_3219(.VSS(VSS),.VDD(VDD),.Y(I11729),.A(g5772));
  NOT NOT1_3220(.VSS(VSS),.VDD(VDD),.Y(g6555),.A(I11729));
  NOT NOT1_3221(.VSS(VSS),.VDD(VDD),.Y(I11732),.A(g6076));
  NOT NOT1_3222(.VSS(VSS),.VDD(VDD),.Y(g6556),.A(I11732));
  NOT NOT1_3223(.VSS(VSS),.VDD(VDD),.Y(I11736),.A(g6076));
  NOT NOT1_3224(.VSS(VSS),.VDD(VDD),.Y(g6562),.A(I11736));
  NOT NOT1_3225(.VSS(VSS),.VDD(VDD),.Y(I11740),.A(g6136));
  NOT NOT1_3226(.VSS(VSS),.VDD(VDD),.Y(g6566),.A(I11740));
  NOT NOT1_3227(.VSS(VSS),.VDD(VDD),.Y(I11744),.A(g6120));
  NOT NOT1_3228(.VSS(VSS),.VDD(VDD),.Y(g6568),.A(I11744));
  NOT NOT1_3229(.VSS(VSS),.VDD(VDD),.Y(I11747),.A(g6123));
  NOT NOT1_3230(.VSS(VSS),.VDD(VDD),.Y(g6569),.A(I11747));
  NOT NOT1_3231(.VSS(VSS),.VDD(VDD),.Y(I11764),.A(g6056));
  NOT NOT1_3232(.VSS(VSS),.VDD(VDD),.Y(g6572),.A(I11764));
  NOT NOT1_3233(.VSS(VSS),.VDD(VDD),.Y(g6573),.A(g5868));
  NOT NOT1_3234(.VSS(VSS),.VDD(VDD),.Y(I11773),.A(g6262));
  NOT NOT1_3235(.VSS(VSS),.VDD(VDD),.Y(g6581),.A(I11773));
  NOT NOT1_3236(.VSS(VSS),.VDD(VDD),.Y(I11778),.A(g6180));
  NOT NOT1_3237(.VSS(VSS),.VDD(VDD),.Y(g6586),.A(I11778));
  NOT NOT1_3238(.VSS(VSS),.VDD(VDD),.Y(I11781),.A(g6284));
  NOT NOT1_3239(.VSS(VSS),.VDD(VDD),.Y(g6587),.A(I11781));
  NOT NOT1_3240(.VSS(VSS),.VDD(VDD),.Y(g6588),.A(g5836));
  NOT NOT1_3241(.VSS(VSS),.VDD(VDD),.Y(g6589),.A(g6083));
  NOT NOT1_3242(.VSS(VSS),.VDD(VDD),.Y(I11787),.A(g6273));
  NOT NOT1_3243(.VSS(VSS),.VDD(VDD),.Y(g6591),.A(I11787));
  NOT NOT1_3244(.VSS(VSS),.VDD(VDD),.Y(I11790),.A(g6282));
  NOT NOT1_3245(.VSS(VSS),.VDD(VDD),.Y(g6592),.A(I11790));
  NOT NOT1_3246(.VSS(VSS),.VDD(VDD),.Y(I11793),.A(g6188));
  NOT NOT1_3247(.VSS(VSS),.VDD(VDD),.Y(g6593),.A(I11793));
  NOT NOT1_3248(.VSS(VSS),.VDD(VDD),.Y(I11796),.A(g6287));
  NOT NOT1_3249(.VSS(VSS),.VDD(VDD),.Y(g6594),.A(I11796));
  NOT NOT1_3250(.VSS(VSS),.VDD(VDD),.Y(g6595),.A(g6083));
  NOT NOT1_3251(.VSS(VSS),.VDD(VDD),.Y(I11800),.A(g6164));
  NOT NOT1_3252(.VSS(VSS),.VDD(VDD),.Y(g6596),.A(I11800));
  NOT NOT1_3253(.VSS(VSS),.VDD(VDD),.Y(I11803),.A(g6280));
  NOT NOT1_3254(.VSS(VSS),.VDD(VDD),.Y(g6597),.A(I11803));
  NOT NOT1_3255(.VSS(VSS),.VDD(VDD),.Y(I11806),.A(g6275));
  NOT NOT1_3256(.VSS(VSS),.VDD(VDD),.Y(g6598),.A(I11806));
  NOT NOT1_3257(.VSS(VSS),.VDD(VDD),.Y(I11809),.A(g6285));
  NOT NOT1_3258(.VSS(VSS),.VDD(VDD),.Y(g6599),.A(I11809));
  NOT NOT1_3259(.VSS(VSS),.VDD(VDD),.Y(g6601),.A(g6083));
  NOT NOT1_3260(.VSS(VSS),.VDD(VDD),.Y(I11815),.A(g6169));
  NOT NOT1_3261(.VSS(VSS),.VDD(VDD),.Y(g6603),.A(I11815));
  NOT NOT1_3262(.VSS(VSS),.VDD(VDD),.Y(I11818),.A(g6276));
  NOT NOT1_3263(.VSS(VSS),.VDD(VDD),.Y(g6604),.A(I11818));
  NOT NOT1_3264(.VSS(VSS),.VDD(VDD),.Y(I11821),.A(g6170));
  NOT NOT1_3265(.VSS(VSS),.VDD(VDD),.Y(g6605),.A(I11821));
  NOT NOT1_3266(.VSS(VSS),.VDD(VDD),.Y(I11824),.A(g6283));
  NOT NOT1_3267(.VSS(VSS),.VDD(VDD),.Y(g6606),.A(I11824));
  NOT NOT1_3268(.VSS(VSS),.VDD(VDD),.Y(I11827),.A(g6231));
  NOT NOT1_3269(.VSS(VSS),.VDD(VDD),.Y(g6607),.A(I11827));
  NOT NOT1_3270(.VSS(VSS),.VDD(VDD),.Y(I11832),.A(g6274));
  NOT NOT1_3271(.VSS(VSS),.VDD(VDD),.Y(g6612),.A(I11832));
  NOT NOT1_3272(.VSS(VSS),.VDD(VDD),.Y(I11835),.A(g6181));
  NOT NOT1_3273(.VSS(VSS),.VDD(VDD),.Y(g6613),.A(I11835));
  NOT NOT1_3274(.VSS(VSS),.VDD(VDD),.Y(I11838),.A(g6281));
  NOT NOT1_3275(.VSS(VSS),.VDD(VDD),.Y(g6614),.A(I11838));
  NOT NOT1_3276(.VSS(VSS),.VDD(VDD),.Y(I11848),.A(g6159));
  NOT NOT1_3277(.VSS(VSS),.VDD(VDD),.Y(g6616),.A(I11848));
  NOT NOT1_3278(.VSS(VSS),.VDD(VDD),.Y(I11851),.A(g6277));
  NOT NOT1_3279(.VSS(VSS),.VDD(VDD),.Y(g6617),.A(I11851));
  NOT NOT1_3280(.VSS(VSS),.VDD(VDD),.Y(g6618),.A(g6003));
  NOT NOT1_3281(.VSS(VSS),.VDD(VDD),.Y(I11855),.A(g5751));
  NOT NOT1_3282(.VSS(VSS),.VDD(VDD),.Y(g6621),.A(I11855));
  NOT NOT1_3283(.VSS(VSS),.VDD(VDD),.Y(I11858),.A(g6165));
  NOT NOT1_3284(.VSS(VSS),.VDD(VDD),.Y(g6622),.A(I11858));
  NOT NOT1_3285(.VSS(VSS),.VDD(VDD),.Y(I11861),.A(g5747));
  NOT NOT1_3286(.VSS(VSS),.VDD(VDD),.Y(g6623),.A(I11861));
  NOT NOT1_3287(.VSS(VSS),.VDD(VDD),.Y(I11864),.A(g5753));
  NOT NOT1_3288(.VSS(VSS),.VDD(VDD),.Y(g6624),.A(I11864));
  NOT NOT1_3289(.VSS(VSS),.VDD(VDD),.Y(I11867),.A(g6286));
  NOT NOT1_3290(.VSS(VSS),.VDD(VDD),.Y(g6625),.A(I11867));
  NOT NOT1_3291(.VSS(VSS),.VDD(VDD),.Y(I11870),.A(g5752));
  NOT NOT1_3292(.VSS(VSS),.VDD(VDD),.Y(g6626),.A(I11870));
  NOT NOT1_3293(.VSS(VSS),.VDD(VDD),.Y(I11880),.A(g5748));
  NOT NOT1_3294(.VSS(VSS),.VDD(VDD),.Y(g6628),.A(I11880));
  NOT NOT1_3295(.VSS(VSS),.VDD(VDD),.Y(I11884),.A(g6091));
  NOT NOT1_3296(.VSS(VSS),.VDD(VDD),.Y(g6630),.A(I11884));
  NOT NOT1_3297(.VSS(VSS),.VDD(VDD),.Y(I11887),.A(g5918));
  NOT NOT1_3298(.VSS(VSS),.VDD(VDD),.Y(g6631),.A(I11887));
  NOT NOT1_3299(.VSS(VSS),.VDD(VDD),.Y(I11890),.A(g6135));
  NOT NOT1_3300(.VSS(VSS),.VDD(VDD),.Y(g6632),.A(I11890));
  NOT NOT1_3301(.VSS(VSS),.VDD(VDD),.Y(I11894),.A(g5956));
  NOT NOT1_3302(.VSS(VSS),.VDD(VDD),.Y(g6634),.A(I11894));
  NOT NOT1_3303(.VSS(VSS),.VDD(VDD),.Y(I11897),.A(g6141));
  NOT NOT1_3304(.VSS(VSS),.VDD(VDD),.Y(g6635),.A(I11897));
  NOT NOT1_3305(.VSS(VSS),.VDD(VDD),.Y(I11900),.A(g5847));
  NOT NOT1_3306(.VSS(VSS),.VDD(VDD),.Y(g6636),.A(I11900));
  NOT NOT1_3307(.VSS(VSS),.VDD(VDD),.Y(I11903),.A(g5939));
  NOT NOT1_3308(.VSS(VSS),.VDD(VDD),.Y(g6637),.A(I11903));
  NOT NOT1_3309(.VSS(VSS),.VDD(VDD),.Y(g6639),.A(g6198));
  NOT NOT1_3310(.VSS(VSS),.VDD(VDD),.Y(I11908),.A(g5918));
  NOT NOT1_3311(.VSS(VSS),.VDD(VDD),.Y(g6640),.A(I11908));
  NOT NOT1_3312(.VSS(VSS),.VDD(VDD),.Y(I11912),.A(g5897));
  NOT NOT1_3313(.VSS(VSS),.VDD(VDD),.Y(g6642),.A(I11912));
  NOT NOT1_3314(.VSS(VSS),.VDD(VDD),.Y(g6644),.A(g6208));
  NOT NOT1_3315(.VSS(VSS),.VDD(VDD),.Y(I11917),.A(g5897));
  NOT NOT1_3316(.VSS(VSS),.VDD(VDD),.Y(g6645),.A(I11917));
  NOT NOT1_3317(.VSS(VSS),.VDD(VDD),.Y(I11920),.A(g5874));
  NOT NOT1_3318(.VSS(VSS),.VDD(VDD),.Y(g6646),.A(I11920));
  NOT NOT1_3319(.VSS(VSS),.VDD(VDD),.Y(I11923),.A(g5939));
  NOT NOT1_3320(.VSS(VSS),.VDD(VDD),.Y(g6647),.A(I11923));
  NOT NOT1_3321(.VSS(VSS),.VDD(VDD),.Y(I11926),.A(g6190));
  NOT NOT1_3322(.VSS(VSS),.VDD(VDD),.Y(g6648),.A(I11926));
  NOT NOT1_3323(.VSS(VSS),.VDD(VDD),.Y(I11929),.A(g6190));
  NOT NOT1_3324(.VSS(VSS),.VDD(VDD),.Y(g6649),.A(I11929));
  NOT NOT1_3325(.VSS(VSS),.VDD(VDD),.Y(g6650),.A(g6213));
  NOT NOT1_3326(.VSS(VSS),.VDD(VDD),.Y(I11933),.A(g5847));
  NOT NOT1_3327(.VSS(VSS),.VDD(VDD),.Y(g6651),.A(I11933));
  NOT NOT1_3328(.VSS(VSS),.VDD(VDD),.Y(I11936),.A(g5918));
  NOT NOT1_3329(.VSS(VSS),.VDD(VDD),.Y(g6652),.A(I11936));
  NOT NOT1_3330(.VSS(VSS),.VDD(VDD),.Y(I11939),.A(g6015));
  NOT NOT1_3331(.VSS(VSS),.VDD(VDD),.Y(g6653),.A(I11939));
  NOT NOT1_3332(.VSS(VSS),.VDD(VDD),.Y(I11942),.A(g6015));
  NOT NOT1_3333(.VSS(VSS),.VDD(VDD),.Y(g6654),.A(I11942));
  NOT NOT1_3334(.VSS(VSS),.VDD(VDD),.Y(I11945),.A(g5874));
  NOT NOT1_3335(.VSS(VSS),.VDD(VDD),.Y(g6655),.A(I11945));
  NOT NOT1_3336(.VSS(VSS),.VDD(VDD),.Y(I11948),.A(g5897));
  NOT NOT1_3337(.VSS(VSS),.VDD(VDD),.Y(g6656),.A(I11948));
  NOT NOT1_3338(.VSS(VSS),.VDD(VDD),.Y(I11951),.A(g5847));
  NOT NOT1_3339(.VSS(VSS),.VDD(VDD),.Y(g6657),.A(I11951));
  NOT NOT1_3340(.VSS(VSS),.VDD(VDD),.Y(g6658),.A(g6224));
  NOT NOT1_3341(.VSS(VSS),.VDD(VDD),.Y(I11955),.A(g5988));
  NOT NOT1_3342(.VSS(VSS),.VDD(VDD),.Y(g6659),.A(I11955));
  NOT NOT1_3343(.VSS(VSS),.VDD(VDD),.Y(I11958),.A(g5874));
  NOT NOT1_3344(.VSS(VSS),.VDD(VDD),.Y(g6660),.A(I11958));
  NOT NOT1_3345(.VSS(VSS),.VDD(VDD),.Y(I11961),.A(g5988));
  NOT NOT1_3346(.VSS(VSS),.VDD(VDD),.Y(g6661),.A(I11961));
  NOT NOT1_3347(.VSS(VSS),.VDD(VDD),.Y(I11964),.A(g5971));
  NOT NOT1_3348(.VSS(VSS),.VDD(VDD),.Y(g6662),.A(I11964));
  NOT NOT1_3349(.VSS(VSS),.VDD(VDD),.Y(I11967),.A(g5971));
  NOT NOT1_3350(.VSS(VSS),.VDD(VDD),.Y(g6663),.A(I11967));
  NOT NOT1_3351(.VSS(VSS),.VDD(VDD),.Y(I11971),.A(g6179));
  NOT NOT1_3352(.VSS(VSS),.VDD(VDD),.Y(g6671),.A(I11971));
  NOT NOT1_3353(.VSS(VSS),.VDD(VDD),.Y(I11974),.A(g5956));
  NOT NOT1_3354(.VSS(VSS),.VDD(VDD),.Y(g6672),.A(I11974));
  NOT NOT1_3355(.VSS(VSS),.VDD(VDD),.Y(I11978),.A(g6186));
  NOT NOT1_3356(.VSS(VSS),.VDD(VDD),.Y(g6674),.A(I11978));
  NOT NOT1_3357(.VSS(VSS),.VDD(VDD),.Y(I11981),.A(g6246));
  NOT NOT1_3358(.VSS(VSS),.VDD(VDD),.Y(g6675),.A(I11981));
  NOT NOT1_3359(.VSS(VSS),.VDD(VDD),.Y(I11984),.A(g6246));
  NOT NOT1_3360(.VSS(VSS),.VDD(VDD),.Y(g6676),.A(I11984));
  NOT NOT1_3361(.VSS(VSS),.VDD(VDD),.Y(I11987),.A(g6278));
  NOT NOT1_3362(.VSS(VSS),.VDD(VDD),.Y(g6677),.A(I11987));
  NOT NOT1_3363(.VSS(VSS),.VDD(VDD),.Y(I11991),.A(g5939));
  NOT NOT1_3364(.VSS(VSS),.VDD(VDD),.Y(g6681),.A(I11991));
  NOT NOT1_3365(.VSS(VSS),.VDD(VDD),.Y(I11994),.A(g6195));
  NOT NOT1_3366(.VSS(VSS),.VDD(VDD),.Y(g6682),.A(I11994));
  NOT NOT1_3367(.VSS(VSS),.VDD(VDD),.Y(g6683),.A(g6237));
  NOT NOT1_3368(.VSS(VSS),.VDD(VDD),.Y(I11998),.A(g5918));
  NOT NOT1_3369(.VSS(VSS),.VDD(VDD),.Y(g6684),.A(I11998));
  NOT NOT1_3370(.VSS(VSS),.VDD(VDD),.Y(I12003),.A(g6202));
  NOT NOT1_3371(.VSS(VSS),.VDD(VDD),.Y(g6687),.A(I12003));
  NOT NOT1_3372(.VSS(VSS),.VDD(VDD),.Y(I12008),.A(g5897));
  NOT NOT1_3373(.VSS(VSS),.VDD(VDD),.Y(g6692),.A(I12008));
  NOT NOT1_3374(.VSS(VSS),.VDD(VDD),.Y(I12011),.A(g5939));
  NOT NOT1_3375(.VSS(VSS),.VDD(VDD),.Y(g6693),.A(I12011));
  NOT NOT1_3376(.VSS(VSS),.VDD(VDD),.Y(I12022),.A(g5874));
  NOT NOT1_3377(.VSS(VSS),.VDD(VDD),.Y(g6696),.A(I12022));
  NOT NOT1_3378(.VSS(VSS),.VDD(VDD),.Y(I12025),.A(g5918));
  NOT NOT1_3379(.VSS(VSS),.VDD(VDD),.Y(g6697),.A(I12025));
  NOT NOT1_3380(.VSS(VSS),.VDD(VDD),.Y(g6700),.A(g6244));
  NOT NOT1_3381(.VSS(VSS),.VDD(VDD),.Y(I12038),.A(g5847));
  NOT NOT1_3382(.VSS(VSS),.VDD(VDD),.Y(g6702),.A(I12038));
  NOT NOT1_3383(.VSS(VSS),.VDD(VDD),.Y(I12041),.A(g5897));
  NOT NOT1_3384(.VSS(VSS),.VDD(VDD),.Y(g6703),.A(I12041));
  NOT NOT1_3385(.VSS(VSS),.VDD(VDD),.Y(I12044),.A(g5847));
  NOT NOT1_3386(.VSS(VSS),.VDD(VDD),.Y(g6704),.A(I12044));
  NOT NOT1_3387(.VSS(VSS),.VDD(VDD),.Y(g6708),.A(g6250));
  NOT NOT1_3388(.VSS(VSS),.VDD(VDD),.Y(I12059),.A(g5874));
  NOT NOT1_3389(.VSS(VSS),.VDD(VDD),.Y(g6711),.A(I12059));
  NOT NOT1_3390(.VSS(VSS),.VDD(VDD),.Y(I12062),.A(g5988));
  NOT NOT1_3391(.VSS(VSS),.VDD(VDD),.Y(g6712),.A(I12062));
  NOT NOT1_3392(.VSS(VSS),.VDD(VDD),.Y(I12065),.A(g5897));
  NOT NOT1_3393(.VSS(VSS),.VDD(VDD),.Y(g6713),.A(I12065));
  NOT NOT1_3394(.VSS(VSS),.VDD(VDD),.Y(I12068),.A(g5847));
  NOT NOT1_3395(.VSS(VSS),.VDD(VDD),.Y(g6714),.A(I12068));
  NOT NOT1_3396(.VSS(VSS),.VDD(VDD),.Y(g6720),.A(g6254));
  NOT NOT1_3397(.VSS(VSS),.VDD(VDD),.Y(g6721),.A(g6257));
  NOT NOT1_3398(.VSS(VSS),.VDD(VDD),.Y(I12085),.A(g5971));
  NOT NOT1_3399(.VSS(VSS),.VDD(VDD),.Y(g6723),.A(I12085));
  NOT NOT1_3400(.VSS(VSS),.VDD(VDD),.Y(I12088),.A(g5874));
  NOT NOT1_3401(.VSS(VSS),.VDD(VDD),.Y(g6724),.A(I12088));
  NOT NOT1_3402(.VSS(VSS),.VDD(VDD),.Y(I12091),.A(g5988));
  NOT NOT1_3403(.VSS(VSS),.VDD(VDD),.Y(g6725),.A(I12091));
  NOT NOT1_3404(.VSS(VSS),.VDD(VDD),.Y(g6729),.A(g6263));
  NOT NOT1_3405(.VSS(VSS),.VDD(VDD),.Y(I12098),.A(g5956));
  NOT NOT1_3406(.VSS(VSS),.VDD(VDD),.Y(g6730),.A(I12098));
  NOT NOT1_3407(.VSS(VSS),.VDD(VDD),.Y(I12101),.A(g5971));
  NOT NOT1_3408(.VSS(VSS),.VDD(VDD),.Y(g6731),.A(I12101));
  NOT NOT1_3409(.VSS(VSS),.VDD(VDD),.Y(I12108),.A(g5939));
  NOT NOT1_3410(.VSS(VSS),.VDD(VDD),.Y(g6736),.A(I12108));
  NOT NOT1_3411(.VSS(VSS),.VDD(VDD),.Y(I12111),.A(g5956));
  NOT NOT1_3412(.VSS(VSS),.VDD(VDD),.Y(g6737),.A(I12111));
  NOT NOT1_3413(.VSS(VSS),.VDD(VDD),.Y(I12117),.A(g5918));
  NOT NOT1_3414(.VSS(VSS),.VDD(VDD),.Y(g6741),.A(I12117));
  NOT NOT1_3415(.VSS(VSS),.VDD(VDD),.Y(I12120),.A(g5939));
  NOT NOT1_3416(.VSS(VSS),.VDD(VDD),.Y(g6742),.A(I12120));
  NOT NOT1_3417(.VSS(VSS),.VDD(VDD),.Y(I12124),.A(g5847));
  NOT NOT1_3418(.VSS(VSS),.VDD(VDD),.Y(g6744),.A(I12124));
  NOT NOT1_3419(.VSS(VSS),.VDD(VDD),.Y(I12128),.A(g5897));
  NOT NOT1_3420(.VSS(VSS),.VDD(VDD),.Y(g6751),.A(I12128));
  NOT NOT1_3421(.VSS(VSS),.VDD(VDD),.Y(I12131),.A(g5918));
  NOT NOT1_3422(.VSS(VSS),.VDD(VDD),.Y(g6752),.A(I12131));
  NOT NOT1_3423(.VSS(VSS),.VDD(VDD),.Y(I12135),.A(g5988));
  NOT NOT1_3424(.VSS(VSS),.VDD(VDD),.Y(g6754),.A(I12135));
  NOT NOT1_3425(.VSS(VSS),.VDD(VDD),.Y(I12138),.A(g5874));
  NOT NOT1_3426(.VSS(VSS),.VDD(VDD),.Y(g6755),.A(I12138));
  NOT NOT1_3427(.VSS(VSS),.VDD(VDD),.Y(I12141),.A(g5897));
  NOT NOT1_3428(.VSS(VSS),.VDD(VDD),.Y(g6756),.A(I12141));
  NOT NOT1_3429(.VSS(VSS),.VDD(VDD),.Y(I12145),.A(g5971));
  NOT NOT1_3430(.VSS(VSS),.VDD(VDD),.Y(g6758),.A(I12145));
  NOT NOT1_3431(.VSS(VSS),.VDD(VDD),.Y(I12148),.A(g5988));
  NOT NOT1_3432(.VSS(VSS),.VDD(VDD),.Y(g6759),.A(I12148));
  NOT NOT1_3433(.VSS(VSS),.VDD(VDD),.Y(I12151),.A(g5847));
  NOT NOT1_3434(.VSS(VSS),.VDD(VDD),.Y(g6760),.A(I12151));
  NOT NOT1_3435(.VSS(VSS),.VDD(VDD),.Y(I12154),.A(g5874));
  NOT NOT1_3436(.VSS(VSS),.VDD(VDD),.Y(g6761),.A(I12154));
  NOT NOT1_3437(.VSS(VSS),.VDD(VDD),.Y(I12158),.A(g5956));
  NOT NOT1_3438(.VSS(VSS),.VDD(VDD),.Y(g6763),.A(I12158));
  NOT NOT1_3439(.VSS(VSS),.VDD(VDD),.Y(I12161),.A(g5971));
  NOT NOT1_3440(.VSS(VSS),.VDD(VDD),.Y(g6764),.A(I12161));
  NOT NOT1_3441(.VSS(VSS),.VDD(VDD),.Y(I12164),.A(g5847));
  NOT NOT1_3442(.VSS(VSS),.VDD(VDD),.Y(g6765),.A(I12164));
  NOT NOT1_3443(.VSS(VSS),.VDD(VDD),.Y(I12167),.A(g5939));
  NOT NOT1_3444(.VSS(VSS),.VDD(VDD),.Y(g6766),.A(I12167));
  NOT NOT1_3445(.VSS(VSS),.VDD(VDD),.Y(I12170),.A(g5956));
  NOT NOT1_3446(.VSS(VSS),.VDD(VDD),.Y(g6767),.A(I12170));
  NOT NOT1_3447(.VSS(VSS),.VDD(VDD),.Y(I12173),.A(g5918));
  NOT NOT1_3448(.VSS(VSS),.VDD(VDD),.Y(g6768),.A(I12173));
  NOT NOT1_3449(.VSS(VSS),.VDD(VDD),.Y(I12176),.A(g5939));
  NOT NOT1_3450(.VSS(VSS),.VDD(VDD),.Y(g6769),.A(I12176));
  NOT NOT1_3451(.VSS(VSS),.VDD(VDD),.Y(I12187),.A(g5897));
  NOT NOT1_3452(.VSS(VSS),.VDD(VDD),.Y(g6772),.A(I12187));
  NOT NOT1_3453(.VSS(VSS),.VDD(VDD),.Y(I12190),.A(g5918));
  NOT NOT1_3454(.VSS(VSS),.VDD(VDD),.Y(g6773),.A(I12190));
  NOT NOT1_3455(.VSS(VSS),.VDD(VDD),.Y(I12193),.A(g6468));
  NOT NOT1_3456(.VSS(VSS),.VDD(VDD),.Y(g6774),.A(I12193));
  NOT NOT1_3457(.VSS(VSS),.VDD(VDD),.Y(I12196),.A(g6471));
  NOT NOT1_3458(.VSS(VSS),.VDD(VDD),.Y(g6775),.A(I12196));
  NOT NOT1_3459(.VSS(VSS),.VDD(VDD),.Y(I12199),.A(g6475));
  NOT NOT1_3460(.VSS(VSS),.VDD(VDD),.Y(g6776),.A(I12199));
  NOT NOT1_3461(.VSS(VSS),.VDD(VDD),.Y(I12202),.A(g6481));
  NOT NOT1_3462(.VSS(VSS),.VDD(VDD),.Y(g6777),.A(I12202));
  NOT NOT1_3463(.VSS(VSS),.VDD(VDD),.Y(I12205),.A(g6488));
  NOT NOT1_3464(.VSS(VSS),.VDD(VDD),.Y(g6778),.A(I12205));
  NOT NOT1_3465(.VSS(VSS),.VDD(VDD),.Y(I12208),.A(g6496));
  NOT NOT1_3466(.VSS(VSS),.VDD(VDD),.Y(g6779),.A(I12208));
  NOT NOT1_3467(.VSS(VSS),.VDD(VDD),.Y(I12211),.A(g6502));
  NOT NOT1_3468(.VSS(VSS),.VDD(VDD),.Y(g6780),.A(I12211));
  NOT NOT1_3469(.VSS(VSS),.VDD(VDD),.Y(I12214),.A(g6507));
  NOT NOT1_3470(.VSS(VSS),.VDD(VDD),.Y(g6781),.A(I12214));
  NOT NOT1_3471(.VSS(VSS),.VDD(VDD),.Y(I12217),.A(g6631));
  NOT NOT1_3472(.VSS(VSS),.VDD(VDD),.Y(g6782),.A(I12217));
  NOT NOT1_3473(.VSS(VSS),.VDD(VDD),.Y(I12220),.A(g6645));
  NOT NOT1_3474(.VSS(VSS),.VDD(VDD),.Y(g6783),.A(I12220));
  NOT NOT1_3475(.VSS(VSS),.VDD(VDD),.Y(I12223),.A(g6655));
  NOT NOT1_3476(.VSS(VSS),.VDD(VDD),.Y(g6784),.A(I12223));
  NOT NOT1_3477(.VSS(VSS),.VDD(VDD),.Y(I12226),.A(g6636));
  NOT NOT1_3478(.VSS(VSS),.VDD(VDD),.Y(g6785),.A(I12226));
  NOT NOT1_3479(.VSS(VSS),.VDD(VDD),.Y(I12229),.A(g6659));
  NOT NOT1_3480(.VSS(VSS),.VDD(VDD),.Y(g6786),.A(I12229));
  NOT NOT1_3481(.VSS(VSS),.VDD(VDD),.Y(I12232),.A(g6662));
  NOT NOT1_3482(.VSS(VSS),.VDD(VDD),.Y(g6787),.A(I12232));
  NOT NOT1_3483(.VSS(VSS),.VDD(VDD),.Y(I12235),.A(g6634));
  NOT NOT1_3484(.VSS(VSS),.VDD(VDD),.Y(g6788),.A(I12235));
  NOT NOT1_3485(.VSS(VSS),.VDD(VDD),.Y(I12238),.A(g6637));
  NOT NOT1_3486(.VSS(VSS),.VDD(VDD),.Y(g6789),.A(I12238));
  NOT NOT1_3487(.VSS(VSS),.VDD(VDD),.Y(I12241),.A(g6640));
  NOT NOT1_3488(.VSS(VSS),.VDD(VDD),.Y(g6790),.A(I12241));
  NOT NOT1_3489(.VSS(VSS),.VDD(VDD),.Y(I12244),.A(g6642));
  NOT NOT1_3490(.VSS(VSS),.VDD(VDD),.Y(g6791),.A(I12244));
  NOT NOT1_3491(.VSS(VSS),.VDD(VDD),.Y(I12247),.A(g6646));
  NOT NOT1_3492(.VSS(VSS),.VDD(VDD),.Y(g6792),.A(I12247));
  NOT NOT1_3493(.VSS(VSS),.VDD(VDD),.Y(I12250),.A(g6651));
  NOT NOT1_3494(.VSS(VSS),.VDD(VDD),.Y(g6793),.A(I12250));
  NOT NOT1_3495(.VSS(VSS),.VDD(VDD),.Y(I12253),.A(g6427));
  NOT NOT1_3496(.VSS(VSS),.VDD(VDD),.Y(g6794),.A(I12253));
  NOT NOT1_3497(.VSS(VSS),.VDD(VDD),.Y(I12256),.A(g6647));
  NOT NOT1_3498(.VSS(VSS),.VDD(VDD),.Y(g6795),.A(I12256));
  NOT NOT1_3499(.VSS(VSS),.VDD(VDD),.Y(I12259),.A(g6652));
  NOT NOT1_3500(.VSS(VSS),.VDD(VDD),.Y(g6796),.A(I12259));
  NOT NOT1_3501(.VSS(VSS),.VDD(VDD),.Y(I12262),.A(g6656));
  NOT NOT1_3502(.VSS(VSS),.VDD(VDD),.Y(g6797),.A(I12262));
  NOT NOT1_3503(.VSS(VSS),.VDD(VDD),.Y(I12265),.A(g6660));
  NOT NOT1_3504(.VSS(VSS),.VDD(VDD),.Y(g6798),.A(I12265));
  NOT NOT1_3505(.VSS(VSS),.VDD(VDD),.Y(I12268),.A(g6661));
  NOT NOT1_3506(.VSS(VSS),.VDD(VDD),.Y(g6799),.A(I12268));
  NOT NOT1_3507(.VSS(VSS),.VDD(VDD),.Y(I12271),.A(g6663));
  NOT NOT1_3508(.VSS(VSS),.VDD(VDD),.Y(g6800),.A(I12271));
  NOT NOT1_3509(.VSS(VSS),.VDD(VDD),.Y(I12274),.A(g6672));
  NOT NOT1_3510(.VSS(VSS),.VDD(VDD),.Y(g6801),.A(I12274));
  NOT NOT1_3511(.VSS(VSS),.VDD(VDD),.Y(I12277),.A(g6681));
  NOT NOT1_3512(.VSS(VSS),.VDD(VDD),.Y(g6802),.A(I12277));
  NOT NOT1_3513(.VSS(VSS),.VDD(VDD),.Y(I12280),.A(g6684));
  NOT NOT1_3514(.VSS(VSS),.VDD(VDD),.Y(g6803),.A(I12280));
  NOT NOT1_3515(.VSS(VSS),.VDD(VDD),.Y(I12283),.A(g6692));
  NOT NOT1_3516(.VSS(VSS),.VDD(VDD),.Y(g6804),.A(I12283));
  NOT NOT1_3517(.VSS(VSS),.VDD(VDD),.Y(I12286),.A(g6696));
  NOT NOT1_3518(.VSS(VSS),.VDD(VDD),.Y(g6805),.A(I12286));
  NOT NOT1_3519(.VSS(VSS),.VDD(VDD),.Y(I12289),.A(g6702));
  NOT NOT1_3520(.VSS(VSS),.VDD(VDD),.Y(g6806),.A(I12289));
  NOT NOT1_3521(.VSS(VSS),.VDD(VDD),.Y(I12292),.A(g6657));
  NOT NOT1_3522(.VSS(VSS),.VDD(VDD),.Y(g6807),.A(I12292));
  NOT NOT1_3523(.VSS(VSS),.VDD(VDD),.Y(I12295),.A(g6693));
  NOT NOT1_3524(.VSS(VSS),.VDD(VDD),.Y(g6808),.A(I12295));
  NOT NOT1_3525(.VSS(VSS),.VDD(VDD),.Y(I12298),.A(g6697));
  NOT NOT1_3526(.VSS(VSS),.VDD(VDD),.Y(g6809),.A(I12298));
  NOT NOT1_3527(.VSS(VSS),.VDD(VDD),.Y(I12301),.A(g6703));
  NOT NOT1_3528(.VSS(VSS),.VDD(VDD),.Y(g6810),.A(I12301));
  NOT NOT1_3529(.VSS(VSS),.VDD(VDD),.Y(I12304),.A(g6711));
  NOT NOT1_3530(.VSS(VSS),.VDD(VDD),.Y(g6811),.A(I12304));
  NOT NOT1_3531(.VSS(VSS),.VDD(VDD),.Y(I12307),.A(g6712));
  NOT NOT1_3532(.VSS(VSS),.VDD(VDD),.Y(g6812),.A(I12307));
  NOT NOT1_3533(.VSS(VSS),.VDD(VDD),.Y(I12310),.A(g6723));
  NOT NOT1_3534(.VSS(VSS),.VDD(VDD),.Y(g6813),.A(I12310));
  NOT NOT1_3535(.VSS(VSS),.VDD(VDD),.Y(I12313),.A(g6730));
  NOT NOT1_3536(.VSS(VSS),.VDD(VDD),.Y(g6814),.A(I12313));
  NOT NOT1_3537(.VSS(VSS),.VDD(VDD),.Y(I12316),.A(g6736));
  NOT NOT1_3538(.VSS(VSS),.VDD(VDD),.Y(g6815),.A(I12316));
  NOT NOT1_3539(.VSS(VSS),.VDD(VDD),.Y(I12319),.A(g6741));
  NOT NOT1_3540(.VSS(VSS),.VDD(VDD),.Y(g6816),.A(I12319));
  NOT NOT1_3541(.VSS(VSS),.VDD(VDD),.Y(I12322),.A(g6751));
  NOT NOT1_3542(.VSS(VSS),.VDD(VDD),.Y(g6817),.A(I12322));
  NOT NOT1_3543(.VSS(VSS),.VDD(VDD),.Y(I12325),.A(g6755));
  NOT NOT1_3544(.VSS(VSS),.VDD(VDD),.Y(g6818),.A(I12325));
  NOT NOT1_3545(.VSS(VSS),.VDD(VDD),.Y(I12328),.A(g6760));
  NOT NOT1_3546(.VSS(VSS),.VDD(VDD),.Y(g6819),.A(I12328));
  NOT NOT1_3547(.VSS(VSS),.VDD(VDD),.Y(I12331),.A(g6704));
  NOT NOT1_3548(.VSS(VSS),.VDD(VDD),.Y(g6820),.A(I12331));
  NOT NOT1_3549(.VSS(VSS),.VDD(VDD),.Y(I12334),.A(g6713));
  NOT NOT1_3550(.VSS(VSS),.VDD(VDD),.Y(g6821),.A(I12334));
  NOT NOT1_3551(.VSS(VSS),.VDD(VDD),.Y(I12337),.A(g6724));
  NOT NOT1_3552(.VSS(VSS),.VDD(VDD),.Y(g6822),.A(I12337));
  NOT NOT1_3553(.VSS(VSS),.VDD(VDD),.Y(I12340),.A(g6725));
  NOT NOT1_3554(.VSS(VSS),.VDD(VDD),.Y(g6823),.A(I12340));
  NOT NOT1_3555(.VSS(VSS),.VDD(VDD),.Y(I12343),.A(g6731));
  NOT NOT1_3556(.VSS(VSS),.VDD(VDD),.Y(g6824),.A(I12343));
  NOT NOT1_3557(.VSS(VSS),.VDD(VDD),.Y(I12346),.A(g6737));
  NOT NOT1_3558(.VSS(VSS),.VDD(VDD),.Y(g6825),.A(I12346));
  NOT NOT1_3559(.VSS(VSS),.VDD(VDD),.Y(I12349),.A(g6742));
  NOT NOT1_3560(.VSS(VSS),.VDD(VDD),.Y(g6826),.A(I12349));
  NOT NOT1_3561(.VSS(VSS),.VDD(VDD),.Y(I12352),.A(g6752));
  NOT NOT1_3562(.VSS(VSS),.VDD(VDD),.Y(g6827),.A(I12352));
  NOT NOT1_3563(.VSS(VSS),.VDD(VDD),.Y(I12355),.A(g6756));
  NOT NOT1_3564(.VSS(VSS),.VDD(VDD),.Y(g6828),.A(I12355));
  NOT NOT1_3565(.VSS(VSS),.VDD(VDD),.Y(I12358),.A(g6761));
  NOT NOT1_3566(.VSS(VSS),.VDD(VDD),.Y(g6829),.A(I12358));
  NOT NOT1_3567(.VSS(VSS),.VDD(VDD),.Y(I12361),.A(g6765));
  NOT NOT1_3568(.VSS(VSS),.VDD(VDD),.Y(g6830),.A(I12361));
  NOT NOT1_3569(.VSS(VSS),.VDD(VDD),.Y(I12364),.A(g6714));
  NOT NOT1_3570(.VSS(VSS),.VDD(VDD),.Y(g6831),.A(I12364));
  NOT NOT1_3571(.VSS(VSS),.VDD(VDD),.Y(I12367),.A(g6754));
  NOT NOT1_3572(.VSS(VSS),.VDD(VDD),.Y(g6832),.A(I12367));
  NOT NOT1_3573(.VSS(VSS),.VDD(VDD),.Y(I12370),.A(g6758));
  NOT NOT1_3574(.VSS(VSS),.VDD(VDD),.Y(g6833),.A(I12370));
  NOT NOT1_3575(.VSS(VSS),.VDD(VDD),.Y(I12373),.A(g6763));
  NOT NOT1_3576(.VSS(VSS),.VDD(VDD),.Y(g6834),.A(I12373));
  NOT NOT1_3577(.VSS(VSS),.VDD(VDD),.Y(I12376),.A(g6766));
  NOT NOT1_3578(.VSS(VSS),.VDD(VDD),.Y(g6835),.A(I12376));
  NOT NOT1_3579(.VSS(VSS),.VDD(VDD),.Y(I12379),.A(g6768));
  NOT NOT1_3580(.VSS(VSS),.VDD(VDD),.Y(g6836),.A(I12379));
  NOT NOT1_3581(.VSS(VSS),.VDD(VDD),.Y(I12382),.A(g6772));
  NOT NOT1_3582(.VSS(VSS),.VDD(VDD),.Y(g6837),.A(I12382));
  NOT NOT1_3583(.VSS(VSS),.VDD(VDD),.Y(I12385),.A(g6397));
  NOT NOT1_3584(.VSS(VSS),.VDD(VDD),.Y(g6838),.A(I12385));
  NOT NOT1_3585(.VSS(VSS),.VDD(VDD),.Y(I12388),.A(g6403));
  NOT NOT1_3586(.VSS(VSS),.VDD(VDD),.Y(g6839),.A(I12388));
  NOT NOT1_3587(.VSS(VSS),.VDD(VDD),.Y(I12391),.A(g6744));
  NOT NOT1_3588(.VSS(VSS),.VDD(VDD),.Y(g6840),.A(I12391));
  NOT NOT1_3589(.VSS(VSS),.VDD(VDD),.Y(I12394),.A(g6759));
  NOT NOT1_3590(.VSS(VSS),.VDD(VDD),.Y(g6841),.A(I12394));
  NOT NOT1_3591(.VSS(VSS),.VDD(VDD),.Y(I12397),.A(g6764));
  NOT NOT1_3592(.VSS(VSS),.VDD(VDD),.Y(g6842),.A(I12397));
  NOT NOT1_3593(.VSS(VSS),.VDD(VDD),.Y(I12400),.A(g6767));
  NOT NOT1_3594(.VSS(VSS),.VDD(VDD),.Y(g6843),.A(I12400));
  NOT NOT1_3595(.VSS(VSS),.VDD(VDD),.Y(I12403),.A(g6769));
  NOT NOT1_3596(.VSS(VSS),.VDD(VDD),.Y(g6844),.A(I12403));
  NOT NOT1_3597(.VSS(VSS),.VDD(VDD),.Y(I12406),.A(g6773));
  NOT NOT1_3598(.VSS(VSS),.VDD(VDD),.Y(g6845),.A(I12406));
  NOT NOT1_3599(.VSS(VSS),.VDD(VDD),.Y(I12409),.A(g6398));
  NOT NOT1_3600(.VSS(VSS),.VDD(VDD),.Y(g6846),.A(I12409));
  NOT NOT1_3601(.VSS(VSS),.VDD(VDD),.Y(I12412),.A(g6404));
  NOT NOT1_3602(.VSS(VSS),.VDD(VDD),.Y(g6847),.A(I12412));
  NOT NOT1_3603(.VSS(VSS),.VDD(VDD),.Y(I12415),.A(g6410));
  NOT NOT1_3604(.VSS(VSS),.VDD(VDD),.Y(g6848),.A(I12415));
  NOT NOT1_3605(.VSS(VSS),.VDD(VDD),.Y(I12418),.A(g6572));
  NOT NOT1_3606(.VSS(VSS),.VDD(VDD),.Y(g6849),.A(I12418));
  NOT NOT1_3607(.VSS(VSS),.VDD(VDD),.Y(I12421),.A(g6486));
  NOT NOT1_3608(.VSS(VSS),.VDD(VDD),.Y(g6850),.A(I12421));
  NOT NOT1_3609(.VSS(VSS),.VDD(VDD),.Y(I12424),.A(g6446));
  NOT NOT1_3610(.VSS(VSS),.VDD(VDD),.Y(g6851),.A(I12424));
  NOT NOT1_3611(.VSS(VSS),.VDD(VDD),.Y(I12427),.A(g6553));
  NOT NOT1_3612(.VSS(VSS),.VDD(VDD),.Y(g6852),.A(I12427));
  NOT NOT1_3613(.VSS(VSS),.VDD(VDD),.Y(I12430),.A(g6432));
  NOT NOT1_3614(.VSS(VSS),.VDD(VDD),.Y(g6853),.A(I12430));
  NOT NOT1_3615(.VSS(VSS),.VDD(VDD),.Y(I12433),.A(g6632));
  NOT NOT1_3616(.VSS(VSS),.VDD(VDD),.Y(g6854),.A(I12433));
  NOT NOT1_3617(.VSS(VSS),.VDD(VDD),.Y(I12436),.A(g6635));
  NOT NOT1_3618(.VSS(VSS),.VDD(VDD),.Y(g6855),.A(I12436));
  NOT NOT1_3619(.VSS(VSS),.VDD(VDD),.Y(I12439),.A(g6566));
  NOT NOT1_3620(.VSS(VSS),.VDD(VDD),.Y(g6856),.A(I12439));
  NOT NOT1_3621(.VSS(VSS),.VDD(VDD),.Y(I12442),.A(g6542));
  NOT NOT1_3622(.VSS(VSS),.VDD(VDD),.Y(g6857),.A(I12442));
  NOT NOT1_3623(.VSS(VSS),.VDD(VDD),.Y(I12445),.A(g6568));
  NOT NOT1_3624(.VSS(VSS),.VDD(VDD),.Y(g6858),.A(I12445));
  NOT NOT1_3625(.VSS(VSS),.VDD(VDD),.Y(I12448),.A(g6569));
  NOT NOT1_3626(.VSS(VSS),.VDD(VDD),.Y(g6859),.A(I12448));
  NOT NOT1_3627(.VSS(VSS),.VDD(VDD),.Y(I12451),.A(g6524));
  NOT NOT1_3628(.VSS(VSS),.VDD(VDD),.Y(g6860),.A(I12451));
  NOT NOT1_3629(.VSS(VSS),.VDD(VDD),.Y(I12454),.A(g6581));
  NOT NOT1_3630(.VSS(VSS),.VDD(VDD),.Y(g6861),.A(I12454));
  NOT NOT1_3631(.VSS(VSS),.VDD(VDD),.Y(I12457),.A(g6671));
  NOT NOT1_3632(.VSS(VSS),.VDD(VDD),.Y(g6862),.A(I12457));
  NOT NOT1_3633(.VSS(VSS),.VDD(VDD),.Y(I12460),.A(g6674));
  NOT NOT1_3634(.VSS(VSS),.VDD(VDD),.Y(g6863),.A(I12460));
  NOT NOT1_3635(.VSS(VSS),.VDD(VDD),.Y(I12463),.A(g6682));
  NOT NOT1_3636(.VSS(VSS),.VDD(VDD),.Y(g6864),.A(I12463));
  NOT NOT1_3637(.VSS(VSS),.VDD(VDD),.Y(I12466),.A(g6687));
  NOT NOT1_3638(.VSS(VSS),.VDD(VDD),.Y(g6865),.A(I12466));
  NOT NOT1_3639(.VSS(VSS),.VDD(VDD),.Y(I12469),.A(g6586));
  NOT NOT1_3640(.VSS(VSS),.VDD(VDD),.Y(g6866),.A(I12469));
  NOT NOT1_3641(.VSS(VSS),.VDD(VDD),.Y(I12472),.A(g6591));
  NOT NOT1_3642(.VSS(VSS),.VDD(VDD),.Y(g6867),.A(I12472));
  NOT NOT1_3643(.VSS(VSS),.VDD(VDD),.Y(I12475),.A(g6596));
  NOT NOT1_3644(.VSS(VSS),.VDD(VDD),.Y(g6868),.A(I12475));
  NOT NOT1_3645(.VSS(VSS),.VDD(VDD),.Y(I12478),.A(g6603));
  NOT NOT1_3646(.VSS(VSS),.VDD(VDD),.Y(g6869),.A(I12478));
  NOT NOT1_3647(.VSS(VSS),.VDD(VDD),.Y(I12481),.A(g6616));
  NOT NOT1_3648(.VSS(VSS),.VDD(VDD),.Y(g6870),.A(I12481));
  NOT NOT1_3649(.VSS(VSS),.VDD(VDD),.Y(I12484),.A(g6621));
  NOT NOT1_3650(.VSS(VSS),.VDD(VDD),.Y(g6871),.A(I12484));
  NOT NOT1_3651(.VSS(VSS),.VDD(VDD),.Y(I12487),.A(g6623));
  NOT NOT1_3652(.VSS(VSS),.VDD(VDD),.Y(g6872),.A(I12487));
  NOT NOT1_3653(.VSS(VSS),.VDD(VDD),.Y(I12490),.A(g6625));
  NOT NOT1_3654(.VSS(VSS),.VDD(VDD),.Y(g6873),.A(I12490));
  NOT NOT1_3655(.VSS(VSS),.VDD(VDD),.Y(I12493),.A(g6587));
  NOT NOT1_3656(.VSS(VSS),.VDD(VDD),.Y(g6874),.A(I12493));
  NOT NOT1_3657(.VSS(VSS),.VDD(VDD),.Y(I12496),.A(g6592));
  NOT NOT1_3658(.VSS(VSS),.VDD(VDD),.Y(g6875),.A(I12496));
  NOT NOT1_3659(.VSS(VSS),.VDD(VDD),.Y(I12499),.A(g6597));
  NOT NOT1_3660(.VSS(VSS),.VDD(VDD),.Y(g6876),.A(I12499));
  NOT NOT1_3661(.VSS(VSS),.VDD(VDD),.Y(I12502),.A(g6604));
  NOT NOT1_3662(.VSS(VSS),.VDD(VDD),.Y(g6877),.A(I12502));
  NOT NOT1_3663(.VSS(VSS),.VDD(VDD),.Y(I12505),.A(g6612));
  NOT NOT1_3664(.VSS(VSS),.VDD(VDD),.Y(g6878),.A(I12505));
  NOT NOT1_3665(.VSS(VSS),.VDD(VDD),.Y(I12508),.A(g6593));
  NOT NOT1_3666(.VSS(VSS),.VDD(VDD),.Y(g6879),.A(I12508));
  NOT NOT1_3667(.VSS(VSS),.VDD(VDD),.Y(I12511),.A(g6598));
  NOT NOT1_3668(.VSS(VSS),.VDD(VDD),.Y(g6880),.A(I12511));
  NOT NOT1_3669(.VSS(VSS),.VDD(VDD),.Y(I12514),.A(g6605));
  NOT NOT1_3670(.VSS(VSS),.VDD(VDD),.Y(g6881),.A(I12514));
  NOT NOT1_3671(.VSS(VSS),.VDD(VDD),.Y(I12517),.A(g6613));
  NOT NOT1_3672(.VSS(VSS),.VDD(VDD),.Y(g6882),.A(I12517));
  NOT NOT1_3673(.VSS(VSS),.VDD(VDD),.Y(I12520),.A(g6622));
  NOT NOT1_3674(.VSS(VSS),.VDD(VDD),.Y(g6883),.A(I12520));
  NOT NOT1_3675(.VSS(VSS),.VDD(VDD),.Y(I12523),.A(g6624));
  NOT NOT1_3676(.VSS(VSS),.VDD(VDD),.Y(g6884),.A(I12523));
  NOT NOT1_3677(.VSS(VSS),.VDD(VDD),.Y(I12526),.A(g6626));
  NOT NOT1_3678(.VSS(VSS),.VDD(VDD),.Y(g6885),.A(I12526));
  NOT NOT1_3679(.VSS(VSS),.VDD(VDD),.Y(I12529),.A(g6628));
  NOT NOT1_3680(.VSS(VSS),.VDD(VDD),.Y(g6886),.A(I12529));
  NOT NOT1_3681(.VSS(VSS),.VDD(VDD),.Y(I12532),.A(g6594));
  NOT NOT1_3682(.VSS(VSS),.VDD(VDD),.Y(g6887),.A(I12532));
  NOT NOT1_3683(.VSS(VSS),.VDD(VDD),.Y(I12535),.A(g6599));
  NOT NOT1_3684(.VSS(VSS),.VDD(VDD),.Y(g6888),.A(I12535));
  NOT NOT1_3685(.VSS(VSS),.VDD(VDD),.Y(I12538),.A(g6606));
  NOT NOT1_3686(.VSS(VSS),.VDD(VDD),.Y(g6889),.A(I12538));
  NOT NOT1_3687(.VSS(VSS),.VDD(VDD),.Y(I12541),.A(g6614));
  NOT NOT1_3688(.VSS(VSS),.VDD(VDD),.Y(g6890),.A(I12541));
  NOT NOT1_3689(.VSS(VSS),.VDD(VDD),.Y(I12544),.A(g6617));
  NOT NOT1_3690(.VSS(VSS),.VDD(VDD),.Y(g6891),.A(I12544));
  NOT NOT1_3691(.VSS(VSS),.VDD(VDD),.Y(I12547),.A(g6708));
  NOT NOT1_3692(.VSS(VSS),.VDD(VDD),.Y(g6892),.A(I12547));
  NOT NOT1_3693(.VSS(VSS),.VDD(VDD),.Y(g6894),.A(g6525));
  NOT NOT1_3694(.VSS(VSS),.VDD(VDD),.Y(I12558),.A(g6449));
  NOT NOT1_3695(.VSS(VSS),.VDD(VDD),.Y(g6895),.A(I12558));
  NOT NOT1_3696(.VSS(VSS),.VDD(VDD),.Y(I12561),.A(g6449));
  NOT NOT1_3697(.VSS(VSS),.VDD(VDD),.Y(g6896),.A(I12561));
  NOT NOT1_3698(.VSS(VSS),.VDD(VDD),.Y(I12564),.A(g6720));
  NOT NOT1_3699(.VSS(VSS),.VDD(VDD),.Y(g6897),.A(I12564));
  NOT NOT1_3700(.VSS(VSS),.VDD(VDD),.Y(I12567),.A(g6721));
  NOT NOT1_3701(.VSS(VSS),.VDD(VDD),.Y(g6898),.A(I12567));
  NOT NOT1_3702(.VSS(VSS),.VDD(VDD),.Y(g6899),.A(g6525));
  NOT NOT1_3703(.VSS(VSS),.VDD(VDD),.Y(I12571),.A(g6729));
  NOT NOT1_3704(.VSS(VSS),.VDD(VDD),.Y(g6900),.A(I12571));
  NOT NOT1_3705(.VSS(VSS),.VDD(VDD),.Y(g6901),.A(g6525));
  NOT NOT1_3706(.VSS(VSS),.VDD(VDD),.Y(I12582),.A(g6745));
  NOT NOT1_3707(.VSS(VSS),.VDD(VDD),.Y(g6903),.A(I12582));
  NOT NOT1_3708(.VSS(VSS),.VDD(VDD),.Y(g6904),.A(g6426));
  NOT NOT1_3709(.VSS(VSS),.VDD(VDD),.Y(I12586),.A(g6643));
  NOT NOT1_3710(.VSS(VSS),.VDD(VDD),.Y(g6905),.A(I12586));
  NOT NOT1_3711(.VSS(VSS),.VDD(VDD),.Y(I12592),.A(g1008));
  NOT NOT1_3712(.VSS(VSS),.VDD(VDD),.Y(g6909),.A(I12592));
  NOT NOT1_3713(.VSS(VSS),.VDD(VDD),.Y(I12609),.A(g6571));
  NOT NOT1_3714(.VSS(VSS),.VDD(VDD),.Y(g6918),.A(I12609));
  NOT NOT1_3715(.VSS(VSS),.VDD(VDD),.Y(g6922),.A(g6525));
  NOT NOT1_3716(.VSS(VSS),.VDD(VDD),.Y(I12629),.A(g6523));
  NOT NOT1_3717(.VSS(VSS),.VDD(VDD),.Y(g6936),.A(I12629));
  NOT NOT1_3718(.VSS(VSS),.VDD(VDD),.Y(I12632),.A(g6514));
  NOT NOT1_3719(.VSS(VSS),.VDD(VDD),.Y(g6937),.A(I12632));
  NOT NOT1_3720(.VSS(VSS),.VDD(VDD),.Y(I12635),.A(g6509));
  NOT NOT1_3721(.VSS(VSS),.VDD(VDD),.Y(g6938),.A(I12635));
  NOT NOT1_3722(.VSS(VSS),.VDD(VDD),.Y(g6939),.A(g6543));
  NOT NOT1_3723(.VSS(VSS),.VDD(VDD),.Y(I12639),.A(g6506));
  NOT NOT1_3724(.VSS(VSS),.VDD(VDD),.Y(g6940),.A(I12639));
  NOT NOT1_3725(.VSS(VSS),.VDD(VDD),.Y(I12643),.A(g6501));
  NOT NOT1_3726(.VSS(VSS),.VDD(VDD),.Y(g6944),.A(I12643));
  NOT NOT1_3727(.VSS(VSS),.VDD(VDD),.Y(I12646),.A(g6493));
  NOT NOT1_3728(.VSS(VSS),.VDD(VDD),.Y(g6945),.A(I12646));
  NOT NOT1_3729(.VSS(VSS),.VDD(VDD),.Y(I12649),.A(g6457));
  NOT NOT1_3730(.VSS(VSS),.VDD(VDD),.Y(g6946),.A(I12649));
  NOT NOT1_3731(.VSS(VSS),.VDD(VDD),.Y(I12652),.A(g6664));
  NOT NOT1_3732(.VSS(VSS),.VDD(VDD),.Y(g6947),.A(I12652));
  NOT NOT1_3733(.VSS(VSS),.VDD(VDD),.Y(I12655),.A(g6458));
  NOT NOT1_3734(.VSS(VSS),.VDD(VDD),.Y(g6948),.A(I12655));
  NOT NOT1_3735(.VSS(VSS),.VDD(VDD),.Y(I12659),.A(g6459));
  NOT NOT1_3736(.VSS(VSS),.VDD(VDD),.Y(g6950),.A(I12659));
  NOT NOT1_3737(.VSS(VSS),.VDD(VDD),.Y(g6953),.A(g6745));
  NOT NOT1_3738(.VSS(VSS),.VDD(VDD),.Y(I12666),.A(g6476));
  NOT NOT1_3739(.VSS(VSS),.VDD(VDD),.Y(g6955),.A(I12666));
  NOT NOT1_3740(.VSS(VSS),.VDD(VDD),.Y(I12669),.A(g6477));
  NOT NOT1_3741(.VSS(VSS),.VDD(VDD),.Y(g6956),.A(I12669));
  NOT NOT1_3742(.VSS(VSS),.VDD(VDD),.Y(I12672),.A(g6473));
  NOT NOT1_3743(.VSS(VSS),.VDD(VDD),.Y(g6957),.A(I12672));
  NOT NOT1_3744(.VSS(VSS),.VDD(VDD),.Y(I12675),.A(g6510));
  NOT NOT1_3745(.VSS(VSS),.VDD(VDD),.Y(g6958),.A(I12675));
  NOT NOT1_3746(.VSS(VSS),.VDD(VDD),.Y(I12678),.A(g6516));
  NOT NOT1_3747(.VSS(VSS),.VDD(VDD),.Y(g6959),.A(I12678));
  NOT NOT1_3748(.VSS(VSS),.VDD(VDD),.Y(I12681),.A(g6469));
  NOT NOT1_3749(.VSS(VSS),.VDD(VDD),.Y(g6960),.A(I12681));
  NOT NOT1_3750(.VSS(VSS),.VDD(VDD),.Y(I12684),.A(g6472));
  NOT NOT1_3751(.VSS(VSS),.VDD(VDD),.Y(g6961),.A(I12684));
  NOT NOT1_3752(.VSS(VSS),.VDD(VDD),.Y(I12687),.A(g6745));
  NOT NOT1_3753(.VSS(VSS),.VDD(VDD),.Y(g6962),.A(I12687));
  NOT NOT1_3754(.VSS(VSS),.VDD(VDD),.Y(I12690),.A(g6467));
  NOT NOT1_3755(.VSS(VSS),.VDD(VDD),.Y(g6963),.A(I12690));
  NOT NOT1_3756(.VSS(VSS),.VDD(VDD),.Y(I12696),.A(g6503));
  NOT NOT1_3757(.VSS(VSS),.VDD(VDD),.Y(g6967),.A(I12696));
  NOT NOT1_3758(.VSS(VSS),.VDD(VDD),.Y(I12699),.A(g6504));
  NOT NOT1_3759(.VSS(VSS),.VDD(VDD),.Y(g6968),.A(I12699));
  NOT NOT1_3760(.VSS(VSS),.VDD(VDD),.Y(I12702),.A(g6497));
  NOT NOT1_3761(.VSS(VSS),.VDD(VDD),.Y(g6969),.A(I12702));
  NOT NOT1_3762(.VSS(VSS),.VDD(VDD),.Y(I12708),.A(g6482));
  NOT NOT1_3763(.VSS(VSS),.VDD(VDD),.Y(g6973),.A(I12708));
  NOT NOT1_3764(.VSS(VSS),.VDD(VDD),.Y(I12712),.A(g6543));
  NOT NOT1_3765(.VSS(VSS),.VDD(VDD),.Y(g6975),.A(I12712));
  NOT NOT1_3766(.VSS(VSS),.VDD(VDD),.Y(g6977),.A(g6664));
  NOT NOT1_3767(.VSS(VSS),.VDD(VDD),.Y(I12717),.A(g6543));
  NOT NOT1_3768(.VSS(VSS),.VDD(VDD),.Y(g6978),.A(I12717));
  NOT NOT1_3769(.VSS(VSS),.VDD(VDD),.Y(I12722),.A(g6611));
  NOT NOT1_3770(.VSS(VSS),.VDD(VDD),.Y(g6983),.A(I12722));
  NOT NOT1_3771(.VSS(VSS),.VDD(VDD),.Y(I12725),.A(g6565));
  NOT NOT1_3772(.VSS(VSS),.VDD(VDD),.Y(g6984),.A(I12725));
  NOT NOT1_3773(.VSS(VSS),.VDD(VDD),.Y(I12731),.A(g6579));
  NOT NOT1_3774(.VSS(VSS),.VDD(VDD),.Y(g6993),.A(I12731));
  NOT NOT1_3775(.VSS(VSS),.VDD(VDD),.Y(I12737),.A(g6460));
  NOT NOT1_3776(.VSS(VSS),.VDD(VDD),.Y(g6997),.A(I12737));
  NOT NOT1_3777(.VSS(VSS),.VDD(VDD),.Y(I12742),.A(g6590));
  NOT NOT1_3778(.VSS(VSS),.VDD(VDD),.Y(g7000),.A(I12742));
  NOT NOT1_3779(.VSS(VSS),.VDD(VDD),.Y(I12748),.A(g6585));
  NOT NOT1_3780(.VSS(VSS),.VDD(VDD),.Y(g7006),.A(I12748));
  NOT NOT1_3781(.VSS(VSS),.VDD(VDD),.Y(I12753),.A(g6445));
  NOT NOT1_3782(.VSS(VSS),.VDD(VDD),.Y(g7009),.A(I12753));
  NOT NOT1_3783(.VSS(VSS),.VDD(VDD),.Y(I12757),.A(g6577));
  NOT NOT1_3784(.VSS(VSS),.VDD(VDD),.Y(g7013),.A(I12757));
  NOT NOT1_3785(.VSS(VSS),.VDD(VDD),.Y(I12760),.A(g6685));
  NOT NOT1_3786(.VSS(VSS),.VDD(VDD),.Y(g7014),.A(I12760));
  NOT NOT1_3787(.VSS(VSS),.VDD(VDD),.Y(I12763),.A(g6686));
  NOT NOT1_3788(.VSS(VSS),.VDD(VDD),.Y(g7015),.A(I12763));
  NOT NOT1_3789(.VSS(VSS),.VDD(VDD),.Y(I12768),.A(g6718));
  NOT NOT1_3790(.VSS(VSS),.VDD(VDD),.Y(g7018),.A(I12768));
  NOT NOT1_3791(.VSS(VSS),.VDD(VDD),.Y(I12771),.A(g6735));
  NOT NOT1_3792(.VSS(VSS),.VDD(VDD),.Y(g7019),.A(I12771));
  NOT NOT1_3793(.VSS(VSS),.VDD(VDD),.Y(I12776),.A(g6739));
  NOT NOT1_3794(.VSS(VSS),.VDD(VDD),.Y(g7022),.A(I12776));
  NOT NOT1_3795(.VSS(VSS),.VDD(VDD),.Y(I12779),.A(g6740));
  NOT NOT1_3796(.VSS(VSS),.VDD(VDD),.Y(g7023),.A(I12779));
  NOT NOT1_3797(.VSS(VSS),.VDD(VDD),.Y(I12782),.A(g6463));
  NOT NOT1_3798(.VSS(VSS),.VDD(VDD),.Y(g7024),.A(I12782));
  NOT NOT1_3799(.VSS(VSS),.VDD(VDD),.Y(g7028),.A(g6525));
  NOT NOT1_3800(.VSS(VSS),.VDD(VDD),.Y(g7032),.A(g6525));
  NOT NOT1_3801(.VSS(VSS),.VDD(VDD),.Y(g7034),.A(g6525));
  NOT NOT1_3802(.VSS(VSS),.VDD(VDD),.Y(g7035),.A(g6543));
  NOT NOT1_3803(.VSS(VSS),.VDD(VDD),.Y(g7037),.A(g6525));
  NOT NOT1_3804(.VSS(VSS),.VDD(VDD),.Y(g7039),.A(g6543));
  NOT NOT1_3805(.VSS(VSS),.VDD(VDD),.Y(g7042),.A(g6543));
  NOT NOT1_3806(.VSS(VSS),.VDD(VDD),.Y(g7043),.A(g6543));
  NOT NOT1_3807(.VSS(VSS),.VDD(VDD),.Y(g7044),.A(g6543));
  NOT NOT1_3808(.VSS(VSS),.VDD(VDD),.Y(g7045),.A(g6490));
  NOT NOT1_3809(.VSS(VSS),.VDD(VDD),.Y(I12806),.A(g6602));
  NOT NOT1_3810(.VSS(VSS),.VDD(VDD),.Y(g7046),.A(I12806));
  NOT NOT1_3811(.VSS(VSS),.VDD(VDD),.Y(g7047),.A(g6498));
  NOT NOT1_3812(.VSS(VSS),.VDD(VDD),.Y(I12810),.A(g6607));
  NOT NOT1_3813(.VSS(VSS),.VDD(VDD),.Y(g7048),.A(I12810));
  NOT NOT1_3814(.VSS(VSS),.VDD(VDD),.Y(I12813),.A(g6607));
  NOT NOT1_3815(.VSS(VSS),.VDD(VDD),.Y(g7049),.A(I12813));
  NOT NOT1_3816(.VSS(VSS),.VDD(VDD),.Y(g7050),.A(g6618));
  NOT NOT1_3817(.VSS(VSS),.VDD(VDD),.Y(g7054),.A(g6511));
  NOT NOT1_3818(.VSS(VSS),.VDD(VDD),.Y(g7055),.A(g6517));
  NOT NOT1_3819(.VSS(VSS),.VDD(VDD),.Y(g7056),.A(g6520));
  NOT NOT1_3820(.VSS(VSS),.VDD(VDD),.Y(g7057),.A(g6644));
  NOT NOT1_3821(.VSS(VSS),.VDD(VDD),.Y(g7058),.A(g6649));
  NOT NOT1_3822(.VSS(VSS),.VDD(VDD),.Y(g7059),.A(g6538));
  NOT NOT1_3823(.VSS(VSS),.VDD(VDD),.Y(g7060),.A(g6654));
  NOT NOT1_3824(.VSS(VSS),.VDD(VDD),.Y(g7061),.A(g6650));
  NOT NOT1_3825(.VSS(VSS),.VDD(VDD),.Y(I12826),.A(g6441));
  NOT NOT1_3826(.VSS(VSS),.VDD(VDD),.Y(g7063),.A(I12826));
  NOT NOT1_3827(.VSS(VSS),.VDD(VDD),.Y(I12829),.A(g6441));
  NOT NOT1_3828(.VSS(VSS),.VDD(VDD),.Y(g7064),.A(I12829));
  NOT NOT1_3829(.VSS(VSS),.VDD(VDD),.Y(I12839),.A(g6630));
  NOT NOT1_3830(.VSS(VSS),.VDD(VDD),.Y(g7066),.A(I12839));
  NOT NOT1_3831(.VSS(VSS),.VDD(VDD),.Y(g7067),.A(g6658));
  NOT NOT1_3832(.VSS(VSS),.VDD(VDD),.Y(g7068),.A(g6556));
  NOT NOT1_3833(.VSS(VSS),.VDD(VDD),.Y(g7070),.A(g6562));
  NOT NOT1_3834(.VSS(VSS),.VDD(VDD),.Y(g7077),.A(g6676));
  NOT NOT1_3835(.VSS(VSS),.VDD(VDD),.Y(g7078),.A(g6683));
  NOT NOT1_3836(.VSS(VSS),.VDD(VDD),.Y(g7090),.A(g6525));
  NOT NOT1_3837(.VSS(VSS),.VDD(VDD),.Y(g7091),.A(g6525));
  NOT NOT1_3838(.VSS(VSS),.VDD(VDD),.Y(I12866),.A(g6483));
  NOT NOT1_3839(.VSS(VSS),.VDD(VDD),.Y(g7092),.A(I12866));
  NOT NOT1_3840(.VSS(VSS),.VDD(VDD),.Y(g7094),.A(g6525));
  NOT NOT1_3841(.VSS(VSS),.VDD(VDD),.Y(I12877),.A(g6700));
  NOT NOT1_3842(.VSS(VSS),.VDD(VDD),.Y(g7095),.A(I12877));
  NOT NOT1_3843(.VSS(VSS),.VDD(VDD),.Y(I12881),.A(g6478));
  NOT NOT1_3844(.VSS(VSS),.VDD(VDD),.Y(g7097),.A(I12881));
  NOT NOT1_3845(.VSS(VSS),.VDD(VDD),.Y(g7098),.A(g6525));
  NOT NOT1_3846(.VSS(VSS),.VDD(VDD),.Y(I12885),.A(g6946));
  NOT NOT1_3847(.VSS(VSS),.VDD(VDD),.Y(g7099),.A(I12885));
  NOT NOT1_3848(.VSS(VSS),.VDD(VDD),.Y(I12888),.A(g6948));
  NOT NOT1_3849(.VSS(VSS),.VDD(VDD),.Y(g7100),.A(I12888));
  NOT NOT1_3850(.VSS(VSS),.VDD(VDD),.Y(I12891),.A(g6950));
  NOT NOT1_3851(.VSS(VSS),.VDD(VDD),.Y(g7101),.A(I12891));
  NOT NOT1_3852(.VSS(VSS),.VDD(VDD),.Y(I12894),.A(g7009));
  NOT NOT1_3853(.VSS(VSS),.VDD(VDD),.Y(g7102),.A(I12894));
  NOT NOT1_3854(.VSS(VSS),.VDD(VDD),.Y(I12897),.A(g6962));
  NOT NOT1_3855(.VSS(VSS),.VDD(VDD),.Y(g7103),.A(I12897));
  NOT NOT1_3856(.VSS(VSS),.VDD(VDD),.Y(I12900),.A(g6947));
  NOT NOT1_3857(.VSS(VSS),.VDD(VDD),.Y(g7104),.A(I12900));
  NOT NOT1_3858(.VSS(VSS),.VDD(VDD),.Y(I12903),.A(g6905));
  NOT NOT1_3859(.VSS(VSS),.VDD(VDD),.Y(g7105),.A(I12903));
  NOT NOT1_3860(.VSS(VSS),.VDD(VDD),.Y(I12906),.A(g6918));
  NOT NOT1_3861(.VSS(VSS),.VDD(VDD),.Y(g7106),.A(I12906));
  NOT NOT1_3862(.VSS(VSS),.VDD(VDD),.Y(I12909),.A(g7046));
  NOT NOT1_3863(.VSS(VSS),.VDD(VDD),.Y(g7107),.A(I12909));
  NOT NOT1_3864(.VSS(VSS),.VDD(VDD),.Y(I12912),.A(g7006));
  NOT NOT1_3865(.VSS(VSS),.VDD(VDD),.Y(g7108),.A(I12912));
  NOT NOT1_3866(.VSS(VSS),.VDD(VDD),.Y(I12915),.A(g7000));
  NOT NOT1_3867(.VSS(VSS),.VDD(VDD),.Y(g7109),.A(I12915));
  NOT NOT1_3868(.VSS(VSS),.VDD(VDD),.Y(I12918),.A(g7013));
  NOT NOT1_3869(.VSS(VSS),.VDD(VDD),.Y(g7110),.A(I12918));
  NOT NOT1_3870(.VSS(VSS),.VDD(VDD),.Y(I12921),.A(g6993));
  NOT NOT1_3871(.VSS(VSS),.VDD(VDD),.Y(g7111),.A(I12921));
  NOT NOT1_3872(.VSS(VSS),.VDD(VDD),.Y(I12924),.A(g6983));
  NOT NOT1_3873(.VSS(VSS),.VDD(VDD),.Y(g7112),.A(I12924));
  NOT NOT1_3874(.VSS(VSS),.VDD(VDD),.Y(I12927),.A(g7014));
  NOT NOT1_3875(.VSS(VSS),.VDD(VDD),.Y(g7113),.A(I12927));
  NOT NOT1_3876(.VSS(VSS),.VDD(VDD),.Y(I12930),.A(g7019));
  NOT NOT1_3877(.VSS(VSS),.VDD(VDD),.Y(g7114),.A(I12930));
  NOT NOT1_3878(.VSS(VSS),.VDD(VDD),.Y(I12933),.A(g7018));
  NOT NOT1_3879(.VSS(VSS),.VDD(VDD),.Y(g7115),.A(I12933));
  NOT NOT1_3880(.VSS(VSS),.VDD(VDD),.Y(I12936),.A(g7015));
  NOT NOT1_3881(.VSS(VSS),.VDD(VDD),.Y(g7116),.A(I12936));
  NOT NOT1_3882(.VSS(VSS),.VDD(VDD),.Y(I12939),.A(g7022));
  NOT NOT1_3883(.VSS(VSS),.VDD(VDD),.Y(g7117),.A(I12939));
  NOT NOT1_3884(.VSS(VSS),.VDD(VDD),.Y(I12942),.A(g7023));
  NOT NOT1_3885(.VSS(VSS),.VDD(VDD),.Y(g7118),.A(I12942));
  NOT NOT1_3886(.VSS(VSS),.VDD(VDD),.Y(I12945),.A(g7066));
  NOT NOT1_3887(.VSS(VSS),.VDD(VDD),.Y(g7119),.A(I12945));
  NOT NOT1_3888(.VSS(VSS),.VDD(VDD),.Y(I12948),.A(g6919));
  NOT NOT1_3889(.VSS(VSS),.VDD(VDD),.Y(g7120),.A(I12948));
  NOT NOT1_3890(.VSS(VSS),.VDD(VDD),.Y(I12958),.A(g6920));
  NOT NOT1_3891(.VSS(VSS),.VDD(VDD),.Y(g7122),.A(I12958));
  NOT NOT1_3892(.VSS(VSS),.VDD(VDD),.Y(I12961),.A(g6921));
  NOT NOT1_3893(.VSS(VSS),.VDD(VDD),.Y(g7123),.A(I12961));
  NOT NOT1_3894(.VSS(VSS),.VDD(VDD),.Y(g7124),.A(g6896));
  NOT NOT1_3895(.VSS(VSS),.VDD(VDD),.Y(I12965),.A(g6924));
  NOT NOT1_3896(.VSS(VSS),.VDD(VDD),.Y(g7125),.A(I12965));
  NOT NOT1_3897(.VSS(VSS),.VDD(VDD),.Y(I12968),.A(g6925));
  NOT NOT1_3898(.VSS(VSS),.VDD(VDD),.Y(g7126),.A(I12968));
  NOT NOT1_3899(.VSS(VSS),.VDD(VDD),.Y(g7127),.A(g6974));
  NOT NOT1_3900(.VSS(VSS),.VDD(VDD),.Y(I12973),.A(g6927));
  NOT NOT1_3901(.VSS(VSS),.VDD(VDD),.Y(g7129),.A(I12973));
  NOT NOT1_3902(.VSS(VSS),.VDD(VDD),.Y(I12976),.A(g6928));
  NOT NOT1_3903(.VSS(VSS),.VDD(VDD),.Y(g7130),.A(I12976));
  NOT NOT1_3904(.VSS(VSS),.VDD(VDD),.Y(g7131),.A(g6976));
  NOT NOT1_3905(.VSS(VSS),.VDD(VDD),.Y(I12980),.A(g6929));
  NOT NOT1_3906(.VSS(VSS),.VDD(VDD),.Y(g7132),.A(I12980));
  NOT NOT1_3907(.VSS(VSS),.VDD(VDD),.Y(I12983),.A(g6930));
  NOT NOT1_3908(.VSS(VSS),.VDD(VDD),.Y(g7133),.A(I12983));
  NOT NOT1_3909(.VSS(VSS),.VDD(VDD),.Y(I12986),.A(g6931));
  NOT NOT1_3910(.VSS(VSS),.VDD(VDD),.Y(g7134),.A(I12986));
  NOT NOT1_3911(.VSS(VSS),.VDD(VDD),.Y(I12989),.A(g6932));
  NOT NOT1_3912(.VSS(VSS),.VDD(VDD),.Y(g7135),.A(I12989));
  NOT NOT1_3913(.VSS(VSS),.VDD(VDD),.Y(I12993),.A(g6933));
  NOT NOT1_3914(.VSS(VSS),.VDD(VDD),.Y(g7137),.A(I12993));
  NOT NOT1_3915(.VSS(VSS),.VDD(VDD),.Y(I12996),.A(g6934));
  NOT NOT1_3916(.VSS(VSS),.VDD(VDD),.Y(g7138),.A(I12996));
  NOT NOT1_3917(.VSS(VSS),.VDD(VDD),.Y(I12999),.A(g7029));
  NOT NOT1_3918(.VSS(VSS),.VDD(VDD),.Y(g7139),.A(I12999));
  NOT NOT1_3919(.VSS(VSS),.VDD(VDD),.Y(I13009),.A(g6935));
  NOT NOT1_3920(.VSS(VSS),.VDD(VDD),.Y(g7141),.A(I13009));
  NOT NOT1_3921(.VSS(VSS),.VDD(VDD),.Y(I13012),.A(g7071));
  NOT NOT1_3922(.VSS(VSS),.VDD(VDD),.Y(g7142),.A(I13012));
  NOT NOT1_3923(.VSS(VSS),.VDD(VDD),.Y(g7143),.A(g6996));
  NOT NOT1_3924(.VSS(VSS),.VDD(VDD),.Y(I13023),.A(g7040));
  NOT NOT1_3925(.VSS(VSS),.VDD(VDD),.Y(g7145),.A(I13023));
  NOT NOT1_3926(.VSS(VSS),.VDD(VDD),.Y(g7146),.A(g6998));
  NOT NOT1_3927(.VSS(VSS),.VDD(VDD),.Y(g7147),.A(g6904));
  NOT NOT1_3928(.VSS(VSS),.VDD(VDD),.Y(I13028),.A(g7087));
  NOT NOT1_3929(.VSS(VSS),.VDD(VDD),.Y(g7148),.A(I13028));
  NOT NOT1_3930(.VSS(VSS),.VDD(VDD),.Y(I13031),.A(g6984));
  NOT NOT1_3931(.VSS(VSS),.VDD(VDD),.Y(g7149),.A(I13031));
  NOT NOT1_3932(.VSS(VSS),.VDD(VDD),.Y(g7150),.A(g6952));
  NOT NOT1_3933(.VSS(VSS),.VDD(VDD),.Y(I13035),.A(g6964));
  NOT NOT1_3934(.VSS(VSS),.VDD(VDD),.Y(g7151),.A(I13035));
  NOT NOT1_3935(.VSS(VSS),.VDD(VDD),.Y(I13039),.A(g6961));
  NOT NOT1_3936(.VSS(VSS),.VDD(VDD),.Y(g7155),.A(I13039));
  NOT NOT1_3937(.VSS(VSS),.VDD(VDD),.Y(I13042),.A(g6963));
  NOT NOT1_3938(.VSS(VSS),.VDD(VDD),.Y(g7156),.A(I13042));
  NOT NOT1_3939(.VSS(VSS),.VDD(VDD),.Y(I13045),.A(g6955));
  NOT NOT1_3940(.VSS(VSS),.VDD(VDD),.Y(g7157),.A(I13045));
  NOT NOT1_3941(.VSS(VSS),.VDD(VDD),.Y(I13048),.A(g6956));
  NOT NOT1_3942(.VSS(VSS),.VDD(VDD),.Y(g7158),.A(I13048));
  NOT NOT1_3943(.VSS(VSS),.VDD(VDD),.Y(I13051),.A(g6967));
  NOT NOT1_3944(.VSS(VSS),.VDD(VDD),.Y(g7159),.A(I13051));
  NOT NOT1_3945(.VSS(VSS),.VDD(VDD),.Y(I13054),.A(g6960));
  NOT NOT1_3946(.VSS(VSS),.VDD(VDD),.Y(g7160),.A(I13054));
  NOT NOT1_3947(.VSS(VSS),.VDD(VDD),.Y(I13057),.A(g6968));
  NOT NOT1_3948(.VSS(VSS),.VDD(VDD),.Y(g7161),.A(I13057));
  NOT NOT1_3949(.VSS(VSS),.VDD(VDD),.Y(I13060),.A(g6959));
  NOT NOT1_3950(.VSS(VSS),.VDD(VDD),.Y(g7162),.A(I13060));
  NOT NOT1_3951(.VSS(VSS),.VDD(VDD),.Y(I13063),.A(g6973));
  NOT NOT1_3952(.VSS(VSS),.VDD(VDD),.Y(g7163),.A(I13063));
  NOT NOT1_3953(.VSS(VSS),.VDD(VDD),.Y(I13066),.A(g6957));
  NOT NOT1_3954(.VSS(VSS),.VDD(VDD),.Y(g7164),.A(I13066));
  NOT NOT1_3955(.VSS(VSS),.VDD(VDD),.Y(I13072),.A(g6969));
  NOT NOT1_3956(.VSS(VSS),.VDD(VDD),.Y(g7168),.A(I13072));
  NOT NOT1_3957(.VSS(VSS),.VDD(VDD),.Y(I13075),.A(g6958));
  NOT NOT1_3958(.VSS(VSS),.VDD(VDD),.Y(g7169),.A(I13075));
  NOT NOT1_3959(.VSS(VSS),.VDD(VDD),.Y(g7171),.A(g7071));
  NOT NOT1_3960(.VSS(VSS),.VDD(VDD),.Y(g7172),.A(g7092));
  NOT NOT1_3961(.VSS(VSS),.VDD(VDD),.Y(g7173),.A(g6980));
  NOT NOT1_3962(.VSS(VSS),.VDD(VDD),.Y(g7174),.A(g7097));
  NOT NOT1_3963(.VSS(VSS),.VDD(VDD),.Y(I13084),.A(g7071));
  NOT NOT1_3964(.VSS(VSS),.VDD(VDD),.Y(g7176),.A(I13084));
  NOT NOT1_3965(.VSS(VSS),.VDD(VDD),.Y(I13088),.A(g7045));
  NOT NOT1_3966(.VSS(VSS),.VDD(VDD),.Y(g7178),.A(I13088));
  NOT NOT1_3967(.VSS(VSS),.VDD(VDD),.Y(I13092),.A(g7047));
  NOT NOT1_3968(.VSS(VSS),.VDD(VDD),.Y(g7180),.A(I13092));
  NOT NOT1_3969(.VSS(VSS),.VDD(VDD),.Y(I13099),.A(g7054));
  NOT NOT1_3970(.VSS(VSS),.VDD(VDD),.Y(g7185),.A(I13099));
  NOT NOT1_3971(.VSS(VSS),.VDD(VDD),.Y(I13103),.A(g7055));
  NOT NOT1_3972(.VSS(VSS),.VDD(VDD),.Y(g7187),.A(I13103));
  NOT NOT1_3973(.VSS(VSS),.VDD(VDD),.Y(I13106),.A(g7056));
  NOT NOT1_3974(.VSS(VSS),.VDD(VDD),.Y(g7188),.A(I13106));
  NOT NOT1_3975(.VSS(VSS),.VDD(VDD),.Y(I13109),.A(g7059));
  NOT NOT1_3976(.VSS(VSS),.VDD(VDD),.Y(g7189),.A(I13109));
  NOT NOT1_3977(.VSS(VSS),.VDD(VDD),.Y(I13112),.A(g7021));
  NOT NOT1_3978(.VSS(VSS),.VDD(VDD),.Y(g7190),.A(I13112));
  NOT NOT1_3979(.VSS(VSS),.VDD(VDD),.Y(I13118),.A(g7068));
  NOT NOT1_3980(.VSS(VSS),.VDD(VDD),.Y(g7194),.A(I13118));
  NOT NOT1_3981(.VSS(VSS),.VDD(VDD),.Y(I13122),.A(g7070));
  NOT NOT1_3982(.VSS(VSS),.VDD(VDD),.Y(g7196),.A(I13122));
  NOT NOT1_3983(.VSS(VSS),.VDD(VDD),.Y(I13126),.A(g6949));
  NOT NOT1_3984(.VSS(VSS),.VDD(VDD),.Y(g7198),.A(I13126));
  NOT NOT1_3985(.VSS(VSS),.VDD(VDD),.Y(I13131),.A(g6951));
  NOT NOT1_3986(.VSS(VSS),.VDD(VDD),.Y(g7205),.A(I13131));
  NOT NOT1_3987(.VSS(VSS),.VDD(VDD),.Y(I13134),.A(g7017));
  NOT NOT1_3988(.VSS(VSS),.VDD(VDD),.Y(g7206),.A(I13134));
  NOT NOT1_3989(.VSS(VSS),.VDD(VDD),.Y(I13137),.A(g7027));
  NOT NOT1_3990(.VSS(VSS),.VDD(VDD),.Y(g7207),.A(I13137));
  NOT NOT1_3991(.VSS(VSS),.VDD(VDD),.Y(I13140),.A(g6954));
  NOT NOT1_3992(.VSS(VSS),.VDD(VDD),.Y(g7208),.A(I13140));
  NOT NOT1_3993(.VSS(VSS),.VDD(VDD),.Y(I13144),.A(g7031));
  NOT NOT1_3994(.VSS(VSS),.VDD(VDD),.Y(g7210),.A(I13144));
  NOT NOT1_3995(.VSS(VSS),.VDD(VDD),.Y(I13147),.A(g7024));
  NOT NOT1_3996(.VSS(VSS),.VDD(VDD),.Y(g7211),.A(I13147));
  NOT NOT1_3997(.VSS(VSS),.VDD(VDD),.Y(I13152),.A(g6966));
  NOT NOT1_3998(.VSS(VSS),.VDD(VDD),.Y(g7216),.A(I13152));
  NOT NOT1_3999(.VSS(VSS),.VDD(VDD),.Y(I13157),.A(g6997));
  NOT NOT1_4000(.VSS(VSS),.VDD(VDD),.Y(g7221),.A(I13157));
  NOT NOT1_4001(.VSS(VSS),.VDD(VDD),.Y(I13161),.A(g7080));
  NOT NOT1_4002(.VSS(VSS),.VDD(VDD),.Y(g7223),.A(I13161));
  NOT NOT1_4003(.VSS(VSS),.VDD(VDD),.Y(I13164),.A(g7086));
  NOT NOT1_4004(.VSS(VSS),.VDD(VDD),.Y(g7224),.A(I13164));
  NOT NOT1_4005(.VSS(VSS),.VDD(VDD),.Y(g7225),.A(g6936));
  NOT NOT1_4006(.VSS(VSS),.VDD(VDD),.Y(g7226),.A(g6937));
  NOT NOT1_4007(.VSS(VSS),.VDD(VDD),.Y(g7229),.A(g6938));
  NOT NOT1_4008(.VSS(VSS),.VDD(VDD),.Y(I13173),.A(g7089));
  NOT NOT1_4009(.VSS(VSS),.VDD(VDD),.Y(g7231),.A(I13173));
  NOT NOT1_4010(.VSS(VSS),.VDD(VDD),.Y(g7233),.A(g6940));
  NOT NOT1_4011(.VSS(VSS),.VDD(VDD),.Y(g7236),.A(g6944));
  NOT NOT1_4012(.VSS(VSS),.VDD(VDD),.Y(g7239),.A(g6945));
  NOT NOT1_4013(.VSS(VSS),.VDD(VDD),.Y(I13185),.A(g7020));
  NOT NOT1_4014(.VSS(VSS),.VDD(VDD),.Y(g7241),.A(I13185));
  NOT NOT1_4015(.VSS(VSS),.VDD(VDD),.Y(I13189),.A(g7002));
  NOT NOT1_4016(.VSS(VSS),.VDD(VDD),.Y(g7243),.A(I13189));
  NOT NOT1_4017(.VSS(VSS),.VDD(VDD),.Y(I13193),.A(g7007));
  NOT NOT1_4018(.VSS(VSS),.VDD(VDD),.Y(g7245),.A(I13193));
  NOT NOT1_4019(.VSS(VSS),.VDD(VDD),.Y(I13196),.A(g7008));
  NOT NOT1_4020(.VSS(VSS),.VDD(VDD),.Y(g7246),.A(I13196));
  NOT NOT1_4021(.VSS(VSS),.VDD(VDD),.Y(I13199),.A(g7025));
  NOT NOT1_4022(.VSS(VSS),.VDD(VDD),.Y(g7247),.A(I13199));
  NOT NOT1_4023(.VSS(VSS),.VDD(VDD),.Y(I13203),.A(g7088));
  NOT NOT1_4024(.VSS(VSS),.VDD(VDD),.Y(g7251),.A(I13203));
  NOT NOT1_4025(.VSS(VSS),.VDD(VDD),.Y(g7253),.A(g7049));
  NOT NOT1_4026(.VSS(VSS),.VDD(VDD),.Y(I13209),.A(g6912));
  NOT NOT1_4027(.VSS(VSS),.VDD(VDD),.Y(g7255),.A(I13209));
  NOT NOT1_4028(.VSS(VSS),.VDD(VDD),.Y(g7256),.A(g7058));
  NOT NOT1_4029(.VSS(VSS),.VDD(VDD),.Y(g7259),.A(g7060));
  NOT NOT1_4030(.VSS(VSS),.VDD(VDD),.Y(g7260),.A(g7064));
  NOT NOT1_4031(.VSS(VSS),.VDD(VDD),.Y(I13225),.A(g7095));
  NOT NOT1_4032(.VSS(VSS),.VDD(VDD),.Y(g7261),.A(I13225));
  NOT NOT1_4033(.VSS(VSS),.VDD(VDD),.Y(I13228),.A(g6892));
  NOT NOT1_4034(.VSS(VSS),.VDD(VDD),.Y(g7262),.A(I13228));
  NOT NOT1_4035(.VSS(VSS),.VDD(VDD),.Y(I13231),.A(g6897));
  NOT NOT1_4036(.VSS(VSS),.VDD(VDD),.Y(g7263),.A(I13231));
  NOT NOT1_4037(.VSS(VSS),.VDD(VDD),.Y(I13234),.A(g6898));
  NOT NOT1_4038(.VSS(VSS),.VDD(VDD),.Y(g7264),.A(I13234));
  NOT NOT1_4039(.VSS(VSS),.VDD(VDD),.Y(g7265),.A(g7077));
  NOT NOT1_4040(.VSS(VSS),.VDD(VDD),.Y(I13238),.A(g6900));
  NOT NOT1_4041(.VSS(VSS),.VDD(VDD),.Y(g7266),.A(I13238));
  NOT NOT1_4042(.VSS(VSS),.VDD(VDD),.Y(I13241),.A(g7030));
  NOT NOT1_4043(.VSS(VSS),.VDD(VDD),.Y(g7267),.A(I13241));
  NOT NOT1_4044(.VSS(VSS),.VDD(VDD),.Y(I13244),.A(g7033));
  NOT NOT1_4045(.VSS(VSS),.VDD(VDD),.Y(g7268),.A(I13244));
  NOT NOT1_4046(.VSS(VSS),.VDD(VDD),.Y(I13247),.A(g6906));
  NOT NOT1_4047(.VSS(VSS),.VDD(VDD),.Y(g7269),.A(I13247));
  NOT NOT1_4048(.VSS(VSS),.VDD(VDD),.Y(I13250),.A(g7036));
  NOT NOT1_4049(.VSS(VSS),.VDD(VDD),.Y(g7270),.A(I13250));
  NOT NOT1_4050(.VSS(VSS),.VDD(VDD),.Y(I13255),.A(g7057));
  NOT NOT1_4051(.VSS(VSS),.VDD(VDD),.Y(g7273),.A(I13255));
  NOT NOT1_4052(.VSS(VSS),.VDD(VDD),.Y(I13258),.A(g6907));
  NOT NOT1_4053(.VSS(VSS),.VDD(VDD),.Y(g7274),.A(I13258));
  NOT NOT1_4054(.VSS(VSS),.VDD(VDD),.Y(I13261),.A(g7041));
  NOT NOT1_4055(.VSS(VSS),.VDD(VDD),.Y(g7275),.A(I13261));
  NOT NOT1_4056(.VSS(VSS),.VDD(VDD),.Y(I13264),.A(g7061));
  NOT NOT1_4057(.VSS(VSS),.VDD(VDD),.Y(g7276),.A(I13264));
  NOT NOT1_4058(.VSS(VSS),.VDD(VDD),.Y(I13267),.A(g6913));
  NOT NOT1_4059(.VSS(VSS),.VDD(VDD),.Y(g7277),.A(I13267));
  NOT NOT1_4060(.VSS(VSS),.VDD(VDD),.Y(I13271),.A(g7067));
  NOT NOT1_4061(.VSS(VSS),.VDD(VDD),.Y(g7279),.A(I13271));
  NOT NOT1_4062(.VSS(VSS),.VDD(VDD),.Y(I13274),.A(g6917));
  NOT NOT1_4063(.VSS(VSS),.VDD(VDD),.Y(g7280),.A(I13274));
  NOT NOT1_4064(.VSS(VSS),.VDD(VDD),.Y(I13277),.A(g7078));
  NOT NOT1_4065(.VSS(VSS),.VDD(VDD),.Y(g7281),.A(I13277));
  NOT NOT1_4066(.VSS(VSS),.VDD(VDD),.Y(I13281),.A(g7155));
  NOT NOT1_4067(.VSS(VSS),.VDD(VDD),.Y(g7283),.A(I13281));
  NOT NOT1_4068(.VSS(VSS),.VDD(VDD),.Y(I13284),.A(g7156));
  NOT NOT1_4069(.VSS(VSS),.VDD(VDD),.Y(g7284),.A(I13284));
  NOT NOT1_4070(.VSS(VSS),.VDD(VDD),.Y(I13287),.A(g7157));
  NOT NOT1_4071(.VSS(VSS),.VDD(VDD),.Y(g7285),.A(I13287));
  NOT NOT1_4072(.VSS(VSS),.VDD(VDD),.Y(I13290),.A(g7158));
  NOT NOT1_4073(.VSS(VSS),.VDD(VDD),.Y(g7286),.A(I13290));
  NOT NOT1_4074(.VSS(VSS),.VDD(VDD),.Y(I13293),.A(g7159));
  NOT NOT1_4075(.VSS(VSS),.VDD(VDD),.Y(g7287),.A(I13293));
  NOT NOT1_4076(.VSS(VSS),.VDD(VDD),.Y(I13296),.A(g7161));
  NOT NOT1_4077(.VSS(VSS),.VDD(VDD),.Y(g7288),.A(I13296));
  NOT NOT1_4078(.VSS(VSS),.VDD(VDD),.Y(I13299),.A(g7163));
  NOT NOT1_4079(.VSS(VSS),.VDD(VDD),.Y(g7289),.A(I13299));
  NOT NOT1_4080(.VSS(VSS),.VDD(VDD),.Y(I13302),.A(g7164));
  NOT NOT1_4081(.VSS(VSS),.VDD(VDD),.Y(g7290),.A(I13302));
  NOT NOT1_4082(.VSS(VSS),.VDD(VDD),.Y(I13305),.A(g7168));
  NOT NOT1_4083(.VSS(VSS),.VDD(VDD),.Y(g7291),.A(I13305));
  NOT NOT1_4084(.VSS(VSS),.VDD(VDD),.Y(I13308),.A(g7169));
  NOT NOT1_4085(.VSS(VSS),.VDD(VDD),.Y(g7292),.A(I13308));
  NOT NOT1_4086(.VSS(VSS),.VDD(VDD),.Y(I13311),.A(g7162));
  NOT NOT1_4087(.VSS(VSS),.VDD(VDD),.Y(g7293),.A(I13311));
  NOT NOT1_4088(.VSS(VSS),.VDD(VDD),.Y(I13314),.A(g7160));
  NOT NOT1_4089(.VSS(VSS),.VDD(VDD),.Y(g7294),.A(I13314));
  NOT NOT1_4090(.VSS(VSS),.VDD(VDD),.Y(I13317),.A(g7211));
  NOT NOT1_4091(.VSS(VSS),.VDD(VDD),.Y(g7295),.A(I13317));
  NOT NOT1_4092(.VSS(VSS),.VDD(VDD),.Y(I13320),.A(g7139));
  NOT NOT1_4093(.VSS(VSS),.VDD(VDD),.Y(g7296),.A(I13320));
  NOT NOT1_4094(.VSS(VSS),.VDD(VDD),.Y(I13323),.A(g7145));
  NOT NOT1_4095(.VSS(VSS),.VDD(VDD),.Y(g7297),.A(I13323));
  NOT NOT1_4096(.VSS(VSS),.VDD(VDD),.Y(I13326),.A(g7176));
  NOT NOT1_4097(.VSS(VSS),.VDD(VDD),.Y(g7298),.A(I13326));
  NOT NOT1_4098(.VSS(VSS),.VDD(VDD),.Y(I13329),.A(g7247));
  NOT NOT1_4099(.VSS(VSS),.VDD(VDD),.Y(g7299),.A(I13329));
  NOT NOT1_4100(.VSS(VSS),.VDD(VDD),.Y(I13332),.A(g7241));
  NOT NOT1_4101(.VSS(VSS),.VDD(VDD),.Y(g7300),.A(I13332));
  NOT NOT1_4102(.VSS(VSS),.VDD(VDD),.Y(I13335),.A(g7206));
  NOT NOT1_4103(.VSS(VSS),.VDD(VDD),.Y(g7301),.A(I13335));
  NOT NOT1_4104(.VSS(VSS),.VDD(VDD),.Y(I13338),.A(g7190));
  NOT NOT1_4105(.VSS(VSS),.VDD(VDD),.Y(g7302),.A(I13338));
  NOT NOT1_4106(.VSS(VSS),.VDD(VDD),.Y(I13341),.A(g7207));
  NOT NOT1_4107(.VSS(VSS),.VDD(VDD),.Y(g7303),.A(I13341));
  NOT NOT1_4108(.VSS(VSS),.VDD(VDD),.Y(I13344),.A(g7210));
  NOT NOT1_4109(.VSS(VSS),.VDD(VDD),.Y(g7304),.A(I13344));
  NOT NOT1_4110(.VSS(VSS),.VDD(VDD),.Y(I13347),.A(g7224));
  NOT NOT1_4111(.VSS(VSS),.VDD(VDD),.Y(g7305),.A(I13347));
  NOT NOT1_4112(.VSS(VSS),.VDD(VDD),.Y(I13350),.A(g7223));
  NOT NOT1_4113(.VSS(VSS),.VDD(VDD),.Y(g7306),.A(I13350));
  NOT NOT1_4114(.VSS(VSS),.VDD(VDD),.Y(I13353),.A(g7231));
  NOT NOT1_4115(.VSS(VSS),.VDD(VDD),.Y(g7307),.A(I13353));
  NOT NOT1_4116(.VSS(VSS),.VDD(VDD),.Y(I13356),.A(g7221));
  NOT NOT1_4117(.VSS(VSS),.VDD(VDD),.Y(g7308),.A(I13356));
  NOT NOT1_4118(.VSS(VSS),.VDD(VDD),.Y(I13359),.A(g7255));
  NOT NOT1_4119(.VSS(VSS),.VDD(VDD),.Y(g7309),.A(I13359));
  NOT NOT1_4120(.VSS(VSS),.VDD(VDD),.Y(I13362),.A(g7265));
  NOT NOT1_4121(.VSS(VSS),.VDD(VDD),.Y(g7310),.A(I13362));
  NOT NOT1_4122(.VSS(VSS),.VDD(VDD),.Y(I13365),.A(g7267));
  NOT NOT1_4123(.VSS(VSS),.VDD(VDD),.Y(g7311),.A(I13365));
  NOT NOT1_4124(.VSS(VSS),.VDD(VDD),.Y(I13369),.A(g7268));
  NOT NOT1_4125(.VSS(VSS),.VDD(VDD),.Y(g7313),.A(I13369));
  NOT NOT1_4126(.VSS(VSS),.VDD(VDD),.Y(I13373),.A(g7270));
  NOT NOT1_4127(.VSS(VSS),.VDD(VDD),.Y(g7315),.A(I13373));
  NOT NOT1_4128(.VSS(VSS),.VDD(VDD),.Y(I13383),.A(g7275));
  NOT NOT1_4129(.VSS(VSS),.VDD(VDD),.Y(g7317),.A(I13383));
  NOT NOT1_4130(.VSS(VSS),.VDD(VDD),.Y(g7319),.A(g7124));
  NOT NOT1_4131(.VSS(VSS),.VDD(VDD),.Y(I13388),.A(g7149));
  NOT NOT1_4132(.VSS(VSS),.VDD(VDD),.Y(g7320),.A(I13388));
  NOT NOT1_4133(.VSS(VSS),.VDD(VDD),.Y(I13403),.A(g7269));
  NOT NOT1_4134(.VSS(VSS),.VDD(VDD),.Y(g7327),.A(I13403));
  NOT NOT1_4135(.VSS(VSS),.VDD(VDD),.Y(I13407),.A(g7271));
  NOT NOT1_4136(.VSS(VSS),.VDD(VDD),.Y(g7329),.A(I13407));
  NOT NOT1_4137(.VSS(VSS),.VDD(VDD),.Y(I13410),.A(g7274));
  NOT NOT1_4138(.VSS(VSS),.VDD(VDD),.Y(g7330),.A(I13410));
  NOT NOT1_4139(.VSS(VSS),.VDD(VDD),.Y(I13413),.A(g7127));
  NOT NOT1_4140(.VSS(VSS),.VDD(VDD),.Y(g7331),.A(I13413));
  NOT NOT1_4141(.VSS(VSS),.VDD(VDD),.Y(I13416),.A(g7165));
  NOT NOT1_4142(.VSS(VSS),.VDD(VDD),.Y(g7332),.A(I13416));
  NOT NOT1_4143(.VSS(VSS),.VDD(VDD),.Y(I13419),.A(g7277));
  NOT NOT1_4144(.VSS(VSS),.VDD(VDD),.Y(g7333),.A(I13419));
  NOT NOT1_4145(.VSS(VSS),.VDD(VDD),.Y(I13422),.A(g7131));
  NOT NOT1_4146(.VSS(VSS),.VDD(VDD),.Y(g7334),.A(I13422));
  NOT NOT1_4147(.VSS(VSS),.VDD(VDD),.Y(I13425),.A(g7166));
  NOT NOT1_4148(.VSS(VSS),.VDD(VDD),.Y(g7335),.A(I13425));
  NOT NOT1_4149(.VSS(VSS),.VDD(VDD),.Y(I13428),.A(g7167));
  NOT NOT1_4150(.VSS(VSS),.VDD(VDD),.Y(g7336),.A(I13428));
  NOT NOT1_4151(.VSS(VSS),.VDD(VDD),.Y(I13432),.A(g7280));
  NOT NOT1_4152(.VSS(VSS),.VDD(VDD),.Y(g7338),.A(I13432));
  NOT NOT1_4153(.VSS(VSS),.VDD(VDD),.Y(I13435),.A(g7170));
  NOT NOT1_4154(.VSS(VSS),.VDD(VDD),.Y(g7339),.A(I13435));
  NOT NOT1_4155(.VSS(VSS),.VDD(VDD),.Y(I13438),.A(g7143));
  NOT NOT1_4156(.VSS(VSS),.VDD(VDD),.Y(g7340),.A(I13438));
  NOT NOT1_4157(.VSS(VSS),.VDD(VDD),.Y(I13441),.A(g7146));
  NOT NOT1_4158(.VSS(VSS),.VDD(VDD),.Y(g7341),.A(I13441));
  NOT NOT1_4159(.VSS(VSS),.VDD(VDD),.Y(I13444),.A(g7282));
  NOT NOT1_4160(.VSS(VSS),.VDD(VDD),.Y(g7342),.A(I13444));
  NOT NOT1_4161(.VSS(VSS),.VDD(VDD),.Y(I13447),.A(g7261));
  NOT NOT1_4162(.VSS(VSS),.VDD(VDD),.Y(g7343),.A(I13447));
  NOT NOT1_4163(.VSS(VSS),.VDD(VDD),.Y(g7344),.A(g7150));
  NOT NOT1_4164(.VSS(VSS),.VDD(VDD),.Y(I13451),.A(g7262));
  NOT NOT1_4165(.VSS(VSS),.VDD(VDD),.Y(g7345),.A(I13451));
  NOT NOT1_4166(.VSS(VSS),.VDD(VDD),.Y(I13454),.A(g7147));
  NOT NOT1_4167(.VSS(VSS),.VDD(VDD),.Y(g7346),.A(I13454));
  NOT NOT1_4168(.VSS(VSS),.VDD(VDD),.Y(I13457),.A(g7120));
  NOT NOT1_4169(.VSS(VSS),.VDD(VDD),.Y(g7347),.A(I13457));
  NOT NOT1_4170(.VSS(VSS),.VDD(VDD),.Y(I13460),.A(g7263));
  NOT NOT1_4171(.VSS(VSS),.VDD(VDD),.Y(g7348),.A(I13460));
  NOT NOT1_4172(.VSS(VSS),.VDD(VDD),.Y(I13463),.A(g7264));
  NOT NOT1_4173(.VSS(VSS),.VDD(VDD),.Y(g7349),.A(I13463));
  NOT NOT1_4174(.VSS(VSS),.VDD(VDD),.Y(I13466),.A(g7122));
  NOT NOT1_4175(.VSS(VSS),.VDD(VDD),.Y(g7350),.A(I13466));
  NOT NOT1_4176(.VSS(VSS),.VDD(VDD),.Y(I13469),.A(g7123));
  NOT NOT1_4177(.VSS(VSS),.VDD(VDD),.Y(g7351),.A(I13469));
  NOT NOT1_4178(.VSS(VSS),.VDD(VDD),.Y(I13472),.A(g7266));
  NOT NOT1_4179(.VSS(VSS),.VDD(VDD),.Y(g7352),.A(I13472));
  NOT NOT1_4180(.VSS(VSS),.VDD(VDD),.Y(I13475),.A(g7125));
  NOT NOT1_4181(.VSS(VSS),.VDD(VDD),.Y(g7353),.A(I13475));
  NOT NOT1_4182(.VSS(VSS),.VDD(VDD),.Y(I13478),.A(g7126));
  NOT NOT1_4183(.VSS(VSS),.VDD(VDD),.Y(g7354),.A(I13478));
  NOT NOT1_4184(.VSS(VSS),.VDD(VDD),.Y(I13481),.A(g7254));
  NOT NOT1_4185(.VSS(VSS),.VDD(VDD),.Y(g7355),.A(I13481));
  NOT NOT1_4186(.VSS(VSS),.VDD(VDD),.Y(I13484),.A(g7128));
  NOT NOT1_4187(.VSS(VSS),.VDD(VDD),.Y(g7356),.A(I13484));
  NOT NOT1_4188(.VSS(VSS),.VDD(VDD),.Y(I13487),.A(g7129));
  NOT NOT1_4189(.VSS(VSS),.VDD(VDD),.Y(g7357),.A(I13487));
  NOT NOT1_4190(.VSS(VSS),.VDD(VDD),.Y(I13490),.A(g7130));
  NOT NOT1_4191(.VSS(VSS),.VDD(VDD),.Y(g7358),.A(I13490));
  NOT NOT1_4192(.VSS(VSS),.VDD(VDD),.Y(I13493),.A(g7132));
  NOT NOT1_4193(.VSS(VSS),.VDD(VDD),.Y(g7359),.A(I13493));
  NOT NOT1_4194(.VSS(VSS),.VDD(VDD),.Y(I13496),.A(g7133));
  NOT NOT1_4195(.VSS(VSS),.VDD(VDD),.Y(g7360),.A(I13496));
  NOT NOT1_4196(.VSS(VSS),.VDD(VDD),.Y(I13499),.A(g7134));
  NOT NOT1_4197(.VSS(VSS),.VDD(VDD),.Y(g7361),.A(I13499));
  NOT NOT1_4198(.VSS(VSS),.VDD(VDD),.Y(I13502),.A(g7135));
  NOT NOT1_4199(.VSS(VSS),.VDD(VDD),.Y(g7362),.A(I13502));
  NOT NOT1_4200(.VSS(VSS),.VDD(VDD),.Y(I13506),.A(g7148));
  NOT NOT1_4201(.VSS(VSS),.VDD(VDD),.Y(g7364),.A(I13506));
  NOT NOT1_4202(.VSS(VSS),.VDD(VDD),.Y(I13509),.A(g7137));
  NOT NOT1_4203(.VSS(VSS),.VDD(VDD),.Y(g7365),.A(I13509));
  NOT NOT1_4204(.VSS(VSS),.VDD(VDD),.Y(I13512),.A(g7138));
  NOT NOT1_4205(.VSS(VSS),.VDD(VDD),.Y(g7366),.A(I13512));
  NOT NOT1_4206(.VSS(VSS),.VDD(VDD),.Y(I13515),.A(g7152));
  NOT NOT1_4207(.VSS(VSS),.VDD(VDD),.Y(g7367),.A(I13515));
  NOT NOT1_4208(.VSS(VSS),.VDD(VDD),.Y(I13518),.A(g7141));
  NOT NOT1_4209(.VSS(VSS),.VDD(VDD),.Y(g7405),.A(I13518));
  NOT NOT1_4210(.VSS(VSS),.VDD(VDD),.Y(g7411),.A(g7202));
  NOT NOT1_4211(.VSS(VSS),.VDD(VDD),.Y(I13524),.A(g7151));
  NOT NOT1_4212(.VSS(VSS),.VDD(VDD),.Y(g7413),.A(I13524));
  NOT NOT1_4213(.VSS(VSS),.VDD(VDD),.Y(I13527),.A(g7217));
  NOT NOT1_4214(.VSS(VSS),.VDD(VDD),.Y(g7414),.A(I13527));
  NOT NOT1_4215(.VSS(VSS),.VDD(VDD),.Y(I13533),.A(g7220));
  NOT NOT1_4216(.VSS(VSS),.VDD(VDD),.Y(g7418),.A(I13533));
  NOT NOT1_4217(.VSS(VSS),.VDD(VDD),.Y(I13537),.A(g7152));
  NOT NOT1_4218(.VSS(VSS),.VDD(VDD),.Y(g7420),.A(I13537));
  NOT NOT1_4219(.VSS(VSS),.VDD(VDD),.Y(I13541),.A(g7209));
  NOT NOT1_4220(.VSS(VSS),.VDD(VDD),.Y(g7422),.A(I13541));
  NOT NOT1_4221(.VSS(VSS),.VDD(VDD),.Y(I13544),.A(g1167));
  NOT NOT1_4222(.VSS(VSS),.VDD(VDD),.Y(g7423),.A(I13544));
  NOT NOT1_4223(.VSS(VSS),.VDD(VDD),.Y(I13547),.A(g1170));
  NOT NOT1_4224(.VSS(VSS),.VDD(VDD),.Y(g7424),.A(I13547));
  NOT NOT1_4225(.VSS(VSS),.VDD(VDD),.Y(I13550),.A(g1173));
  NOT NOT1_4226(.VSS(VSS),.VDD(VDD),.Y(g7425),.A(I13550));
  NOT NOT1_4227(.VSS(VSS),.VDD(VDD),.Y(I13559),.A(g7177));
  NOT NOT1_4228(.VSS(VSS),.VDD(VDD),.Y(g7432),.A(I13559));
  NOT NOT1_4229(.VSS(VSS),.VDD(VDD),.Y(I13562),.A(g7179));
  NOT NOT1_4230(.VSS(VSS),.VDD(VDD),.Y(g7433),.A(I13562));
  NOT NOT1_4231(.VSS(VSS),.VDD(VDD),.Y(I13565),.A(g7181));
  NOT NOT1_4232(.VSS(VSS),.VDD(VDD),.Y(g7434),.A(I13565));
  NOT NOT1_4233(.VSS(VSS),.VDD(VDD),.Y(I13570),.A(g7198));
  NOT NOT1_4234(.VSS(VSS),.VDD(VDD),.Y(g7437),.A(I13570));
  NOT NOT1_4235(.VSS(VSS),.VDD(VDD),.Y(I13574),.A(g7205));
  NOT NOT1_4236(.VSS(VSS),.VDD(VDD),.Y(g7439),.A(I13574));
  NOT NOT1_4237(.VSS(VSS),.VDD(VDD),.Y(I13577),.A(g7186));
  NOT NOT1_4238(.VSS(VSS),.VDD(VDD),.Y(g7440),.A(I13577));
  NOT NOT1_4239(.VSS(VSS),.VDD(VDD),.Y(I13580),.A(g7208));
  NOT NOT1_4240(.VSS(VSS),.VDD(VDD),.Y(g7441),.A(I13580));
  NOT NOT1_4241(.VSS(VSS),.VDD(VDD),.Y(I13583),.A(g7252));
  NOT NOT1_4242(.VSS(VSS),.VDD(VDD),.Y(g7442),.A(I13583));
  NOT NOT1_4243(.VSS(VSS),.VDD(VDD),.Y(I13595),.A(g7216));
  NOT NOT1_4244(.VSS(VSS),.VDD(VDD),.Y(g7446),.A(I13595));
  NOT NOT1_4245(.VSS(VSS),.VDD(VDD),.Y(I13605),.A(g7197));
  NOT NOT1_4246(.VSS(VSS),.VDD(VDD),.Y(g7448),.A(I13605));
  NOT NOT1_4247(.VSS(VSS),.VDD(VDD),.Y(I13610),.A(g7227));
  NOT NOT1_4248(.VSS(VSS),.VDD(VDD),.Y(g7454),.A(I13610));
  NOT NOT1_4249(.VSS(VSS),.VDD(VDD),.Y(I13613),.A(g7273));
  NOT NOT1_4250(.VSS(VSS),.VDD(VDD),.Y(g7455),.A(I13613));
  NOT NOT1_4251(.VSS(VSS),.VDD(VDD),.Y(g7456),.A(g7174));
  NOT NOT1_4252(.VSS(VSS),.VDD(VDD),.Y(I13617),.A(g7276));
  NOT NOT1_4253(.VSS(VSS),.VDD(VDD),.Y(g7459),.A(I13617));
  NOT NOT1_4254(.VSS(VSS),.VDD(VDD),.Y(g7460),.A(g7172));
  NOT NOT1_4255(.VSS(VSS),.VDD(VDD),.Y(g7463),.A(g7239));
  NOT NOT1_4256(.VSS(VSS),.VDD(VDD),.Y(I13622),.A(g7279));
  NOT NOT1_4257(.VSS(VSS),.VDD(VDD),.Y(g7466),.A(I13622));
  NOT NOT1_4258(.VSS(VSS),.VDD(VDD),.Y(g7467),.A(g7236));
  NOT NOT1_4259(.VSS(VSS),.VDD(VDD),.Y(g7470),.A(g7253));
  NOT NOT1_4260(.VSS(VSS),.VDD(VDD),.Y(g7471),.A(g7233));
  NOT NOT1_4261(.VSS(VSS),.VDD(VDD),.Y(I13628),.A(g7248));
  NOT NOT1_4262(.VSS(VSS),.VDD(VDD),.Y(g7474),.A(I13628));
  NOT NOT1_4263(.VSS(VSS),.VDD(VDD),.Y(I13631),.A(g7248));
  NOT NOT1_4264(.VSS(VSS),.VDD(VDD),.Y(g7475),.A(I13631));
  NOT NOT1_4265(.VSS(VSS),.VDD(VDD),.Y(g7476),.A(g7229));
  NOT NOT1_4266(.VSS(VSS),.VDD(VDD),.Y(I13635),.A(g7243));
  NOT NOT1_4267(.VSS(VSS),.VDD(VDD),.Y(g7479),.A(I13635));
  NOT NOT1_4268(.VSS(VSS),.VDD(VDD),.Y(g7483),.A(g7226));
  NOT NOT1_4269(.VSS(VSS),.VDD(VDD),.Y(I13646),.A(g7245));
  NOT NOT1_4270(.VSS(VSS),.VDD(VDD),.Y(g7486),.A(I13646));
  NOT NOT1_4271(.VSS(VSS),.VDD(VDD),.Y(I13649),.A(g7281));
  NOT NOT1_4272(.VSS(VSS),.VDD(VDD),.Y(g7487),.A(I13649));
  NOT NOT1_4273(.VSS(VSS),.VDD(VDD),.Y(g7488),.A(g7225));
  NOT NOT1_4274(.VSS(VSS),.VDD(VDD),.Y(I13653),.A(g7246));
  NOT NOT1_4275(.VSS(VSS),.VDD(VDD),.Y(g7491),.A(I13653));
  NOT NOT1_4276(.VSS(VSS),.VDD(VDD),.Y(I13656),.A(g7228));
  NOT NOT1_4277(.VSS(VSS),.VDD(VDD),.Y(g7492),.A(I13656));
  NOT NOT1_4278(.VSS(VSS),.VDD(VDD),.Y(I13659),.A(g7232));
  NOT NOT1_4279(.VSS(VSS),.VDD(VDD),.Y(g7493),.A(I13659));
  NOT NOT1_4280(.VSS(VSS),.VDD(VDD),.Y(g7494),.A(g7260));
  NOT NOT1_4281(.VSS(VSS),.VDD(VDD),.Y(I13663),.A(g7235));
  NOT NOT1_4282(.VSS(VSS),.VDD(VDD),.Y(g7495),.A(I13663));
  NOT NOT1_4283(.VSS(VSS),.VDD(VDD),.Y(I13666),.A(g7238));
  NOT NOT1_4284(.VSS(VSS),.VDD(VDD),.Y(g7496),.A(I13666));
  NOT NOT1_4285(.VSS(VSS),.VDD(VDD),.Y(I13669),.A(g7240));
  NOT NOT1_4286(.VSS(VSS),.VDD(VDD),.Y(g7497),.A(I13669));
  NOT NOT1_4287(.VSS(VSS),.VDD(VDD),.Y(I13672),.A(g7242));
  NOT NOT1_4288(.VSS(VSS),.VDD(VDD),.Y(g7498),.A(I13672));
  NOT NOT1_4289(.VSS(VSS),.VDD(VDD),.Y(g7499),.A(g7258));
  NOT NOT1_4290(.VSS(VSS),.VDD(VDD),.Y(I13676),.A(g7256));
  NOT NOT1_4291(.VSS(VSS),.VDD(VDD),.Y(g7500),.A(I13676));
  NOT NOT1_4292(.VSS(VSS),.VDD(VDD),.Y(I13679),.A(g7259));
  NOT NOT1_4293(.VSS(VSS),.VDD(VDD),.Y(g7501),.A(I13679));
  NOT NOT1_4294(.VSS(VSS),.VDD(VDD),.Y(I13682),.A(g7251));
  NOT NOT1_4295(.VSS(VSS),.VDD(VDD),.Y(g7502),.A(I13682));
  NOT NOT1_4296(.VSS(VSS),.VDD(VDD),.Y(I13692),.A(g7343));
  NOT NOT1_4297(.VSS(VSS),.VDD(VDD),.Y(g7504),.A(I13692));
  NOT NOT1_4298(.VSS(VSS),.VDD(VDD),.Y(I13695),.A(g7345));
  NOT NOT1_4299(.VSS(VSS),.VDD(VDD),.Y(g7505),.A(I13695));
  NOT NOT1_4300(.VSS(VSS),.VDD(VDD),.Y(I13698),.A(g7348));
  NOT NOT1_4301(.VSS(VSS),.VDD(VDD),.Y(g7506),.A(I13698));
  NOT NOT1_4302(.VSS(VSS),.VDD(VDD),.Y(I13701),.A(g7349));
  NOT NOT1_4303(.VSS(VSS),.VDD(VDD),.Y(g7507),.A(I13701));
  NOT NOT1_4304(.VSS(VSS),.VDD(VDD),.Y(I13704),.A(g7352));
  NOT NOT1_4305(.VSS(VSS),.VDD(VDD),.Y(g7508),.A(I13704));
  NOT NOT1_4306(.VSS(VSS),.VDD(VDD),.Y(I13707),.A(g7420));
  NOT NOT1_4307(.VSS(VSS),.VDD(VDD),.Y(g7509),.A(I13707));
  NOT NOT1_4308(.VSS(VSS),.VDD(VDD),.Y(I13710),.A(g7340));
  NOT NOT1_4309(.VSS(VSS),.VDD(VDD),.Y(g7510),.A(I13710));
  NOT NOT1_4310(.VSS(VSS),.VDD(VDD),.Y(I13713),.A(g7341));
  NOT NOT1_4311(.VSS(VSS),.VDD(VDD),.Y(g7511),.A(I13713));
  NOT NOT1_4312(.VSS(VSS),.VDD(VDD),.Y(I13716),.A(g7331));
  NOT NOT1_4313(.VSS(VSS),.VDD(VDD),.Y(g7512),.A(I13716));
  NOT NOT1_4314(.VSS(VSS),.VDD(VDD),.Y(I13719),.A(g7334));
  NOT NOT1_4315(.VSS(VSS),.VDD(VDD),.Y(g7513),.A(I13719));
  NOT NOT1_4316(.VSS(VSS),.VDD(VDD),.Y(I13722),.A(g7442));
  NOT NOT1_4317(.VSS(VSS),.VDD(VDD),.Y(g7514),.A(I13722));
  NOT NOT1_4318(.VSS(VSS),.VDD(VDD),.Y(I13725),.A(g7437));
  NOT NOT1_4319(.VSS(VSS),.VDD(VDD),.Y(g7515),.A(I13725));
  NOT NOT1_4320(.VSS(VSS),.VDD(VDD),.Y(I13728),.A(g7439));
  NOT NOT1_4321(.VSS(VSS),.VDD(VDD),.Y(g7516),.A(I13728));
  NOT NOT1_4322(.VSS(VSS),.VDD(VDD),.Y(I13731),.A(g7441));
  NOT NOT1_4323(.VSS(VSS),.VDD(VDD),.Y(g7517),.A(I13731));
  NOT NOT1_4324(.VSS(VSS),.VDD(VDD),.Y(I13734),.A(g7422));
  NOT NOT1_4325(.VSS(VSS),.VDD(VDD),.Y(g7518),.A(I13734));
  NOT NOT1_4326(.VSS(VSS),.VDD(VDD),.Y(I13737),.A(g7446));
  NOT NOT1_4327(.VSS(VSS),.VDD(VDD),.Y(g7519),.A(I13737));
  NOT NOT1_4328(.VSS(VSS),.VDD(VDD),.Y(I13740),.A(g7364));
  NOT NOT1_4329(.VSS(VSS),.VDD(VDD),.Y(g7520),.A(I13740));
  NOT NOT1_4330(.VSS(VSS),.VDD(VDD),.Y(I13743),.A(g7454));
  NOT NOT1_4331(.VSS(VSS),.VDD(VDD),.Y(g7521),.A(I13743));
  NOT NOT1_4332(.VSS(VSS),.VDD(VDD),.Y(I13746),.A(g7311));
  NOT NOT1_4333(.VSS(VSS),.VDD(VDD),.Y(g7522),.A(I13746));
  NOT NOT1_4334(.VSS(VSS),.VDD(VDD),.Y(I13749),.A(g7313));
  NOT NOT1_4335(.VSS(VSS),.VDD(VDD),.Y(g7523),.A(I13749));
  NOT NOT1_4336(.VSS(VSS),.VDD(VDD),.Y(I13752),.A(g7315));
  NOT NOT1_4337(.VSS(VSS),.VDD(VDD),.Y(g7524),.A(I13752));
  NOT NOT1_4338(.VSS(VSS),.VDD(VDD),.Y(I13755),.A(g7317));
  NOT NOT1_4339(.VSS(VSS),.VDD(VDD),.Y(g7525),.A(I13755));
  NOT NOT1_4340(.VSS(VSS),.VDD(VDD),.Y(I13758),.A(g7414));
  NOT NOT1_4341(.VSS(VSS),.VDD(VDD),.Y(g7526),.A(I13758));
  NOT NOT1_4342(.VSS(VSS),.VDD(VDD),.Y(I13761),.A(g7418));
  NOT NOT1_4343(.VSS(VSS),.VDD(VDD),.Y(g7527),.A(I13761));
  NOT NOT1_4344(.VSS(VSS),.VDD(VDD),.Y(I13764),.A(g7479));
  NOT NOT1_4345(.VSS(VSS),.VDD(VDD),.Y(g7528),.A(I13764));
  NOT NOT1_4346(.VSS(VSS),.VDD(VDD),.Y(I13767),.A(g7486));
  NOT NOT1_4347(.VSS(VSS),.VDD(VDD),.Y(g7529),.A(I13767));
  NOT NOT1_4348(.VSS(VSS),.VDD(VDD),.Y(I13770),.A(g7491));
  NOT NOT1_4349(.VSS(VSS),.VDD(VDD),.Y(g7530),.A(I13770));
  NOT NOT1_4350(.VSS(VSS),.VDD(VDD),.Y(I13773),.A(g7496));
  NOT NOT1_4351(.VSS(VSS),.VDD(VDD),.Y(g7531),.A(I13773));
  NOT NOT1_4352(.VSS(VSS),.VDD(VDD),.Y(I13776),.A(g7497));
  NOT NOT1_4353(.VSS(VSS),.VDD(VDD),.Y(g7532),.A(I13776));
  NOT NOT1_4354(.VSS(VSS),.VDD(VDD),.Y(I13779),.A(g7406));
  NOT NOT1_4355(.VSS(VSS),.VDD(VDD),.Y(g7533),.A(I13779));
  NOT NOT1_4356(.VSS(VSS),.VDD(VDD),.Y(I13782),.A(g7498));
  NOT NOT1_4357(.VSS(VSS),.VDD(VDD),.Y(g7534),.A(I13782));
  NOT NOT1_4358(.VSS(VSS),.VDD(VDD),.Y(I13794),.A(g7346));
  NOT NOT1_4359(.VSS(VSS),.VDD(VDD),.Y(g7538),.A(I13794));
  NOT NOT1_4360(.VSS(VSS),.VDD(VDD),.Y(I13797),.A(g7502));
  NOT NOT1_4361(.VSS(VSS),.VDD(VDD),.Y(g7539),.A(I13797));
  NOT NOT1_4362(.VSS(VSS),.VDD(VDD),.Y(I13807),.A(g7320));
  NOT NOT1_4363(.VSS(VSS),.VDD(VDD),.Y(g7541),.A(I13807));
  NOT NOT1_4364(.VSS(VSS),.VDD(VDD),.Y(I13810),.A(g7312));
  NOT NOT1_4365(.VSS(VSS),.VDD(VDD),.Y(g7542),.A(I13810));
  NOT NOT1_4366(.VSS(VSS),.VDD(VDD),.Y(I13813),.A(g7314));
  NOT NOT1_4367(.VSS(VSS),.VDD(VDD),.Y(g7543),.A(I13813));
  NOT NOT1_4368(.VSS(VSS),.VDD(VDD),.Y(I13816),.A(g7455));
  NOT NOT1_4369(.VSS(VSS),.VDD(VDD),.Y(g7544),.A(I13816));
  NOT NOT1_4370(.VSS(VSS),.VDD(VDD),.Y(I13819),.A(g7426));
  NOT NOT1_4371(.VSS(VSS),.VDD(VDD),.Y(g7545),.A(I13819));
  NOT NOT1_4372(.VSS(VSS),.VDD(VDD),.Y(I13822),.A(g7459));
  NOT NOT1_4373(.VSS(VSS),.VDD(VDD),.Y(g7546),.A(I13822));
  NOT NOT1_4374(.VSS(VSS),.VDD(VDD),.Y(I13825),.A(g7318));
  NOT NOT1_4375(.VSS(VSS),.VDD(VDD),.Y(g7547),.A(I13825));
  NOT NOT1_4376(.VSS(VSS),.VDD(VDD),.Y(I13828),.A(g7321));
  NOT NOT1_4377(.VSS(VSS),.VDD(VDD),.Y(g7548),.A(I13828));
  NOT NOT1_4378(.VSS(VSS),.VDD(VDD),.Y(I13831),.A(g7322));
  NOT NOT1_4379(.VSS(VSS),.VDD(VDD),.Y(g7549),.A(I13831));
  NOT NOT1_4380(.VSS(VSS),.VDD(VDD),.Y(I13834),.A(g7466));
  NOT NOT1_4381(.VSS(VSS),.VDD(VDD),.Y(g7550),.A(I13834));
  NOT NOT1_4382(.VSS(VSS),.VDD(VDD),.Y(I13837),.A(g7324));
  NOT NOT1_4383(.VSS(VSS),.VDD(VDD),.Y(g7551),.A(I13837));
  NOT NOT1_4384(.VSS(VSS),.VDD(VDD),.Y(I13843),.A(g7326));
  NOT NOT1_4385(.VSS(VSS),.VDD(VDD),.Y(g7555),.A(I13843));
  NOT NOT1_4386(.VSS(VSS),.VDD(VDD),.Y(I13846),.A(g7487));
  NOT NOT1_4387(.VSS(VSS),.VDD(VDD),.Y(g7556),.A(I13846));
  NOT NOT1_4388(.VSS(VSS),.VDD(VDD),.Y(I13850),.A(g7328));
  NOT NOT1_4389(.VSS(VSS),.VDD(VDD),.Y(g7558),.A(I13850));
  NOT NOT1_4390(.VSS(VSS),.VDD(VDD),.Y(I13854),.A(g7327));
  NOT NOT1_4391(.VSS(VSS),.VDD(VDD),.Y(g7560),.A(I13854));
  NOT NOT1_4392(.VSS(VSS),.VDD(VDD),.Y(I13858),.A(g7329));
  NOT NOT1_4393(.VSS(VSS),.VDD(VDD),.Y(g7562),.A(I13858));
  NOT NOT1_4394(.VSS(VSS),.VDD(VDD),.Y(I13861),.A(g7330));
  NOT NOT1_4395(.VSS(VSS),.VDD(VDD),.Y(g7563),.A(I13861));
  NOT NOT1_4396(.VSS(VSS),.VDD(VDD),.Y(I13865),.A(g7333));
  NOT NOT1_4397(.VSS(VSS),.VDD(VDD),.Y(g7565),.A(I13865));
  NOT NOT1_4398(.VSS(VSS),.VDD(VDD),.Y(I13869),.A(g7338));
  NOT NOT1_4399(.VSS(VSS),.VDD(VDD),.Y(g7574),.A(I13869));
  NOT NOT1_4400(.VSS(VSS),.VDD(VDD),.Y(I13873),.A(g7342));
  NOT NOT1_4401(.VSS(VSS),.VDD(VDD),.Y(g7576),.A(I13873));
  NOT NOT1_4402(.VSS(VSS),.VDD(VDD),.Y(I13876),.A(g7347));
  NOT NOT1_4403(.VSS(VSS),.VDD(VDD),.Y(g7577),.A(I13876));
  NOT NOT1_4404(.VSS(VSS),.VDD(VDD),.Y(I13879),.A(g7332));
  NOT NOT1_4405(.VSS(VSS),.VDD(VDD),.Y(g7578),.A(I13879));
  NOT NOT1_4406(.VSS(VSS),.VDD(VDD),.Y(I13882),.A(g7350));
  NOT NOT1_4407(.VSS(VSS),.VDD(VDD),.Y(g7579),.A(I13882));
  NOT NOT1_4408(.VSS(VSS),.VDD(VDD),.Y(I13885),.A(g7351));
  NOT NOT1_4409(.VSS(VSS),.VDD(VDD),.Y(g7580),.A(I13885));
  NOT NOT1_4410(.VSS(VSS),.VDD(VDD),.Y(I13888),.A(g7335));
  NOT NOT1_4411(.VSS(VSS),.VDD(VDD),.Y(g7581),.A(I13888));
  NOT NOT1_4412(.VSS(VSS),.VDD(VDD),.Y(I13891),.A(g7336));
  NOT NOT1_4413(.VSS(VSS),.VDD(VDD),.Y(g7582),.A(I13891));
  NOT NOT1_4414(.VSS(VSS),.VDD(VDD),.Y(I13894),.A(g7353));
  NOT NOT1_4415(.VSS(VSS),.VDD(VDD),.Y(g7583),.A(I13894));
  NOT NOT1_4416(.VSS(VSS),.VDD(VDD),.Y(I13897),.A(g7354));
  NOT NOT1_4417(.VSS(VSS),.VDD(VDD),.Y(g7584),.A(I13897));
  NOT NOT1_4418(.VSS(VSS),.VDD(VDD),.Y(I13900),.A(g7356));
  NOT NOT1_4419(.VSS(VSS),.VDD(VDD),.Y(g7585),.A(I13900));
  NOT NOT1_4420(.VSS(VSS),.VDD(VDD),.Y(I13903),.A(g7357));
  NOT NOT1_4421(.VSS(VSS),.VDD(VDD),.Y(g7586),.A(I13903));
  NOT NOT1_4422(.VSS(VSS),.VDD(VDD),.Y(I13906),.A(g7358));
  NOT NOT1_4423(.VSS(VSS),.VDD(VDD),.Y(g7587),.A(I13906));
  NOT NOT1_4424(.VSS(VSS),.VDD(VDD),.Y(I13909),.A(g7339));
  NOT NOT1_4425(.VSS(VSS),.VDD(VDD),.Y(g7588),.A(I13909));
  NOT NOT1_4426(.VSS(VSS),.VDD(VDD),.Y(I13912),.A(g7359));
  NOT NOT1_4427(.VSS(VSS),.VDD(VDD),.Y(g7589),.A(I13912));
  NOT NOT1_4428(.VSS(VSS),.VDD(VDD),.Y(I13915),.A(g7360));
  NOT NOT1_4429(.VSS(VSS),.VDD(VDD),.Y(g7590),.A(I13915));
  NOT NOT1_4430(.VSS(VSS),.VDD(VDD),.Y(I13918),.A(g7361));
  NOT NOT1_4431(.VSS(VSS),.VDD(VDD),.Y(g7591),.A(I13918));
  NOT NOT1_4432(.VSS(VSS),.VDD(VDD),.Y(I13921),.A(g7362));
  NOT NOT1_4433(.VSS(VSS),.VDD(VDD),.Y(g7592),.A(I13921));
  NOT NOT1_4434(.VSS(VSS),.VDD(VDD),.Y(I13924),.A(g7365));
  NOT NOT1_4435(.VSS(VSS),.VDD(VDD),.Y(g7593),.A(I13924));
  NOT NOT1_4436(.VSS(VSS),.VDD(VDD),.Y(I13927),.A(g7366));
  NOT NOT1_4437(.VSS(VSS),.VDD(VDD),.Y(g7594),.A(I13927));
  NOT NOT1_4438(.VSS(VSS),.VDD(VDD),.Y(I13930),.A(g7405));
  NOT NOT1_4439(.VSS(VSS),.VDD(VDD),.Y(g7595),.A(I13930));
  NOT NOT1_4440(.VSS(VSS),.VDD(VDD),.Y(g7599),.A(g7450));
  NOT NOT1_4441(.VSS(VSS),.VDD(VDD),.Y(g7601),.A(g7450));
  NOT NOT1_4442(.VSS(VSS),.VDD(VDD),.Y(I13940),.A(g7355));
  NOT NOT1_4443(.VSS(VSS),.VDD(VDD),.Y(g7603),.A(I13940));
  NOT NOT1_4444(.VSS(VSS),.VDD(VDD),.Y(g7610),.A(g7450));
  NOT NOT1_4445(.VSS(VSS),.VDD(VDD),.Y(I13956),.A(g7499));
  NOT NOT1_4446(.VSS(VSS),.VDD(VDD),.Y(g7627),.A(I13956));
  NOT NOT1_4447(.VSS(VSS),.VDD(VDD),.Y(I13962),.A(g7413));
  NOT NOT1_4448(.VSS(VSS),.VDD(VDD),.Y(g7633),.A(I13962));
  NOT NOT1_4449(.VSS(VSS),.VDD(VDD),.Y(I13979),.A(g7415));
  NOT NOT1_4450(.VSS(VSS),.VDD(VDD),.Y(g7686),.A(I13979));
  NOT NOT1_4451(.VSS(VSS),.VDD(VDD),.Y(g7688),.A(g7406));
  NOT NOT1_4452(.VSS(VSS),.VDD(VDD),.Y(I13997),.A(g7432));
  NOT NOT1_4453(.VSS(VSS),.VDD(VDD),.Y(g7702),.A(I13997));
  NOT NOT1_4454(.VSS(VSS),.VDD(VDD),.Y(I14001),.A(g7433));
  NOT NOT1_4455(.VSS(VSS),.VDD(VDD),.Y(g7704),.A(I14001));
  NOT NOT1_4456(.VSS(VSS),.VDD(VDD),.Y(I14005),.A(g7434));
  NOT NOT1_4457(.VSS(VSS),.VDD(VDD),.Y(g7708),.A(I14005));
  NOT NOT1_4458(.VSS(VSS),.VDD(VDD),.Y(I14009),.A(g7436));
  NOT NOT1_4459(.VSS(VSS),.VDD(VDD),.Y(g7710),.A(I14009));
  NOT NOT1_4460(.VSS(VSS),.VDD(VDD),.Y(I14012),.A(g7438));
  NOT NOT1_4461(.VSS(VSS),.VDD(VDD),.Y(g7711),.A(I14012));
  NOT NOT1_4462(.VSS(VSS),.VDD(VDD),.Y(I14015),.A(g7440));
  NOT NOT1_4463(.VSS(VSS),.VDD(VDD),.Y(g7712),.A(I14015));
  NOT NOT1_4464(.VSS(VSS),.VDD(VDD),.Y(I14019),.A(g7480));
  NOT NOT1_4465(.VSS(VSS),.VDD(VDD),.Y(g7714),.A(I14019));
  NOT NOT1_4466(.VSS(VSS),.VDD(VDD),.Y(I14022),.A(g7443));
  NOT NOT1_4467(.VSS(VSS),.VDD(VDD),.Y(g7715),.A(I14022));
  NOT NOT1_4468(.VSS(VSS),.VDD(VDD),.Y(I14025),.A(g7500));
  NOT NOT1_4469(.VSS(VSS),.VDD(VDD),.Y(g7716),.A(I14025));
  NOT NOT1_4470(.VSS(VSS),.VDD(VDD),.Y(I14028),.A(g7501));
  NOT NOT1_4471(.VSS(VSS),.VDD(VDD),.Y(g7717),.A(I14028));
  NOT NOT1_4472(.VSS(VSS),.VDD(VDD),.Y(I14031),.A(g7448));
  NOT NOT1_4473(.VSS(VSS),.VDD(VDD),.Y(g7718),.A(I14031));
  NOT NOT1_4474(.VSS(VSS),.VDD(VDD),.Y(g7719),.A(g7475));
  NOT NOT1_4475(.VSS(VSS),.VDD(VDD),.Y(I14035),.A(g7310));
  NOT NOT1_4476(.VSS(VSS),.VDD(VDD),.Y(g7720),.A(I14035));
  NOT NOT1_4477(.VSS(VSS),.VDD(VDD),.Y(g7721),.A(g7344));
  NOT NOT1_4478(.VSS(VSS),.VDD(VDD),.Y(I14039),.A(g7449));
  NOT NOT1_4479(.VSS(VSS),.VDD(VDD),.Y(g7722),.A(I14039));
  NOT NOT1_4480(.VSS(VSS),.VDD(VDD),.Y(I14042),.A(g7470));
  NOT NOT1_4481(.VSS(VSS),.VDD(VDD),.Y(g7723),.A(I14042));
  NOT NOT1_4482(.VSS(VSS),.VDD(VDD),.Y(I14046),.A(g7492));
  NOT NOT1_4483(.VSS(VSS),.VDD(VDD),.Y(g7725),.A(I14046));
  NOT NOT1_4484(.VSS(VSS),.VDD(VDD),.Y(I14049),.A(g7493));
  NOT NOT1_4485(.VSS(VSS),.VDD(VDD),.Y(g7726),.A(I14049));
  NOT NOT1_4486(.VSS(VSS),.VDD(VDD),.Y(I14052),.A(g7494));
  NOT NOT1_4487(.VSS(VSS),.VDD(VDD),.Y(g7727),.A(I14052));
  NOT NOT1_4488(.VSS(VSS),.VDD(VDD),.Y(I14055),.A(g7495));
  NOT NOT1_4489(.VSS(VSS),.VDD(VDD),.Y(g7728),.A(I14055));
  NOT NOT1_4490(.VSS(VSS),.VDD(VDD),.Y(I14058),.A(g7544));
  NOT NOT1_4491(.VSS(VSS),.VDD(VDD),.Y(g7729),.A(I14058));
  NOT NOT1_4492(.VSS(VSS),.VDD(VDD),.Y(I14061),.A(g7546));
  NOT NOT1_4493(.VSS(VSS),.VDD(VDD),.Y(g7730),.A(I14061));
  NOT NOT1_4494(.VSS(VSS),.VDD(VDD),.Y(I14064),.A(g7556));
  NOT NOT1_4495(.VSS(VSS),.VDD(VDD),.Y(g7731),.A(I14064));
  NOT NOT1_4496(.VSS(VSS),.VDD(VDD),.Y(I14067),.A(g7550));
  NOT NOT1_4497(.VSS(VSS),.VDD(VDD),.Y(g7732),.A(I14067));
  NOT NOT1_4498(.VSS(VSS),.VDD(VDD),.Y(I14070),.A(g7714));
  NOT NOT1_4499(.VSS(VSS),.VDD(VDD),.Y(g7733),.A(I14070));
  NOT NOT1_4500(.VSS(VSS),.VDD(VDD),.Y(I14073),.A(g7627));
  NOT NOT1_4501(.VSS(VSS),.VDD(VDD),.Y(g7734),.A(I14073));
  NOT NOT1_4502(.VSS(VSS),.VDD(VDD),.Y(I14076),.A(g7577));
  NOT NOT1_4503(.VSS(VSS),.VDD(VDD),.Y(g7735),.A(I14076));
  NOT NOT1_4504(.VSS(VSS),.VDD(VDD),.Y(I14079),.A(g7579));
  NOT NOT1_4505(.VSS(VSS),.VDD(VDD),.Y(g7736),.A(I14079));
  NOT NOT1_4506(.VSS(VSS),.VDD(VDD),.Y(I14082),.A(g7539));
  NOT NOT1_4507(.VSS(VSS),.VDD(VDD),.Y(g7737),.A(I14082));
  NOT NOT1_4508(.VSS(VSS),.VDD(VDD),.Y(I14085),.A(g7583));
  NOT NOT1_4509(.VSS(VSS),.VDD(VDD),.Y(g7738),.A(I14085));
  NOT NOT1_4510(.VSS(VSS),.VDD(VDD),.Y(I14088),.A(g7585));
  NOT NOT1_4511(.VSS(VSS),.VDD(VDD),.Y(g7739),.A(I14088));
  NOT NOT1_4512(.VSS(VSS),.VDD(VDD),.Y(I14091),.A(g7589));
  NOT NOT1_4513(.VSS(VSS),.VDD(VDD),.Y(g7740),.A(I14091));
  NOT NOT1_4514(.VSS(VSS),.VDD(VDD),.Y(I14094),.A(g7593));
  NOT NOT1_4515(.VSS(VSS),.VDD(VDD),.Y(g7741),.A(I14094));
  NOT NOT1_4516(.VSS(VSS),.VDD(VDD),.Y(I14097),.A(g7595));
  NOT NOT1_4517(.VSS(VSS),.VDD(VDD),.Y(g7742),.A(I14097));
  NOT NOT1_4518(.VSS(VSS),.VDD(VDD),.Y(I14100),.A(g7580));
  NOT NOT1_4519(.VSS(VSS),.VDD(VDD),.Y(g7743),.A(I14100));
  NOT NOT1_4520(.VSS(VSS),.VDD(VDD),.Y(I14103),.A(g7584));
  NOT NOT1_4521(.VSS(VSS),.VDD(VDD),.Y(g7744),.A(I14103));
  NOT NOT1_4522(.VSS(VSS),.VDD(VDD),.Y(I14106),.A(g7586));
  NOT NOT1_4523(.VSS(VSS),.VDD(VDD),.Y(g7745),.A(I14106));
  NOT NOT1_4524(.VSS(VSS),.VDD(VDD),.Y(I14109),.A(g7590));
  NOT NOT1_4525(.VSS(VSS),.VDD(VDD),.Y(g7746),.A(I14109));
  NOT NOT1_4526(.VSS(VSS),.VDD(VDD),.Y(I14112),.A(g7560));
  NOT NOT1_4527(.VSS(VSS),.VDD(VDD),.Y(g7747),.A(I14112));
  NOT NOT1_4528(.VSS(VSS),.VDD(VDD),.Y(I14115),.A(g7563));
  NOT NOT1_4529(.VSS(VSS),.VDD(VDD),.Y(g7748),.A(I14115));
  NOT NOT1_4530(.VSS(VSS),.VDD(VDD),.Y(I14118),.A(g7565));
  NOT NOT1_4531(.VSS(VSS),.VDD(VDD),.Y(g7749),.A(I14118));
  NOT NOT1_4532(.VSS(VSS),.VDD(VDD),.Y(I14121),.A(g7587));
  NOT NOT1_4533(.VSS(VSS),.VDD(VDD),.Y(g7750),.A(I14121));
  NOT NOT1_4534(.VSS(VSS),.VDD(VDD),.Y(I14124),.A(g7591));
  NOT NOT1_4535(.VSS(VSS),.VDD(VDD),.Y(g7751),.A(I14124));
  NOT NOT1_4536(.VSS(VSS),.VDD(VDD),.Y(I14127),.A(g7594));
  NOT NOT1_4537(.VSS(VSS),.VDD(VDD),.Y(g7752),.A(I14127));
  NOT NOT1_4538(.VSS(VSS),.VDD(VDD),.Y(I14130),.A(g7592));
  NOT NOT1_4539(.VSS(VSS),.VDD(VDD),.Y(g7753),.A(I14130));
  NOT NOT1_4540(.VSS(VSS),.VDD(VDD),.Y(I14133),.A(g7574));
  NOT NOT1_4541(.VSS(VSS),.VDD(VDD),.Y(g7754),.A(I14133));
  NOT NOT1_4542(.VSS(VSS),.VDD(VDD),.Y(I14136),.A(g7633));
  NOT NOT1_4543(.VSS(VSS),.VDD(VDD),.Y(g7755),.A(I14136));
  NOT NOT1_4544(.VSS(VSS),.VDD(VDD),.Y(I14139),.A(g7548));
  NOT NOT1_4545(.VSS(VSS),.VDD(VDD),.Y(g7756),.A(I14139));
  NOT NOT1_4546(.VSS(VSS),.VDD(VDD),.Y(I14142),.A(g7551));
  NOT NOT1_4547(.VSS(VSS),.VDD(VDD),.Y(g7757),.A(I14142));
  NOT NOT1_4548(.VSS(VSS),.VDD(VDD),.Y(I14145),.A(g7542));
  NOT NOT1_4549(.VSS(VSS),.VDD(VDD),.Y(g7758),.A(I14145));
  NOT NOT1_4550(.VSS(VSS),.VDD(VDD),.Y(I14148),.A(g7543));
  NOT NOT1_4551(.VSS(VSS),.VDD(VDD),.Y(g7759),.A(I14148));
  NOT NOT1_4552(.VSS(VSS),.VDD(VDD),.Y(I14151),.A(g7555));
  NOT NOT1_4553(.VSS(VSS),.VDD(VDD),.Y(g7760),.A(I14151));
  NOT NOT1_4554(.VSS(VSS),.VDD(VDD),.Y(I14154),.A(g7558));
  NOT NOT1_4555(.VSS(VSS),.VDD(VDD),.Y(g7761),.A(I14154));
  NOT NOT1_4556(.VSS(VSS),.VDD(VDD),.Y(I14157),.A(g7547));
  NOT NOT1_4557(.VSS(VSS),.VDD(VDD),.Y(g7762),.A(I14157));
  NOT NOT1_4558(.VSS(VSS),.VDD(VDD),.Y(I14160),.A(g7549));
  NOT NOT1_4559(.VSS(VSS),.VDD(VDD),.Y(g7763),.A(I14160));
  NOT NOT1_4560(.VSS(VSS),.VDD(VDD),.Y(I14163),.A(g7533));
  NOT NOT1_4561(.VSS(VSS),.VDD(VDD),.Y(g7764),.A(I14163));
  NOT NOT1_4562(.VSS(VSS),.VDD(VDD),.Y(I14166),.A(g7702));
  NOT NOT1_4563(.VSS(VSS),.VDD(VDD),.Y(g7765),.A(I14166));
  NOT NOT1_4564(.VSS(VSS),.VDD(VDD),.Y(I14169),.A(g7715));
  NOT NOT1_4565(.VSS(VSS),.VDD(VDD),.Y(g7766),.A(I14169));
  NOT NOT1_4566(.VSS(VSS),.VDD(VDD),.Y(I14172),.A(g7545));
  NOT NOT1_4567(.VSS(VSS),.VDD(VDD),.Y(g7767),.A(I14172));
  NOT NOT1_4568(.VSS(VSS),.VDD(VDD),.Y(I14175),.A(g7718));
  NOT NOT1_4569(.VSS(VSS),.VDD(VDD),.Y(g7768),.A(I14175));
  NOT NOT1_4570(.VSS(VSS),.VDD(VDD),.Y(I14178),.A(g7562));
  NOT NOT1_4571(.VSS(VSS),.VDD(VDD),.Y(g7769),.A(I14178));
  NOT NOT1_4572(.VSS(VSS),.VDD(VDD),.Y(I14181),.A(g7725));
  NOT NOT1_4573(.VSS(VSS),.VDD(VDD),.Y(g7770),.A(I14181));
  NOT NOT1_4574(.VSS(VSS),.VDD(VDD),.Y(I14184),.A(g7726));
  NOT NOT1_4575(.VSS(VSS),.VDD(VDD),.Y(g7771),.A(I14184));
  NOT NOT1_4576(.VSS(VSS),.VDD(VDD),.Y(I14187),.A(g7728));
  NOT NOT1_4577(.VSS(VSS),.VDD(VDD),.Y(g7772),.A(I14187));
  NOT NOT1_4578(.VSS(VSS),.VDD(VDD),.Y(I14190),.A(g7531));
  NOT NOT1_4579(.VSS(VSS),.VDD(VDD),.Y(g7773),.A(I14190));
  NOT NOT1_4580(.VSS(VSS),.VDD(VDD),.Y(I14193),.A(g7532));
  NOT NOT1_4581(.VSS(VSS),.VDD(VDD),.Y(g7774),.A(I14193));
  NOT NOT1_4582(.VSS(VSS),.VDD(VDD),.Y(I14196),.A(g7534));
  NOT NOT1_4583(.VSS(VSS),.VDD(VDD),.Y(g7775),.A(I14196));
  NOT NOT1_4584(.VSS(VSS),.VDD(VDD),.Y(I14199),.A(g7704));
  NOT NOT1_4585(.VSS(VSS),.VDD(VDD),.Y(g7776),.A(I14199));
  NOT NOT1_4586(.VSS(VSS),.VDD(VDD),.Y(I14202),.A(g7708));
  NOT NOT1_4587(.VSS(VSS),.VDD(VDD),.Y(g7777),.A(I14202));
  NOT NOT1_4588(.VSS(VSS),.VDD(VDD),.Y(I14205),.A(g7710));
  NOT NOT1_4589(.VSS(VSS),.VDD(VDD),.Y(g7778),.A(I14205));
  NOT NOT1_4590(.VSS(VSS),.VDD(VDD),.Y(I14208),.A(g7711));
  NOT NOT1_4591(.VSS(VSS),.VDD(VDD),.Y(g7779),.A(I14208));
  NOT NOT1_4592(.VSS(VSS),.VDD(VDD),.Y(I14211),.A(g7712));
  NOT NOT1_4593(.VSS(VSS),.VDD(VDD),.Y(g7780),.A(I14211));
  NOT NOT1_4594(.VSS(VSS),.VDD(VDD),.Y(I14214),.A(g7576));
  NOT NOT1_4595(.VSS(VSS),.VDD(VDD),.Y(g7781),.A(I14214));
  NOT NOT1_4596(.VSS(VSS),.VDD(VDD),.Y(I14224),.A(g7722));
  NOT NOT1_4597(.VSS(VSS),.VDD(VDD),.Y(g7789),.A(I14224));
  NOT NOT1_4598(.VSS(VSS),.VDD(VDD),.Y(I14227),.A(g7552));
  NOT NOT1_4599(.VSS(VSS),.VDD(VDD),.Y(g7790),.A(I14227));
  NOT NOT1_4600(.VSS(VSS),.VDD(VDD),.Y(I14231),.A(g7566));
  NOT NOT1_4601(.VSS(VSS),.VDD(VDD),.Y(g7792),.A(I14231));
  NOT NOT1_4602(.VSS(VSS),.VDD(VDD),.Y(I14234),.A(g7614));
  NOT NOT1_4603(.VSS(VSS),.VDD(VDD),.Y(g7793),.A(I14234));
  NOT NOT1_4604(.VSS(VSS),.VDD(VDD),.Y(I14238),.A(g7608));
  NOT NOT1_4605(.VSS(VSS),.VDD(VDD),.Y(g7811),.A(I14238));
  NOT NOT1_4606(.VSS(VSS),.VDD(VDD),.Y(I14251),.A(g7541));
  NOT NOT1_4607(.VSS(VSS),.VDD(VDD),.Y(g7829),.A(I14251));
  NOT NOT1_4608(.VSS(VSS),.VDD(VDD),.Y(I14257),.A(g7716));
  NOT NOT1_4609(.VSS(VSS),.VDD(VDD),.Y(g7835),.A(I14257));
  NOT NOT1_4610(.VSS(VSS),.VDD(VDD),.Y(I14260),.A(g7717));
  NOT NOT1_4611(.VSS(VSS),.VDD(VDD),.Y(g7836),.A(I14260));
  NOT NOT1_4612(.VSS(VSS),.VDD(VDD),.Y(I14264),.A(g7698));
  NOT NOT1_4613(.VSS(VSS),.VDD(VDD),.Y(g7838),.A(I14264));
  NOT NOT1_4614(.VSS(VSS),.VDD(VDD),.Y(I14267),.A(g7695));
  NOT NOT1_4615(.VSS(VSS),.VDD(VDD),.Y(g7855),.A(I14267));
  NOT NOT1_4616(.VSS(VSS),.VDD(VDD),.Y(I14270),.A(g7703));
  NOT NOT1_4617(.VSS(VSS),.VDD(VDD),.Y(g7870),.A(I14270));
  NOT NOT1_4618(.VSS(VSS),.VDD(VDD),.Y(I14273),.A(g7631));
  NOT NOT1_4619(.VSS(VSS),.VDD(VDD),.Y(g7887),.A(I14273));
  NOT NOT1_4620(.VSS(VSS),.VDD(VDD),.Y(I14276),.A(g7720));
  NOT NOT1_4621(.VSS(VSS),.VDD(VDD),.Y(g7904),.A(I14276));
  NOT NOT1_4622(.VSS(VSS),.VDD(VDD),.Y(I14279),.A(g7700));
  NOT NOT1_4623(.VSS(VSS),.VDD(VDD),.Y(g7905),.A(I14279));
  NOT NOT1_4624(.VSS(VSS),.VDD(VDD),.Y(I14282),.A(g7709));
  NOT NOT1_4625(.VSS(VSS),.VDD(VDD),.Y(g7920),.A(I14282));
  NOT NOT1_4626(.VSS(VSS),.VDD(VDD),.Y(I14285),.A(g7625));
  NOT NOT1_4627(.VSS(VSS),.VDD(VDD),.Y(g7937),.A(I14285));
  NOT NOT1_4628(.VSS(VSS),.VDD(VDD),.Y(I14288),.A(g7705));
  NOT NOT1_4629(.VSS(VSS),.VDD(VDD),.Y(g7951),.A(I14288));
  NOT NOT1_4630(.VSS(VSS),.VDD(VDD),.Y(I14291),.A(g7680));
  NOT NOT1_4631(.VSS(VSS),.VDD(VDD),.Y(g7966),.A(I14291));
  NOT NOT1_4632(.VSS(VSS),.VDD(VDD),.Y(I14294),.A(g7553));
  NOT NOT1_4633(.VSS(VSS),.VDD(VDD),.Y(g7983),.A(I14294));
  NOT NOT1_4634(.VSS(VSS),.VDD(VDD),.Y(g7992),.A(g7557));
  NOT NOT1_4635(.VSS(VSS),.VDD(VDD),.Y(I14298),.A(g7678));
  NOT NOT1_4636(.VSS(VSS),.VDD(VDD),.Y(g7993),.A(I14298));
  NOT NOT1_4637(.VSS(VSS),.VDD(VDD),.Y(g8008),.A(g7559));
  NOT NOT1_4638(.VSS(VSS),.VDD(VDD),.Y(I14305),.A(g7537));
  NOT NOT1_4639(.VSS(VSS),.VDD(VDD),.Y(g8012),.A(I14305));
  NOT NOT1_4640(.VSS(VSS),.VDD(VDD),.Y(g8013),.A(g7561));
  NOT NOT1_4641(.VSS(VSS),.VDD(VDD),.Y(g8014),.A(g7564));
  NOT NOT1_4642(.VSS(VSS),.VDD(VDD),.Y(g8015),.A(g7689));
  NOT NOT1_4643(.VSS(VSS),.VDD(VDD),.Y(I14311),.A(g7566));
  NOT NOT1_4644(.VSS(VSS),.VDD(VDD),.Y(g8016),.A(I14311));
  NOT NOT1_4645(.VSS(VSS),.VDD(VDD),.Y(g8017),.A(g7692));
  NOT NOT1_4646(.VSS(VSS),.VDD(VDD),.Y(I14315),.A(g7676));
  NOT NOT1_4647(.VSS(VSS),.VDD(VDD),.Y(g8018),.A(I14315));
  NOT NOT1_4648(.VSS(VSS),.VDD(VDD),.Y(I14318),.A(g7657));
  NOT NOT1_4649(.VSS(VSS),.VDD(VDD),.Y(g8029),.A(I14318));
  NOT NOT1_4650(.VSS(VSS),.VDD(VDD),.Y(g8038),.A(g7694));
  NOT NOT1_4651(.VSS(VSS),.VDD(VDD),.Y(g8039),.A(g7696));
  NOT NOT1_4652(.VSS(VSS),.VDD(VDD),.Y(g8040),.A(g7699));
  NOT NOT1_4653(.VSS(VSS),.VDD(VDD),.Y(g8041),.A(g7701));
  NOT NOT1_4654(.VSS(VSS),.VDD(VDD),.Y(I14325),.A(g7713));
  NOT NOT1_4655(.VSS(VSS),.VDD(VDD),.Y(g8042),.A(I14325));
  NOT NOT1_4656(.VSS(VSS),.VDD(VDD),.Y(I14330),.A(g7538));
  NOT NOT1_4657(.VSS(VSS),.VDD(VDD),.Y(g8061),.A(I14330));
  NOT NOT1_4658(.VSS(VSS),.VDD(VDD),.Y(I14334),.A(g7578));
  NOT NOT1_4659(.VSS(VSS),.VDD(VDD),.Y(g8063),.A(I14334));
  NOT NOT1_4660(.VSS(VSS),.VDD(VDD),.Y(I14338),.A(g7581));
  NOT NOT1_4661(.VSS(VSS),.VDD(VDD),.Y(g8065),.A(I14338));
  NOT NOT1_4662(.VSS(VSS),.VDD(VDD),.Y(I14342),.A(g7582));
  NOT NOT1_4663(.VSS(VSS),.VDD(VDD),.Y(g8067),.A(I14342));
  NOT NOT1_4664(.VSS(VSS),.VDD(VDD),.Y(I14349),.A(g7588));
  NOT NOT1_4665(.VSS(VSS),.VDD(VDD),.Y(g8072),.A(I14349));
  NOT NOT1_4666(.VSS(VSS),.VDD(VDD),.Y(I14370),.A(g7603));
  NOT NOT1_4667(.VSS(VSS),.VDD(VDD),.Y(g8093),.A(I14370));
  NOT NOT1_4668(.VSS(VSS),.VDD(VDD),.Y(g8094),.A(g7705));
  NOT NOT1_4669(.VSS(VSS),.VDD(VDD),.Y(I14374),.A(g7693));
  NOT NOT1_4670(.VSS(VSS),.VDD(VDD),.Y(g8111),.A(I14374));
  NOT NOT1_4671(.VSS(VSS),.VDD(VDD),.Y(I14378),.A(g7691));
  NOT NOT1_4672(.VSS(VSS),.VDD(VDD),.Y(g8131),.A(I14378));
  NOT NOT1_4673(.VSS(VSS),.VDD(VDD),.Y(I14381),.A(g7596));
  NOT NOT1_4674(.VSS(VSS),.VDD(VDD),.Y(g8145),.A(I14381));
  NOT NOT1_4675(.VSS(VSS),.VDD(VDD),.Y(I14388),.A(g7605));
  NOT NOT1_4676(.VSS(VSS),.VDD(VDD),.Y(g8152),.A(I14388));
  NOT NOT1_4677(.VSS(VSS),.VDD(VDD),.Y(I14394),.A(g7536));
  NOT NOT1_4678(.VSS(VSS),.VDD(VDD),.Y(g8156),.A(I14394));
  NOT NOT1_4679(.VSS(VSS),.VDD(VDD),.Y(I14397),.A(g7686));
  NOT NOT1_4680(.VSS(VSS),.VDD(VDD),.Y(g8172),.A(I14397));
  NOT NOT1_4681(.VSS(VSS),.VDD(VDD),.Y(I14400),.A(g7677));
  NOT NOT1_4682(.VSS(VSS),.VDD(VDD),.Y(g8173),.A(I14400));
  NOT NOT1_4683(.VSS(VSS),.VDD(VDD),.Y(I14403),.A(g7679));
  NOT NOT1_4684(.VSS(VSS),.VDD(VDD),.Y(g8174),.A(I14403));
  NOT NOT1_4685(.VSS(VSS),.VDD(VDD),.Y(I14406),.A(g7681));
  NOT NOT1_4686(.VSS(VSS),.VDD(VDD),.Y(g8175),.A(I14406));
  NOT NOT1_4687(.VSS(VSS),.VDD(VDD),.Y(I14410),.A(g7697));
  NOT NOT1_4688(.VSS(VSS),.VDD(VDD),.Y(g8177),.A(I14410));
  NOT NOT1_4689(.VSS(VSS),.VDD(VDD),.Y(I14413),.A(g7723));
  NOT NOT1_4690(.VSS(VSS),.VDD(VDD),.Y(g8178),.A(I14413));
  NOT NOT1_4691(.VSS(VSS),.VDD(VDD),.Y(I14416),.A(g7727));
  NOT NOT1_4692(.VSS(VSS),.VDD(VDD),.Y(g8179),.A(I14416));
  NOT NOT1_4693(.VSS(VSS),.VDD(VDD),.Y(g8180),.A(g7719));
  NOT NOT1_4694(.VSS(VSS),.VDD(VDD),.Y(I14420),.A(g7554));
  NOT NOT1_4695(.VSS(VSS),.VDD(VDD),.Y(g8181),.A(I14420));
  NOT NOT1_4696(.VSS(VSS),.VDD(VDD),.Y(g8198),.A(g7721));
  NOT NOT1_4697(.VSS(VSS),.VDD(VDD),.Y(I14424),.A(g7652));
  NOT NOT1_4698(.VSS(VSS),.VDD(VDD),.Y(g8199),.A(I14424));
  NOT NOT1_4699(.VSS(VSS),.VDD(VDD),.Y(I14427),.A(g7835));
  NOT NOT1_4700(.VSS(VSS),.VDD(VDD),.Y(g8216),.A(I14427));
  NOT NOT1_4701(.VSS(VSS),.VDD(VDD),.Y(I14430),.A(g7836));
  NOT NOT1_4702(.VSS(VSS),.VDD(VDD),.Y(g8217),.A(I14430));
  NOT NOT1_4703(.VSS(VSS),.VDD(VDD),.Y(I14433),.A(g8061));
  NOT NOT1_4704(.VSS(VSS),.VDD(VDD),.Y(g8218),.A(I14433));
  NOT NOT1_4705(.VSS(VSS),.VDD(VDD),.Y(I14436),.A(g7904));
  NOT NOT1_4706(.VSS(VSS),.VDD(VDD),.Y(g8219),.A(I14436));
  NOT NOT1_4707(.VSS(VSS),.VDD(VDD),.Y(I14439),.A(g8063));
  NOT NOT1_4708(.VSS(VSS),.VDD(VDD),.Y(g8220),.A(I14439));
  NOT NOT1_4709(.VSS(VSS),.VDD(VDD),.Y(I14442),.A(g8065));
  NOT NOT1_4710(.VSS(VSS),.VDD(VDD),.Y(g8221),.A(I14442));
  NOT NOT1_4711(.VSS(VSS),.VDD(VDD),.Y(I14445),.A(g8067));
  NOT NOT1_4712(.VSS(VSS),.VDD(VDD),.Y(g8222),.A(I14445));
  NOT NOT1_4713(.VSS(VSS),.VDD(VDD),.Y(I14448),.A(g7792));
  NOT NOT1_4714(.VSS(VSS),.VDD(VDD),.Y(g8223),.A(I14448));
  NOT NOT1_4715(.VSS(VSS),.VDD(VDD),.Y(I14451),.A(g8172));
  NOT NOT1_4716(.VSS(VSS),.VDD(VDD),.Y(g8224),.A(I14451));
  NOT NOT1_4717(.VSS(VSS),.VDD(VDD),.Y(I14454),.A(g8177));
  NOT NOT1_4718(.VSS(VSS),.VDD(VDD),.Y(g8225),.A(I14454));
  NOT NOT1_4719(.VSS(VSS),.VDD(VDD),.Y(I14457),.A(g8093));
  NOT NOT1_4720(.VSS(VSS),.VDD(VDD),.Y(g8226),.A(I14457));
  NOT NOT1_4721(.VSS(VSS),.VDD(VDD),.Y(I14460),.A(g7789));
  NOT NOT1_4722(.VSS(VSS),.VDD(VDD),.Y(g8227),.A(I14460));
  NOT NOT1_4723(.VSS(VSS),.VDD(VDD),.Y(I14463),.A(g8072));
  NOT NOT1_4724(.VSS(VSS),.VDD(VDD),.Y(g8228),.A(I14463));
  NOT NOT1_4725(.VSS(VSS),.VDD(VDD),.Y(I14489),.A(g7829));
  NOT NOT1_4726(.VSS(VSS),.VDD(VDD),.Y(g8234),.A(I14489));
  NOT NOT1_4727(.VSS(VSS),.VDD(VDD),.Y(I14492),.A(g7829));
  NOT NOT1_4728(.VSS(VSS),.VDD(VDD),.Y(g8235),.A(I14492));
  NOT NOT1_4729(.VSS(VSS),.VDD(VDD),.Y(I14531),.A(g8178));
  NOT NOT1_4730(.VSS(VSS),.VDD(VDD),.Y(g8284),.A(I14531));
  NOT NOT1_4731(.VSS(VSS),.VDD(VDD),.Y(I14573),.A(g8179));
  NOT NOT1_4732(.VSS(VSS),.VDD(VDD),.Y(g8324),.A(I14573));
  NOT NOT1_4733(.VSS(VSS),.VDD(VDD),.Y(g8342),.A(g8008));
  NOT NOT1_4734(.VSS(VSS),.VDD(VDD),.Y(g8363),.A(g7992));
  NOT NOT1_4735(.VSS(VSS),.VDD(VDD),.Y(I14603),.A(g7827));
  NOT NOT1_4736(.VSS(VSS),.VDD(VDD),.Y(g8381),.A(I14603));
  NOT NOT1_4737(.VSS(VSS),.VDD(VDD),.Y(g8386),.A(g8014));
  NOT NOT1_4738(.VSS(VSS),.VDD(VDD),.Y(I14614),.A(g7832));
  NOT NOT1_4739(.VSS(VSS),.VDD(VDD),.Y(g8406),.A(I14614));
  NOT NOT1_4740(.VSS(VSS),.VDD(VDD),.Y(g8407),.A(g8013));
  NOT NOT1_4741(.VSS(VSS),.VDD(VDD),.Y(g8421),.A(g8017));
  NOT NOT1_4742(.VSS(VSS),.VDD(VDD),.Y(I14623),.A(g7833));
  NOT NOT1_4743(.VSS(VSS),.VDD(VDD),.Y(g8442),.A(I14623));
  NOT NOT1_4744(.VSS(VSS),.VDD(VDD),.Y(g8443),.A(g8015));
  NOT NOT1_4745(.VSS(VSS),.VDD(VDD),.Y(g8463),.A(g8094));
  NOT NOT1_4746(.VSS(VSS),.VDD(VDD),.Y(g8464),.A(g8039));
  NOT NOT1_4747(.VSS(VSS),.VDD(VDD),.Y(I14637),.A(g8012));
  NOT NOT1_4748(.VSS(VSS),.VDD(VDD),.Y(g8481),.A(I14637));
  NOT NOT1_4749(.VSS(VSS),.VDD(VDD),.Y(g8482),.A(g8094));
  NOT NOT1_4750(.VSS(VSS),.VDD(VDD),.Y(g8483),.A(g8038));
  NOT NOT1_4751(.VSS(VSS),.VDD(VDD),.Y(g8493),.A(g8041));
  NOT NOT1_4752(.VSS(VSS),.VDD(VDD),.Y(I14643),.A(g7837));
  NOT NOT1_4753(.VSS(VSS),.VDD(VDD),.Y(g8510),.A(I14643));
  NOT NOT1_4754(.VSS(VSS),.VDD(VDD),.Y(I14646),.A(g7790));
  NOT NOT1_4755(.VSS(VSS),.VDD(VDD),.Y(g8511),.A(I14646));
  NOT NOT1_4756(.VSS(VSS),.VDD(VDD),.Y(g8512),.A(g8094));
  NOT NOT1_4757(.VSS(VSS),.VDD(VDD),.Y(g8514),.A(g8040));
  NOT NOT1_4758(.VSS(VSS),.VDD(VDD),.Y(g8524),.A(g7855));
  NOT NOT1_4759(.VSS(VSS),.VDD(VDD),.Y(g8541),.A(g8094));
  NOT NOT1_4760(.VSS(VSS),.VDD(VDD),.Y(I14657),.A(g7782));
  NOT NOT1_4761(.VSS(VSS),.VDD(VDD),.Y(g8544),.A(I14657));
  NOT NOT1_4762(.VSS(VSS),.VDD(VDD),.Y(g8545),.A(g7905));
  NOT NOT1_4763(.VSS(VSS),.VDD(VDD),.Y(g8562),.A(g8094));
  NOT NOT1_4764(.VSS(VSS),.VDD(VDD),.Y(I14662),.A(g7783));
  NOT NOT1_4765(.VSS(VSS),.VDD(VDD),.Y(g8563),.A(I14662));
  NOT NOT1_4766(.VSS(VSS),.VDD(VDD),.Y(g8564),.A(g7951));
  NOT NOT1_4767(.VSS(VSS),.VDD(VDD),.Y(g8581),.A(g8094));
  NOT NOT1_4768(.VSS(VSS),.VDD(VDD),.Y(g8582),.A(g8094));
  NOT NOT1_4769(.VSS(VSS),.VDD(VDD),.Y(I14668),.A(g7787));
  NOT NOT1_4770(.VSS(VSS),.VDD(VDD),.Y(g8583),.A(I14668));
  NOT NOT1_4771(.VSS(VSS),.VDD(VDD),.Y(g8585),.A(g7993));
  NOT NOT1_4772(.VSS(VSS),.VDD(VDD),.Y(g8602),.A(g8094));
  NOT NOT1_4773(.VSS(VSS),.VDD(VDD),.Y(I14674),.A(g7788));
  NOT NOT1_4774(.VSS(VSS),.VDD(VDD),.Y(g8603),.A(I14674));
  NOT NOT1_4775(.VSS(VSS),.VDD(VDD),.Y(I14677),.A(g7791));
  NOT NOT1_4776(.VSS(VSS),.VDD(VDD),.Y(g8604),.A(I14677));
  NOT NOT1_4777(.VSS(VSS),.VDD(VDD),.Y(I14680),.A(g7810));
  NOT NOT1_4778(.VSS(VSS),.VDD(VDD),.Y(g8605),.A(I14680));
  NOT NOT1_4779(.VSS(VSS),.VDD(VDD),.Y(I14683),.A(g7825));
  NOT NOT1_4780(.VSS(VSS),.VDD(VDD),.Y(g8606),.A(I14683));
  NOT NOT1_4781(.VSS(VSS),.VDD(VDD),.Y(I14687),.A(g7826));
  NOT NOT1_4782(.VSS(VSS),.VDD(VDD),.Y(g8608),.A(I14687));
  NOT NOT1_4783(.VSS(VSS),.VDD(VDD),.Y(I14695),.A(g8016));
  NOT NOT1_4784(.VSS(VSS),.VDD(VDD),.Y(g8619),.A(I14695));
  NOT NOT1_4785(.VSS(VSS),.VDD(VDD),.Y(I14709),.A(g8198));
  NOT NOT1_4786(.VSS(VSS),.VDD(VDD),.Y(g8631),.A(I14709));
  NOT NOT1_4787(.VSS(VSS),.VDD(VDD),.Y(I14712),.A(g8059));
  NOT NOT1_4788(.VSS(VSS),.VDD(VDD),.Y(g8632),.A(I14712));
  NOT NOT1_4789(.VSS(VSS),.VDD(VDD),.Y(I14718),.A(g8068));
  NOT NOT1_4790(.VSS(VSS),.VDD(VDD),.Y(g8636),.A(I14718));
  NOT NOT1_4791(.VSS(VSS),.VDD(VDD),.Y(I14722),.A(g8076));
  NOT NOT1_4792(.VSS(VSS),.VDD(VDD),.Y(g8638),.A(I14722));
  NOT NOT1_4793(.VSS(VSS),.VDD(VDD),.Y(I14725),.A(g8145));
  NOT NOT1_4794(.VSS(VSS),.VDD(VDD),.Y(g8639),.A(I14725));
  NOT NOT1_4795(.VSS(VSS),.VDD(VDD),.Y(I14728),.A(g8152));
  NOT NOT1_4796(.VSS(VSS),.VDD(VDD),.Y(g8640),.A(I14728));
  NOT NOT1_4797(.VSS(VSS),.VDD(VDD),.Y(I14732),.A(g8155));
  NOT NOT1_4798(.VSS(VSS),.VDD(VDD),.Y(g8642),.A(I14732));
  NOT NOT1_4799(.VSS(VSS),.VDD(VDD),.Y(I14739),.A(g8173));
  NOT NOT1_4800(.VSS(VSS),.VDD(VDD),.Y(g8647),.A(I14739));
  NOT NOT1_4801(.VSS(VSS),.VDD(VDD),.Y(I14743),.A(g8174));
  NOT NOT1_4802(.VSS(VSS),.VDD(VDD),.Y(g8649),.A(I14743));
  NOT NOT1_4803(.VSS(VSS),.VDD(VDD),.Y(I14747),.A(g8175));
  NOT NOT1_4804(.VSS(VSS),.VDD(VDD),.Y(g8651),.A(I14747));
  NOT NOT1_4805(.VSS(VSS),.VDD(VDD),.Y(I14763),.A(g7834));
  NOT NOT1_4806(.VSS(VSS),.VDD(VDD),.Y(g8657),.A(I14763));
  NOT NOT1_4807(.VSS(VSS),.VDD(VDD),.Y(I14777),.A(g8511));
  NOT NOT1_4808(.VSS(VSS),.VDD(VDD),.Y(g8661),.A(I14777));
  NOT NOT1_4809(.VSS(VSS),.VDD(VDD),.Y(I14780),.A(g8284));
  NOT NOT1_4810(.VSS(VSS),.VDD(VDD),.Y(g8662),.A(I14780));
  NOT NOT1_4811(.VSS(VSS),.VDD(VDD),.Y(I14783),.A(g8324));
  NOT NOT1_4812(.VSS(VSS),.VDD(VDD),.Y(g8663),.A(I14783));
  NOT NOT1_4813(.VSS(VSS),.VDD(VDD),.Y(I14786),.A(g8606));
  NOT NOT1_4814(.VSS(VSS),.VDD(VDD),.Y(g8664),.A(I14786));
  NOT NOT1_4815(.VSS(VSS),.VDD(VDD),.Y(I14789),.A(g8544));
  NOT NOT1_4816(.VSS(VSS),.VDD(VDD),.Y(g8665),.A(I14789));
  NOT NOT1_4817(.VSS(VSS),.VDD(VDD),.Y(I14792),.A(g8583));
  NOT NOT1_4818(.VSS(VSS),.VDD(VDD),.Y(g8666),.A(I14792));
  NOT NOT1_4819(.VSS(VSS),.VDD(VDD),.Y(I14795),.A(g8604));
  NOT NOT1_4820(.VSS(VSS),.VDD(VDD),.Y(g8667),.A(I14795));
  NOT NOT1_4821(.VSS(VSS),.VDD(VDD),.Y(I14798),.A(g8605));
  NOT NOT1_4822(.VSS(VSS),.VDD(VDD),.Y(g8668),.A(I14798));
  NOT NOT1_4823(.VSS(VSS),.VDD(VDD),.Y(I14801),.A(g8608));
  NOT NOT1_4824(.VSS(VSS),.VDD(VDD),.Y(g8669),.A(I14801));
  NOT NOT1_4825(.VSS(VSS),.VDD(VDD),.Y(I14804),.A(g8563));
  NOT NOT1_4826(.VSS(VSS),.VDD(VDD),.Y(g8670),.A(I14804));
  NOT NOT1_4827(.VSS(VSS),.VDD(VDD),.Y(I14807),.A(g8603));
  NOT NOT1_4828(.VSS(VSS),.VDD(VDD),.Y(g8671),.A(I14807));
  NOT NOT1_4829(.VSS(VSS),.VDD(VDD),.Y(I14810),.A(g8481));
  NOT NOT1_4830(.VSS(VSS),.VDD(VDD),.Y(g8672),.A(I14810));
  NOT NOT1_4831(.VSS(VSS),.VDD(VDD),.Y(I14813),.A(g8640));
  NOT NOT1_4832(.VSS(VSS),.VDD(VDD),.Y(g8673),.A(I14813));
  NOT NOT1_4833(.VSS(VSS),.VDD(VDD),.Y(I14816),.A(g8642));
  NOT NOT1_4834(.VSS(VSS),.VDD(VDD),.Y(g8674),.A(I14816));
  NOT NOT1_4835(.VSS(VSS),.VDD(VDD),.Y(I14819),.A(g8647));
  NOT NOT1_4836(.VSS(VSS),.VDD(VDD),.Y(g8675),.A(I14819));
  NOT NOT1_4837(.VSS(VSS),.VDD(VDD),.Y(I14822),.A(g8649));
  NOT NOT1_4838(.VSS(VSS),.VDD(VDD),.Y(g8676),.A(I14822));
  NOT NOT1_4839(.VSS(VSS),.VDD(VDD),.Y(I14825),.A(g8651));
  NOT NOT1_4840(.VSS(VSS),.VDD(VDD),.Y(g8677),.A(I14825));
  NOT NOT1_4841(.VSS(VSS),.VDD(VDD),.Y(I14828),.A(g8639));
  NOT NOT1_4842(.VSS(VSS),.VDD(VDD),.Y(g8678),.A(I14828));
  NOT NOT1_4843(.VSS(VSS),.VDD(VDD),.Y(I14844),.A(g8641));
  NOT NOT1_4844(.VSS(VSS),.VDD(VDD),.Y(g8682),.A(I14844));
  NOT NOT1_4845(.VSS(VSS),.VDD(VDD),.Y(g8683),.A(g8235));
  NOT NOT1_4846(.VSS(VSS),.VDD(VDD),.Y(I14848),.A(g8625));
  NOT NOT1_4847(.VSS(VSS),.VDD(VDD),.Y(g8684),.A(I14848));
  NOT NOT1_4848(.VSS(VSS),.VDD(VDD),.Y(I14851),.A(g8630));
  NOT NOT1_4849(.VSS(VSS),.VDD(VDD),.Y(g8685),.A(I14851));
  NOT NOT1_4850(.VSS(VSS),.VDD(VDD),.Y(I14857),.A(g8657));
  NOT NOT1_4851(.VSS(VSS),.VDD(VDD),.Y(g8689),.A(I14857));
  NOT NOT1_4852(.VSS(VSS),.VDD(VDD),.Y(I14904),.A(g8629));
  NOT NOT1_4853(.VSS(VSS),.VDD(VDD),.Y(g8734),.A(I14904));
  NOT NOT1_4854(.VSS(VSS),.VDD(VDD),.Y(g8743),.A(g8524));
  NOT NOT1_4855(.VSS(VSS),.VDD(VDD),.Y(g8746),.A(g8524));
  NOT NOT1_4856(.VSS(VSS),.VDD(VDD),.Y(g8747),.A(g8545));
  NOT NOT1_4857(.VSS(VSS),.VDD(VDD),.Y(g8750),.A(g8524));
  NOT NOT1_4858(.VSS(VSS),.VDD(VDD),.Y(g8751),.A(g8545));
  NOT NOT1_4859(.VSS(VSS),.VDD(VDD),.Y(g8752),.A(g8564));
  NOT NOT1_4860(.VSS(VSS),.VDD(VDD),.Y(I14925),.A(g8381));
  NOT NOT1_4861(.VSS(VSS),.VDD(VDD),.Y(g8753),.A(I14925));
  NOT NOT1_4862(.VSS(VSS),.VDD(VDD),.Y(g8754),.A(g8524));
  NOT NOT1_4863(.VSS(VSS),.VDD(VDD),.Y(g8755),.A(g8545));
  NOT NOT1_4864(.VSS(VSS),.VDD(VDD),.Y(g8756),.A(g8564));
  NOT NOT1_4865(.VSS(VSS),.VDD(VDD),.Y(g8757),.A(g8585));
  NOT NOT1_4866(.VSS(VSS),.VDD(VDD),.Y(g8759),.A(g8524));
  NOT NOT1_4867(.VSS(VSS),.VDD(VDD),.Y(g8760),.A(g8545));
  NOT NOT1_4868(.VSS(VSS),.VDD(VDD),.Y(g8761),.A(g8564));
  NOT NOT1_4869(.VSS(VSS),.VDD(VDD),.Y(g8762),.A(g8585));
  NOT NOT1_4870(.VSS(VSS),.VDD(VDD),.Y(g8765),.A(g8524));
  NOT NOT1_4871(.VSS(VSS),.VDD(VDD),.Y(g8766),.A(g8545));
  NOT NOT1_4872(.VSS(VSS),.VDD(VDD),.Y(g8767),.A(g8564));
  NOT NOT1_4873(.VSS(VSS),.VDD(VDD),.Y(g8768),.A(g8585));
  NOT NOT1_4874(.VSS(VSS),.VDD(VDD),.Y(g8770),.A(g8545));
  NOT NOT1_4875(.VSS(VSS),.VDD(VDD),.Y(g8771),.A(g8564));
  NOT NOT1_4876(.VSS(VSS),.VDD(VDD),.Y(g8772),.A(g8585));
  NOT NOT1_4877(.VSS(VSS),.VDD(VDD),.Y(I14964),.A(g8406));
  NOT NOT1_4878(.VSS(VSS),.VDD(VDD),.Y(g8774),.A(I14964));
  NOT NOT1_4879(.VSS(VSS),.VDD(VDD),.Y(g8775),.A(g8564));
  NOT NOT1_4880(.VSS(VSS),.VDD(VDD),.Y(g8776),.A(g8585));
  NOT NOT1_4881(.VSS(VSS),.VDD(VDD),.Y(I14974),.A(g8442));
  NOT NOT1_4882(.VSS(VSS),.VDD(VDD),.Y(g8778),.A(I14974));
  NOT NOT1_4883(.VSS(VSS),.VDD(VDD),.Y(g8780),.A(g8524));
  NOT NOT1_4884(.VSS(VSS),.VDD(VDD),.Y(g8781),.A(g8585));
  NOT NOT1_4885(.VSS(VSS),.VDD(VDD),.Y(g8783),.A(g8524));
  NOT NOT1_4886(.VSS(VSS),.VDD(VDD),.Y(g8784),.A(g8545));
  NOT NOT1_4887(.VSS(VSS),.VDD(VDD),.Y(g8786),.A(g8545));
  NOT NOT1_4888(.VSS(VSS),.VDD(VDD),.Y(g8787),.A(g8564));
  NOT NOT1_4889(.VSS(VSS),.VDD(VDD),.Y(g8789),.A(g8564));
  NOT NOT1_4890(.VSS(VSS),.VDD(VDD),.Y(g8790),.A(g8585));
  NOT NOT1_4891(.VSS(VSS),.VDD(VDD),.Y(g8791),.A(g8585));
  NOT NOT1_4892(.VSS(VSS),.VDD(VDD),.Y(I14996),.A(g8510));
  NOT NOT1_4893(.VSS(VSS),.VDD(VDD),.Y(g8792),.A(I14996));
  NOT NOT1_4894(.VSS(VSS),.VDD(VDD),.Y(I15003),.A(g8633));
  NOT NOT1_4895(.VSS(VSS),.VDD(VDD),.Y(g8797),.A(I15003));
  NOT NOT1_4896(.VSS(VSS),.VDD(VDD),.Y(I15007),.A(g8627));
  NOT NOT1_4897(.VSS(VSS),.VDD(VDD),.Y(g8799),.A(I15007));
  NOT NOT1_4898(.VSS(VSS),.VDD(VDD),.Y(I15010),.A(g8584));
  NOT NOT1_4899(.VSS(VSS),.VDD(VDD),.Y(g8800),.A(I15010));
  NOT NOT1_4900(.VSS(VSS),.VDD(VDD),.Y(I15014),.A(g8607));
  NOT NOT1_4901(.VSS(VSS),.VDD(VDD),.Y(g8802),.A(I15014));
  NOT NOT1_4902(.VSS(VSS),.VDD(VDD),.Y(I15062),.A(g8632));
  NOT NOT1_4903(.VSS(VSS),.VDD(VDD),.Y(g8808),.A(I15062));
  NOT NOT1_4904(.VSS(VSS),.VDD(VDD),.Y(I15065),.A(g8636));
  NOT NOT1_4905(.VSS(VSS),.VDD(VDD),.Y(g8809),.A(I15065));
  NOT NOT1_4906(.VSS(VSS),.VDD(VDD),.Y(I15068),.A(g8638));
  NOT NOT1_4907(.VSS(VSS),.VDD(VDD),.Y(g8810),.A(I15068));
  NOT NOT1_4908(.VSS(VSS),.VDD(VDD),.Y(I15160),.A(g8631));
  NOT NOT1_4909(.VSS(VSS),.VDD(VDD),.Y(g8856),.A(I15160));
  NOT NOT1_4910(.VSS(VSS),.VDD(VDD),.Y(I15178),.A(g8753));
  NOT NOT1_4911(.VSS(VSS),.VDD(VDD),.Y(g8864),.A(I15178));
  NOT NOT1_4912(.VSS(VSS),.VDD(VDD),.Y(I15181),.A(g8734));
  NOT NOT1_4913(.VSS(VSS),.VDD(VDD),.Y(g8865),.A(I15181));
  NOT NOT1_4914(.VSS(VSS),.VDD(VDD),.Y(I15184),.A(g8684));
  NOT NOT1_4915(.VSS(VSS),.VDD(VDD),.Y(g8866),.A(I15184));
  NOT NOT1_4916(.VSS(VSS),.VDD(VDD),.Y(I15187),.A(g8682));
  NOT NOT1_4917(.VSS(VSS),.VDD(VDD),.Y(g8867),.A(I15187));
  NOT NOT1_4918(.VSS(VSS),.VDD(VDD),.Y(I15190),.A(g8685));
  NOT NOT1_4919(.VSS(VSS),.VDD(VDD),.Y(g8868),.A(I15190));
  NOT NOT1_4920(.VSS(VSS),.VDD(VDD),.Y(I15193),.A(g8774));
  NOT NOT1_4921(.VSS(VSS),.VDD(VDD),.Y(g8869),.A(I15193));
  NOT NOT1_4922(.VSS(VSS),.VDD(VDD),.Y(I15196),.A(g8778));
  NOT NOT1_4923(.VSS(VSS),.VDD(VDD),.Y(g8870),.A(I15196));
  NOT NOT1_4924(.VSS(VSS),.VDD(VDD),.Y(I15199),.A(g8792));
  NOT NOT1_4925(.VSS(VSS),.VDD(VDD),.Y(g8871),.A(I15199));
  NOT NOT1_4926(.VSS(VSS),.VDD(VDD),.Y(I15202),.A(g8797));
  NOT NOT1_4927(.VSS(VSS),.VDD(VDD),.Y(g8872),.A(I15202));
  NOT NOT1_4928(.VSS(VSS),.VDD(VDD),.Y(I15205),.A(g8809));
  NOT NOT1_4929(.VSS(VSS),.VDD(VDD),.Y(g8873),.A(I15205));
  NOT NOT1_4930(.VSS(VSS),.VDD(VDD),.Y(I15208),.A(g8810));
  NOT NOT1_4931(.VSS(VSS),.VDD(VDD),.Y(g8874),.A(I15208));
  NOT NOT1_4932(.VSS(VSS),.VDD(VDD),.Y(I15211),.A(g8808));
  NOT NOT1_4933(.VSS(VSS),.VDD(VDD),.Y(g8875),.A(I15211));
  NOT NOT1_4934(.VSS(VSS),.VDD(VDD),.Y(I15218),.A(g8801));
  NOT NOT1_4935(.VSS(VSS),.VDD(VDD),.Y(g8880),.A(I15218));
  NOT NOT1_4936(.VSS(VSS),.VDD(VDD),.Y(g8881),.A(g8683));
  NOT NOT1_4937(.VSS(VSS),.VDD(VDD),.Y(I15222),.A(g8834));
  NOT NOT1_4938(.VSS(VSS),.VDD(VDD),.Y(g8882),.A(I15222));
  NOT NOT1_4939(.VSS(VSS),.VDD(VDD),.Y(I15225),.A(g8689));
  NOT NOT1_4940(.VSS(VSS),.VDD(VDD),.Y(g8883),.A(I15225));
  NOT NOT1_4941(.VSS(VSS),.VDD(VDD),.Y(I15308),.A(g8799));
  NOT NOT1_4942(.VSS(VSS),.VDD(VDD),.Y(g8898),.A(I15308));
  NOT NOT1_4943(.VSS(VSS),.VDD(VDD),.Y(I15315),.A(g8738));
  NOT NOT1_4944(.VSS(VSS),.VDD(VDD),.Y(g8903),.A(I15315));
  NOT NOT1_4945(.VSS(VSS),.VDD(VDD),.Y(I15324),.A(g8779));
  NOT NOT1_4946(.VSS(VSS),.VDD(VDD),.Y(g8910),.A(I15324));
  NOT NOT1_4947(.VSS(VSS),.VDD(VDD),.Y(I15329),.A(g8793));
  NOT NOT1_4948(.VSS(VSS),.VDD(VDD),.Y(g8913),.A(I15329));
  NOT NOT1_4949(.VSS(VSS),.VDD(VDD),.Y(I15334),.A(g8800));
  NOT NOT1_4950(.VSS(VSS),.VDD(VDD),.Y(g8916),.A(I15334));
  NOT NOT1_4951(.VSS(VSS),.VDD(VDD),.Y(I15337),.A(g8802));
  NOT NOT1_4952(.VSS(VSS),.VDD(VDD),.Y(g8917),.A(I15337));
  NOT NOT1_4953(.VSS(VSS),.VDD(VDD),.Y(I15340),.A(g8856));
  NOT NOT1_4954(.VSS(VSS),.VDD(VDD),.Y(g8918),.A(I15340));
  NOT NOT1_4955(.VSS(VSS),.VDD(VDD),.Y(I15379),.A(g8882));
  NOT NOT1_4956(.VSS(VSS),.VDD(VDD),.Y(g8955),.A(I15379));
  NOT NOT1_4957(.VSS(VSS),.VDD(VDD),.Y(I15382),.A(g8883));
  NOT NOT1_4958(.VSS(VSS),.VDD(VDD),.Y(g8956),.A(I15382));
  NOT NOT1_4959(.VSS(VSS),.VDD(VDD),.Y(I15385),.A(g8880));
  NOT NOT1_4960(.VSS(VSS),.VDD(VDD),.Y(g8957),.A(I15385));
  NOT NOT1_4961(.VSS(VSS),.VDD(VDD),.Y(I15388),.A(g8898));
  NOT NOT1_4962(.VSS(VSS),.VDD(VDD),.Y(g8958),.A(I15388));
  NOT NOT1_4963(.VSS(VSS),.VDD(VDD),.Y(I15391),.A(g8917));
  NOT NOT1_4964(.VSS(VSS),.VDD(VDD),.Y(g8959),.A(I15391));
  NOT NOT1_4965(.VSS(VSS),.VDD(VDD),.Y(I15394),.A(g8916));
  NOT NOT1_4966(.VSS(VSS),.VDD(VDD),.Y(g8960),.A(I15394));
  NOT NOT1_4967(.VSS(VSS),.VDD(VDD),.Y(I15405),.A(g8902));
  NOT NOT1_4968(.VSS(VSS),.VDD(VDD),.Y(g8967),.A(I15405));
  NOT NOT1_4969(.VSS(VSS),.VDD(VDD),.Y(I15408),.A(g8896));
  NOT NOT1_4970(.VSS(VSS),.VDD(VDD),.Y(g8968),.A(I15408));
  NOT NOT1_4971(.VSS(VSS),.VDD(VDD),.Y(I15411),.A(g8897));
  NOT NOT1_4972(.VSS(VSS),.VDD(VDD),.Y(g8969),.A(I15411));
  NOT NOT1_4973(.VSS(VSS),.VDD(VDD),.Y(I15414),.A(g8900));
  NOT NOT1_4974(.VSS(VSS),.VDD(VDD),.Y(g8970),.A(I15414));
  NOT NOT1_4975(.VSS(VSS),.VDD(VDD),.Y(I15417),.A(g8893));
  NOT NOT1_4976(.VSS(VSS),.VDD(VDD),.Y(g8971),.A(I15417));
  NOT NOT1_4977(.VSS(VSS),.VDD(VDD),.Y(I15420),.A(g8881));
  NOT NOT1_4978(.VSS(VSS),.VDD(VDD),.Y(g8972),.A(I15420));
  NOT NOT1_4979(.VSS(VSS),.VDD(VDD),.Y(I15423),.A(g8894));
  NOT NOT1_4980(.VSS(VSS),.VDD(VDD),.Y(g8973),.A(I15423));
  NOT NOT1_4981(.VSS(VSS),.VDD(VDD),.Y(I15426),.A(g8895));
  NOT NOT1_4982(.VSS(VSS),.VDD(VDD),.Y(g8974),.A(I15426));
  NOT NOT1_4983(.VSS(VSS),.VDD(VDD),.Y(I15429),.A(g8899));
  NOT NOT1_4984(.VSS(VSS),.VDD(VDD),.Y(g8975),.A(I15429));
  NOT NOT1_4985(.VSS(VSS),.VDD(VDD),.Y(I15433),.A(g8911));
  NOT NOT1_4986(.VSS(VSS),.VDD(VDD),.Y(g8977),.A(I15433));
  NOT NOT1_4987(.VSS(VSS),.VDD(VDD),.Y(I15475),.A(g8901));
  NOT NOT1_4988(.VSS(VSS),.VDD(VDD),.Y(g9017),.A(I15475));
  NOT NOT1_4989(.VSS(VSS),.VDD(VDD),.Y(I15478),.A(g8910));
  NOT NOT1_4990(.VSS(VSS),.VDD(VDD),.Y(g9018),.A(I15478));
  NOT NOT1_4991(.VSS(VSS),.VDD(VDD),.Y(I15481),.A(g8913));
  NOT NOT1_4992(.VSS(VSS),.VDD(VDD),.Y(g9019),.A(I15481));
  NOT NOT1_4993(.VSS(VSS),.VDD(VDD),.Y(I15484),.A(g8918));
  NOT NOT1_4994(.VSS(VSS),.VDD(VDD),.Y(g9020),.A(I15484));
  NOT NOT1_4995(.VSS(VSS),.VDD(VDD),.Y(I15492),.A(g8971));
  NOT NOT1_4996(.VSS(VSS),.VDD(VDD),.Y(g9026),.A(I15492));
  NOT NOT1_4997(.VSS(VSS),.VDD(VDD),.Y(I15495),.A(g8973));
  NOT NOT1_4998(.VSS(VSS),.VDD(VDD),.Y(g9027),.A(I15495));
  NOT NOT1_4999(.VSS(VSS),.VDD(VDD),.Y(I15498),.A(g8974));
  NOT NOT1_5000(.VSS(VSS),.VDD(VDD),.Y(g9028),.A(I15498));
  NOT NOT1_5001(.VSS(VSS),.VDD(VDD),.Y(I15501),.A(g8975));
  NOT NOT1_5002(.VSS(VSS),.VDD(VDD),.Y(g9029),.A(I15501));
  NOT NOT1_5003(.VSS(VSS),.VDD(VDD),.Y(I15504),.A(g8967));
  NOT NOT1_5004(.VSS(VSS),.VDD(VDD),.Y(g9030),.A(I15504));
  NOT NOT1_5005(.VSS(VSS),.VDD(VDD),.Y(I15507),.A(g8968));
  NOT NOT1_5006(.VSS(VSS),.VDD(VDD),.Y(g9031),.A(I15507));
  NOT NOT1_5007(.VSS(VSS),.VDD(VDD),.Y(I15510),.A(g8969));
  NOT NOT1_5008(.VSS(VSS),.VDD(VDD),.Y(g9032),.A(I15510));
  NOT NOT1_5009(.VSS(VSS),.VDD(VDD),.Y(I15513),.A(g8970));
  NOT NOT1_5010(.VSS(VSS),.VDD(VDD),.Y(g9033),.A(I15513));
  NOT NOT1_5011(.VSS(VSS),.VDD(VDD),.Y(I15516),.A(g8977));
  NOT NOT1_5012(.VSS(VSS),.VDD(VDD),.Y(g9034),.A(I15516));
  NOT NOT1_5013(.VSS(VSS),.VDD(VDD),.Y(I15519),.A(g9019));
  NOT NOT1_5014(.VSS(VSS),.VDD(VDD),.Y(g9035),.A(I15519));
  NOT NOT1_5015(.VSS(VSS),.VDD(VDD),.Y(I15522),.A(g9018));
  NOT NOT1_5016(.VSS(VSS),.VDD(VDD),.Y(g9036),.A(I15522));
  NOT NOT1_5017(.VSS(VSS),.VDD(VDD),.Y(I15527),.A(g9020));
  NOT NOT1_5018(.VSS(VSS),.VDD(VDD),.Y(g9039),.A(I15527));
  NOT NOT1_5019(.VSS(VSS),.VDD(VDD),.Y(I15530),.A(g8972));
  NOT NOT1_5020(.VSS(VSS),.VDD(VDD),.Y(g9042),.A(I15530));
  NOT NOT1_5021(.VSS(VSS),.VDD(VDD),.Y(I15533),.A(g9002));
  NOT NOT1_5022(.VSS(VSS),.VDD(VDD),.Y(g9043),.A(I15533));
  NOT NOT1_5023(.VSS(VSS),.VDD(VDD),.Y(I15536),.A(g9004));
  NOT NOT1_5024(.VSS(VSS),.VDD(VDD),.Y(g9044),.A(I15536));
  NOT NOT1_5025(.VSS(VSS),.VDD(VDD),.Y(I15539),.A(g9005));
  NOT NOT1_5026(.VSS(VSS),.VDD(VDD),.Y(g9045),.A(I15539));
  NOT NOT1_5027(.VSS(VSS),.VDD(VDD),.Y(I15543),.A(g9006));
  NOT NOT1_5028(.VSS(VSS),.VDD(VDD),.Y(g9047),.A(I15543));
  NOT NOT1_5029(.VSS(VSS),.VDD(VDD),.Y(I15546),.A(g9007));
  NOT NOT1_5030(.VSS(VSS),.VDD(VDD),.Y(g9048),.A(I15546));
  NOT NOT1_5031(.VSS(VSS),.VDD(VDD),.Y(I15550),.A(g9008));
  NOT NOT1_5032(.VSS(VSS),.VDD(VDD),.Y(g9050),.A(I15550));
  NOT NOT1_5033(.VSS(VSS),.VDD(VDD),.Y(I15553),.A(g9009));
  NOT NOT1_5034(.VSS(VSS),.VDD(VDD),.Y(g9051),.A(I15553));
  NOT NOT1_5035(.VSS(VSS),.VDD(VDD),.Y(I15557),.A(g9010));
  NOT NOT1_5036(.VSS(VSS),.VDD(VDD),.Y(g9053),.A(I15557));
  NOT NOT1_5037(.VSS(VSS),.VDD(VDD),.Y(I15562),.A(g8979));
  NOT NOT1_5038(.VSS(VSS),.VDD(VDD),.Y(g9056),.A(I15562));
  NOT NOT1_5039(.VSS(VSS),.VDD(VDD),.Y(I15565),.A(g8980));
  NOT NOT1_5040(.VSS(VSS),.VDD(VDD),.Y(g9057),.A(I15565));
  NOT NOT1_5041(.VSS(VSS),.VDD(VDD),.Y(I15568),.A(g8981));
  NOT NOT1_5042(.VSS(VSS),.VDD(VDD),.Y(g9058),.A(I15568));
  NOT NOT1_5043(.VSS(VSS),.VDD(VDD),.Y(I15571),.A(g8982));
  NOT NOT1_5044(.VSS(VSS),.VDD(VDD),.Y(g9059),.A(I15571));
  NOT NOT1_5045(.VSS(VSS),.VDD(VDD),.Y(I15574),.A(g8983));
  NOT NOT1_5046(.VSS(VSS),.VDD(VDD),.Y(g9060),.A(I15574));
  NOT NOT1_5047(.VSS(VSS),.VDD(VDD),.Y(I15577),.A(g8984));
  NOT NOT1_5048(.VSS(VSS),.VDD(VDD),.Y(g9061),.A(I15577));
  NOT NOT1_5049(.VSS(VSS),.VDD(VDD),.Y(I15580),.A(g8985));
  NOT NOT1_5050(.VSS(VSS),.VDD(VDD),.Y(g9062),.A(I15580));
  NOT NOT1_5051(.VSS(VSS),.VDD(VDD),.Y(I15583),.A(g8986));
  NOT NOT1_5052(.VSS(VSS),.VDD(VDD),.Y(g9063),.A(I15583));
  NOT NOT1_5053(.VSS(VSS),.VDD(VDD),.Y(I15586),.A(g8987));
  NOT NOT1_5054(.VSS(VSS),.VDD(VDD),.Y(g9064),.A(I15586));
  NOT NOT1_5055(.VSS(VSS),.VDD(VDD),.Y(I15589),.A(g8988));
  NOT NOT1_5056(.VSS(VSS),.VDD(VDD),.Y(g9065),.A(I15589));
  NOT NOT1_5057(.VSS(VSS),.VDD(VDD),.Y(I15592),.A(g8989));
  NOT NOT1_5058(.VSS(VSS),.VDD(VDD),.Y(g9066),.A(I15592));
  NOT NOT1_5059(.VSS(VSS),.VDD(VDD),.Y(I15595),.A(g8990));
  NOT NOT1_5060(.VSS(VSS),.VDD(VDD),.Y(g9067),.A(I15595));
  NOT NOT1_5061(.VSS(VSS),.VDD(VDD),.Y(I15598),.A(g8991));
  NOT NOT1_5062(.VSS(VSS),.VDD(VDD),.Y(g9068),.A(I15598));
  NOT NOT1_5063(.VSS(VSS),.VDD(VDD),.Y(I15601),.A(g8992));
  NOT NOT1_5064(.VSS(VSS),.VDD(VDD),.Y(g9069),.A(I15601));
  NOT NOT1_5065(.VSS(VSS),.VDD(VDD),.Y(I15604),.A(g8993));
  NOT NOT1_5066(.VSS(VSS),.VDD(VDD),.Y(g9070),.A(I15604));
  NOT NOT1_5067(.VSS(VSS),.VDD(VDD),.Y(I15607),.A(g8994));
  NOT NOT1_5068(.VSS(VSS),.VDD(VDD),.Y(g9071),.A(I15607));
  NOT NOT1_5069(.VSS(VSS),.VDD(VDD),.Y(I15610),.A(g8995));
  NOT NOT1_5070(.VSS(VSS),.VDD(VDD),.Y(g9072),.A(I15610));
  NOT NOT1_5071(.VSS(VSS),.VDD(VDD),.Y(I15613),.A(g8996));
  NOT NOT1_5072(.VSS(VSS),.VDD(VDD),.Y(g9073),.A(I15613));
  NOT NOT1_5073(.VSS(VSS),.VDD(VDD),.Y(I15616),.A(g8997));
  NOT NOT1_5074(.VSS(VSS),.VDD(VDD),.Y(g9074),.A(I15616));
  NOT NOT1_5075(.VSS(VSS),.VDD(VDD),.Y(I15619),.A(g8998));
  NOT NOT1_5076(.VSS(VSS),.VDD(VDD),.Y(g9075),.A(I15619));
  NOT NOT1_5077(.VSS(VSS),.VDD(VDD),.Y(I15622),.A(g8999));
  NOT NOT1_5078(.VSS(VSS),.VDD(VDD),.Y(g9076),.A(I15622));
  NOT NOT1_5079(.VSS(VSS),.VDD(VDD),.Y(I15625),.A(g9000));
  NOT NOT1_5080(.VSS(VSS),.VDD(VDD),.Y(g9077),.A(I15625));
  NOT NOT1_5081(.VSS(VSS),.VDD(VDD),.Y(I15628),.A(g9001));
  NOT NOT1_5082(.VSS(VSS),.VDD(VDD),.Y(g9078),.A(I15628));
  NOT NOT1_5083(.VSS(VSS),.VDD(VDD),.Y(I15631),.A(g9003));
  NOT NOT1_5084(.VSS(VSS),.VDD(VDD),.Y(g9079),.A(I15631));
  NOT NOT1_5085(.VSS(VSS),.VDD(VDD),.Y(I15635),.A(g8976));
  NOT NOT1_5086(.VSS(VSS),.VDD(VDD),.Y(g9081),.A(I15635));
  NOT NOT1_5087(.VSS(VSS),.VDD(VDD),.Y(I15638),.A(g8978));
  NOT NOT1_5088(.VSS(VSS),.VDD(VDD),.Y(g9082),.A(I15638));
  NOT NOT1_5089(.VSS(VSS),.VDD(VDD),.Y(I15641),.A(g9017));
  NOT NOT1_5090(.VSS(VSS),.VDD(VDD),.Y(g9083),.A(I15641));
  NOT NOT1_5091(.VSS(VSS),.VDD(VDD),.Y(I15645),.A(g9043));
  NOT NOT1_5092(.VSS(VSS),.VDD(VDD),.Y(g9085),.A(I15645));
  NOT NOT1_5093(.VSS(VSS),.VDD(VDD),.Y(I15648),.A(g9044));
  NOT NOT1_5094(.VSS(VSS),.VDD(VDD),.Y(g9086),.A(I15648));
  NOT NOT1_5095(.VSS(VSS),.VDD(VDD),.Y(I15651),.A(g9056));
  NOT NOT1_5096(.VSS(VSS),.VDD(VDD),.Y(g9087),.A(I15651));
  NOT NOT1_5097(.VSS(VSS),.VDD(VDD),.Y(I15654),.A(g9057));
  NOT NOT1_5098(.VSS(VSS),.VDD(VDD),.Y(g9088),.A(I15654));
  NOT NOT1_5099(.VSS(VSS),.VDD(VDD),.Y(I15657),.A(g9059));
  NOT NOT1_5100(.VSS(VSS),.VDD(VDD),.Y(g9089),.A(I15657));
  NOT NOT1_5101(.VSS(VSS),.VDD(VDD),.Y(I15660),.A(g9062));
  NOT NOT1_5102(.VSS(VSS),.VDD(VDD),.Y(g9090),.A(I15660));
  NOT NOT1_5103(.VSS(VSS),.VDD(VDD),.Y(I15663),.A(g9066));
  NOT NOT1_5104(.VSS(VSS),.VDD(VDD),.Y(g9091),.A(I15663));
  NOT NOT1_5105(.VSS(VSS),.VDD(VDD),.Y(I15666),.A(g9070));
  NOT NOT1_5106(.VSS(VSS),.VDD(VDD),.Y(g9092),.A(I15666));
  NOT NOT1_5107(.VSS(VSS),.VDD(VDD),.Y(I15669),.A(g9045));
  NOT NOT1_5108(.VSS(VSS),.VDD(VDD),.Y(g9093),.A(I15669));
  NOT NOT1_5109(.VSS(VSS),.VDD(VDD),.Y(I15672),.A(g9047));
  NOT NOT1_5110(.VSS(VSS),.VDD(VDD),.Y(g9094),.A(I15672));
  NOT NOT1_5111(.VSS(VSS),.VDD(VDD),.Y(I15675),.A(g9058));
  NOT NOT1_5112(.VSS(VSS),.VDD(VDD),.Y(g9095),.A(I15675));
  NOT NOT1_5113(.VSS(VSS),.VDD(VDD),.Y(I15678),.A(g9060));
  NOT NOT1_5114(.VSS(VSS),.VDD(VDD),.Y(g9096),.A(I15678));
  NOT NOT1_5115(.VSS(VSS),.VDD(VDD),.Y(I15681),.A(g9063));
  NOT NOT1_5116(.VSS(VSS),.VDD(VDD),.Y(g9097),.A(I15681));
  NOT NOT1_5117(.VSS(VSS),.VDD(VDD),.Y(I15684),.A(g9067));
  NOT NOT1_5118(.VSS(VSS),.VDD(VDD),.Y(g9098),.A(I15684));
  NOT NOT1_5119(.VSS(VSS),.VDD(VDD),.Y(I15687),.A(g9071));
  NOT NOT1_5120(.VSS(VSS),.VDD(VDD),.Y(g9099),.A(I15687));
  NOT NOT1_5121(.VSS(VSS),.VDD(VDD),.Y(I15690),.A(g9074));
  NOT NOT1_5122(.VSS(VSS),.VDD(VDD),.Y(g9100),.A(I15690));
  NOT NOT1_5123(.VSS(VSS),.VDD(VDD),.Y(I15693),.A(g9048));
  NOT NOT1_5124(.VSS(VSS),.VDD(VDD),.Y(g9101),.A(I15693));
  NOT NOT1_5125(.VSS(VSS),.VDD(VDD),.Y(I15696),.A(g9050));
  NOT NOT1_5126(.VSS(VSS),.VDD(VDD),.Y(g9102),.A(I15696));
  NOT NOT1_5127(.VSS(VSS),.VDD(VDD),.Y(I15699),.A(g9061));
  NOT NOT1_5128(.VSS(VSS),.VDD(VDD),.Y(g9103),.A(I15699));
  NOT NOT1_5129(.VSS(VSS),.VDD(VDD),.Y(I15702),.A(g9064));
  NOT NOT1_5130(.VSS(VSS),.VDD(VDD),.Y(g9104),.A(I15702));
  NOT NOT1_5131(.VSS(VSS),.VDD(VDD),.Y(I15705),.A(g9068));
  NOT NOT1_5132(.VSS(VSS),.VDD(VDD),.Y(g9105),.A(I15705));
  NOT NOT1_5133(.VSS(VSS),.VDD(VDD),.Y(I15708),.A(g9072));
  NOT NOT1_5134(.VSS(VSS),.VDD(VDD),.Y(g9106),.A(I15708));
  NOT NOT1_5135(.VSS(VSS),.VDD(VDD),.Y(I15711),.A(g9075));
  NOT NOT1_5136(.VSS(VSS),.VDD(VDD),.Y(g9107),.A(I15711));
  NOT NOT1_5137(.VSS(VSS),.VDD(VDD),.Y(I15714),.A(g9077));
  NOT NOT1_5138(.VSS(VSS),.VDD(VDD),.Y(g9108),.A(I15714));
  NOT NOT1_5139(.VSS(VSS),.VDD(VDD),.Y(I15717),.A(g9051));
  NOT NOT1_5140(.VSS(VSS),.VDD(VDD),.Y(g9109),.A(I15717));
  NOT NOT1_5141(.VSS(VSS),.VDD(VDD),.Y(I15720),.A(g9053));
  NOT NOT1_5142(.VSS(VSS),.VDD(VDD),.Y(g9110),.A(I15720));
  NOT NOT1_5143(.VSS(VSS),.VDD(VDD),.Y(I15723),.A(g9065));
  NOT NOT1_5144(.VSS(VSS),.VDD(VDD),.Y(g9111),.A(I15723));
  NOT NOT1_5145(.VSS(VSS),.VDD(VDD),.Y(I15726),.A(g9069));
  NOT NOT1_5146(.VSS(VSS),.VDD(VDD),.Y(g9112),.A(I15726));
  NOT NOT1_5147(.VSS(VSS),.VDD(VDD),.Y(I15729),.A(g9073));
  NOT NOT1_5148(.VSS(VSS),.VDD(VDD),.Y(g9113),.A(I15729));
  NOT NOT1_5149(.VSS(VSS),.VDD(VDD),.Y(I15732),.A(g9076));
  NOT NOT1_5150(.VSS(VSS),.VDD(VDD),.Y(g9114),.A(I15732));
  NOT NOT1_5151(.VSS(VSS),.VDD(VDD),.Y(I15735),.A(g9078));
  NOT NOT1_5152(.VSS(VSS),.VDD(VDD),.Y(g9115),.A(I15735));
  NOT NOT1_5153(.VSS(VSS),.VDD(VDD),.Y(I15738),.A(g9079));
  NOT NOT1_5154(.VSS(VSS),.VDD(VDD),.Y(g9116),.A(I15738));
  NOT NOT1_5155(.VSS(VSS),.VDD(VDD),.Y(I15741),.A(g9083));
  NOT NOT1_5156(.VSS(VSS),.VDD(VDD),.Y(g9117),.A(I15741));
  NOT NOT1_5157(.VSS(VSS),.VDD(VDD),.Y(I15747),.A(g9042));
  NOT NOT1_5158(.VSS(VSS),.VDD(VDD),.Y(g9121),.A(I15747));
  NOT NOT1_5159(.VSS(VSS),.VDD(VDD),.Y(I15753),.A(g9080));
  NOT NOT1_5160(.VSS(VSS),.VDD(VDD),.Y(g9125),.A(I15753));
  NOT NOT1_5161(.VSS(VSS),.VDD(VDD),.Y(I15756),.A(g9081));
  NOT NOT1_5162(.VSS(VSS),.VDD(VDD),.Y(g9126),.A(I15756));
  NOT NOT1_5163(.VSS(VSS),.VDD(VDD),.Y(I15759),.A(g9082));
  NOT NOT1_5164(.VSS(VSS),.VDD(VDD),.Y(g9127),.A(I15759));
  NOT NOT1_5165(.VSS(VSS),.VDD(VDD),.Y(I15762),.A(g9039));
  NOT NOT1_5166(.VSS(VSS),.VDD(VDD),.Y(g9128),.A(I15762));
  NOT NOT1_5167(.VSS(VSS),.VDD(VDD),.Y(I15765),.A(g9039));
  NOT NOT1_5168(.VSS(VSS),.VDD(VDD),.Y(g9129),.A(I15765));
  NOT NOT1_5169(.VSS(VSS),.VDD(VDD),.Y(I15770),.A(g9121));
  NOT NOT1_5170(.VSS(VSS),.VDD(VDD),.Y(g9132),.A(I15770));
  NOT NOT1_5171(.VSS(VSS),.VDD(VDD),.Y(I15773),.A(g9126));
  NOT NOT1_5172(.VSS(VSS),.VDD(VDD),.Y(g9133),.A(I15773));
  NOT NOT1_5173(.VSS(VSS),.VDD(VDD),.Y(I15776),.A(g9127));
  NOT NOT1_5174(.VSS(VSS),.VDD(VDD),.Y(g9134),.A(I15776));
  NOT NOT1_5175(.VSS(VSS),.VDD(VDD),.Y(I15784),.A(g9125));
  NOT NOT1_5176(.VSS(VSS),.VDD(VDD),.Y(g9140),.A(I15784));
  NOT NOT1_5177(.VSS(VSS),.VDD(VDD),.Y(g9141),.A(g9129));
  NOT NOT1_5178(.VSS(VSS),.VDD(VDD),.Y(I15791),.A(g9140));
  NOT NOT1_5179(.VSS(VSS),.VDD(VDD),.Y(g9145),.A(I15791));
  NOT NOT1_5180(.VSS(VSS),.VDD(VDD),.Y(g9157),.A(g9141));
  NOT NOT1_5181(.VSS(VSS),.VDD(VDD),.Y(I15803),.A(g9148));
  NOT NOT1_5182(.VSS(VSS),.VDD(VDD),.Y(g9161),.A(I15803));
  NOT NOT1_5183(.VSS(VSS),.VDD(VDD),.Y(I15811),.A(g9151));
  NOT NOT1_5184(.VSS(VSS),.VDD(VDD),.Y(g9177),.A(I15811));
  NOT NOT1_5185(.VSS(VSS),.VDD(VDD),.Y(I15814),.A(g9154));
  NOT NOT1_5186(.VSS(VSS),.VDD(VDD),.Y(g9178),.A(I15814));
  NOT NOT1_5187(.VSS(VSS),.VDD(VDD),.Y(I15824),.A(g9157));
  NOT NOT1_5188(.VSS(VSS),.VDD(VDD),.Y(g9180),.A(I15824));
  NOT NOT1_5189(.VSS(VSS),.VDD(VDD),.Y(g9181),.A(g9177));
  NOT NOT1_5190(.VSS(VSS),.VDD(VDD),.Y(g9182),.A(g9178));
  NOT NOT1_5191(.VSS(VSS),.VDD(VDD),.Y(g9183),.A(g9161));
  NOT NOT1_5192(.VSS(VSS),.VDD(VDD),.Y(I15830),.A(g9180));
  NOT NOT1_5193(.VSS(VSS),.VDD(VDD),.Y(g9184),.A(I15830));
  NOT NOT1_5194(.VSS(VSS),.VDD(VDD),.Y(I15833),.A(g9162));
  NOT NOT1_5195(.VSS(VSS),.VDD(VDD),.Y(g9185),.A(I15833));
  NOT NOT1_5196(.VSS(VSS),.VDD(VDD),.Y(I15836),.A(g9165));
  NOT NOT1_5197(.VSS(VSS),.VDD(VDD),.Y(g9186),.A(I15836));
  NOT NOT1_5198(.VSS(VSS),.VDD(VDD),.Y(I15839),.A(g9168));
  NOT NOT1_5199(.VSS(VSS),.VDD(VDD),.Y(g9187),.A(I15839));
  NOT NOT1_5200(.VSS(VSS),.VDD(VDD),.Y(I15842),.A(g9171));
  NOT NOT1_5201(.VSS(VSS),.VDD(VDD),.Y(g9188),.A(I15842));
  NOT NOT1_5202(.VSS(VSS),.VDD(VDD),.Y(I15845),.A(g9174));
  NOT NOT1_5203(.VSS(VSS),.VDD(VDD),.Y(g9189),.A(I15845));
  NOT NOT1_5204(.VSS(VSS),.VDD(VDD),.Y(g9193),.A(g9181));
  NOT NOT1_5205(.VSS(VSS),.VDD(VDD),.Y(g9194),.A(g9182));
  NOT NOT1_5206(.VSS(VSS),.VDD(VDD),.Y(I15871),.A(g9184));
  NOT NOT1_5207(.VSS(VSS),.VDD(VDD),.Y(g9195),.A(I15871));
  NOT NOT1_5208(.VSS(VSS),.VDD(VDD),.Y(g9196),.A(g9185));
  NOT NOT1_5209(.VSS(VSS),.VDD(VDD),.Y(g9197),.A(g9186));
  NOT NOT1_5210(.VSS(VSS),.VDD(VDD),.Y(g9198),.A(g9187));
  NOT NOT1_5211(.VSS(VSS),.VDD(VDD),.Y(g9199),.A(g9188));
  NOT NOT1_5212(.VSS(VSS),.VDD(VDD),.Y(g9200),.A(g9189));
  NOT NOT1_5213(.VSS(VSS),.VDD(VDD),.Y(g9201),.A(g9183));
  NOT NOT1_5214(.VSS(VSS),.VDD(VDD),.Y(I15894),.A(g9195));
  NOT NOT1_5215(.VSS(VSS),.VDD(VDD),.Y(g9204),.A(I15894));
  NOT NOT1_5216(.VSS(VSS),.VDD(VDD),.Y(g9206),.A(g9196));
  NOT NOT1_5217(.VSS(VSS),.VDD(VDD),.Y(g9207),.A(g9197));
  NOT NOT1_5218(.VSS(VSS),.VDD(VDD),.Y(g9208),.A(g9198));
  NOT NOT1_5219(.VSS(VSS),.VDD(VDD),.Y(g9209),.A(g9199));
  NOT NOT1_5220(.VSS(VSS),.VDD(VDD),.Y(g9210),.A(g9200));
  NOT NOT1_5221(.VSS(VSS),.VDD(VDD),.Y(I15909),.A(g9201));
  NOT NOT1_5222(.VSS(VSS),.VDD(VDD),.Y(g9211),.A(I15909));
  NOT NOT1_5223(.VSS(VSS),.VDD(VDD),.Y(I15912),.A(g9193));
  NOT NOT1_5224(.VSS(VSS),.VDD(VDD),.Y(g9212),.A(I15912));
  NOT NOT1_5225(.VSS(VSS),.VDD(VDD),.Y(I15915),.A(g9194));
  NOT NOT1_5226(.VSS(VSS),.VDD(VDD),.Y(g9213),.A(I15915));
  NOT NOT1_5227(.VSS(VSS),.VDD(VDD),.Y(I15918),.A(g9211));
  NOT NOT1_5228(.VSS(VSS),.VDD(VDD),.Y(g9214),.A(I15918));
  NOT NOT1_5229(.VSS(VSS),.VDD(VDD),.Y(I15921),.A(g9206));
  NOT NOT1_5230(.VSS(VSS),.VDD(VDD),.Y(g9215),.A(I15921));
  NOT NOT1_5231(.VSS(VSS),.VDD(VDD),.Y(I15924),.A(g9207));
  NOT NOT1_5232(.VSS(VSS),.VDD(VDD),.Y(g9216),.A(I15924));
  NOT NOT1_5233(.VSS(VSS),.VDD(VDD),.Y(I15927),.A(g9208));
  NOT NOT1_5234(.VSS(VSS),.VDD(VDD),.Y(g9217),.A(I15927));
  NOT NOT1_5235(.VSS(VSS),.VDD(VDD),.Y(I15930),.A(g9209));
  NOT NOT1_5236(.VSS(VSS),.VDD(VDD),.Y(g9218),.A(I15930));
  NOT NOT1_5237(.VSS(VSS),.VDD(VDD),.Y(I15933),.A(g9210));
  NOT NOT1_5238(.VSS(VSS),.VDD(VDD),.Y(g9219),.A(I15933));
  NOT NOT1_5239(.VSS(VSS),.VDD(VDD),.Y(g9220),.A(g9205));
  NOT NOT1_5240(.VSS(VSS),.VDD(VDD),.Y(I15937),.A(g9212));
  NOT NOT1_5241(.VSS(VSS),.VDD(VDD),.Y(g9221),.A(I15937));
  NOT NOT1_5242(.VSS(VSS),.VDD(VDD),.Y(I15940),.A(g9213));
  NOT NOT1_5243(.VSS(VSS),.VDD(VDD),.Y(g9222),.A(I15940));
  NOT NOT1_5244(.VSS(VSS),.VDD(VDD),.Y(I15943),.A(g9214));
  NOT NOT1_5245(.VSS(VSS),.VDD(VDD),.Y(g9223),.A(I15943));
  NOT NOT1_5246(.VSS(VSS),.VDD(VDD),.Y(I15947),.A(g9221));
  NOT NOT1_5247(.VSS(VSS),.VDD(VDD),.Y(g9227),.A(I15947));
  NOT NOT1_5248(.VSS(VSS),.VDD(VDD),.Y(I15950),.A(g9222));
  NOT NOT1_5249(.VSS(VSS),.VDD(VDD),.Y(g9230),.A(I15950));
  NOT NOT1_5250(.VSS(VSS),.VDD(VDD),.Y(I15953),.A(g9215));
  NOT NOT1_5251(.VSS(VSS),.VDD(VDD),.Y(g9233),.A(I15953));
  NOT NOT1_5252(.VSS(VSS),.VDD(VDD),.Y(I15956),.A(g9216));
  NOT NOT1_5253(.VSS(VSS),.VDD(VDD),.Y(g9234),.A(I15956));
  NOT NOT1_5254(.VSS(VSS),.VDD(VDD),.Y(I15959),.A(g9217));
  NOT NOT1_5255(.VSS(VSS),.VDD(VDD),.Y(g9235),.A(I15959));
  NOT NOT1_5256(.VSS(VSS),.VDD(VDD),.Y(I15962),.A(g9218));
  NOT NOT1_5257(.VSS(VSS),.VDD(VDD),.Y(g9236),.A(I15962));
  NOT NOT1_5258(.VSS(VSS),.VDD(VDD),.Y(I15965),.A(g9219));
  NOT NOT1_5259(.VSS(VSS),.VDD(VDD),.Y(g9237),.A(I15965));
  NOT NOT1_5260(.VSS(VSS),.VDD(VDD),.Y(I15971),.A(g9233));
  NOT NOT1_5261(.VSS(VSS),.VDD(VDD),.Y(g9241),.A(I15971));
  NOT NOT1_5262(.VSS(VSS),.VDD(VDD),.Y(I15974),.A(g9234));
  NOT NOT1_5263(.VSS(VSS),.VDD(VDD),.Y(g9244),.A(I15974));
  NOT NOT1_5264(.VSS(VSS),.VDD(VDD),.Y(I15978),.A(g9235));
  NOT NOT1_5265(.VSS(VSS),.VDD(VDD),.Y(g9248),.A(I15978));
  NOT NOT1_5266(.VSS(VSS),.VDD(VDD),.Y(I15982),.A(g9236));
  NOT NOT1_5267(.VSS(VSS),.VDD(VDD),.Y(g9252),.A(I15982));
  NOT NOT1_5268(.VSS(VSS),.VDD(VDD),.Y(I15985),.A(g9237));
  NOT NOT1_5269(.VSS(VSS),.VDD(VDD),.Y(g9255),.A(I15985));
  NOT NOT1_5270(.VSS(VSS),.VDD(VDD),.Y(I15990),.A(g9239));
  NOT NOT1_5271(.VSS(VSS),.VDD(VDD),.Y(g9260),.A(I15990));
  NOT NOT1_5272(.VSS(VSS),.VDD(VDD),.Y(I16006),.A(g9261));
  NOT NOT1_5273(.VSS(VSS),.VDD(VDD),.Y(g9280),.A(I16006));
  NOT NOT1_5274(.VSS(VSS),.VDD(VDD),.Y(I16009),.A(g9261));
  NOT NOT1_5275(.VSS(VSS),.VDD(VDD),.Y(g9281),.A(I16009));
  NOT NOT1_5276(.VSS(VSS),.VDD(VDD),.Y(I16017),.A(g9264));
  NOT NOT1_5277(.VSS(VSS),.VDD(VDD),.Y(g9297),.A(I16017));
  NOT NOT1_5278(.VSS(VSS),.VDD(VDD),.Y(I16020),.A(g9264));
  NOT NOT1_5279(.VSS(VSS),.VDD(VDD),.Y(g9298),.A(I16020));
  NOT NOT1_5280(.VSS(VSS),.VDD(VDD),.Y(I16023),.A(g9267));
  NOT NOT1_5281(.VSS(VSS),.VDD(VDD),.Y(g9299),.A(I16023));
  NOT NOT1_5282(.VSS(VSS),.VDD(VDD),.Y(I16026),.A(g9267));
  NOT NOT1_5283(.VSS(VSS),.VDD(VDD),.Y(g9300),.A(I16026));
  NOT NOT1_5284(.VSS(VSS),.VDD(VDD),.Y(g9301),.A(g9260));
  NOT NOT1_5285(.VSS(VSS),.VDD(VDD),.Y(g9302),.A(g9281));
  NOT NOT1_5286(.VSS(VSS),.VDD(VDD),.Y(g9303),.A(g9301));
  NOT NOT1_5287(.VSS(VSS),.VDD(VDD),.Y(g9304),.A(g9298));
  NOT NOT1_5288(.VSS(VSS),.VDD(VDD),.Y(I16033),.A(g9282));
  NOT NOT1_5289(.VSS(VSS),.VDD(VDD),.Y(g9305),.A(I16033));
  NOT NOT1_5290(.VSS(VSS),.VDD(VDD),.Y(I16036),.A(g9282));
  NOT NOT1_5291(.VSS(VSS),.VDD(VDD),.Y(g9306),.A(I16036));
  NOT NOT1_5292(.VSS(VSS),.VDD(VDD),.Y(g9307),.A(g9300));
  NOT NOT1_5293(.VSS(VSS),.VDD(VDD),.Y(I16040),.A(g9285));
  NOT NOT1_5294(.VSS(VSS),.VDD(VDD),.Y(g9308),.A(I16040));
  NOT NOT1_5295(.VSS(VSS),.VDD(VDD),.Y(I16043),.A(g9285));
  NOT NOT1_5296(.VSS(VSS),.VDD(VDD),.Y(g9309),.A(I16043));
  NOT NOT1_5297(.VSS(VSS),.VDD(VDD),.Y(I16046),.A(g9288));
  NOT NOT1_5298(.VSS(VSS),.VDD(VDD),.Y(g9310),.A(I16046));
  NOT NOT1_5299(.VSS(VSS),.VDD(VDD),.Y(I16049),.A(g9288));
  NOT NOT1_5300(.VSS(VSS),.VDD(VDD),.Y(g9311),.A(I16049));
  NOT NOT1_5301(.VSS(VSS),.VDD(VDD),.Y(I16052),.A(g9291));
  NOT NOT1_5302(.VSS(VSS),.VDD(VDD),.Y(g9312),.A(I16052));
  NOT NOT1_5303(.VSS(VSS),.VDD(VDD),.Y(I16055),.A(g9291));
  NOT NOT1_5304(.VSS(VSS),.VDD(VDD),.Y(g9313),.A(I16055));
  NOT NOT1_5305(.VSS(VSS),.VDD(VDD),.Y(I16058),.A(g9294));
  NOT NOT1_5306(.VSS(VSS),.VDD(VDD),.Y(g9314),.A(I16058));
  NOT NOT1_5307(.VSS(VSS),.VDD(VDD),.Y(I16061),.A(g9294));
  NOT NOT1_5308(.VSS(VSS),.VDD(VDD),.Y(g9315),.A(I16061));
  NOT NOT1_5309(.VSS(VSS),.VDD(VDD),.Y(g9316),.A(g9302));
  NOT NOT1_5310(.VSS(VSS),.VDD(VDD),.Y(g9317),.A(g9306));
  NOT NOT1_5311(.VSS(VSS),.VDD(VDD),.Y(g9318),.A(g9304));
  NOT NOT1_5312(.VSS(VSS),.VDD(VDD),.Y(g9319),.A(g9309));
  NOT NOT1_5313(.VSS(VSS),.VDD(VDD),.Y(g9320),.A(g9307));
  NOT NOT1_5314(.VSS(VSS),.VDD(VDD),.Y(g9321),.A(g9311));
  NOT NOT1_5315(.VSS(VSS),.VDD(VDD),.Y(g9322),.A(g9313));
  NOT NOT1_5316(.VSS(VSS),.VDD(VDD),.Y(g9323),.A(g9315));
  NOT NOT1_5317(.VSS(VSS),.VDD(VDD),.Y(I16072),.A(g9303));
  NOT NOT1_5318(.VSS(VSS),.VDD(VDD),.Y(g9324),.A(I16072));
  NOT NOT1_5319(.VSS(VSS),.VDD(VDD),.Y(g9329),.A(g9317));
  NOT NOT1_5320(.VSS(VSS),.VDD(VDD),.Y(g9330),.A(g9319));
  NOT NOT1_5321(.VSS(VSS),.VDD(VDD),.Y(g9331),.A(g9321));
  NOT NOT1_5322(.VSS(VSS),.VDD(VDD),.Y(g9332),.A(g9322));
  NOT NOT1_5323(.VSS(VSS),.VDD(VDD),.Y(g9333),.A(g9323));
  NOT NOT1_5324(.VSS(VSS),.VDD(VDD),.Y(I16084),.A(g9324));
  NOT NOT1_5325(.VSS(VSS),.VDD(VDD),.Y(g9336),.A(I16084));
  NOT NOT1_5326(.VSS(VSS),.VDD(VDD),.Y(I16090),.A(g9336));
  NOT NOT1_5327(.VSS(VSS),.VDD(VDD),.Y(g9340),.A(I16090));
  NOT NOT1_5328(.VSS(VSS),.VDD(VDD),.Y(I16100),.A(g9338));
  NOT NOT1_5329(.VSS(VSS),.VDD(VDD),.Y(g9350),.A(I16100));
  NOT NOT1_5330(.VSS(VSS),.VDD(VDD),.Y(I16103),.A(g9339));
  NOT NOT1_5331(.VSS(VSS),.VDD(VDD),.Y(g9351),.A(I16103));
  NOT NOT1_5332(.VSS(VSS),.VDD(VDD),.Y(I16107),.A(g9337));
  NOT NOT1_5333(.VSS(VSS),.VDD(VDD),.Y(g9353),.A(I16107));
  NOT NOT1_5334(.VSS(VSS),.VDD(VDD),.Y(I16116),.A(g9350));
  NOT NOT1_5335(.VSS(VSS),.VDD(VDD),.Y(g9360),.A(I16116));
  NOT NOT1_5336(.VSS(VSS),.VDD(VDD),.Y(I16119),.A(g9351));
  NOT NOT1_5337(.VSS(VSS),.VDD(VDD),.Y(g9361),.A(I16119));
  NOT NOT1_5338(.VSS(VSS),.VDD(VDD),.Y(I16122),.A(g9353));
  NOT NOT1_5339(.VSS(VSS),.VDD(VDD),.Y(g9362),.A(I16122));
  NOT NOT1_5340(.VSS(VSS),.VDD(VDD),.Y(I16126),.A(g9354));
  NOT NOT1_5341(.VSS(VSS),.VDD(VDD),.Y(g9366),.A(I16126));
  NOT NOT1_5342(.VSS(VSS),.VDD(VDD),.Y(I16129),.A(g9355));
  NOT NOT1_5343(.VSS(VSS),.VDD(VDD),.Y(g9367),.A(I16129));
  NOT NOT1_5344(.VSS(VSS),.VDD(VDD),.Y(I16132),.A(g9356));
  NOT NOT1_5345(.VSS(VSS),.VDD(VDD),.Y(g9368),.A(I16132));
  NOT NOT1_5346(.VSS(VSS),.VDD(VDD),.Y(I16135),.A(g9357));
  NOT NOT1_5347(.VSS(VSS),.VDD(VDD),.Y(g9369),.A(I16135));
  NOT NOT1_5348(.VSS(VSS),.VDD(VDD),.Y(I16138),.A(g9358));
  NOT NOT1_5349(.VSS(VSS),.VDD(VDD),.Y(g9370),.A(I16138));
  NOT NOT1_5350(.VSS(VSS),.VDD(VDD),.Y(I16142),.A(g9366));
  NOT NOT1_5351(.VSS(VSS),.VDD(VDD),.Y(g9372),.A(I16142));
  NOT NOT1_5352(.VSS(VSS),.VDD(VDD),.Y(I16145),.A(g9367));
  NOT NOT1_5353(.VSS(VSS),.VDD(VDD),.Y(g9373),.A(I16145));
  NOT NOT1_5354(.VSS(VSS),.VDD(VDD),.Y(I16148),.A(g9368));
  NOT NOT1_5355(.VSS(VSS),.VDD(VDD),.Y(g9374),.A(I16148));
  NOT NOT1_5356(.VSS(VSS),.VDD(VDD),.Y(I16151),.A(g9369));
  NOT NOT1_5357(.VSS(VSS),.VDD(VDD),.Y(g9375),.A(I16151));
  NOT NOT1_5358(.VSS(VSS),.VDD(VDD),.Y(I16154),.A(g9370));
  NOT NOT1_5359(.VSS(VSS),.VDD(VDD),.Y(g9376),.A(I16154));
  NOT NOT1_5360(.VSS(VSS),.VDD(VDD),.Y(I16158),.A(g9363));
  NOT NOT1_5361(.VSS(VSS),.VDD(VDD),.Y(g9378),.A(I16158));
  NOT NOT1_5362(.VSS(VSS),.VDD(VDD),.Y(I16161),.A(g9363));
  NOT NOT1_5363(.VSS(VSS),.VDD(VDD),.Y(g9379),.A(I16161));
  NOT NOT1_5364(.VSS(VSS),.VDD(VDD),.Y(g9380),.A(g9379));
  NOT NOT1_5365(.VSS(VSS),.VDD(VDD),.Y(I16165),.A(g9377));
  NOT NOT1_5366(.VSS(VSS),.VDD(VDD),.Y(g9381),.A(I16165));
  NOT NOT1_5367(.VSS(VSS),.VDD(VDD),.Y(I16168),.A(g9381));
  NOT NOT1_5368(.VSS(VSS),.VDD(VDD),.Y(g9382),.A(I16168));
  NOT NOT1_5369(.VSS(VSS),.VDD(VDD),.Y(g9383),.A(g9380));
  NOT NOT1_5370(.VSS(VSS),.VDD(VDD),.Y(I16173),.A(g9382));
  NOT NOT1_5371(.VSS(VSS),.VDD(VDD),.Y(g9385),.A(I16173));
  NOT NOT1_5372(.VSS(VSS),.VDD(VDD),.Y(I16176),.A(g9385));
  NOT NOT1_5373(.VSS(VSS),.VDD(VDD),.Y(g9386),.A(I16176));
  NOT NOT1_5374(.VSS(VSS),.VDD(VDD),.Y(I16180),.A(g9387));
  NOT NOT1_5375(.VSS(VSS),.VDD(VDD),.Y(g9388),.A(I16180));
  NOT NOT1_5376(.VSS(VSS),.VDD(VDD),.Y(I16183),.A(g9388));
  NOT NOT1_5377(.VSS(VSS),.VDD(VDD),.Y(g9389),.A(I16183));
//
  AND2 AND2_0(.VSS(VSS),.VDD(VDD),.Y(g1714),.A(g1454),.B(g1450));
  AND2 AND2_1(.VSS(VSS),.VDD(VDD),.Y(g1725),.A(g1409),.B(g1416));
  AND2 AND2_2(.VSS(VSS),.VDD(VDD),.Y(g1728),.A(g1432),.B(g1439));
  AND2 AND2_3(.VSS(VSS),.VDD(VDD),.Y(g1733),.A(g1489),.B(g1481));
  AND2 AND2_4(.VSS(VSS),.VDD(VDD),.Y(g1739),.A(g803),.B(g799));
  AND2 AND2_5(.VSS(VSS),.VDD(VDD),.Y(g1753),.A(g819),.B(g815));
  AND2 AND2_6(.VSS(VSS),.VDD(VDD),.Y(g1834),.A(g933),.B(g929));
  AND2 AND2_7(.VSS(VSS),.VDD(VDD),.Y(g1844),.A(g792),.B(g795));
  AND2 AND2_8(.VSS(VSS),.VDD(VDD),.Y(g1898),.A(g959),.B(g955));
  AND2 AND2_9(.VSS(VSS),.VDD(VDD),.Y(g1913),.A(g1528),.B(g1532));
  AND2 AND2_10(.VSS(VSS),.VDD(VDD),.Y(g1919),.A(g1098),.B(g1087));
  AND2 AND2_11(.VSS(VSS),.VDD(VDD),.Y(g2386),.A(g1130),.B(g1092));
  AND2 AND2_12(.VSS(VSS),.VDD(VDD),.Y(g2768),.A(g1597),.B(g973));
  AND2 AND2_13(.VSS(VSS),.VDD(VDD),.Y(g2781),.A(g1600),.B(g976));
  AND2 AND2_14(.VSS(VSS),.VDD(VDD),.Y(g2827),.A(g1889),.B(g1690));
  AND2 AND2_15(.VSS(VSS),.VDD(VDD),.Y(g2889),.A(g1612),.B(g1077));
  AND2 AND2_16(.VSS(VSS),.VDD(VDD),.Y(g2912),.A(g1080),.B(g1945));
  AND2 AND2_17(.VSS(VSS),.VDD(VDD),.Y(g2935),.A(g1612),.B(g1077));
  AND2 AND2_18(.VSS(VSS),.VDD(VDD),.Y(g2949),.A(g822),.B(g1753));
  AND2 AND2_19(.VSS(VSS),.VDD(VDD),.Y(g2952),.A(g2474),.B(g2215));
  AND2 AND2_20(.VSS(VSS),.VDD(VDD),.Y(g2972),.A(g2397),.B(g2407));
  AND2 AND2_21(.VSS(VSS),.VDD(VDD),.Y(g2979),.A(g1494),.B(g1733));
  AND2 AND2_22(.VSS(VSS),.VDD(VDD),.Y(g2986),.A(g806),.B(g1739));
  AND2 AND2_23(.VSS(VSS),.VDD(VDD),.Y(g3002),.A(g871),.B(g1834));
  AND2 AND2_24(.VSS(VSS),.VDD(VDD),.Y(g3049),.A(g2274),.B(g1844));
  AND2 AND2_25(.VSS(VSS),.VDD(VDD),.Y(g3081),.A(g1682),.B(g1616));
  AND2 AND2_26(.VSS(VSS),.VDD(VDD),.Y(g3094),.A(g945),.B(g1898));
  AND2 AND2_27(.VSS(VSS),.VDD(VDD),.Y(g3188),.A(g2298),.B(g2316));
  AND2 AND2_28(.VSS(VSS),.VDD(VDD),.Y(g3190),.A(g1658),.B(g2424));
  AND2 AND2_29(.VSS(VSS),.VDD(VDD),.Y(g3222),.A(g1537),.B(g1913));
  AND2 AND2_30(.VSS(VSS),.VDD(VDD),.Y(g3226),.A(g1102),.B(g1919));
  AND2 AND2_31(.VSS(VSS),.VDD(VDD),.Y(g3229),.A(g1728),.B(g2015));
  AND4 AND4_0(.VSS(VSS),.VDD(VDD),.Y(g3258),.A(g2298),.B(g2316),.C(g2334),.D(g2354));
  AND2 AND2_32(.VSS(VSS),.VDD(VDD),.Y(g3259),.A(g1976),.B(g1960));
  AND3 AND3_0(.VSS(VSS),.VDD(VDD),.Y(g3313),.A(g2334),.B(g2316),.C(g2298));
  AND3 AND3_1(.VSS(VSS),.VDD(VDD),.Y(g3429),.A(g1454),.B(g1838),.C(g1444));
  AND2 AND2_33(.VSS(VSS),.VDD(VDD),.Y(g3466),.A(g936),.B(g2557));
  AND2 AND2_34(.VSS(VSS),.VDD(VDD),.Y(g3509),.A(g1637),.B(g1616));
  AND2 AND2_35(.VSS(VSS),.VDD(VDD),.Y(g3614),.A(g1134),.B(g2386));
  AND2 AND2_36(.VSS(VSS),.VDD(VDD),.Y(g3984),.A(g2403),.B(g3085));
  AND2 AND2_37(.VSS(VSS),.VDD(VDD),.Y(g4038),.A(g825),.B(g2949));
  AND2 AND2_38(.VSS(VSS),.VDD(VDD),.Y(g4047),.A(g1272),.B(g3503));
  AND2 AND2_39(.VSS(VSS),.VDD(VDD),.Y(g4048),.A(g1288),.B(g3513));
  AND2 AND2_40(.VSS(VSS),.VDD(VDD),.Y(g4049),.A(g141),.B(g3514));
  AND2 AND2_41(.VSS(VSS),.VDD(VDD),.Y(g4052),.A(g1276),.B(g3522));
  AND2 AND2_42(.VSS(VSS),.VDD(VDD),.Y(g4053),.A(g1292),.B(g3523));
  AND2 AND2_43(.VSS(VSS),.VDD(VDD),.Y(g4054),.A(g3767),.B(g2424));
  AND2 AND2_44(.VSS(VSS),.VDD(VDD),.Y(g4058),.A(g3656),.B(g2407));
  AND2 AND2_45(.VSS(VSS),.VDD(VDD),.Y(g4059),.A(g1499),.B(g2979));
  AND2 AND2_46(.VSS(VSS),.VDD(VDD),.Y(g4062),.A(g809),.B(g2986));
  AND2 AND2_47(.VSS(VSS),.VDD(VDD),.Y(g4066),.A(g1280),.B(g3532));
  AND2 AND2_48(.VSS(VSS),.VDD(VDD),.Y(g4067),.A(g133),.B(g3539));
  AND2 AND2_49(.VSS(VSS),.VDD(VDD),.Y(g4068),.A(g121),.B(g3540));
  AND2 AND2_50(.VSS(VSS),.VDD(VDD),.Y(g4073),.A(g1300),.B(g3567));
  AND2 AND2_51(.VSS(VSS),.VDD(VDD),.Y(g4074),.A(g137),.B(g3573));
  AND2 AND2_52(.VSS(VSS),.VDD(VDD),.Y(g4077),.A(g1284),.B(g3582));
  AND4 AND4_1(.VSS(VSS),.VDD(VDD),.Y(g4078),.A(g3753),.B(g3732),.C(g3712),.D(g3700));
  AND2 AND2_53(.VSS(VSS),.VDD(VDD),.Y(g4082),.A(g1296),.B(g3604));
  AND2 AND2_54(.VSS(VSS),.VDD(VDD),.Y(g4083),.A(g125),.B(g3610));
  AND2 AND2_55(.VSS(VSS),.VDD(VDD),.Y(g4086),.A(g103),.B(g3629));
  AND2 AND2_56(.VSS(VSS),.VDD(VDD),.Y(g4091),.A(g129),.B(g3639));
  AND2 AND2_57(.VSS(VSS),.VDD(VDD),.Y(g4097),.A(g2624),.B(g2614));
  AND2 AND2_58(.VSS(VSS),.VDD(VDD),.Y(g4098),.A(g985),.B(g3790));
  AND2 AND2_59(.VSS(VSS),.VDD(VDD),.Y(g4099),.A(g117),.B(g3647));
  AND2 AND2_60(.VSS(VSS),.VDD(VDD),.Y(g4100),.A(g113),.B(g3648));
  AND2 AND2_61(.VSS(VSS),.VDD(VDD),.Y(g4101),.A(g108),.B(g3649));
  AND2 AND2_62(.VSS(VSS),.VDD(VDD),.Y(g4107),.A(g2625),.B(g2615));
  AND2 AND2_63(.VSS(VSS),.VDD(VDD),.Y(g4108),.A(g782),.B(g3655));
  AND2 AND2_64(.VSS(VSS),.VDD(VDD),.Y(g4109),.A(g990),.B(g3790));
  AND2 AND2_65(.VSS(VSS),.VDD(VDD),.Y(g4117),.A(g2626),.B(g2616));
  AND2 AND2_66(.VSS(VSS),.VDD(VDD),.Y(g4118),.A(g995),.B(g3790));
  AND2 AND2_67(.VSS(VSS),.VDD(VDD),.Y(g4123),.A(g2627),.B(g2617));
  AND2 AND2_68(.VSS(VSS),.VDD(VDD),.Y(g4124),.A(g2641),.B(g2640));
  AND2 AND2_69(.VSS(VSS),.VDD(VDD),.Y(g4127),.A(g2628),.B(g2618));
  AND2 AND2_70(.VSS(VSS),.VDD(VDD),.Y(g4128),.A(g98),.B(g3693));
  AND2 AND2_71(.VSS(VSS),.VDD(VDD),.Y(g4129),.A(g2629),.B(g2621));
  AND2 AND2_72(.VSS(VSS),.VDD(VDD),.Y(g4131),.A(g2630),.B(g2622));
  AND2 AND2_73(.VSS(VSS),.VDD(VDD),.Y(g4132),.A(g2637),.B(g2633));
  AND2 AND2_74(.VSS(VSS),.VDD(VDD),.Y(g4133),.A(g2631),.B(g2623));
  AND4 AND4_2(.VSS(VSS),.VDD(VDD),.Y(I7994),.A(g3430),.B(g3398),.C(g3359),.D(g3341));
  AND4 AND4_3(.VSS(VSS),.VDD(VDD),.Y(I7995),.A(g2074),.B(g3287),.C(g2020),.D(g3238));
  AND2 AND2_75(.VSS(VSS),.VDD(VDD),.Y(g4135),.A(I7994),.B(I7995));
  AND2 AND2_76(.VSS(VSS),.VDD(VDD),.Y(g4138),.A(g2638),.B(g2634));
  AND4 AND4_4(.VSS(VSS),.VDD(VDD),.Y(I8000),.A(g3430),.B(g3398),.C(g3359),.D(g3341));
  AND4 AND4_5(.VSS(VSS),.VDD(VDD),.Y(I8001),.A(g2074),.B(g3287),.C(g2020),.D(g1987));
  AND2 AND2_77(.VSS(VSS),.VDD(VDD),.Y(g4139),.A(I8000),.B(I8001));
  AND4 AND4_6(.VSS(VSS),.VDD(VDD),.Y(I8005),.A(g3430),.B(g3398),.C(g3359),.D(g2106));
  AND4 AND4_7(.VSS(VSS),.VDD(VDD),.Y(I8006),.A(g2074),.B(g3287),.C(g2020),.D(g3238));
  AND2 AND2_78(.VSS(VSS),.VDD(VDD),.Y(g4142),.A(I8005),.B(I8006));
  AND2 AND2_79(.VSS(VSS),.VDD(VDD),.Y(g4145),.A(g2639),.B(g2635));
  AND4 AND4_8(.VSS(VSS),.VDD(VDD),.Y(I8014),.A(g3430),.B(g3398),.C(g3359),.D(g3341));
  AND4 AND4_9(.VSS(VSS),.VDD(VDD),.Y(I8015),.A(g2074),.B(g2057),.C(g3264),.D(g3238));
  AND2 AND2_80(.VSS(VSS),.VDD(VDD),.Y(g4147),.A(I8014),.B(I8015));
  AND4 AND4_10(.VSS(VSS),.VDD(VDD),.Y(I8019),.A(g3430),.B(g3398),.C(g3359),.D(g2106));
  AND4 AND4_11(.VSS(VSS),.VDD(VDD),.Y(I8020),.A(g2074),.B(g3287),.C(g2020),.D(g1987));
  AND2 AND2_81(.VSS(VSS),.VDD(VDD),.Y(g4150),.A(I8019),.B(I8020));
  AND2 AND2_82(.VSS(VSS),.VDD(VDD),.Y(g4154),.A(g1098),.B(g3495));
  AND4 AND4_12(.VSS(VSS),.VDD(VDD),.Y(I8028),.A(g3430),.B(g3398),.C(g3359),.D(g3341));
  AND4 AND4_13(.VSS(VSS),.VDD(VDD),.Y(I8029),.A(g2074),.B(g2057),.C(g3264),.D(g1987));
  AND2 AND2_83(.VSS(VSS),.VDD(VDD),.Y(g4155),.A(I8028),.B(I8029));
  AND4 AND4_14(.VSS(VSS),.VDD(VDD),.Y(I8033),.A(g3430),.B(g3398),.C(g3359),.D(g2106));
  AND4 AND4_15(.VSS(VSS),.VDD(VDD),.Y(I8034),.A(g2074),.B(g2057),.C(g3264),.D(g3238));
  AND2 AND2_84(.VSS(VSS),.VDD(VDD),.Y(g4158),.A(I8033),.B(I8034));
  AND2 AND2_85(.VSS(VSS),.VDD(VDD),.Y(g4159),.A(g1102),.B(g3498));
  AND4 AND4_16(.VSS(VSS),.VDD(VDD),.Y(I8040),.A(g3430),.B(g3398),.C(g3359),.D(g3341));
  AND4 AND4_17(.VSS(VSS),.VDD(VDD),.Y(I8041),.A(g2074),.B(g2057),.C(g2020),.D(g3238));
  AND2 AND2_86(.VSS(VSS),.VDD(VDD),.Y(g4163),.A(I8040),.B(I8041));
  AND4 AND4_18(.VSS(VSS),.VDD(VDD),.Y(I8045),.A(g3430),.B(g3398),.C(g3359),.D(g2106));
  AND4 AND4_19(.VSS(VSS),.VDD(VDD),.Y(I8046),.A(g2074),.B(g2057),.C(g3264),.D(g1987));
  AND2 AND2_87(.VSS(VSS),.VDD(VDD),.Y(g4166),.A(I8045),.B(I8046));
  AND2 AND2_88(.VSS(VSS),.VDD(VDD),.Y(g4167),.A(g2783),.B(g1616));
  AND2 AND2_89(.VSS(VSS),.VDD(VDD),.Y(g4168),.A(g1106),.B(g3500));
  AND4 AND4_20(.VSS(VSS),.VDD(VDD),.Y(I8052),.A(g2162),.B(g2149),.C(g2137),.D(g2106));
  AND4 AND4_21(.VSS(VSS),.VDD(VDD),.Y(I8053),.A(g3316),.B(g3287),.C(g3264),.D(g3238));
  AND2 AND2_90(.VSS(VSS),.VDD(VDD),.Y(g4169),.A(I8052),.B(I8053));
  AND4 AND4_22(.VSS(VSS),.VDD(VDD),.Y(I8057),.A(g3430),.B(g3398),.C(g3359),.D(g3341));
  AND4 AND4_23(.VSS(VSS),.VDD(VDD),.Y(I8058),.A(g2074),.B(g2057),.C(g2020),.D(g1987));
  AND2 AND2_91(.VSS(VSS),.VDD(VDD),.Y(g4172),.A(I8057),.B(I8058));
  AND2 AND2_92(.VSS(VSS),.VDD(VDD),.Y(g4175),.A(g1110),.B(g3502));
  AND4 AND4_24(.VSS(VSS),.VDD(VDD),.Y(I8063),.A(g2162),.B(g2149),.C(g2137),.D(g2106));
  AND4 AND4_25(.VSS(VSS),.VDD(VDD),.Y(I8064),.A(g3316),.B(g3287),.C(g3264),.D(g1987));
  AND2 AND2_93(.VSS(VSS),.VDD(VDD),.Y(g4176),.A(I8063),.B(I8064));
  AND2 AND2_94(.VSS(VSS),.VDD(VDD),.Y(g4180),.A(g1114),.B(g3511));
  AND2 AND2_95(.VSS(VSS),.VDD(VDD),.Y(g4181),.A(g1142),.B(g3512));
  AND4 AND4_26(.VSS(VSS),.VDD(VDD),.Y(I8071),.A(g2162),.B(g2149),.C(g2137),.D(g2106));
  AND4 AND4_27(.VSS(VSS),.VDD(VDD),.Y(I8072),.A(g3316),.B(g3287),.C(g2020),.D(g3238));
  AND2 AND2_96(.VSS(VSS),.VDD(VDD),.Y(g4182),.A(I8071),.B(I8072));
  AND2 AND2_97(.VSS(VSS),.VDD(VDD),.Y(g4185),.A(g2636),.B(g2632));
  AND2 AND2_98(.VSS(VSS),.VDD(VDD),.Y(g4186),.A(g1118),.B(g3520));
  AND4 AND4_28(.VSS(VSS),.VDD(VDD),.Y(I8078),.A(g2162),.B(g2149),.C(g2137),.D(g2106));
  AND4 AND4_29(.VSS(VSS),.VDD(VDD),.Y(I8079),.A(g3316),.B(g3287),.C(g2020),.D(g1987));
  AND2 AND2_99(.VSS(VSS),.VDD(VDD),.Y(g4187),.A(I8078),.B(I8079));
  AND2 AND2_100(.VSS(VSS),.VDD(VDD),.Y(g4190),.A(g1122),.B(g3527));
  AND2 AND2_101(.VSS(VSS),.VDD(VDD),.Y(g4192),.A(g1126),.B(g3531));
  AND2 AND2_102(.VSS(VSS),.VDD(VDD),.Y(g4193),.A(g145),.B(g2727));
  AND4 AND4_30(.VSS(VSS),.VDD(VDD),.Y(I8089),.A(g2162),.B(g2149),.C(g2137),.D(g2106));
  AND4 AND4_31(.VSS(VSS),.VDD(VDD),.Y(I8090),.A(g3316),.B(g2057),.C(g2020),.D(g3238));
  AND2 AND2_103(.VSS(VSS),.VDD(VDD),.Y(g4194),.A(I8089),.B(I8090));
  AND2 AND2_104(.VSS(VSS),.VDD(VDD),.Y(g4199),.A(g93),.B(g2769));
  AND4 AND4_32(.VSS(VSS),.VDD(VDD),.Y(I8108),.A(g2162),.B(g2149),.C(g2137),.D(g2106));
  AND4 AND4_33(.VSS(VSS),.VDD(VDD),.Y(I8109),.A(g2074),.B(g3287),.C(g3264),.D(g3238));
  AND2 AND2_105(.VSS(VSS),.VDD(VDD),.Y(g4201),.A(I8108),.B(I8109));
  AND4 AND4_34(.VSS(VSS),.VDD(VDD),.Y(I8114),.A(g2162),.B(g2149),.C(g2137),.D(g2106));
  AND4 AND4_35(.VSS(VSS),.VDD(VDD),.Y(I8115),.A(g2074),.B(g3287),.C(g3264),.D(g1987));
  AND2 AND2_106(.VSS(VSS),.VDD(VDD),.Y(g4216),.A(I8114),.B(I8115));
  AND4 AND4_36(.VSS(VSS),.VDD(VDD),.Y(g4220),.A(g3533),.B(g3549),.C(g3568),.D(g3583));
  AND3 AND3_2(.VSS(VSS),.VDD(VDD),.Y(I8127),.A(g2699),.B(g2674),.C(g2677));
  AND3 AND3_3(.VSS(VSS),.VDD(VDD),.Y(g4224),.A(g2680),.B(g2683),.C(I8127));
  AND4 AND4_37(.VSS(VSS),.VDD(VDD),.Y(g4225),.A(g2686),.B(g2689),.C(g2692),.D(g2695));
  AND3 AND3_4(.VSS(VSS),.VDD(VDD),.Y(I8143),.A(g2674),.B(g2677),.C(g2680));
  AND3 AND3_5(.VSS(VSS),.VDD(VDD),.Y(g4230),.A(g2683),.B(g3491),.C(I8143));
  AND2 AND2_107(.VSS(VSS),.VDD(VDD),.Y(g4236),.A(g3260),.B(g3221));
  AND3 AND3_6(.VSS(VSS),.VDD(VDD),.Y(I8157),.A(g2686),.B(g2689),.C(g2692));
  AND3 AND3_7(.VSS(VSS),.VDD(VDD),.Y(g4238),.A(g2695),.B(g2698),.C(I8157));
  AND2 AND2_108(.VSS(VSS),.VDD(VDD),.Y(g4239),.A(g1541),.B(g3222));
  AND2 AND2_109(.VSS(VSS),.VDD(VDD),.Y(g4246),.A(g1106),.B(g3226));
  AND3 AND3_8(.VSS(VSS),.VDD(VDD),.Y(g4254),.A(g3583),.B(g3568),.C(g3549));
  AND4 AND4_38(.VSS(VSS),.VDD(VDD),.Y(I8186),.A(g3778),.B(g3549),.C(g3568),.D(g3583));
  AND4 AND4_39(.VSS(VSS),.VDD(VDD),.Y(g4255),.A(g3605),.B(g3644),.C(g3635),.D(I8186));
  AND2 AND2_110(.VSS(VSS),.VDD(VDD),.Y(g4268),.A(g2216),.B(g2655));
  AND3 AND3_9(.VSS(VSS),.VDD(VDD),.Y(I8209),.A(g2298),.B(g2316),.C(g2334));
  AND3 AND3_10(.VSS(VSS),.VDD(VDD),.Y(g4269),.A(g2354),.B(g3563),.C(I8209));
  AND2 AND2_111(.VSS(VSS),.VDD(VDD),.Y(g4271),.A(g3666),.B(g3684));
  AND2 AND2_112(.VSS(VSS),.VDD(VDD),.Y(g4272),.A(g3233),.B(g3286));
  AND2 AND2_113(.VSS(VSS),.VDD(VDD),.Y(g4276),.A(g2216),.B(g2618));
  AND2 AND2_114(.VSS(VSS),.VDD(VDD),.Y(g4282),.A(g3549),.B(g3568));
  AND2 AND2_115(.VSS(VSS),.VDD(VDD),.Y(g4284),.A(g3260),.B(g3314));
  AND3 AND3_11(.VSS(VSS),.VDD(VDD),.Y(I8237),.A(g2298),.B(g2316),.C(g2354));
  AND4 AND4_40(.VSS(VSS),.VDD(VDD),.Y(g4287),.A(g3563),.B(g2334),.C(g3579),.D(I8237));
  AND4 AND4_41(.VSS(VSS),.VDD(VDD),.Y(I8240),.A(g2298),.B(g2316),.C(g2334),.D(g2354));
  AND4 AND4_42(.VSS(VSS),.VDD(VDD),.Y(g4288),.A(g3563),.B(g3579),.C(g3603),.D(I8240));
  AND2 AND2_116(.VSS(VSS),.VDD(VDD),.Y(g4299),.A(g3233),.B(g3358));
  AND3 AND3_12(.VSS(VSS),.VDD(VDD),.Y(g4302),.A(g3086),.B(g3659),.C(g3124));
  AND2 AND2_117(.VSS(VSS),.VDD(VDD),.Y(g4304),.A(g2784),.B(g3779));
  AND4 AND4_43(.VSS(VSS),.VDD(VDD),.Y(g4312),.A(g3666),.B(g3684),.C(g3694),.D(g3707));
  AND3 AND3_13(.VSS(VSS),.VDD(VDD),.Y(g4314),.A(g3694),.B(g3684),.C(g3666));
  AND3 AND3_14(.VSS(VSS),.VDD(VDD),.Y(I8288),.A(g3666),.B(g3684),.C(g3694));
  AND3 AND3_15(.VSS(VSS),.VDD(VDD),.Y(g4315),.A(g3707),.B(g3728),.C(I8288));
  AND4 AND4_44(.VSS(VSS),.VDD(VDD),.Y(g4317),.A(g878),.B(g3086),.C(g1857),.D(g3659));
  AND3 AND3_16(.VSS(VSS),.VDD(VDD),.Y(I8296),.A(g3666),.B(g3684),.C(g3707));
  AND4 AND4_45(.VSS(VSS),.VDD(VDD),.Y(g4319),.A(g3728),.B(g3694),.C(g3750),.D(I8296));
  AND4 AND4_46(.VSS(VSS),.VDD(VDD),.Y(I8299),.A(g3666),.B(g3684),.C(g3694),.D(g3707));
  AND4 AND4_47(.VSS(VSS),.VDD(VDD),.Y(g4320),.A(g3728),.B(g3750),.C(g3768),.D(I8299));
  AND2 AND2_118(.VSS(VSS),.VDD(VDD),.Y(g4327),.A(g2959),.B(g1867));
  AND2 AND2_119(.VSS(VSS),.VDD(VDD),.Y(g4333),.A(g1087),.B(g2782));
  AND2 AND2_120(.VSS(VSS),.VDD(VDD),.Y(g4334),.A(g225),.B(g3097));
  AND2 AND2_121(.VSS(VSS),.VDD(VDD),.Y(g4342),.A(g228),.B(g3097));
  AND2 AND2_122(.VSS(VSS),.VDD(VDD),.Y(g4343),.A(g306),.B(g3131));
  AND2 AND2_123(.VSS(VSS),.VDD(VDD),.Y(g4351),.A(g309),.B(g3131));
  AND2 AND2_124(.VSS(VSS),.VDD(VDD),.Y(g4352),.A(g387),.B(g3160));
  AND2 AND2_125(.VSS(VSS),.VDD(VDD),.Y(g4355),.A(g390),.B(g3160));
  AND2 AND2_126(.VSS(VSS),.VDD(VDD),.Y(g4356),.A(g468),.B(g3192));
  AND2 AND2_127(.VSS(VSS),.VDD(VDD),.Y(g4361),.A(g471),.B(g3192));
  AND2 AND2_128(.VSS(VSS),.VDD(VDD),.Y(g4365),.A(g237),.B(g3097));
  AND2 AND2_129(.VSS(VSS),.VDD(VDD),.Y(g4366),.A(g216),.B(g3097));
  AND2 AND2_130(.VSS(VSS),.VDD(VDD),.Y(g4367),.A(g240),.B(g3097));
  AND2 AND2_131(.VSS(VSS),.VDD(VDD),.Y(g4368),.A(g318),.B(g3131));
  AND2 AND2_132(.VSS(VSS),.VDD(VDD),.Y(g4369),.A(g580),.B(g2845));
  AND2 AND2_133(.VSS(VSS),.VDD(VDD),.Y(g4375),.A(g219),.B(g3097));
  AND2 AND2_134(.VSS(VSS),.VDD(VDD),.Y(g4376),.A(g243),.B(g3097));
  AND2 AND2_135(.VSS(VSS),.VDD(VDD),.Y(g4377),.A(g297),.B(g3131));
  AND2 AND2_136(.VSS(VSS),.VDD(VDD),.Y(g4378),.A(g321),.B(g3131));
  AND2 AND2_137(.VSS(VSS),.VDD(VDD),.Y(g4379),.A(g399),.B(g3160));
  AND2 AND2_138(.VSS(VSS),.VDD(VDD),.Y(g4380),.A(g584),.B(g2845));
  AND2 AND2_139(.VSS(VSS),.VDD(VDD),.Y(g4383),.A(g222),.B(g3097));
  AND2 AND2_140(.VSS(VSS),.VDD(VDD),.Y(g4384),.A(g246),.B(g3097));
  AND2 AND2_141(.VSS(VSS),.VDD(VDD),.Y(g4385),.A(g300),.B(g3131));
  AND2 AND2_142(.VSS(VSS),.VDD(VDD),.Y(g4386),.A(g324),.B(g3131));
  AND2 AND2_143(.VSS(VSS),.VDD(VDD),.Y(g4387),.A(g378),.B(g3160));
  AND2 AND2_144(.VSS(VSS),.VDD(VDD),.Y(g4388),.A(g402),.B(g3160));
  AND2 AND2_145(.VSS(VSS),.VDD(VDD),.Y(g4389),.A(g480),.B(g3192));
  AND2 AND2_146(.VSS(VSS),.VDD(VDD),.Y(g4390),.A(g560),.B(g2845));
  AND2 AND2_147(.VSS(VSS),.VDD(VDD),.Y(g4391),.A(g249),.B(g3097));
  AND2 AND2_148(.VSS(VSS),.VDD(VDD),.Y(g4392),.A(g303),.B(g3131));
  AND2 AND2_149(.VSS(VSS),.VDD(VDD),.Y(g4393),.A(g327),.B(g3131));
  AND2 AND2_150(.VSS(VSS),.VDD(VDD),.Y(g4394),.A(g381),.B(g3160));
  AND2 AND2_151(.VSS(VSS),.VDD(VDD),.Y(g4395),.A(g405),.B(g3160));
  AND2 AND2_152(.VSS(VSS),.VDD(VDD),.Y(g4396),.A(g459),.B(g3192));
  AND2 AND2_153(.VSS(VSS),.VDD(VDD),.Y(g4397),.A(g483),.B(g3192));
  AND2 AND2_154(.VSS(VSS),.VDD(VDD),.Y(g4398),.A(g567),.B(g2845));
  AND2 AND2_155(.VSS(VSS),.VDD(VDD),.Y(g4400),.A(g1138),.B(g3614));
  AND4 AND4_48(.VSS(VSS),.VDD(VDD),.Y(I8400),.A(g3430),.B(g3398),.C(g3359),.D(g3341));
  AND4 AND4_49(.VSS(VSS),.VDD(VDD),.Y(I8401),.A(g3316),.B(g3287),.C(g3264),.D(g3238));
  AND2 AND2_156(.VSS(VSS),.VDD(VDD),.Y(g4403),.A(I8400),.B(I8401));
  AND2 AND2_157(.VSS(VSS),.VDD(VDD),.Y(g4407),.A(g252),.B(g3097));
  AND2 AND2_158(.VSS(VSS),.VDD(VDD),.Y(g4408),.A(g330),.B(g3131));
  AND2 AND2_159(.VSS(VSS),.VDD(VDD),.Y(g4409),.A(g384),.B(g3160));
  AND2 AND2_160(.VSS(VSS),.VDD(VDD),.Y(g4410),.A(g408),.B(g3160));
  AND2 AND2_161(.VSS(VSS),.VDD(VDD),.Y(g4411),.A(g462),.B(g3192));
  AND2 AND2_162(.VSS(VSS),.VDD(VDD),.Y(g4412),.A(g486),.B(g3192));
  AND4 AND4_50(.VSS(VSS),.VDD(VDD),.Y(I8412),.A(g3430),.B(g3398),.C(g3359),.D(g3341));
  AND4 AND4_51(.VSS(VSS),.VDD(VDD),.Y(I8413),.A(g3316),.B(g3287),.C(g3264),.D(g1987));
  AND2 AND2_163(.VSS(VSS),.VDD(VDD),.Y(g4414),.A(I8412),.B(I8413));
  AND4 AND4_52(.VSS(VSS),.VDD(VDD),.Y(I8417),.A(g3430),.B(g3398),.C(g3359),.D(g2106));
  AND4 AND4_53(.VSS(VSS),.VDD(VDD),.Y(I8418),.A(g3316),.B(g3287),.C(g3264),.D(g3238));
  AND2 AND2_164(.VSS(VSS),.VDD(VDD),.Y(g4417),.A(I8417),.B(I8418));
  AND2 AND2_165(.VSS(VSS),.VDD(VDD),.Y(g4420),.A(g275),.B(g3097));
  AND2 AND2_166(.VSS(VSS),.VDD(VDD),.Y(g4421),.A(g333),.B(g3131));
  AND2 AND2_167(.VSS(VSS),.VDD(VDD),.Y(g4422),.A(g411),.B(g3160));
  AND2 AND2_168(.VSS(VSS),.VDD(VDD),.Y(g4423),.A(g465),.B(g3192));
  AND2 AND2_169(.VSS(VSS),.VDD(VDD),.Y(g4424),.A(g489),.B(g3192));
  AND2 AND2_170(.VSS(VSS),.VDD(VDD),.Y(g4425),.A(g536),.B(g2845));
  AND4 AND4_54(.VSS(VSS),.VDD(VDD),.Y(I8431),.A(g3430),.B(g3398),.C(g3359),.D(g3341));
  AND4 AND4_55(.VSS(VSS),.VDD(VDD),.Y(I8432),.A(g3316),.B(g3287),.C(g2020),.D(g3238));
  AND2 AND2_171(.VSS(VSS),.VDD(VDD),.Y(g4427),.A(I8431),.B(I8432));
  AND4 AND4_56(.VSS(VSS),.VDD(VDD),.Y(I8436),.A(g3430),.B(g3398),.C(g3359),.D(g2106));
  AND4 AND4_57(.VSS(VSS),.VDD(VDD),.Y(I8437),.A(g3316),.B(g3287),.C(g3264),.D(g1987));
  AND2 AND2_172(.VSS(VSS),.VDD(VDD),.Y(g4430),.A(I8436),.B(I8437));
  AND2 AND2_173(.VSS(VSS),.VDD(VDD),.Y(g4433),.A(g278),.B(g3097));
  AND2 AND2_174(.VSS(VSS),.VDD(VDD),.Y(g4434),.A(g356),.B(g3131));
  AND2 AND2_175(.VSS(VSS),.VDD(VDD),.Y(g4435),.A(g414),.B(g3160));
  AND2 AND2_176(.VSS(VSS),.VDD(VDD),.Y(g4436),.A(g492),.B(g3192));
  AND2 AND2_177(.VSS(VSS),.VDD(VDD),.Y(g4437),.A(g540),.B(g2845));
  AND4 AND4_58(.VSS(VSS),.VDD(VDD),.Y(I8455),.A(g3430),.B(g3398),.C(g3359),.D(g3341));
  AND4 AND4_59(.VSS(VSS),.VDD(VDD),.Y(I8456),.A(g3316),.B(g3287),.C(g2020),.D(g1987));
  AND2 AND2_178(.VSS(VSS),.VDD(VDD),.Y(g4445),.A(I8455),.B(I8456));
  AND4 AND4_60(.VSS(VSS),.VDD(VDD),.Y(I8460),.A(g3430),.B(g3398),.C(g3359),.D(g2106));
  AND4 AND4_61(.VSS(VSS),.VDD(VDD),.Y(I8461),.A(g3316),.B(g3287),.C(g2020),.D(g3238));
  AND2 AND2_179(.VSS(VSS),.VDD(VDD),.Y(g4448),.A(I8460),.B(I8461));
  AND2 AND2_180(.VSS(VSS),.VDD(VDD),.Y(g4451),.A(g359),.B(g3131));
  AND2 AND2_181(.VSS(VSS),.VDD(VDD),.Y(g4452),.A(g437),.B(g3160));
  AND2 AND2_182(.VSS(VSS),.VDD(VDD),.Y(g4453),.A(g495),.B(g3192));
  AND2 AND2_183(.VSS(VSS),.VDD(VDD),.Y(g4454),.A(g544),.B(g2845));
  AND4 AND4_62(.VSS(VSS),.VDD(VDD),.Y(I8490),.A(g3430),.B(g3398),.C(g3359),.D(g3341));
  AND4 AND4_63(.VSS(VSS),.VDD(VDD),.Y(I8491),.A(g3316),.B(g2057),.C(g3264),.D(g3238));
  AND2 AND2_184(.VSS(VSS),.VDD(VDD),.Y(g4466),.A(I8490),.B(I8491));
  AND4 AND4_64(.VSS(VSS),.VDD(VDD),.Y(I8495),.A(g3430),.B(g3398),.C(g3359),.D(g2106));
  AND4 AND4_65(.VSS(VSS),.VDD(VDD),.Y(I8496),.A(g3316),.B(g3287),.C(g2020),.D(g1987));
  AND2 AND2_185(.VSS(VSS),.VDD(VDD),.Y(g4469),.A(I8495),.B(I8496));
  AND2 AND2_186(.VSS(VSS),.VDD(VDD),.Y(g4472),.A(g440),.B(g3160));
  AND2 AND2_187(.VSS(VSS),.VDD(VDD),.Y(g4473),.A(g518),.B(g3192));
  AND4 AND4_66(.VSS(VSS),.VDD(VDD),.Y(I8523),.A(g3430),.B(g3398),.C(g3359),.D(g3341));
  AND4 AND4_67(.VSS(VSS),.VDD(VDD),.Y(I8524),.A(g3316),.B(g2057),.C(g3264),.D(g1987));
  AND2 AND2_188(.VSS(VSS),.VDD(VDD),.Y(g4483),.A(I8523),.B(I8524));
  AND4 AND4_68(.VSS(VSS),.VDD(VDD),.Y(I8528),.A(g3430),.B(g3398),.C(g3359),.D(g2106));
  AND4 AND4_69(.VSS(VSS),.VDD(VDD),.Y(I8529),.A(g3316),.B(g2057),.C(g3264),.D(g3238));
  AND2 AND2_189(.VSS(VSS),.VDD(VDD),.Y(g4486),.A(I8528),.B(I8529));
  AND2 AND2_190(.VSS(VSS),.VDD(VDD),.Y(g4490),.A(g521),.B(g3192));
  AND2 AND2_191(.VSS(VSS),.VDD(VDD),.Y(g4491),.A(g557),.B(g2845));
  AND4 AND4_70(.VSS(VSS),.VDD(VDD),.Y(I8546),.A(g3430),.B(g3398),.C(g3359),.D(g3341));
  AND4 AND4_71(.VSS(VSS),.VDD(VDD),.Y(I8547),.A(g3316),.B(g2057),.C(g2020),.D(g3238));
  AND2 AND2_192(.VSS(VSS),.VDD(VDD),.Y(g4494),.A(I8546),.B(I8547));
  AND4 AND4_72(.VSS(VSS),.VDD(VDD),.Y(I8551),.A(g3430),.B(g3398),.C(g3359),.D(g2106));
  AND4 AND4_73(.VSS(VSS),.VDD(VDD),.Y(I8552),.A(g3316),.B(g2057),.C(g3264),.D(g1987));
  AND2 AND2_193(.VSS(VSS),.VDD(VDD),.Y(g4497),.A(I8551),.B(I8552));
  AND4 AND4_74(.VSS(VSS),.VDD(VDD),.Y(I8568),.A(g3430),.B(g3398),.C(g3359),.D(g3341));
  AND4 AND4_75(.VSS(VSS),.VDD(VDD),.Y(I8569),.A(g3316),.B(g2057),.C(g2020),.D(g1987));
  AND2 AND2_194(.VSS(VSS),.VDD(VDD),.Y(g4504),.A(I8568),.B(I8569));
  AND4 AND4_76(.VSS(VSS),.VDD(VDD),.Y(I8573),.A(g3430),.B(g3398),.C(g3359),.D(g2106));
  AND4 AND4_77(.VSS(VSS),.VDD(VDD),.Y(I8574),.A(g3316),.B(g2057),.C(g2020),.D(g3238));
  AND2 AND2_195(.VSS(VSS),.VDD(VDD),.Y(g4507),.A(I8573),.B(I8574));
  AND4 AND4_78(.VSS(VSS),.VDD(VDD),.Y(I8588),.A(g3430),.B(g3398),.C(g3359),.D(g3341));
  AND4 AND4_79(.VSS(VSS),.VDD(VDD),.Y(I8589),.A(g2074),.B(g3287),.C(g3264),.D(g3238));
  AND2 AND2_196(.VSS(VSS),.VDD(VDD),.Y(g4514),.A(I8588),.B(I8589));
  AND4 AND4_80(.VSS(VSS),.VDD(VDD),.Y(I8593),.A(g3430),.B(g3398),.C(g3359),.D(g2106));
  AND4 AND4_81(.VSS(VSS),.VDD(VDD),.Y(I8594),.A(g3316),.B(g2057),.C(g2020),.D(g1987));
  AND2 AND2_197(.VSS(VSS),.VDD(VDD),.Y(g4517),.A(I8593),.B(I8594));
  AND2 AND2_198(.VSS(VSS),.VDD(VDD),.Y(g4526),.A(g2642),.B(g741));
  AND4 AND4_82(.VSS(VSS),.VDD(VDD),.Y(I8612),.A(g3430),.B(g3398),.C(g3359),.D(g3341));
  AND4 AND4_83(.VSS(VSS),.VDD(VDD),.Y(I8613),.A(g2074),.B(g3287),.C(g3264),.D(g1987));
  AND2 AND2_199(.VSS(VSS),.VDD(VDD),.Y(g4529),.A(I8612),.B(I8613));
  AND4 AND4_84(.VSS(VSS),.VDD(VDD),.Y(I8617),.A(g3430),.B(g3398),.C(g3359),.D(g2106));
  AND4 AND4_85(.VSS(VSS),.VDD(VDD),.Y(I8618),.A(g2074),.B(g3287),.C(g3264),.D(g3238));
  AND2 AND2_200(.VSS(VSS),.VDD(VDD),.Y(g4532),.A(I8617),.B(I8618));
  AND2 AND2_201(.VSS(VSS),.VDD(VDD),.Y(g4546),.A(g2643),.B(g746));
  AND4 AND4_86(.VSS(VSS),.VDD(VDD),.Y(I8642),.A(g3430),.B(g3398),.C(g3359),.D(g2106));
  AND4 AND4_87(.VSS(VSS),.VDD(VDD),.Y(I8643),.A(g2074),.B(g3287),.C(g3264),.D(g1987));
  AND2 AND2_202(.VSS(VSS),.VDD(VDD),.Y(g4549),.A(I8642),.B(I8643));
  AND2 AND2_203(.VSS(VSS),.VDD(VDD),.Y(g4681),.A(g4255),.B(g3533));
  AND2 AND2_204(.VSS(VSS),.VDD(VDD),.Y(g4690),.A(g4081),.B(g3078));
  AND2 AND2_205(.VSS(VSS),.VDD(VDD),.Y(g4691),.A(g4219),.B(g1690));
  AND2 AND2_206(.VSS(VSS),.VDD(VDD),.Y(g4699),.A(g1557),.B(g4276));
  AND2 AND2_207(.VSS(VSS),.VDD(VDD),.Y(g4702),.A(g4243),.B(g1690));
  AND2 AND2_208(.VSS(VSS),.VDD(VDD),.Y(g4705),.A(g190),.B(g3986));
  AND2 AND2_209(.VSS(VSS),.VDD(VDD),.Y(g4707),.A(g812),.B(g4062));
  AND2 AND2_210(.VSS(VSS),.VDD(VDD),.Y(g4711),.A(g190),.B(g4072));
  AND2 AND2_211(.VSS(VSS),.VDD(VDD),.Y(g4712),.A(g1179),.B(g4276));
  AND2 AND2_212(.VSS(VSS),.VDD(VDD),.Y(g4720),.A(g190),.B(g4055));
  AND2 AND2_213(.VSS(VSS),.VDD(VDD),.Y(g4724),.A(g828),.B(g4038));
  AND2 AND2_214(.VSS(VSS),.VDD(VDD),.Y(g4728),.A(g190),.B(g4179));
  AND2 AND2_215(.VSS(VSS),.VDD(VDD),.Y(g4729),.A(g1504),.B(g4059));
  AND2 AND2_216(.VSS(VSS),.VDD(VDD),.Y(g4740),.A(g2242),.B(g4275));
  AND2 AND2_217(.VSS(VSS),.VDD(VDD),.Y(g4743),.A(g3518),.B(g4286));
  AND2 AND2_218(.VSS(VSS),.VDD(VDD),.Y(g4744),.A(g3525),.B(g4296));
  AND2 AND2_219(.VSS(VSS),.VDD(VDD),.Y(g4778),.A(g4169),.B(g1760));
  AND2 AND2_220(.VSS(VSS),.VDD(VDD),.Y(g4779),.A(g4176),.B(g1760));
  AND2 AND2_221(.VSS(VSS),.VDD(VDD),.Y(g4781),.A(g4182),.B(g1760));
  AND2 AND2_222(.VSS(VSS),.VDD(VDD),.Y(g4782),.A(g4187),.B(g1760));
  AND2 AND2_223(.VSS(VSS),.VDD(VDD),.Y(g4783),.A(g948),.B(g4527));
  AND2 AND2_224(.VSS(VSS),.VDD(VDD),.Y(g4785),.A(g1678),.B(g4202));
  AND2 AND2_225(.VSS(VSS),.VDD(VDD),.Y(g4787),.A(g953),.B(g4547));
  AND2 AND2_226(.VSS(VSS),.VDD(VDD),.Y(g4789),.A(g2751),.B(g4202));
  AND2 AND2_227(.VSS(VSS),.VDD(VDD),.Y(g4791),.A(g949),.B(g4562));
  AND2 AND2_228(.VSS(VSS),.VDD(VDD),.Y(g4793),.A(g3887),.B(g4202));
  AND2 AND2_229(.VSS(VSS),.VDD(VDD),.Y(g4794),.A(g954),.B(g4574));
  AND2 AND2_230(.VSS(VSS),.VDD(VDD),.Y(g4796),.A(g950),.B(g4584));
  AND2 AND2_231(.VSS(VSS),.VDD(VDD),.Y(g4797),.A(g3893),.B(g1616));
  AND2 AND2_232(.VSS(VSS),.VDD(VDD),.Y(g4798),.A(g4216),.B(g1760));
  AND2 AND2_233(.VSS(VSS),.VDD(VDD),.Y(g4799),.A(g951),.B(g4596));
  AND2 AND2_234(.VSS(VSS),.VDD(VDD),.Y(g4804),.A(g952),.B(g3876));
  AND2 AND2_235(.VSS(VSS),.VDD(VDD),.Y(g4814),.A(g150),.B(g4265));
  AND3 AND3_17(.VSS(VSS),.VDD(VDD),.Y(I9166),.A(g4041),.B(g2595),.C(g2584));
  AND3 AND3_18(.VSS(VSS),.VDD(VDD),.Y(g4819),.A(g2573),.B(g2562),.C(I9166));
  AND3 AND3_19(.VSS(VSS),.VDD(VDD),.Y(g4823),.A(g4238),.B(g4230),.C(g174));
  AND2 AND2_236(.VSS(VSS),.VDD(VDD),.Y(g4825),.A(g4228),.B(g1964));
  AND2 AND2_237(.VSS(VSS),.VDD(VDD),.Y(g4826),.A(g1545),.B(g4239));
  AND2 AND2_238(.VSS(VSS),.VDD(VDD),.Y(g4830),.A(g4288),.B(g3723));
  AND2 AND2_239(.VSS(VSS),.VDD(VDD),.Y(g4832),.A(g1110),.B(g4246));
  AND3 AND3_20(.VSS(VSS),.VDD(VDD),.Y(I9202),.A(g2605),.B(g4044),.C(g2584));
  AND3 AND3_21(.VSS(VSS),.VDD(VDD),.Y(g4837),.A(g2573),.B(g2562),.C(I9202));
  AND2 AND2_240(.VSS(VSS),.VDD(VDD),.Y(g4838),.A(g4517),.B(g1760));
  AND2 AND2_241(.VSS(VSS),.VDD(VDD),.Y(g4840),.A(g4235),.B(g1980));
  AND2 AND2_242(.VSS(VSS),.VDD(VDD),.Y(g4868),.A(g4227),.B(g4160));
  AND3 AND3_22(.VSS(VSS),.VDD(VDD),.Y(g4872),.A(g1924),.B(g4225),.C(g4224));
  AND4 AND4_88(.VSS(VSS),.VDD(VDD),.Y(g4877),.A(g3746),.B(g3723),.C(g4288),.D(g3764));
  AND3 AND3_23(.VSS(VSS),.VDD(VDD),.Y(I9222),.A(g4041),.B(g4044),.C(g2584));
  AND3 AND3_24(.VSS(VSS),.VDD(VDD),.Y(g4878),.A(g2573),.B(g2562),.C(I9222));
  AND3 AND3_25(.VSS(VSS),.VDD(VDD),.Y(g4883),.A(g3746),.B(g3723),.C(g4288));
  AND3 AND3_26(.VSS(VSS),.VDD(VDD),.Y(I9261),.A(g3777),.B(g3764),.C(g3746));
  AND3 AND3_27(.VSS(VSS),.VDD(VDD),.Y(g4901),.A(g3723),.B(g4288),.C(I9261));
  AND4 AND4_89(.VSS(VSS),.VDD(VDD),.Y(g4902),.A(g4304),.B(g2770),.C(g2746),.D(g2728));
  AND2 AND2_243(.VSS(VSS),.VDD(VDD),.Y(g4906),.A(g4320),.B(g2728));
  AND4 AND4_90(.VSS(VSS),.VDD(VDD),.Y(g4933),.A(g2746),.B(g2728),.C(g4320),.D(g2770));
  AND2 AND2_244(.VSS(VSS),.VDD(VDD),.Y(g4936),.A(g214),.B(g3888));
  AND2 AND2_245(.VSS(VSS),.VDD(VDD),.Y(g4937),.A(g3086),.B(g4309));
  AND2 AND2_246(.VSS(VSS),.VDD(VDD),.Y(g4955),.A(g215),.B(g3891));
  AND2 AND2_247(.VSS(VSS),.VDD(VDD),.Y(g4956),.A(g295),.B(g3892));
  AND3 AND3_28(.VSS(VSS),.VDD(VDD),.Y(g4957),.A(g2746),.B(g2728),.C(g4320));
  AND2 AND2_248(.VSS(VSS),.VDD(VDD),.Y(g4958),.A(g296),.B(g3897));
  AND2 AND2_249(.VSS(VSS),.VDD(VDD),.Y(g4959),.A(g376),.B(g3898));
  AND2 AND2_250(.VSS(VSS),.VDD(VDD),.Y(g4961),.A(g377),.B(g3904));
  AND2 AND2_251(.VSS(VSS),.VDD(VDD),.Y(g4962),.A(g457),.B(g3905));
  AND2 AND2_252(.VSS(VSS),.VDD(VDD),.Y(g4968),.A(g4403),.B(g1760));
  AND2 AND2_253(.VSS(VSS),.VDD(VDD),.Y(g4969),.A(g4362),.B(g2216));
  AND2 AND2_254(.VSS(VSS),.VDD(VDD),.Y(g5001),.A(g458),.B(g3912));
  AND3 AND3_29(.VSS(VSS),.VDD(VDD),.Y(I9330),.A(g2784),.B(g2770),.C(g2746));
  AND3 AND3_30(.VSS(VSS),.VDD(VDD),.Y(g5005),.A(g2728),.B(g4320),.C(I9330));
  AND2 AND2_255(.VSS(VSS),.VDD(VDD),.Y(g5008),.A(g231),.B(g3920));
  AND2 AND2_256(.VSS(VSS),.VDD(VDD),.Y(g5017),.A(g211),.B(g3928));
  AND2 AND2_257(.VSS(VSS),.VDD(VDD),.Y(g5018),.A(g232),.B(g3930));
  AND2 AND2_258(.VSS(VSS),.VDD(VDD),.Y(g5019),.A(g312),.B(g3933));
  AND2 AND2_259(.VSS(VSS),.VDD(VDD),.Y(g5020),.A(g579),.B(g3937));
  AND2 AND2_260(.VSS(VSS),.VDD(VDD),.Y(g5029),.A(g212),.B(g3945));
  AND2 AND2_261(.VSS(VSS),.VDD(VDD),.Y(g5030),.A(g233),.B(g3946));
  AND2 AND2_262(.VSS(VSS),.VDD(VDD),.Y(g5031),.A(g292),.B(g3948));
  AND2 AND2_263(.VSS(VSS),.VDD(VDD),.Y(g5032),.A(g313),.B(g3950));
  AND2 AND2_264(.VSS(VSS),.VDD(VDD),.Y(g5033),.A(g393),.B(g3953));
  AND2 AND2_265(.VSS(VSS),.VDD(VDD),.Y(g5034),.A(g583),.B(g3956));
  AND2 AND2_266(.VSS(VSS),.VDD(VDD),.Y(g5043),.A(g213),.B(g3958));
  AND2 AND2_267(.VSS(VSS),.VDD(VDD),.Y(g5044),.A(g234),.B(g3959));
  AND2 AND2_268(.VSS(VSS),.VDD(VDD),.Y(g5045),.A(g293),.B(g3961));
  AND2 AND2_269(.VSS(VSS),.VDD(VDD),.Y(g5046),.A(g314),.B(g3962));
  AND2 AND2_270(.VSS(VSS),.VDD(VDD),.Y(g5047),.A(g373),.B(g3964));
  AND2 AND2_271(.VSS(VSS),.VDD(VDD),.Y(g5048),.A(g394),.B(g3966));
  AND2 AND2_272(.VSS(VSS),.VDD(VDD),.Y(g5049),.A(g474),.B(g3969));
  AND2 AND2_273(.VSS(VSS),.VDD(VDD),.Y(g5050),.A(g587),.B(g3970));
  AND2 AND2_274(.VSS(VSS),.VDD(VDD),.Y(g5062),.A(g235),.B(g3973));
  AND2 AND2_275(.VSS(VSS),.VDD(VDD),.Y(g5063),.A(g294),.B(g3974));
  AND2 AND2_276(.VSS(VSS),.VDD(VDD),.Y(g5064),.A(g315),.B(g3975));
  AND2 AND2_277(.VSS(VSS),.VDD(VDD),.Y(g5065),.A(g374),.B(g3977));
  AND2 AND2_278(.VSS(VSS),.VDD(VDD),.Y(g5066),.A(g395),.B(g3978));
  AND2 AND2_279(.VSS(VSS),.VDD(VDD),.Y(g5067),.A(g454),.B(g3980));
  AND2 AND2_280(.VSS(VSS),.VDD(VDD),.Y(g5068),.A(g475),.B(g3982));
  AND2 AND2_281(.VSS(VSS),.VDD(VDD),.Y(g5069),.A(g566),.B(g3983));
  AND2 AND2_282(.VSS(VSS),.VDD(VDD),.Y(g5077),.A(g236),.B(g3988));
  AND2 AND2_283(.VSS(VSS),.VDD(VDD),.Y(g5078),.A(g316),.B(g3989));
  AND2 AND2_284(.VSS(VSS),.VDD(VDD),.Y(g5079),.A(g375),.B(g3990));
  AND2 AND2_285(.VSS(VSS),.VDD(VDD),.Y(g5080),.A(g396),.B(g3991));
  AND2 AND2_286(.VSS(VSS),.VDD(VDD),.Y(g5081),.A(g455),.B(g3993));
  AND2 AND2_287(.VSS(VSS),.VDD(VDD),.Y(g5082),.A(g476),.B(g3994));
  AND2 AND2_288(.VSS(VSS),.VDD(VDD),.Y(g5089),.A(g273),.B(g3998));
  AND2 AND2_289(.VSS(VSS),.VDD(VDD),.Y(g5090),.A(g317),.B(g4000));
  AND2 AND2_290(.VSS(VSS),.VDD(VDD),.Y(g5091),.A(g397),.B(g4001));
  AND2 AND2_291(.VSS(VSS),.VDD(VDD),.Y(g5092),.A(g456),.B(g4002));
  AND2 AND2_292(.VSS(VSS),.VDD(VDD),.Y(g5093),.A(g477),.B(g4003));
  AND2 AND2_293(.VSS(VSS),.VDD(VDD),.Y(g5094),.A(g535),.B(g4004));
  AND2 AND2_294(.VSS(VSS),.VDD(VDD),.Y(g5096),.A(g1149),.B(g4400));
  AND2 AND2_295(.VSS(VSS),.VDD(VDD),.Y(g5104),.A(g274),.B(g4010));
  AND2 AND2_296(.VSS(VSS),.VDD(VDD),.Y(g5105),.A(g354),.B(g4013));
  AND2 AND2_297(.VSS(VSS),.VDD(VDD),.Y(g5106),.A(g398),.B(g4015));
  AND2 AND2_298(.VSS(VSS),.VDD(VDD),.Y(g5107),.A(g478),.B(g4016));
  AND2 AND2_299(.VSS(VSS),.VDD(VDD),.Y(g5108),.A(g539),.B(g4017));
  AND2 AND2_300(.VSS(VSS),.VDD(VDD),.Y(g5116),.A(g355),.B(g4021));
  AND2 AND2_301(.VSS(VSS),.VDD(VDD),.Y(g5117),.A(g435),.B(g4024));
  AND2 AND2_302(.VSS(VSS),.VDD(VDD),.Y(g5118),.A(g479),.B(g4026));
  AND2 AND2_303(.VSS(VSS),.VDD(VDD),.Y(g5119),.A(g543),.B(g4027));
  AND2 AND2_304(.VSS(VSS),.VDD(VDD),.Y(g5122),.A(g436),.B(g4030));
  AND2 AND2_305(.VSS(VSS),.VDD(VDD),.Y(g5123),.A(g516),.B(g4033));
  AND2 AND2_306(.VSS(VSS),.VDD(VDD),.Y(g5125),.A(g517),.B(g4036));
  AND2 AND2_307(.VSS(VSS),.VDD(VDD),.Y(g5126),.A(g556),.B(g4037));
  AND4 AND4_91(.VSS(VSS),.VDD(VDD),.Y(I9534),.A(g3019),.B(g3029),.C(g3038),.D(g3052));
  AND4 AND4_92(.VSS(VSS),.VDD(VDD),.Y(I9535),.A(g3062),.B(g2712),.C(g4253),.D(g2752));
  AND2 AND2_308(.VSS(VSS),.VDD(VDD),.Y(g5132),.A(I9534),.B(I9535));
  AND2 AND2_309(.VSS(VSS),.VDD(VDD),.Y(g5142),.A(g1677),.B(g4202));
  AND2 AND2_310(.VSS(VSS),.VDD(VDD),.Y(g5287),.A(g786),.B(g4724));
  AND2 AND2_311(.VSS(VSS),.VDD(VDD),.Y(g5298),.A(g1912),.B(g4814));
  AND2 AND2_312(.VSS(VSS),.VDD(VDD),.Y(g5313),.A(g4820),.B(g2407));
  AND2 AND2_313(.VSS(VSS),.VDD(VDD),.Y(g5314),.A(g1509),.B(g4729));
  AND2 AND2_314(.VSS(VSS),.VDD(VDD),.Y(g5334),.A(g4887),.B(g2424));
  AND2 AND2_315(.VSS(VSS),.VDD(VDD),.Y(g5425),.A(g1528),.B(g4916));
  AND2 AND2_316(.VSS(VSS),.VDD(VDD),.Y(g5428),.A(g775),.B(g4707));
  AND2 AND2_317(.VSS(VSS),.VDD(VDD),.Y(g5432),.A(g1537),.B(g4921));
  AND2 AND2_318(.VSS(VSS),.VDD(VDD),.Y(g5436),.A(g1541),.B(g4926));
  AND2 AND2_319(.VSS(VSS),.VDD(VDD),.Y(g5438),.A(g1545),.B(g4932));
  AND2 AND2_320(.VSS(VSS),.VDD(VDD),.Y(g5441),.A(g4870),.B(g3497));
  AND2 AND2_321(.VSS(VSS),.VDD(VDD),.Y(g5442),.A(g4679),.B(g4202));
  AND2 AND2_322(.VSS(VSS),.VDD(VDD),.Y(g5443),.A(g1549),.B(g4935));
  AND2 AND2_323(.VSS(VSS),.VDD(VDD),.Y(g5452),.A(g4876),.B(g3499));
  AND2 AND2_324(.VSS(VSS),.VDD(VDD),.Y(g5458),.A(g4686),.B(g1616));
  AND2 AND2_325(.VSS(VSS),.VDD(VDD),.Y(g5475),.A(g3801),.B(g5022));
  AND2 AND2_326(.VSS(VSS),.VDD(VDD),.Y(g5479),.A(g5141),.B(g5037));
  AND2 AND2_327(.VSS(VSS),.VDD(VDD),.Y(g5484),.A(g1037),.B(g5096));
  AND2 AND2_328(.VSS(VSS),.VDD(VDD),.Y(g5489),.A(g4912),.B(g5053));
  AND2 AND2_329(.VSS(VSS),.VDD(VDD),.Y(g5513),.A(g4889),.B(g5071));
  AND2 AND2_330(.VSS(VSS),.VDD(VDD),.Y(g5547),.A(g4814),.B(g1819));
  AND2 AND2_331(.VSS(VSS),.VDD(VDD),.Y(g5548),.A(g1549),.B(g4826));
  AND2 AND2_332(.VSS(VSS),.VDD(VDD),.Y(g5552),.A(g1114),.B(g4832));
  AND2 AND2_333(.VSS(VSS),.VDD(VDD),.Y(g5560),.A(g3390),.B(g5036));
  AND2 AND2_334(.VSS(VSS),.VDD(VDD),.Y(g5563),.A(g3390),.B(g5070));
  AND2 AND2_335(.VSS(VSS),.VDD(VDD),.Y(g5570),.A(g1759),.B(g4841));
  AND2 AND2_336(.VSS(VSS),.VDD(VDD),.Y(g5573),.A(g3011),.B(g4841));
  AND2 AND2_337(.VSS(VSS),.VDD(VDD),.Y(g5579),.A(g4090),.B(g4841));
  AND2 AND2_338(.VSS(VSS),.VDD(VDD),.Y(g5583),.A(g1775),.B(g4969));
  AND2 AND2_339(.VSS(VSS),.VDD(VDD),.Y(g5585),.A(g4741),.B(g4841));
  AND2 AND2_340(.VSS(VSS),.VDD(VDD),.Y(g5588),.A(g3028),.B(g4969));
  AND2 AND2_341(.VSS(VSS),.VDD(VDD),.Y(g5593),.A(g4110),.B(g4969));
  AND2 AND2_342(.VSS(VSS),.VDD(VDD),.Y(g5599),.A(g4745),.B(g4969));
  AND2 AND2_343(.VSS(VSS),.VDD(VDD),.Y(g5624),.A(g5140),.B(g2794));
  AND2 AND2_344(.VSS(VSS),.VDD(VDD),.Y(g5699),.A(g1667),.B(g4841));
  AND2 AND2_345(.VSS(VSS),.VDD(VDD),.Y(g5700),.A(g1638),.B(g4969));
  AND2 AND2_346(.VSS(VSS),.VDD(VDD),.Y(g5714),.A(g1532),.B(g4733));
  AND2 AND2_347(.VSS(VSS),.VDD(VDD),.Y(g5765),.A(g1695),.B(g5428));
  AND2 AND2_348(.VSS(VSS),.VDD(VDD),.Y(g5767),.A(g5344),.B(g3079));
  AND2 AND2_349(.VSS(VSS),.VDD(VDD),.Y(g5783),.A(g1897),.B(g5287));
  AND2 AND2_350(.VSS(VSS),.VDD(VDD),.Y(g5817),.A(g5395),.B(g3091));
  AND2 AND2_351(.VSS(VSS),.VDD(VDD),.Y(g5894),.A(g1118),.B(g5552));
  AND2 AND2_352(.VSS(VSS),.VDD(VDD),.Y(g5937),.A(g5562),.B(g2407));
  AND2 AND2_353(.VSS(VSS),.VDD(VDD),.Y(g5969),.A(g5564),.B(g2424));
  AND2 AND2_354(.VSS(VSS),.VDD(VDD),.Y(g5970),.A(g5605),.B(g2424));
  AND2 AND2_355(.VSS(VSS),.VDD(VDD),.Y(g5984),.A(g1041),.B(g5484));
  AND2 AND2_356(.VSS(VSS),.VDD(VDD),.Y(g6001),.A(g5540),.B(g2407));
  AND2 AND2_357(.VSS(VSS),.VDD(VDD),.Y(g6002),.A(g5539),.B(g2407));
  AND3 AND3_31(.VSS(VSS),.VDD(VDD),.Y(I10597),.A(g3769),.B(g3754),.C(g3735));
  AND3 AND3_32(.VSS(VSS),.VDD(VDD),.Y(g6003),.A(g3716),.B(g5633),.C(I10597));
  AND2 AND2_358(.VSS(VSS),.VDD(VDD),.Y(g6005),.A(g5557),.B(g2407));
  AND2 AND2_359(.VSS(VSS),.VDD(VDD),.Y(g6006),.A(g5575),.B(g2424));
  AND2 AND2_360(.VSS(VSS),.VDD(VDD),.Y(g6013),.A(g5589),.B(g2424));
  AND2 AND2_361(.VSS(VSS),.VDD(VDD),.Y(g6021),.A(g5594),.B(g2424));
  AND2 AND2_362(.VSS(VSS),.VDD(VDD),.Y(g6022),.A(g5595),.B(g2424));
  AND2 AND2_363(.VSS(VSS),.VDD(VDD),.Y(g6039),.A(g1037),.B(g5574));
  AND2 AND2_364(.VSS(VSS),.VDD(VDD),.Y(g6040),.A(g1462),.B(g5578));
  AND2 AND2_365(.VSS(VSS),.VDD(VDD),.Y(g6041),.A(g5189),.B(g4969));
  AND2 AND2_366(.VSS(VSS),.VDD(VDD),.Y(g6042),.A(g1041),.B(g5581));
  AND2 AND2_367(.VSS(VSS),.VDD(VDD),.Y(g6043),.A(g1069),.B(g5582));
  AND2 AND2_368(.VSS(VSS),.VDD(VDD),.Y(g6044),.A(g1467),.B(g5584));
  AND2 AND2_369(.VSS(VSS),.VDD(VDD),.Y(g6045),.A(g1472),.B(g5591));
  AND2 AND2_370(.VSS(VSS),.VDD(VDD),.Y(g6046),.A(g1073),.B(g5592));
  AND2 AND2_371(.VSS(VSS),.VDD(VDD),.Y(g6047),.A(g1477),.B(g5596));
  AND2 AND2_372(.VSS(VSS),.VDD(VDD),.Y(g6049),.A(g1045),.B(g5597));
  AND2 AND2_373(.VSS(VSS),.VDD(VDD),.Y(g6052),.A(g1049),.B(g5604));
  AND2 AND2_374(.VSS(VSS),.VDD(VDD),.Y(g6053),.A(g1053),.B(g5608));
  AND2 AND2_375(.VSS(VSS),.VDD(VDD),.Y(g6054),.A(g1057),.B(g5611));
  AND2 AND2_376(.VSS(VSS),.VDD(VDD),.Y(g6055),.A(g5239),.B(g4202));
  AND3 AND3_33(.VSS(VSS),.VDD(VDD),.Y(g6056),.A(g3760),.B(g5286),.C(g1695));
  AND2 AND2_377(.VSS(VSS),.VDD(VDD),.Y(g6057),.A(g1061),.B(g5617));
  AND2 AND2_378(.VSS(VSS),.VDD(VDD),.Y(g6058),.A(g5561),.B(g3501));
  AND2 AND2_379(.VSS(VSS),.VDD(VDD),.Y(g6060),.A(g1065),.B(g5623));
  AND2 AND2_380(.VSS(VSS),.VDD(VDD),.Y(g6061),.A(g5257),.B(g1616));
  AND2 AND2_381(.VSS(VSS),.VDD(VDD),.Y(g6091),.A(g5712),.B(g5038));
  AND2 AND2_382(.VSS(VSS),.VDD(VDD),.Y(g6098),.A(g5681),.B(g1247));
  AND2 AND2_383(.VSS(VSS),.VDD(VDD),.Y(g6105),.A(g5618),.B(g2817));
  AND2 AND2_384(.VSS(VSS),.VDD(VDD),.Y(g6107),.A(g5478),.B(g1849));
  AND2 AND2_385(.VSS(VSS),.VDD(VDD),.Y(g6109),.A(g5453),.B(g5335));
  AND3 AND3_34(.VSS(VSS),.VDD(VDD),.Y(g6112),.A(g5673),.B(g4841),.C(g5541));
  AND2 AND2_386(.VSS(VSS),.VDD(VDD),.Y(g6125),.A(g5548),.B(g4202));
  AND2 AND2_387(.VSS(VSS),.VDD(VDD),.Y(g6145),.A(g1489),.B(g5705));
  AND2 AND2_388(.VSS(VSS),.VDD(VDD),.Y(g6151),.A(g1494),.B(g5709));
  AND2 AND2_389(.VSS(VSS),.VDD(VDD),.Y(g6154),.A(g1499),.B(g5713));
  AND2 AND2_390(.VSS(VSS),.VDD(VDD),.Y(g6157),.A(g1130),.B(g5717));
  AND2 AND2_391(.VSS(VSS),.VDD(VDD),.Y(g6160),.A(g1504),.B(g5718));
  AND2 AND2_392(.VSS(VSS),.VDD(VDD),.Y(g6162),.A(g1134),.B(g5724));
  AND2 AND2_393(.VSS(VSS),.VDD(VDD),.Y(g6166),.A(g1509),.B(g5725));
  AND2 AND2_394(.VSS(VSS),.VDD(VDD),.Y(g6168),.A(g1138),.B(g5191));
  AND2 AND2_395(.VSS(VSS),.VDD(VDD),.Y(g6171),.A(g5363),.B(g4841));
  AND2 AND2_396(.VSS(VSS),.VDD(VDD),.Y(g6172),.A(g1514),.B(g5192));
  AND2 AND2_397(.VSS(VSS),.VDD(VDD),.Y(g6175),.A(g4332),.B(g5614));
  AND2 AND2_398(.VSS(VSS),.VDD(VDD),.Y(g6176),.A(g1149),.B(g5198));
  AND2 AND2_399(.VSS(VSS),.VDD(VDD),.Y(g6182),.A(g1519),.B(g5199));
  AND2 AND2_400(.VSS(VSS),.VDD(VDD),.Y(g6196),.A(g4927),.B(g5615));
  AND2 AND2_401(.VSS(VSS),.VDD(VDD),.Y(g6204),.A(g5542),.B(g5294));
  AND2 AND2_402(.VSS(VSS),.VDD(VDD),.Y(g6239),.A(g1514),.B(g5314));
  AND2 AND2_403(.VSS(VSS),.VDD(VDD),.Y(g6266),.A(g1481),.B(g5285));
  AND2 AND2_404(.VSS(VSS),.VDD(VDD),.Y(g6268),.A(g1092),.B(g5309));
  AND2 AND2_405(.VSS(VSS),.VDD(VDD),.Y(g6394),.A(g5988),.B(g5494));
  AND2 AND2_406(.VSS(VSS),.VDD(VDD),.Y(g6395),.A(g2157),.B(g6007));
  AND2 AND2_407(.VSS(VSS),.VDD(VDD),.Y(g6396),.A(g661),.B(g6008));
  AND2 AND2_408(.VSS(VSS),.VDD(VDD),.Y(g6399),.A(g5971),.B(g5494));
  AND2 AND2_409(.VSS(VSS),.VDD(VDD),.Y(g6400),.A(g150),.B(g6011));
  AND2 AND2_410(.VSS(VSS),.VDD(VDD),.Y(g6401),.A(g5971),.B(g5367));
  AND2 AND2_411(.VSS(VSS),.VDD(VDD),.Y(g6402),.A(g665),.B(g6012));
  AND2 AND2_412(.VSS(VSS),.VDD(VDD),.Y(g6405),.A(g5956),.B(g5494));
  AND2 AND2_413(.VSS(VSS),.VDD(VDD),.Y(g6406),.A(g154),.B(g6018));
  AND2 AND2_414(.VSS(VSS),.VDD(VDD),.Y(g6407),.A(g5956),.B(g5367));
  AND2 AND2_415(.VSS(VSS),.VDD(VDD),.Y(g6408),.A(g669),.B(g6019));
  AND2 AND2_416(.VSS(VSS),.VDD(VDD),.Y(g6409),.A(g706),.B(g6020));
  AND2 AND2_417(.VSS(VSS),.VDD(VDD),.Y(g6411),.A(g5918),.B(g5494));
  AND2 AND2_418(.VSS(VSS),.VDD(VDD),.Y(g6412),.A(g158),.B(g6024));
  AND2 AND2_419(.VSS(VSS),.VDD(VDD),.Y(g6413),.A(g5939),.B(g5367));
  AND2 AND2_420(.VSS(VSS),.VDD(VDD),.Y(g6414),.A(g673),.B(g6025));
  AND2 AND2_421(.VSS(VSS),.VDD(VDD),.Y(g6415),.A(g5988),.B(g5367));
  AND2 AND2_422(.VSS(VSS),.VDD(VDD),.Y(g6416),.A(g710),.B(g6026));
  AND2 AND2_423(.VSS(VSS),.VDD(VDD),.Y(g6417),.A(g718),.B(g6027));
  AND2 AND2_424(.VSS(VSS),.VDD(VDD),.Y(g6418),.A(g5897),.B(g5494));
  AND2 AND2_425(.VSS(VSS),.VDD(VDD),.Y(g6419),.A(g162),.B(g6032));
  AND2 AND2_426(.VSS(VSS),.VDD(VDD),.Y(g6420),.A(g5918),.B(g5367));
  AND2 AND2_427(.VSS(VSS),.VDD(VDD),.Y(g6421),.A(g5847),.B(g5384));
  AND2 AND2_428(.VSS(VSS),.VDD(VDD),.Y(g6422),.A(g714),.B(g6033));
  AND2 AND2_429(.VSS(VSS),.VDD(VDD),.Y(g6423),.A(g5897),.B(g5384));
  AND2 AND2_430(.VSS(VSS),.VDD(VDD),.Y(g6428),.A(g5874),.B(g5494));
  AND2 AND2_431(.VSS(VSS),.VDD(VDD),.Y(g6429),.A(g168),.B(g6035));
  AND2 AND2_432(.VSS(VSS),.VDD(VDD),.Y(g6430),.A(g5874),.B(g5384));
  AND2 AND2_433(.VSS(VSS),.VDD(VDD),.Y(g6431),.A(g5847),.B(g5494));
  AND2 AND2_434(.VSS(VSS),.VDD(VDD),.Y(g6433),.A(g778),.B(g6134));
  AND2 AND2_435(.VSS(VSS),.VDD(VDD),.Y(g6434),.A(g855),.B(g6048));
  AND2 AND2_436(.VSS(VSS),.VDD(VDD),.Y(g6437),.A(g859),.B(g6050));
  AND2 AND2_437(.VSS(VSS),.VDD(VDD),.Y(g6438),.A(g4829),.B(g6051));
  AND2 AND2_438(.VSS(VSS),.VDD(VDD),.Y(g6439),.A(g789),.B(g6150));
  AND2 AND2_439(.VSS(VSS),.VDD(VDD),.Y(g6444),.A(g1676),.B(g6125));
  AND2 AND2_440(.VSS(VSS),.VDD(VDD),.Y(g6447),.A(g734),.B(g6073));
  AND2 AND2_441(.VSS(VSS),.VDD(VDD),.Y(g6448),.A(g5918),.B(g5384));
  AND2 AND2_442(.VSS(VSS),.VDD(VDD),.Y(g6456),.A(g6116),.B(g2407));
  AND2 AND2_443(.VSS(VSS),.VDD(VDD),.Y(g6460),.A(g6178),.B(g2424));
  AND2 AND2_444(.VSS(VSS),.VDD(VDD),.Y(g6462),.A(g6215),.B(g2424));
  AND2 AND2_445(.VSS(VSS),.VDD(VDD),.Y(g6464),.A(g6177),.B(g2424));
  AND2 AND2_446(.VSS(VSS),.VDD(VDD),.Y(g6474),.A(g6203),.B(g2424));
  AND2 AND2_447(.VSS(VSS),.VDD(VDD),.Y(g6487),.A(g5750),.B(g4969));
  AND2 AND2_448(.VSS(VSS),.VDD(VDD),.Y(g6541),.A(g6144),.B(g3510));
  AND2 AND2_449(.VSS(VSS),.VDD(VDD),.Y(g6554),.A(g5762),.B(g1616));
  AND2 AND2_450(.VSS(VSS),.VDD(VDD),.Y(g6567),.A(g6265),.B(g2424));
  AND2 AND2_451(.VSS(VSS),.VDD(VDD),.Y(g6574),.A(g1045),.B(g5984));
  AND2 AND2_452(.VSS(VSS),.VDD(VDD),.Y(g6577),.A(g6142),.B(g4160));
  AND2 AND2_453(.VSS(VSS),.VDD(VDD),.Y(g6578),.A(g6218),.B(g3913));
  AND2 AND2_454(.VSS(VSS),.VDD(VDD),.Y(g6582),.A(g1122),.B(g5894));
  AND2 AND2_455(.VSS(VSS),.VDD(VDD),.Y(g6611),.A(g3390),.B(g6249));
  AND2 AND2_456(.VSS(VSS),.VDD(VDD),.Y(g6629),.A(g6023),.B(g4841));
  AND2 AND2_457(.VSS(VSS),.VDD(VDD),.Y(g6633),.A(g5526),.B(g5987));
  AND2 AND2_458(.VSS(VSS),.VDD(VDD),.Y(g6638),.A(g174),.B(g5755));
  AND2 AND2_459(.VSS(VSS),.VDD(VDD),.Y(g6641),.A(g5939),.B(g5494));
  AND2 AND2_460(.VSS(VSS),.VDD(VDD),.Y(g6643),.A(g1860),.B(g5868));
  AND2 AND2_461(.VSS(VSS),.VDD(VDD),.Y(g6689),.A(g1519),.B(g6239));
  AND2 AND2_462(.VSS(VSS),.VDD(VDD),.Y(g6715),.A(g677),.B(g5843));
  AND2 AND2_463(.VSS(VSS),.VDD(VDD),.Y(g6726),.A(g5897),.B(g5367));
  AND2 AND2_464(.VSS(VSS),.VDD(VDD),.Y(g6727),.A(g681),.B(g5846));
  AND2 AND2_465(.VSS(VSS),.VDD(VDD),.Y(g6732),.A(g5874),.B(g5367));
  AND2 AND2_466(.VSS(VSS),.VDD(VDD),.Y(g6733),.A(g685),.B(g5873));
  AND2 AND2_467(.VSS(VSS),.VDD(VDD),.Y(g6738),.A(g5847),.B(g5367));
  AND2 AND2_468(.VSS(VSS),.VDD(VDD),.Y(g6743),.A(g730),.B(g5916));
  AND2 AND2_469(.VSS(VSS),.VDD(VDD),.Y(g6745),.A(g1872),.B(g6198));
  AND2 AND2_470(.VSS(VSS),.VDD(VDD),.Y(g6753),.A(g5939),.B(g5384));
  AND2 AND2_471(.VSS(VSS),.VDD(VDD),.Y(g6757),.A(g5874),.B(g5412));
  AND2 AND2_472(.VSS(VSS),.VDD(VDD),.Y(g6762),.A(g5847),.B(g5412));
  AND2 AND2_473(.VSS(VSS),.VDD(VDD),.Y(g6771),.A(g146),.B(g6004));
  AND2 AND2_474(.VSS(VSS),.VDD(VDD),.Y(g6908),.A(g6478),.B(g5246));
  AND2 AND2_475(.VSS(VSS),.VDD(VDD),.Y(g6914),.A(g6483),.B(g5246));
  AND2 AND2_476(.VSS(VSS),.VDD(VDD),.Y(g6915),.A(g6493),.B(g5246));
  AND2 AND2_477(.VSS(VSS),.VDD(VDD),.Y(g6916),.A(g727),.B(g6515));
  AND2 AND2_478(.VSS(VSS),.VDD(VDD),.Y(g6923),.A(g6570),.B(g5612));
  AND2 AND2_479(.VSS(VSS),.VDD(VDD),.Y(g6941),.A(g1126),.B(g6582));
  AND2 AND2_480(.VSS(VSS),.VDD(VDD),.Y(g6949),.A(g5483),.B(g6589));
  AND2 AND2_481(.VSS(VSS),.VDD(VDD),.Y(g6951),.A(g5511),.B(g6595));
  AND2 AND2_482(.VSS(VSS),.VDD(VDD),.Y(g6954),.A(g5518),.B(g6601));
  AND2 AND2_483(.VSS(VSS),.VDD(VDD),.Y(g6965),.A(g55),.B(g6489));
  AND2 AND2_484(.VSS(VSS),.VDD(VDD),.Y(g6966),.A(g6580),.B(g5580));
  AND2 AND2_485(.VSS(VSS),.VDD(VDD),.Y(g6970),.A(g5035),.B(g6490));
  AND2 AND2_486(.VSS(VSS),.VDD(VDD),.Y(g6971),.A(g6424),.B(g4969));
  AND2 AND2_487(.VSS(VSS),.VDD(VDD),.Y(g6972),.A(g5661),.B(g6498));
  AND2 AND2_488(.VSS(VSS),.VDD(VDD),.Y(g6974),.A(g3613),.B(g6505));
  AND2 AND2_489(.VSS(VSS),.VDD(VDD),.Y(g6976),.A(g4399),.B(g6508));
  AND2 AND2_490(.VSS(VSS),.VDD(VDD),.Y(g6979),.A(g5095),.B(g6511));
  AND2 AND2_491(.VSS(VSS),.VDD(VDD),.Y(g6990),.A(g799),.B(g6517));
  AND2 AND2_492(.VSS(VSS),.VDD(VDD),.Y(g6991),.A(g5689),.B(g6520));
  AND2 AND2_493(.VSS(VSS),.VDD(VDD),.Y(g6992),.A(g6610),.B(g3519));
  AND2 AND2_494(.VSS(VSS),.VDD(VDD),.Y(g6994),.A(g3658),.B(g6538));
  AND2 AND2_495(.VSS(VSS),.VDD(VDD),.Y(g6995),.A(g6435),.B(g1616));
  AND2 AND2_496(.VSS(VSS),.VDD(VDD),.Y(g6996),.A(g3678),.B(g6552));
  AND2 AND2_497(.VSS(VSS),.VDD(VDD),.Y(g6998),.A(g4474),.B(g6555));
  AND2 AND2_498(.VSS(VSS),.VDD(VDD),.Y(g6999),.A(g815),.B(g6556));
  AND2 AND2_499(.VSS(VSS),.VDD(VDD),.Y(g7001),.A(g3722),.B(g6562));
  AND2 AND2_500(.VSS(VSS),.VDD(VDD),.Y(g7002),.A(g6770),.B(g5054));
  AND2 AND2_501(.VSS(VSS),.VDD(VDD),.Y(g7003),.A(g1462),.B(g6689));
  AND2 AND2_502(.VSS(VSS),.VDD(VDD),.Y(g7007),.A(g6627),.B(g5072));
  AND2 AND2_503(.VSS(VSS),.VDD(VDD),.Y(g7008),.A(g6615),.B(g5083));
  AND2 AND2_504(.VSS(VSS),.VDD(VDD),.Y(g7010),.A(g1049),.B(g6574));
  AND2 AND2_505(.VSS(VSS),.VDD(VDD),.Y(g7017),.A(g3390),.B(g6706));
  AND2 AND2_506(.VSS(VSS),.VDD(VDD),.Y(g7021),.A(g3390),.B(g6673));
  AND2 AND2_507(.VSS(VSS),.VDD(VDD),.Y(g7027),.A(g3390),.B(g6698));
  AND2 AND2_508(.VSS(VSS),.VDD(VDD),.Y(g7030),.A(g6705),.B(g5723));
  AND2 AND2_509(.VSS(VSS),.VDD(VDD),.Y(g7031),.A(g3390),.B(g6717));
  AND2 AND2_510(.VSS(VSS),.VDD(VDD),.Y(g7033),.A(g6716),.B(g5190));
  AND2 AND2_511(.VSS(VSS),.VDD(VDD),.Y(g7036),.A(g6728),.B(g5197));
  AND2 AND2_512(.VSS(VSS),.VDD(VDD),.Y(g7038),.A(g6466),.B(g4841));
  AND2 AND2_513(.VSS(VSS),.VDD(VDD),.Y(g7041),.A(g6734),.B(g5206));
  AND2 AND2_514(.VSS(VSS),.VDD(VDD),.Y(g7071),.A(g6639),.B(g1872));
  AND2 AND2_515(.VSS(VSS),.VDD(VDD),.Y(g7079),.A(g4259),.B(g6677));
  AND2 AND2_516(.VSS(VSS),.VDD(VDD),.Y(g7087),.A(g6440),.B(g5311));
  AND2 AND2_517(.VSS(VSS),.VDD(VDD),.Y(g7096),.A(g6677),.B(g5101));
  AND2 AND2_518(.VSS(VSS),.VDD(VDD),.Y(g7128),.A(g6926),.B(g3047));
  AND2 AND2_519(.VSS(VSS),.VDD(VDD),.Y(g7136),.A(g4057),.B(g6953));
  AND2 AND2_520(.VSS(VSS),.VDD(VDD),.Y(g7175),.A(g6893),.B(g4841));
  AND2 AND2_521(.VSS(VSS),.VDD(VDD),.Y(g7177),.A(g7016),.B(g5586));
  AND2 AND2_522(.VSS(VSS),.VDD(VDD),.Y(g7179),.A(g6121),.B(g7035));
  AND2 AND2_523(.VSS(VSS),.VDD(VDD),.Y(g7181),.A(g6124),.B(g7039));
  AND2 AND2_524(.VSS(VSS),.VDD(VDD),.Y(g7182),.A(g6902),.B(g4969));
  AND2 AND2_525(.VSS(VSS),.VDD(VDD),.Y(g7183),.A(g6132),.B(g7042));
  AND2 AND2_526(.VSS(VSS),.VDD(VDD),.Y(g7184),.A(g6138),.B(g7043));
  AND2 AND2_527(.VSS(VSS),.VDD(VDD),.Y(g7186),.A(g6600),.B(g7044));
  AND2 AND2_528(.VSS(VSS),.VDD(VDD),.Y(g7192),.A(g7026),.B(g3526));
  AND2 AND2_529(.VSS(VSS),.VDD(VDD),.Y(g7193),.A(g6911),.B(g1616));
  AND2 AND2_530(.VSS(VSS),.VDD(VDD),.Y(g7195),.A(g6984),.B(g4226));
  AND2 AND2_531(.VSS(VSS),.VDD(VDD),.Y(g7197),.A(g7093),.B(g5055));
  AND2 AND2_532(.VSS(VSS),.VDD(VDD),.Y(g7199),.A(g1467),.B(g7003));
  AND2 AND2_533(.VSS(VSS),.VDD(VDD),.Y(g7212),.A(g1053),.B(g7010));
  AND2 AND2_534(.VSS(VSS),.VDD(VDD),.Y(g7215),.A(g6111),.B(g6984));
  AND2 AND2_535(.VSS(VSS),.VDD(VDD),.Y(g7217),.A(g1142),.B(g6941));
  AND2 AND2_536(.VSS(VSS),.VDD(VDD),.Y(g7228),.A(g6688),.B(g7090));
  AND2 AND2_537(.VSS(VSS),.VDD(VDD),.Y(g7232),.A(g6694),.B(g7091));
  AND2 AND2_538(.VSS(VSS),.VDD(VDD),.Y(g7235),.A(g6699),.B(g7094));
  AND2 AND2_539(.VSS(VSS),.VDD(VDD),.Y(g7238),.A(g6707),.B(g7098));
  AND2 AND2_540(.VSS(VSS),.VDD(VDD),.Y(g7240),.A(g6719),.B(g6894));
  AND2 AND2_541(.VSS(VSS),.VDD(VDD),.Y(g7242),.A(g7081),.B(g6899));
  AND2 AND2_542(.VSS(VSS),.VDD(VDD),.Y(g7252),.A(g3591),.B(g6977));
  AND2 AND2_543(.VSS(VSS),.VDD(VDD),.Y(g7271),.A(g6436),.B(g6922));
  AND2 AND2_544(.VSS(VSS),.VDD(VDD),.Y(g7278),.A(g6965),.B(g1745));
  AND2 AND2_545(.VSS(VSS),.VDD(VDD),.Y(g7282),.A(g5830),.B(g6939));
  AND2 AND2_546(.VSS(VSS),.VDD(VDD),.Y(g7323),.A(g4065),.B(g7171));
  AND2 AND2_547(.VSS(VSS),.VDD(VDD),.Y(g7412),.A(g7121),.B(g4841));
  AND2 AND2_548(.VSS(VSS),.VDD(VDD),.Y(g7415),.A(g7222),.B(g5603));
  AND2 AND2_549(.VSS(VSS),.VDD(VDD),.Y(g7416),.A(g7140),.B(g4969));
  AND2 AND2_550(.VSS(VSS),.VDD(VDD),.Y(g7417),.A(g7144),.B(g1616));
  AND2 AND2_551(.VSS(VSS),.VDD(VDD),.Y(g7419),.A(g7230),.B(g3530));
  AND2 AND2_552(.VSS(VSS),.VDD(VDD),.Y(g7427),.A(g1472),.B(g7199));
  AND2 AND2_553(.VSS(VSS),.VDD(VDD),.Y(g7429),.A(g1057),.B(g7212));
  AND2 AND2_554(.VSS(VSS),.VDD(VDD),.Y(g7449),.A(g7272),.B(g6901));
  AND2 AND2_555(.VSS(VSS),.VDD(VDD),.Y(g7536),.A(g4414),.B(g7367));
  AND2 AND2_556(.VSS(VSS),.VDD(VDD),.Y(g7537),.A(g7363),.B(g7411));
  AND2 AND2_557(.VSS(VSS),.VDD(VDD),.Y(g7552),.A(g7319),.B(g5749));
  AND2 AND2_558(.VSS(VSS),.VDD(VDD),.Y(g7553),.A(g7367),.B(g4135));
  AND2 AND2_559(.VSS(VSS),.VDD(VDD),.Y(g7554),.A(g7367),.B(g4139));
  AND2 AND2_560(.VSS(VSS),.VDD(VDD),.Y(g7557),.A(g7367),.B(g4147));
  AND2 AND2_561(.VSS(VSS),.VDD(VDD),.Y(g7559),.A(g7367),.B(g4155));
  AND2 AND2_562(.VSS(VSS),.VDD(VDD),.Y(g7561),.A(g7367),.B(g4163));
  AND2 AND2_563(.VSS(VSS),.VDD(VDD),.Y(g7564),.A(g7367),.B(g4172));
  AND2 AND2_564(.VSS(VSS),.VDD(VDD),.Y(g7596),.A(g7428),.B(g7028));
  AND2 AND2_565(.VSS(VSS),.VDD(VDD),.Y(g7597),.A(g7316),.B(g4841));
  AND2 AND2_566(.VSS(VSS),.VDD(VDD),.Y(g7598),.A(g7483),.B(g3466));
  AND2 AND2_567(.VSS(VSS),.VDD(VDD),.Y(g7600),.A(g7460),.B(g3466));
  AND2 AND2_568(.VSS(VSS),.VDD(VDD),.Y(g7602),.A(g7476),.B(g3466));
  AND2 AND2_569(.VSS(VSS),.VDD(VDD),.Y(g7604),.A(g7456),.B(g3466));
  AND2 AND2_570(.VSS(VSS),.VDD(VDD),.Y(g7605),.A(g7435),.B(g5607));
  AND2 AND2_571(.VSS(VSS),.VDD(VDD),.Y(g7606),.A(g7471),.B(g3466));
  AND2 AND2_572(.VSS(VSS),.VDD(VDD),.Y(g7607),.A(g7325),.B(g4969));
  AND2 AND2_573(.VSS(VSS),.VDD(VDD),.Y(g7608),.A(g7367),.B(g4169));
  AND2 AND2_574(.VSS(VSS),.VDD(VDD),.Y(g7609),.A(g7467),.B(g3466));
  AND2 AND2_575(.VSS(VSS),.VDD(VDD),.Y(g7611),.A(g7367),.B(g4507));
  AND2 AND2_576(.VSS(VSS),.VDD(VDD),.Y(g7614),.A(g7367),.B(g4176));
  AND2 AND2_577(.VSS(VSS),.VDD(VDD),.Y(g7615),.A(g7488),.B(g3466));
  AND2 AND2_578(.VSS(VSS),.VDD(VDD),.Y(g7616),.A(g7367),.B(g4517));
  AND2 AND2_579(.VSS(VSS),.VDD(VDD),.Y(g7625),.A(g7367),.B(g4182));
  AND2 AND2_580(.VSS(VSS),.VDD(VDD),.Y(g7626),.A(g7463),.B(g3466));
  AND2 AND2_581(.VSS(VSS),.VDD(VDD),.Y(g7628),.A(g7367),.B(g4532));
  AND2 AND2_582(.VSS(VSS),.VDD(VDD),.Y(g7631),.A(g7367),.B(g4187));
  AND2 AND2_583(.VSS(VSS),.VDD(VDD),.Y(g7632),.A(g7445),.B(g3548));
  AND2 AND2_584(.VSS(VSS),.VDD(VDD),.Y(g7634),.A(g7367),.B(g4549));
  AND2 AND2_585(.VSS(VSS),.VDD(VDD),.Y(g7652),.A(g7367),.B(g4194));
  AND2 AND2_586(.VSS(VSS),.VDD(VDD),.Y(g7653),.A(g7480),.B(g5754));
  AND2 AND2_587(.VSS(VSS),.VDD(VDD),.Y(g7654),.A(g7367),.B(g4142));
  AND2 AND2_588(.VSS(VSS),.VDD(VDD),.Y(g7657),.A(g7367),.B(g4201));
  AND2 AND2_589(.VSS(VSS),.VDD(VDD),.Y(g7658),.A(g7367),.B(g4150));
  AND2 AND2_590(.VSS(VSS),.VDD(VDD),.Y(g7676),.A(g7367),.B(g4216));
  AND2 AND2_591(.VSS(VSS),.VDD(VDD),.Y(g7677),.A(g7503),.B(g5073));
  AND2 AND2_592(.VSS(VSS),.VDD(VDD),.Y(g7678),.A(g7367),.B(g4158));
  AND2 AND2_593(.VSS(VSS),.VDD(VDD),.Y(g7679),.A(g7447),.B(g5084));
  AND2 AND2_594(.VSS(VSS),.VDD(VDD),.Y(g7680),.A(g7367),.B(g4166));
  AND2 AND2_595(.VSS(VSS),.VDD(VDD),.Y(g7681),.A(g7444),.B(g5099));
  AND2 AND2_596(.VSS(VSS),.VDD(VDD),.Y(g7683),.A(g1061),.B(g7429));
  AND2 AND2_597(.VSS(VSS),.VDD(VDD),.Y(g7689),.A(g7367),.B(g4417));
  AND2 AND2_598(.VSS(VSS),.VDD(VDD),.Y(g7691),.A(g7367),.B(g4427));
  AND2 AND2_599(.VSS(VSS),.VDD(VDD),.Y(g7692),.A(g7367),.B(g4430));
  AND2 AND2_600(.VSS(VSS),.VDD(VDD),.Y(g7693),.A(g7367),.B(g4445));
  AND2 AND2_601(.VSS(VSS),.VDD(VDD),.Y(g7694),.A(g7367),.B(g4448));
  AND2 AND2_602(.VSS(VSS),.VDD(VDD),.Y(g7695),.A(g7367),.B(g4466));
  AND2 AND2_603(.VSS(VSS),.VDD(VDD),.Y(g7696),.A(g7367),.B(g4469));
  AND2 AND2_604(.VSS(VSS),.VDD(VDD),.Y(g7698),.A(g7367),.B(g4483));
  AND2 AND2_605(.VSS(VSS),.VDD(VDD),.Y(g7699),.A(g7367),.B(g4486));
  AND2 AND2_606(.VSS(VSS),.VDD(VDD),.Y(g7700),.A(g7367),.B(g4494));
  AND2 AND2_607(.VSS(VSS),.VDD(VDD),.Y(g7701),.A(g7367),.B(g4497));
  AND2 AND2_608(.VSS(VSS),.VDD(VDD),.Y(g7703),.A(g7367),.B(g4504));
  AND2 AND2_609(.VSS(VSS),.VDD(VDD),.Y(g7705),.A(g7367),.B(g4514));
  AND2 AND2_610(.VSS(VSS),.VDD(VDD),.Y(g7709),.A(g7367),.B(g4529));
  AND2 AND2_611(.VSS(VSS),.VDD(VDD),.Y(g7713),.A(g4403),.B(g7367));
  AND2 AND2_612(.VSS(VSS),.VDD(VDD),.Y(g7724),.A(g7337),.B(g5938));
  AND2 AND2_613(.VSS(VSS),.VDD(VDD),.Y(g7827),.A(g7575),.B(g7173));
  AND2 AND2_614(.VSS(VSS),.VDD(VDD),.Y(g7832),.A(g5343),.B(g7599));
  AND2 AND2_615(.VSS(VSS),.VDD(VDD),.Y(g7833),.A(g6461),.B(g7601));
  AND2 AND2_616(.VSS(VSS),.VDD(VDD),.Y(g7837),.A(g6470),.B(g7610));
  AND2 AND2_617(.VSS(VSS),.VDD(VDD),.Y(g8059),.A(g7682),.B(g7032));
  AND2 AND2_618(.VSS(VSS),.VDD(VDD),.Y(g8060),.A(g7535),.B(g4841));
  AND2 AND2_619(.VSS(VSS),.VDD(VDD),.Y(g8062),.A(g7476),.B(g7634));
  AND2 AND2_620(.VSS(VSS),.VDD(VDD),.Y(g8064),.A(g7483),.B(g7634));
  AND2 AND2_621(.VSS(VSS),.VDD(VDD),.Y(g8066),.A(g7488),.B(g7634));
  AND2 AND2_622(.VSS(VSS),.VDD(VDD),.Y(g8068),.A(g7687),.B(g5610));
  AND2 AND2_623(.VSS(VSS),.VDD(VDD),.Y(g8069),.A(g7456),.B(g7634));
  AND2 AND2_624(.VSS(VSS),.VDD(VDD),.Y(g8070),.A(g863),.B(g7616));
  AND2 AND2_625(.VSS(VSS),.VDD(VDD),.Y(g8071),.A(g7540),.B(g4969));
  AND2 AND2_626(.VSS(VSS),.VDD(VDD),.Y(g8074),.A(g855),.B(g7616));
  AND2 AND2_627(.VSS(VSS),.VDD(VDD),.Y(g8075),.A(g7460),.B(g7634));
  AND2 AND2_628(.VSS(VSS),.VDD(VDD),.Y(g8076),.A(g7690),.B(g3521));
  AND2 AND2_629(.VSS(VSS),.VDD(VDD),.Y(g8077),.A(g859),.B(g7616));
  AND2 AND2_630(.VSS(VSS),.VDD(VDD),.Y(g8078),.A(g7463),.B(g7634));
  AND2 AND2_631(.VSS(VSS),.VDD(VDD),.Y(g8079),.A(g831),.B(g7658));
  AND2 AND2_632(.VSS(VSS),.VDD(VDD),.Y(g8080),.A(g7467),.B(g7634));
  AND2 AND2_633(.VSS(VSS),.VDD(VDD),.Y(g8081),.A(g834),.B(g7658));
  AND2 AND2_634(.VSS(VSS),.VDD(VDD),.Y(g8087),.A(g7471),.B(g7634));
  AND2 AND2_635(.VSS(VSS),.VDD(VDD),.Y(g8088),.A(g837),.B(g7658));
  AND2 AND2_636(.VSS(VSS),.VDD(VDD),.Y(g8089),.A(g840),.B(g7658));
  AND2 AND2_637(.VSS(VSS),.VDD(VDD),.Y(g8090),.A(g843),.B(g7658));
  AND2 AND2_638(.VSS(VSS),.VDD(VDD),.Y(g8147),.A(g1065),.B(g7683));
  AND2 AND2_639(.VSS(VSS),.VDD(VDD),.Y(g8150),.A(g846),.B(g7658));
  AND2 AND2_640(.VSS(VSS),.VDD(VDD),.Y(g8151),.A(g849),.B(g7658));
  AND2 AND2_641(.VSS(VSS),.VDD(VDD),.Y(g8153),.A(g852),.B(g7658));
  AND2 AND2_642(.VSS(VSS),.VDD(VDD),.Y(g8229),.A(g8180),.B(g5680));
  AND2 AND2_643(.VSS(VSS),.VDD(VDD),.Y(g8237),.A(g89),.B(g8131));
  AND2 AND2_644(.VSS(VSS),.VDD(VDD),.Y(g8238),.A(g100),.B(g8131));
  AND2 AND2_645(.VSS(VSS),.VDD(VDD),.Y(g8256),.A(g95),.B(g8131));
  AND2 AND2_646(.VSS(VSS),.VDD(VDD),.Y(g8257),.A(g146),.B(g8042));
  AND2 AND2_647(.VSS(VSS),.VDD(VDD),.Y(g8258),.A(g142),.B(g8111));
  AND2 AND2_648(.VSS(VSS),.VDD(VDD),.Y(g8259),.A(g4538),.B(g7855));
  AND2 AND2_649(.VSS(VSS),.VDD(VDD),.Y(g8260),.A(g138),.B(g8111));
  AND2 AND2_650(.VSS(VSS),.VDD(VDD),.Y(g8261),.A(g174),.B(g8042));
  AND2 AND2_651(.VSS(VSS),.VDD(VDD),.Y(g8262),.A(g4554),.B(g7855));
  AND2 AND2_652(.VSS(VSS),.VDD(VDD),.Y(g8263),.A(g4555),.B(g7905));
  AND2 AND2_653(.VSS(VSS),.VDD(VDD),.Y(g8264),.A(g105),.B(g8131));
  AND2 AND2_654(.VSS(VSS),.VDD(VDD),.Y(g8265),.A(g134),.B(g8111));
  AND2 AND2_655(.VSS(VSS),.VDD(VDD),.Y(g8266),.A(g2157),.B(g8042));
  AND2 AND2_656(.VSS(VSS),.VDD(VDD),.Y(g8267),.A(g154),.B(g8042));
  AND2 AND2_657(.VSS(VSS),.VDD(VDD),.Y(g8268),.A(g4568),.B(g7905));
  AND2 AND2_658(.VSS(VSS),.VDD(VDD),.Y(g8269),.A(g4569),.B(g7951));
  AND2 AND2_659(.VSS(VSS),.VDD(VDD),.Y(g8270),.A(g110),.B(g8131));
  AND2 AND2_660(.VSS(VSS),.VDD(VDD),.Y(g8271),.A(g130),.B(g8111));
  AND2 AND2_661(.VSS(VSS),.VDD(VDD),.Y(g8272),.A(g158),.B(g8042));
  AND2 AND2_662(.VSS(VSS),.VDD(VDD),.Y(g8273),.A(g185),.B(g8156));
  AND2 AND2_663(.VSS(VSS),.VDD(VDD),.Y(g8274),.A(g4580),.B(g7951));
  AND2 AND2_664(.VSS(VSS),.VDD(VDD),.Y(g8275),.A(g4581),.B(g7993));
  AND2 AND2_665(.VSS(VSS),.VDD(VDD),.Y(g8276),.A(g150),.B(g8042));
  AND2 AND2_666(.VSS(VSS),.VDD(VDD),.Y(g8277),.A(g162),.B(g8042));
  AND2 AND2_667(.VSS(VSS),.VDD(VDD),.Y(g8278),.A(g4589),.B(g7993));
  AND2 AND2_668(.VSS(VSS),.VDD(VDD),.Y(g8280),.A(g114),.B(g8111));
  AND2 AND2_669(.VSS(VSS),.VDD(VDD),.Y(g8281),.A(g168),.B(g8042));
  AND2 AND2_670(.VSS(VSS),.VDD(VDD),.Y(g8282),.A(g179),.B(g8156));
  AND2 AND2_671(.VSS(VSS),.VDD(VDD),.Y(g8283),.A(g267),.B(g7838));
  AND2 AND2_672(.VSS(VSS),.VDD(VDD),.Y(g8285),.A(g118),.B(g8111));
  AND2 AND2_673(.VSS(VSS),.VDD(VDD),.Y(g8286),.A(g180),.B(g8156));
  AND2 AND2_674(.VSS(VSS),.VDD(VDD),.Y(g8287),.A(g4500),.B(g7855));
  AND2 AND2_675(.VSS(VSS),.VDD(VDD),.Y(g8288),.A(g270),.B(g7838));
  AND2 AND2_676(.VSS(VSS),.VDD(VDD),.Y(g8289),.A(g348),.B(g7870));
  AND2 AND2_677(.VSS(VSS),.VDD(VDD),.Y(g8290),.A(g588),.B(g8181));
  AND2 AND2_678(.VSS(VSS),.VDD(VDD),.Y(g8291),.A(g122),.B(g8111));
  AND2 AND2_679(.VSS(VSS),.VDD(VDD),.Y(g8292),.A(g181),.B(g8156));
  AND2 AND2_680(.VSS(VSS),.VDD(VDD),.Y(g8293),.A(g4510),.B(g7855));
  AND2 AND2_681(.VSS(VSS),.VDD(VDD),.Y(g8294),.A(g281),.B(g7838));
  AND2 AND2_682(.VSS(VSS),.VDD(VDD),.Y(g8295),.A(g4512),.B(g7905));
  AND2 AND2_683(.VSS(VSS),.VDD(VDD),.Y(g8296),.A(g351),.B(g7870));
  AND2 AND2_684(.VSS(VSS),.VDD(VDD),.Y(g8297),.A(g429),.B(g7920));
  AND2 AND2_685(.VSS(VSS),.VDD(VDD),.Y(g8298),.A(g553),.B(g8181));
  AND2 AND2_686(.VSS(VSS),.VDD(VDD),.Y(g8299),.A(g591),.B(g8181));
  AND2 AND2_687(.VSS(VSS),.VDD(VDD),.Y(g8300),.A(g126),.B(g8111));
  AND2 AND2_688(.VSS(VSS),.VDD(VDD),.Y(g8301),.A(g182),.B(g8156));
  AND2 AND2_689(.VSS(VSS),.VDD(VDD),.Y(g8302),.A(g4521),.B(g7855));
  AND2 AND2_690(.VSS(VSS),.VDD(VDD),.Y(g8303),.A(g284),.B(g7838));
  AND2 AND2_691(.VSS(VSS),.VDD(VDD),.Y(g8304),.A(g4523),.B(g7905));
  AND2 AND2_692(.VSS(VSS),.VDD(VDD),.Y(g8305),.A(g362),.B(g7870));
  AND2 AND2_693(.VSS(VSS),.VDD(VDD),.Y(g8306),.A(g4525),.B(g7951));
  AND2 AND2_694(.VSS(VSS),.VDD(VDD),.Y(g8307),.A(g432),.B(g7920));
  AND2 AND2_695(.VSS(VSS),.VDD(VDD),.Y(g8308),.A(g510),.B(g7966));
  AND2 AND2_696(.VSS(VSS),.VDD(VDD),.Y(g8309),.A(g550),.B(g8181));
  AND2 AND2_697(.VSS(VSS),.VDD(VDD),.Y(g8310),.A(g573),.B(g8181));
  AND2 AND2_698(.VSS(VSS),.VDD(VDD),.Y(g8311),.A(g4540),.B(g7905));
  AND2 AND2_699(.VSS(VSS),.VDD(VDD),.Y(g8312),.A(g365),.B(g7870));
  AND2 AND2_700(.VSS(VSS),.VDD(VDD),.Y(g8313),.A(g4542),.B(g7951));
  AND2 AND2_701(.VSS(VSS),.VDD(VDD),.Y(g8314),.A(g443),.B(g7920));
  AND2 AND2_702(.VSS(VSS),.VDD(VDD),.Y(g8315),.A(g4544),.B(g7993));
  AND2 AND2_703(.VSS(VSS),.VDD(VDD),.Y(g8316),.A(g513),.B(g7966));
  AND2 AND2_704(.VSS(VSS),.VDD(VDD),.Y(g8317),.A(g547),.B(g8181));
  AND2 AND2_705(.VSS(VSS),.VDD(VDD),.Y(g8318),.A(g183),.B(g8156));
  AND2 AND2_706(.VSS(VSS),.VDD(VDD),.Y(g8319),.A(g255),.B(g7838));
  AND2 AND2_707(.VSS(VSS),.VDD(VDD),.Y(g8320),.A(g4557),.B(g7951));
  AND2 AND2_708(.VSS(VSS),.VDD(VDD),.Y(g8321),.A(g446),.B(g7920));
  AND2 AND2_709(.VSS(VSS),.VDD(VDD),.Y(g8322),.A(g4559),.B(g7993));
  AND2 AND2_710(.VSS(VSS),.VDD(VDD),.Y(g8323),.A(g524),.B(g7966));
  AND2 AND2_711(.VSS(VSS),.VDD(VDD),.Y(g8325),.A(g184),.B(g8156));
  AND2 AND2_712(.VSS(VSS),.VDD(VDD),.Y(g8326),.A(g258),.B(g7838));
  AND2 AND2_713(.VSS(VSS),.VDD(VDD),.Y(g8327),.A(g336),.B(g7870));
  AND2 AND2_714(.VSS(VSS),.VDD(VDD),.Y(g8328),.A(g4571),.B(g7993));
  AND2 AND2_715(.VSS(VSS),.VDD(VDD),.Y(g8329),.A(g527),.B(g7966));
  AND2 AND2_716(.VSS(VSS),.VDD(VDD),.Y(g8330),.A(g261),.B(g7838));
  AND2 AND2_717(.VSS(VSS),.VDD(VDD),.Y(g8331),.A(g339),.B(g7870));
  AND2 AND2_718(.VSS(VSS),.VDD(VDD),.Y(g8332),.A(g417),.B(g7920));
  AND2 AND2_719(.VSS(VSS),.VDD(VDD),.Y(g8333),.A(g563),.B(g8181));
  AND2 AND2_720(.VSS(VSS),.VDD(VDD),.Y(g8334),.A(g264),.B(g7838));
  AND2 AND2_721(.VSS(VSS),.VDD(VDD),.Y(g8335),.A(g342),.B(g7870));
  AND2 AND2_722(.VSS(VSS),.VDD(VDD),.Y(g8336),.A(g420),.B(g7920));
  AND2 AND2_723(.VSS(VSS),.VDD(VDD),.Y(g8337),.A(g498),.B(g7966));
  AND2 AND2_724(.VSS(VSS),.VDD(VDD),.Y(g8338),.A(g570),.B(g8181));
  AND2 AND2_725(.VSS(VSS),.VDD(VDD),.Y(g8339),.A(g345),.B(g7870));
  AND2 AND2_726(.VSS(VSS),.VDD(VDD),.Y(g8340),.A(g423),.B(g7920));
  AND2 AND2_727(.VSS(VSS),.VDD(VDD),.Y(g8341),.A(g501),.B(g7966));
  AND2 AND2_728(.VSS(VSS),.VDD(VDD),.Y(g8359),.A(g642),.B(g7793));
  AND2 AND2_729(.VSS(VSS),.VDD(VDD),.Y(g8361),.A(g426),.B(g7920));
  AND2 AND2_730(.VSS(VSS),.VDD(VDD),.Y(g8362),.A(g504),.B(g7966));
  AND2 AND2_731(.VSS(VSS),.VDD(VDD),.Y(g8377),.A(g507),.B(g7966));
  AND2 AND2_732(.VSS(VSS),.VDD(VDD),.Y(g8378),.A(g677),.B(g7887));
  AND2 AND2_733(.VSS(VSS),.VDD(VDD),.Y(g8379),.A(g691),.B(g7793));
  AND2 AND2_734(.VSS(VSS),.VDD(VDD),.Y(g8380),.A(g681),.B(g7887));
  AND2 AND2_735(.VSS(VSS),.VDD(VDD),.Y(g8382),.A(g685),.B(g7887));
  AND2 AND2_736(.VSS(VSS),.VDD(VDD),.Y(g8383),.A(g730),.B(g7937));
  AND2 AND2_737(.VSS(VSS),.VDD(VDD),.Y(g8384),.A(g636),.B(g7793));
  AND2 AND2_738(.VSS(VSS),.VDD(VDD),.Y(g8385),.A(g695),.B(g7811));
  AND2 AND2_739(.VSS(VSS),.VDD(VDD),.Y(g8403),.A(g639),.B(g7793));
  AND2 AND2_740(.VSS(VSS),.VDD(VDD),.Y(g8404),.A(g710),.B(g7937));
  AND2 AND2_741(.VSS(VSS),.VDD(VDD),.Y(g8405),.A(g741),.B(g8018));
  AND2 AND2_742(.VSS(VSS),.VDD(VDD),.Y(g8438),.A(g649),.B(g7793));
  AND2 AND2_743(.VSS(VSS),.VDD(VDD),.Y(g8439),.A(g699),.B(g7811));
  AND2 AND2_744(.VSS(VSS),.VDD(VDD),.Y(g8440),.A(g714),.B(g7937));
  AND2 AND2_745(.VSS(VSS),.VDD(VDD),.Y(g8441),.A(g746),.B(g8018));
  AND2 AND2_746(.VSS(VSS),.VDD(VDD),.Y(g8455),.A(g652),.B(g7793));
  AND2 AND2_747(.VSS(VSS),.VDD(VDD),.Y(g8456),.A(g703),.B(g7811));
  AND2 AND2_748(.VSS(VSS),.VDD(VDD),.Y(g8457),.A(g724),.B(g7811));
  AND2 AND2_749(.VSS(VSS),.VDD(VDD),.Y(g8458),.A(g756),.B(g8199));
  AND2 AND2_750(.VSS(VSS),.VDD(VDD),.Y(g8459),.A(g655),.B(g7793));
  AND2 AND2_751(.VSS(VSS),.VDD(VDD),.Y(g8460),.A(g757),.B(g8199));
  AND2 AND2_752(.VSS(VSS),.VDD(VDD),.Y(g8461),.A(g658),.B(g7793));
  AND2 AND2_753(.VSS(VSS),.VDD(VDD),.Y(g8462),.A(g49),.B(g8199));
  AND2 AND2_754(.VSS(VSS),.VDD(VDD),.Y(g8513),.A(g718),.B(g7937));
  AND2 AND2_755(.VSS(VSS),.VDD(VDD),.Y(g8542),.A(g661),.B(g7887));
  AND2 AND2_756(.VSS(VSS),.VDD(VDD),.Y(g8543),.A(g706),.B(g7887));
  AND2 AND2_757(.VSS(VSS),.VDD(VDD),.Y(g8584),.A(g8146),.B(g7034));
  AND2 AND2_758(.VSS(VSS),.VDD(VDD),.Y(g8607),.A(g8154),.B(g5616));
  AND2 AND2_759(.VSS(VSS),.VDD(VDD),.Y(g8609),.A(g7828),.B(g4969));
  AND2 AND2_760(.VSS(VSS),.VDD(VDD),.Y(g8610),.A(g665),.B(g7887));
  AND2 AND2_761(.VSS(VSS),.VDD(VDD),.Y(g8611),.A(g669),.B(g7887));
  AND2 AND2_762(.VSS(VSS),.VDD(VDD),.Y(g8612),.A(g673),.B(g7887));
  AND2 AND2_763(.VSS(VSS),.VDD(VDD),.Y(g8620),.A(g751),.B(g8199));
  AND2 AND2_764(.VSS(VSS),.VDD(VDD),.Y(g8621),.A(g734),.B(g7937));
  AND2 AND2_765(.VSS(VSS),.VDD(VDD),.Y(g8622),.A(g738),.B(g7811));
  AND2 AND2_766(.VSS(VSS),.VDD(VDD),.Y(g8623),.A(g755),.B(g8199));
  AND2 AND2_767(.VSS(VSS),.VDD(VDD),.Y(g8624),.A(g754),.B(g8199));
  AND2 AND2_768(.VSS(VSS),.VDD(VDD),.Y(g8626),.A(g752),.B(g8199));
  AND2 AND2_769(.VSS(VSS),.VDD(VDD),.Y(g8628),.A(g753),.B(g8199));
  AND2 AND2_770(.VSS(VSS),.VDD(VDD),.Y(g8643),.A(g547),.B(g8094));
  AND2 AND2_771(.VSS(VSS),.VDD(VDD),.Y(g8645),.A(g550),.B(g8094));
  AND2 AND2_772(.VSS(VSS),.VDD(VDD),.Y(g8646),.A(g553),.B(g8094));
  AND2 AND2_773(.VSS(VSS),.VDD(VDD),.Y(g8648),.A(g588),.B(g8094));
  AND2 AND2_774(.VSS(VSS),.VDD(VDD),.Y(g8650),.A(g591),.B(g8094));
  AND2 AND2_775(.VSS(VSS),.VDD(VDD),.Y(g8652),.A(g563),.B(g8094));
  AND2 AND2_776(.VSS(VSS),.VDD(VDD),.Y(g8653),.A(g573),.B(g8094));
  AND2 AND2_777(.VSS(VSS),.VDD(VDD),.Y(g8654),.A(g570),.B(g8094));
  AND2 AND2_778(.VSS(VSS),.VDD(VDD),.Y(g8660),.A(g1069),.B(g8147));
  AND2 AND2_779(.VSS(VSS),.VDD(VDD),.Y(g8686),.A(g3819),.B(g8342));
  AND2 AND2_780(.VSS(VSS),.VDD(VDD),.Y(g8687),.A(g3488),.B(g8363));
  AND2 AND2_781(.VSS(VSS),.VDD(VDD),.Y(g8688),.A(g3812),.B(g8342));
  AND2 AND2_782(.VSS(VSS),.VDD(VDD),.Y(g8690),.A(g3485),.B(g8363));
  AND2 AND2_783(.VSS(VSS),.VDD(VDD),.Y(g8691),.A(g3805),.B(g8342));
  AND2 AND2_784(.VSS(VSS),.VDD(VDD),.Y(g8692),.A(g3462),.B(g8363));
  AND2 AND2_785(.VSS(VSS),.VDD(VDD),.Y(g8693),.A(g3798),.B(g8342));
  AND2 AND2_786(.VSS(VSS),.VDD(VDD),.Y(g8695),.A(g2709),.B(g8363));
  AND2 AND2_787(.VSS(VSS),.VDD(VDD),.Y(g8696),.A(g3743),.B(g8342));
  AND2 AND2_788(.VSS(VSS),.VDD(VDD),.Y(g8697),.A(g3761),.B(g8342));
  AND2 AND2_789(.VSS(VSS),.VDD(VDD),.Y(g8698),.A(g3774),.B(g8342));
  AND2 AND2_790(.VSS(VSS),.VDD(VDD),.Y(g8700),.A(g3784),.B(g8342));
  AND2 AND2_791(.VSS(VSS),.VDD(VDD),.Y(g8701),.A(g2700),.B(g8363));
  AND2 AND2_792(.VSS(VSS),.VDD(VDD),.Y(g8702),.A(g2837),.B(g8386));
  AND2 AND2_793(.VSS(VSS),.VDD(VDD),.Y(g8703),.A(g3574),.B(g8407));
  AND2 AND2_794(.VSS(VSS),.VDD(VDD),.Y(g8704),.A(g2829),.B(g8386));
  AND2 AND2_795(.VSS(VSS),.VDD(VDD),.Y(g8705),.A(g2798),.B(g8421));
  AND2 AND2_796(.VSS(VSS),.VDD(VDD),.Y(g8708),.A(g3557),.B(g8407));
  AND2 AND2_797(.VSS(VSS),.VDD(VDD),.Y(g8709),.A(g2818),.B(g8386));
  AND2 AND2_798(.VSS(VSS),.VDD(VDD),.Y(g8710),.A(g2790),.B(g8421));
  AND2 AND2_799(.VSS(VSS),.VDD(VDD),.Y(g8711),.A(g3542),.B(g8407));
  AND2 AND2_800(.VSS(VSS),.VDD(VDD),.Y(g8712),.A(g2804),.B(g8386));
  AND2 AND2_801(.VSS(VSS),.VDD(VDD),.Y(g8713),.A(g2777),.B(g8421));
  AND2 AND2_802(.VSS(VSS),.VDD(VDD),.Y(g8714),.A(g2873),.B(g8407));
  AND2 AND2_803(.VSS(VSS),.VDD(VDD),.Y(g8715),.A(g2761),.B(g8386));
  AND2 AND2_804(.VSS(VSS),.VDD(VDD),.Y(g8716),.A(g3506),.B(g8443));
  AND2 AND2_805(.VSS(VSS),.VDD(VDD),.Y(g8717),.A(g2764),.B(g8421));
  AND2 AND2_806(.VSS(VSS),.VDD(VDD),.Y(g8718),.A(g2774),.B(g8386));
  AND2 AND2_807(.VSS(VSS),.VDD(VDD),.Y(g8719),.A(g2821),.B(g8443));
  AND2 AND2_808(.VSS(VSS),.VDD(VDD),.Y(g8720),.A(g3825),.B(g8421));
  AND2 AND2_809(.VSS(VSS),.VDD(VDD),.Y(g8721),.A(g2703),.B(g8464));
  AND2 AND2_810(.VSS(VSS),.VDD(VDD),.Y(g8722),.A(g2787),.B(g8386));
  AND2 AND2_811(.VSS(VSS),.VDD(VDD),.Y(g8723),.A(g2706),.B(g8421));
  AND2 AND2_812(.VSS(VSS),.VDD(VDD),.Y(g8724),.A(g3822),.B(g8464));
  AND2 AND2_813(.VSS(VSS),.VDD(VDD),.Y(g8725),.A(g3008),.B(g8493));
  AND2 AND2_814(.VSS(VSS),.VDD(VDD),.Y(g8726),.A(g2795),.B(g8386));
  AND2 AND2_815(.VSS(VSS),.VDD(VDD),.Y(g8727),.A(g2724),.B(g8421));
  AND2 AND2_816(.VSS(VSS),.VDD(VDD),.Y(g8728),.A(g3815),.B(g8464));
  AND2 AND2_817(.VSS(VSS),.VDD(VDD),.Y(g8729),.A(g2999),.B(g8493));
  AND2 AND2_818(.VSS(VSS),.VDD(VDD),.Y(g8730),.A(g2863),.B(g8407));
  AND2 AND2_819(.VSS(VSS),.VDD(VDD),.Y(g8731),.A(g2743),.B(g8421));
  AND2 AND2_820(.VSS(VSS),.VDD(VDD),.Y(g8732),.A(g3808),.B(g8464));
  AND2 AND2_821(.VSS(VSS),.VDD(VDD),.Y(g8733),.A(g2996),.B(g8493));
  AND2 AND2_822(.VSS(VSS),.VDD(VDD),.Y(g8735),.A(g2807),.B(g8443));
  AND2 AND2_823(.VSS(VSS),.VDD(VDD),.Y(g8736),.A(g3771),.B(g8464));
  AND2 AND2_824(.VSS(VSS),.VDD(VDD),.Y(g8737),.A(g2992),.B(g8493));
  AND2 AND2_825(.VSS(VSS),.VDD(VDD),.Y(g8738),.A(g8619),.B(g3338));
  AND2 AND2_826(.VSS(VSS),.VDD(VDD),.Y(g8739),.A(g3780),.B(g8464));
  AND2 AND2_827(.VSS(VSS),.VDD(VDD),.Y(g8740),.A(g2966),.B(g8493));
  AND2 AND2_828(.VSS(VSS),.VDD(VDD),.Y(g8741),.A(g3787),.B(g8464));
  AND2 AND2_829(.VSS(VSS),.VDD(VDD),.Y(g8742),.A(g2973),.B(g8493));
  AND2 AND2_830(.VSS(VSS),.VDD(VDD),.Y(g8744),.A(g3802),.B(g8464));
  AND2 AND2_831(.VSS(VSS),.VDD(VDD),.Y(g8745),.A(g2982),.B(g8493));
  AND2 AND2_832(.VSS(VSS),.VDD(VDD),.Y(g8748),.A(g2721),.B(g8483));
  AND2 AND2_833(.VSS(VSS),.VDD(VDD),.Y(g8749),.A(g2989),.B(g8493));
  AND2 AND2_834(.VSS(VSS),.VDD(VDD),.Y(g8764),.A(g8231),.B(g4969));
  AND2 AND2_835(.VSS(VSS),.VDD(VDD),.Y(g8779),.A(g8634),.B(g7037));
  AND2 AND2_836(.VSS(VSS),.VDD(VDD),.Y(g8793),.A(g8637),.B(g5622));
  AND2 AND2_837(.VSS(VSS),.VDD(VDD),.Y(g8813),.A(g255),.B(g8524));
  AND2 AND2_838(.VSS(VSS),.VDD(VDD),.Y(g8814),.A(g3880),.B(g8463));
  AND2 AND2_839(.VSS(VSS),.VDD(VDD),.Y(g8815),.A(g258),.B(g8524));
  AND2 AND2_840(.VSS(VSS),.VDD(VDD),.Y(g8816),.A(g336),.B(g8545));
  AND2 AND2_841(.VSS(VSS),.VDD(VDD),.Y(g8817),.A(g4545),.B(g8482));
  AND2 AND2_842(.VSS(VSS),.VDD(VDD),.Y(g8820),.A(g261),.B(g8524));
  AND2 AND2_843(.VSS(VSS),.VDD(VDD),.Y(g8821),.A(g339),.B(g8545));
  AND2 AND2_844(.VSS(VSS),.VDD(VDD),.Y(g8822),.A(g417),.B(g8564));
  AND2 AND2_845(.VSS(VSS),.VDD(VDD),.Y(g8823),.A(g4561),.B(g8512));
  AND2 AND2_846(.VSS(VSS),.VDD(VDD),.Y(g8824),.A(g264),.B(g8524));
  AND2 AND2_847(.VSS(VSS),.VDD(VDD),.Y(g8825),.A(g342),.B(g8545));
  AND2 AND2_848(.VSS(VSS),.VDD(VDD),.Y(g8826),.A(g420),.B(g8564));
  AND2 AND2_849(.VSS(VSS),.VDD(VDD),.Y(g8827),.A(g498),.B(g8585));
  AND2 AND2_850(.VSS(VSS),.VDD(VDD),.Y(g8828),.A(g4573),.B(g8541));
  AND2 AND2_851(.VSS(VSS),.VDD(VDD),.Y(g8829),.A(g267),.B(g8524));
  AND2 AND2_852(.VSS(VSS),.VDD(VDD),.Y(g8830),.A(g345),.B(g8545));
  AND2 AND2_853(.VSS(VSS),.VDD(VDD),.Y(g8831),.A(g423),.B(g8564));
  AND2 AND2_854(.VSS(VSS),.VDD(VDD),.Y(g8832),.A(g501),.B(g8585));
  AND2 AND2_855(.VSS(VSS),.VDD(VDD),.Y(g8833),.A(g4583),.B(g8562));
  AND2 AND2_856(.VSS(VSS),.VDD(VDD),.Y(g8835),.A(g270),.B(g8524));
  AND2 AND2_857(.VSS(VSS),.VDD(VDD),.Y(g8836),.A(g348),.B(g8545));
  AND2 AND2_858(.VSS(VSS),.VDD(VDD),.Y(g8837),.A(g426),.B(g8564));
  AND2 AND2_859(.VSS(VSS),.VDD(VDD),.Y(g8838),.A(g504),.B(g8585));
  AND2 AND2_860(.VSS(VSS),.VDD(VDD),.Y(g8839),.A(g4050),.B(g8581));
  AND2 AND2_861(.VSS(VSS),.VDD(VDD),.Y(g8840),.A(g4590),.B(g8582));
  AND2 AND2_862(.VSS(VSS),.VDD(VDD),.Y(g8841),.A(g351),.B(g8545));
  AND2 AND2_863(.VSS(VSS),.VDD(VDD),.Y(g8842),.A(g429),.B(g8564));
  AND2 AND2_864(.VSS(VSS),.VDD(VDD),.Y(g8843),.A(g507),.B(g8585));
  AND2 AND2_865(.VSS(VSS),.VDD(VDD),.Y(g8844),.A(g4056),.B(g8602));
  AND2 AND2_866(.VSS(VSS),.VDD(VDD),.Y(g8845),.A(g432),.B(g8564));
  AND2 AND2_867(.VSS(VSS),.VDD(VDD),.Y(g8846),.A(g510),.B(g8585));
  AND2 AND2_868(.VSS(VSS),.VDD(VDD),.Y(g8848),.A(g281),.B(g8524));
  AND2 AND2_869(.VSS(VSS),.VDD(VDD),.Y(g8849),.A(g513),.B(g8585));
  AND2 AND2_870(.VSS(VSS),.VDD(VDD),.Y(g8851),.A(g284),.B(g8524));
  AND2 AND2_871(.VSS(VSS),.VDD(VDD),.Y(g8852),.A(g362),.B(g8545));
  AND2 AND2_872(.VSS(VSS),.VDD(VDD),.Y(g8853),.A(g365),.B(g8545));
  AND2 AND2_873(.VSS(VSS),.VDD(VDD),.Y(g8854),.A(g443),.B(g8564));
  AND2 AND2_874(.VSS(VSS),.VDD(VDD),.Y(g8857),.A(g446),.B(g8564));
  AND2 AND2_875(.VSS(VSS),.VDD(VDD),.Y(g8858),.A(g524),.B(g8585));
  AND2 AND2_876(.VSS(VSS),.VDD(VDD),.Y(g8860),.A(g527),.B(g8585));
  AND2 AND2_877(.VSS(VSS),.VDD(VDD),.Y(g8876),.A(g8769),.B(g6102));
  AND2 AND2_878(.VSS(VSS),.VDD(VDD),.Y(g8877),.A(g8773),.B(g6104));
  AND2 AND2_879(.VSS(VSS),.VDD(VDD),.Y(g8878),.A(g8777),.B(g6106));
  AND2 AND2_880(.VSS(VSS),.VDD(VDD),.Y(g8879),.A(g8782),.B(g6108));
  AND2 AND2_881(.VSS(VSS),.VDD(VDD),.Y(g8892),.A(g8681),.B(g4969));
  AND2 AND2_882(.VSS(VSS),.VDD(VDD),.Y(g8901),.A(g8804),.B(g5631));
  AND2 AND2_883(.VSS(VSS),.VDD(VDD),.Y(g8911),.A(g8798),.B(g7688));
  AND2 AND2_884(.VSS(VSS),.VDD(VDD),.Y(g8912),.A(g8796),.B(g8239));
  AND2 AND2_885(.VSS(VSS),.VDD(VDD),.Y(g8914),.A(g8795),.B(g8239));
  AND2 AND2_886(.VSS(VSS),.VDD(VDD),.Y(g8915),.A(g8794),.B(g8239));
  AND2 AND2_887(.VSS(VSS),.VDD(VDD),.Y(g8919),.A(g4567),.B(g8743));
  AND2 AND2_888(.VSS(VSS),.VDD(VDD),.Y(g8920),.A(g4578),.B(g8746));
  AND2 AND2_889(.VSS(VSS),.VDD(VDD),.Y(g8921),.A(g4579),.B(g8747));
  AND2 AND2_890(.VSS(VSS),.VDD(VDD),.Y(g8922),.A(g4586),.B(g8750));
  AND2 AND2_891(.VSS(VSS),.VDD(VDD),.Y(g8923),.A(g4587),.B(g8751));
  AND2 AND2_892(.VSS(VSS),.VDD(VDD),.Y(g8924),.A(g4588),.B(g8752));
  AND2 AND2_893(.VSS(VSS),.VDD(VDD),.Y(g8925),.A(g4592),.B(g8754));
  AND2 AND2_894(.VSS(VSS),.VDD(VDD),.Y(g8926),.A(g4593),.B(g8755));
  AND2 AND2_895(.VSS(VSS),.VDD(VDD),.Y(g8927),.A(g4594),.B(g8756));
  AND2 AND2_896(.VSS(VSS),.VDD(VDD),.Y(g8928),.A(g4595),.B(g8757));
  AND2 AND2_897(.VSS(VSS),.VDD(VDD),.Y(g8929),.A(g3865),.B(g8759));
  AND2 AND2_898(.VSS(VSS),.VDD(VDD),.Y(g8930),.A(g3866),.B(g8760));
  AND2 AND2_899(.VSS(VSS),.VDD(VDD),.Y(g8931),.A(g3867),.B(g8761));
  AND2 AND2_900(.VSS(VSS),.VDD(VDD),.Y(g8932),.A(g3868),.B(g8762));
  AND2 AND2_901(.VSS(VSS),.VDD(VDD),.Y(g8933),.A(g4511),.B(g8765));
  AND2 AND2_902(.VSS(VSS),.VDD(VDD),.Y(g8934),.A(g3873),.B(g8766));
  AND2 AND2_903(.VSS(VSS),.VDD(VDD),.Y(g8935),.A(g3874),.B(g8767));
  AND2 AND2_904(.VSS(VSS),.VDD(VDD),.Y(g8936),.A(g3875),.B(g8768));
  AND2 AND2_905(.VSS(VSS),.VDD(VDD),.Y(g8937),.A(g4524),.B(g8770));
  AND2 AND2_906(.VSS(VSS),.VDD(VDD),.Y(g8938),.A(g3878),.B(g8771));
  AND2 AND2_907(.VSS(VSS),.VDD(VDD),.Y(g8939),.A(g3879),.B(g8772));
  AND2 AND2_908(.VSS(VSS),.VDD(VDD),.Y(g8940),.A(g4543),.B(g8775));
  AND2 AND2_909(.VSS(VSS),.VDD(VDD),.Y(g8941),.A(g3882),.B(g8776));
  AND2 AND2_910(.VSS(VSS),.VDD(VDD),.Y(g8942),.A(g4522),.B(g8780));
  AND2 AND2_911(.VSS(VSS),.VDD(VDD),.Y(g8943),.A(g4560),.B(g8781));
  AND2 AND2_912(.VSS(VSS),.VDD(VDD),.Y(g8944),.A(g4539),.B(g8783));
  AND2 AND2_913(.VSS(VSS),.VDD(VDD),.Y(g8945),.A(g4541),.B(g8784));
  AND2 AND2_914(.VSS(VSS),.VDD(VDD),.Y(g8946),.A(g4556),.B(g8786));
  AND2 AND2_915(.VSS(VSS),.VDD(VDD),.Y(g8947),.A(g4558),.B(g8787));
  AND2 AND2_916(.VSS(VSS),.VDD(VDD),.Y(g8948),.A(g4570),.B(g8789));
  AND2 AND2_917(.VSS(VSS),.VDD(VDD),.Y(g8949),.A(g4572),.B(g8790));
  AND2 AND2_918(.VSS(VSS),.VDD(VDD),.Y(g8950),.A(g4582),.B(g8791));
  AND2 AND2_919(.VSS(VSS),.VDD(VDD),.Y(g8951),.A(g8785),.B(g6072));
  AND2 AND2_920(.VSS(VSS),.VDD(VDD),.Y(g8952),.A(g8788),.B(g6075));
  AND2 AND2_921(.VSS(VSS),.VDD(VDD),.Y(g8953),.A(g8758),.B(g6093));
  AND2 AND2_922(.VSS(VSS),.VDD(VDD),.Y(g8954),.A(g8763),.B(g6097));
  AND2 AND2_923(.VSS(VSS),.VDD(VDD),.Y(g8961),.A(g8885),.B(g5317));
  AND2 AND2_924(.VSS(VSS),.VDD(VDD),.Y(g8962),.A(g8890),.B(g5317));
  AND2 AND2_925(.VSS(VSS),.VDD(VDD),.Y(g8963),.A(g8891),.B(g5317));
  AND2 AND2_926(.VSS(VSS),.VDD(VDD),.Y(g8976),.A(g8903),.B(g6588));
  AND2 AND2_927(.VSS(VSS),.VDD(VDD),.Y(g8978),.A(g8909),.B(g5587));
  AND2 AND2_928(.VSS(VSS),.VDD(VDD),.Y(g9012),.A(g8908),.B(g8239));
  AND2 AND2_929(.VSS(VSS),.VDD(VDD),.Y(g9013),.A(g8907),.B(g8239));
  AND2 AND2_930(.VSS(VSS),.VDD(VDD),.Y(g9014),.A(g8906),.B(g8239));
  AND2 AND2_931(.VSS(VSS),.VDD(VDD),.Y(g9015),.A(g8905),.B(g8239));
  AND2 AND2_932(.VSS(VSS),.VDD(VDD),.Y(g9016),.A(g8904),.B(g8239));
  AND2 AND2_933(.VSS(VSS),.VDD(VDD),.Y(g9021),.A(g8886),.B(g5317));
  AND2 AND2_934(.VSS(VSS),.VDD(VDD),.Y(g9022),.A(g8887),.B(g5317));
  AND2 AND2_935(.VSS(VSS),.VDD(VDD),.Y(g9023),.A(g8888),.B(g5317));
  AND2 AND2_936(.VSS(VSS),.VDD(VDD),.Y(g9024),.A(g8884),.B(g5317));
  AND2 AND2_937(.VSS(VSS),.VDD(VDD),.Y(g9025),.A(g8889),.B(g5317));
  AND2 AND2_938(.VSS(VSS),.VDD(VDD),.Y(g9037),.A(g8965),.B(g5345));
  AND2 AND2_939(.VSS(VSS),.VDD(VDD),.Y(g9038),.A(g8966),.B(g5345));
  AND2 AND2_940(.VSS(VSS),.VDD(VDD),.Y(g9080),.A(g9011),.B(g5598));
  AND2 AND2_941(.VSS(VSS),.VDD(VDD),.Y(g9084),.A(g8964),.B(g5345));
  AND2 AND2_942(.VSS(VSS),.VDD(VDD),.Y(g9118),.A(g9046),.B(g5345));
  AND2 AND2_943(.VSS(VSS),.VDD(VDD),.Y(g9119),.A(g9049),.B(g5345));
  AND2 AND2_944(.VSS(VSS),.VDD(VDD),.Y(g9120),.A(g9052),.B(g5345));
  AND2 AND2_945(.VSS(VSS),.VDD(VDD),.Y(g9130),.A(g9054),.B(g5345));
  AND2 AND2_946(.VSS(VSS),.VDD(VDD),.Y(g9131),.A(g9055),.B(g5345));
  AND2 AND2_947(.VSS(VSS),.VDD(VDD),.Y(g9142),.A(g9124),.B(g6059));
  AND2 AND2_948(.VSS(VSS),.VDD(VDD),.Y(g9143),.A(g9122),.B(g6089));
  AND2 AND2_949(.VSS(VSS),.VDD(VDD),.Y(g9144),.A(g9123),.B(g6096));
  AND2 AND2_950(.VSS(VSS),.VDD(VDD),.Y(g9146),.A(g9135),.B(g6101));
  AND2 AND2_951(.VSS(VSS),.VDD(VDD),.Y(g9147),.A(g9136),.B(g6103));
  AND2 AND2_952(.VSS(VSS),.VDD(VDD),.Y(g9158),.A(g9137),.B(g6070));
  AND2 AND2_953(.VSS(VSS),.VDD(VDD),.Y(g9159),.A(g9138),.B(g6074));
  AND2 AND2_954(.VSS(VSS),.VDD(VDD),.Y(g9160),.A(g9139),.B(g6092));
  AND2 AND2_955(.VSS(VSS),.VDD(VDD),.Y(g9226),.A(g9220),.B(g5403));
  AND2 AND2_956(.VSS(VSS),.VDD(VDD),.Y(g9238),.A(g4748),.B(g9223));
  AND2 AND2_957(.VSS(VSS),.VDD(VDD),.Y(g9240),.A(g9223),.B(g5261));
  AND2 AND2_958(.VSS(VSS),.VDD(VDD),.Y(g9247),.A(g4748),.B(g9227));
  AND2 AND2_959(.VSS(VSS),.VDD(VDD),.Y(g9251),.A(g4748),.B(g9230));
  AND2 AND2_960(.VSS(VSS),.VDD(VDD),.Y(g9258),.A(g9227),.B(g5628));
  AND2 AND2_961(.VSS(VSS),.VDD(VDD),.Y(g9259),.A(g9230),.B(g5639));
  AND2 AND2_962(.VSS(VSS),.VDD(VDD),.Y(g9270),.A(g4748),.B(g9241));
  AND2 AND2_963(.VSS(VSS),.VDD(VDD),.Y(g9271),.A(g4748),.B(g9244));
  AND2 AND2_964(.VSS(VSS),.VDD(VDD),.Y(g9272),.A(g4748),.B(g9248));
  AND2 AND2_965(.VSS(VSS),.VDD(VDD),.Y(g9273),.A(g4748),.B(g9252));
  AND2 AND2_966(.VSS(VSS),.VDD(VDD),.Y(g9274),.A(g4748),.B(g9255));
  AND2 AND2_967(.VSS(VSS),.VDD(VDD),.Y(g9275),.A(g9241),.B(g5645));
  AND2 AND2_968(.VSS(VSS),.VDD(VDD),.Y(g9276),.A(g9244),.B(g5649));
  AND2 AND2_969(.VSS(VSS),.VDD(VDD),.Y(g9277),.A(g9248),.B(g5654));
  AND2 AND2_970(.VSS(VSS),.VDD(VDD),.Y(g9278),.A(g9252),.B(g5658));
  AND2 AND2_971(.VSS(VSS),.VDD(VDD),.Y(g9279),.A(g9255),.B(g5665));
  AND2 AND2_972(.VSS(VSS),.VDD(VDD),.Y(g9327),.A(g9316),.B(g5757));
  AND2 AND2_973(.VSS(VSS),.VDD(VDD),.Y(g9328),.A(g9324),.B(g6465));
  AND2 AND2_974(.VSS(VSS),.VDD(VDD),.Y(g9334),.A(g9318),.B(g6205));
  AND2 AND2_975(.VSS(VSS),.VDD(VDD),.Y(g9335),.A(g9320),.B(g6206));
  AND2 AND2_976(.VSS(VSS),.VDD(VDD),.Y(g9343),.A(g9328),.B(g1738));
  AND2 AND2_977(.VSS(VSS),.VDD(VDD),.Y(g9344),.A(g9329),.B(g6211));
  AND2 AND2_978(.VSS(VSS),.VDD(VDD),.Y(g9345),.A(g9330),.B(g6217));
  AND2 AND2_979(.VSS(VSS),.VDD(VDD),.Y(g9346),.A(g9331),.B(g6222));
  AND2 AND2_980(.VSS(VSS),.VDD(VDD),.Y(g9347),.A(g9332),.B(g6226));
  AND2 AND2_981(.VSS(VSS),.VDD(VDD),.Y(g9348),.A(g9333),.B(g6229));
  AND2 AND2_982(.VSS(VSS),.VDD(VDD),.Y(g9349),.A(g9340),.B(g5690));
  AND2 AND2_983(.VSS(VSS),.VDD(VDD),.Y(g9359),.A(g4748),.B(g9340));
  AND2 AND2_984(.VSS(VSS),.VDD(VDD),.Y(g9371),.A(g9352),.B(g5917));
  AND2 AND2_985(.VSS(VSS),.VDD(VDD),.Y(g9384),.A(g9383),.B(g6245));
//
  OR3 OR3_0(.VSS(VSS),.VDD(VDD),.Y(g1690),.A(g1021),.B(g1025),.C(g1018));
  OR4 OR4_0(.VSS(VSS),.VDD(VDD),.Y(I5757),.A(g969),.B(g970),.C(g966),.D(g963));
  OR4 OR4_1(.VSS(VSS),.VDD(VDD),.Y(g1872),.A(g971),.B(g962),.C(g972),.D(I5757));
  OR2 OR2_0(.VSS(VSS),.VDD(VDD),.Y(g1955),.A(g1189),.B(g16));
  OR2 OR2_1(.VSS(VSS),.VDD(VDD),.Y(g2043),.A(g1263),.B(g1257));
  OR4 OR4_2(.VSS(VSS),.VDD(VDD),.Y(g2206),.A(g1363),.B(g1364),.C(g1365),.D(g1366));
  OR4 OR4_3(.VSS(VSS),.VDD(VDD),.Y(g2213),.A(g1367),.B(g1368),.C(g1369),.D(g1370));
  OR4 OR4_4(.VSS(VSS),.VDD(VDD),.Y(g2214),.A(g1376),.B(g1377),.C(g1378),.D(g1379));
  OR4 OR4_5(.VSS(VSS),.VDD(VDD),.Y(g2229),.A(g1371),.B(g1372),.C(g1373),.D(g1374));
  OR4 OR4_6(.VSS(VSS),.VDD(VDD),.Y(g2230),.A(g1380),.B(g1381),.C(g1382),.D(g1383));
  OR4 OR4_7(.VSS(VSS),.VDD(VDD),.Y(g2262),.A(g1384),.B(g1385),.C(g1386),.D(g1387));
  OR4 OR4_8(.VSS(VSS),.VDD(VDD),.Y(I6208),.A(g891),.B(g896),.C(g901),.D(g906));
  OR4 OR4_9(.VSS(VSS),.VDD(VDD),.Y(I6209),.A(g911),.B(g916),.C(g921),.D(g883));
  OR2 OR2_2(.VSS(VSS),.VDD(VDD),.Y(g2368),.A(I6208),.B(I6209));
  OR2 OR2_3(.VSS(VSS),.VDD(VDD),.Y(g2845),.A(g1877),.B(g576));
  OR2 OR2_4(.VSS(VSS),.VDD(VDD),.Y(g3097),.A(g1746),.B(g287));
  OR2 OR2_5(.VSS(VSS),.VDD(VDD),.Y(g3131),.A(g1749),.B(g368));
  OR2 OR2_6(.VSS(VSS),.VDD(VDD),.Y(g3160),.A(g1751),.B(g449));
  OR2 OR2_7(.VSS(VSS),.VDD(VDD),.Y(g3192),.A(g1756),.B(g530));
  OR2 OR2_8(.VSS(VSS),.VDD(VDD),.Y(g3339),.A(g1424),.B(g2014));
  OR2 OR2_9(.VSS(VSS),.VDD(VDD),.Y(g3541),.A(g1663),.B(g1421));
  OR4 OR4_10(.VSS(VSS),.VDD(VDD),.Y(I7232),.A(g2367),.B(g2352),.C(g2378),.D(g2330));
  OR4 OR4_11(.VSS(VSS),.VDD(VDD),.Y(I7233),.A(g2315),.B(g2385),.C(g2294),.D(g2395));
  OR2 OR2_10(.VSS(VSS),.VDD(VDD),.Y(g3760),.A(I7232),.B(I7233));
  OR2 OR2_11(.VSS(VSS),.VDD(VDD),.Y(g3986),.A(g202),.B(g3129));
  OR2 OR2_12(.VSS(VSS),.VDD(VDD),.Y(g4055),.A(g187),.B(g3012));
  OR2 OR2_13(.VSS(VSS),.VDD(VDD),.Y(g4072),.A(g196),.B(g2995));
  OR2 OR2_14(.VSS(VSS),.VDD(VDD),.Y(g4179),.A(g207),.B(g3083));
  OR2 OR2_15(.VSS(VSS),.VDD(VDD),.Y(g4249),.A(g3617),.B(g1639));
  OR2 OR2_16(.VSS(VSS),.VDD(VDD),.Y(g4264),.A(g2490),.B(g3315));
  OR4 OR4_12(.VSS(VSS),.VDD(VDD),.Y(I8224),.A(g3019),.B(g3029),.C(g3038),.D(g3052));
  OR4 OR4_13(.VSS(VSS),.VDD(VDD),.Y(I8225),.A(g3062),.B(g2712),.C(g2734),.D(g2752));
  OR2 OR2_17(.VSS(VSS),.VDD(VDD),.Y(g4280),.A(I8224),.B(I8225));
  OR2 OR2_18(.VSS(VSS),.VDD(VDD),.Y(g4283),.A(g3587),.B(g2665));
  OR2 OR2_19(.VSS(VSS),.VDD(VDD),.Y(g4295),.A(g2828),.B(g2668));
  OR2 OR2_20(.VSS(VSS),.VDD(VDD),.Y(g4297),.A(g3617),.B(g3602));
  OR2 OR2_21(.VSS(VSS),.VDD(VDD),.Y(g4364),.A(g2952),.B(g1725));
  OR3 OR3_1(.VSS(VSS),.VDD(VDD),.Y(I8363),.A(g2655),.B(g1163),.C(g1160));
  OR4 OR4_14(.VSS(VSS),.VDD(VDD),.Y(g4374),.A(g1182),.B(g1186),.C(g1179),.D(I8363));
  OR2 OR2_22(.VSS(VSS),.VDD(VDD),.Y(g4413),.A(g2371),.B(g3285));
  OR2 OR2_23(.VSS(VSS),.VDD(VDD),.Y(g4688),.A(g4193),.B(g3190));
  OR3 OR3_2(.VSS(VSS),.VDD(VDD),.Y(I9029),.A(g4504),.B(g4494),.C(g4430));
  OR4 OR4_15(.VSS(VSS),.VDD(VDD),.Y(g4727),.A(g4417),.B(g4172),.C(g4163),.D(I9029));
  OR3 OR3_3(.VSS(VSS),.VDD(VDD),.Y(I9038),.A(g4507),.B(g4497),.C(g4486));
  OR3 OR3_4(.VSS(VSS),.VDD(VDD),.Y(g4734),.A(g4469),.B(g4448),.C(I9038));
  OR3 OR3_5(.VSS(VSS),.VDD(VDD),.Y(I9041),.A(g4483),.B(g4466),.C(g4445));
  OR4 OR4_16(.VSS(VSS),.VDD(VDD),.Y(g4735),.A(g4427),.B(g4414),.C(g4403),.D(I9041));
  OR3 OR3_6(.VSS(VSS),.VDD(VDD),.Y(I9044),.A(g4150),.B(g4142),.C(g4549));
  OR3 OR3_7(.VSS(VSS),.VDD(VDD),.Y(g4736),.A(g4532),.B(g4517),.C(I9044));
  OR3 OR3_8(.VSS(VSS),.VDD(VDD),.Y(I9047),.A(g4155),.B(g4147),.C(g4139));
  OR4 OR4_17(.VSS(VSS),.VDD(VDD),.Y(g4737),.A(g4135),.B(g4529),.C(g4514),.D(I9047));
  OR2 OR2_24(.VSS(VSS),.VDD(VDD),.Y(g4747),.A(g3984),.B(g2912));
  OR3 OR3_9(.VSS(VSS),.VDD(VDD),.Y(I9099),.A(g4127),.B(g4123),.C(g4117));
  OR4 OR4_18(.VSS(VSS),.VDD(VDD),.Y(g4786),.A(g4107),.B(g4097),.C(g4124),.D(I9099));
  OR4 OR4_19(.VSS(VSS),.VDD(VDD),.Y(I9107),.A(g4133),.B(g4145),.C(g4138),.D(g4132));
  OR4 OR4_20(.VSS(VSS),.VDD(VDD),.Y(g4790),.A(g4185),.B(g4131),.C(g4129),.D(I9107));
  OR2 OR2_25(.VSS(VSS),.VDD(VDD),.Y(g4812),.A(g2490),.B(g4237));
  OR2 OR2_26(.VSS(VSS),.VDD(VDD),.Y(g4829),.A(g863),.B(g4051));
  OR2 OR2_27(.VSS(VSS),.VDD(VDD),.Y(g4870),.A(g4154),.B(g3081));
  OR2 OR2_28(.VSS(VSS),.VDD(VDD),.Y(g4876),.A(g4159),.B(g4167));
  OR2 OR2_29(.VSS(VSS),.VDD(VDD),.Y(g4927),.A(g4318),.B(g1590));
  OR2 OR2_30(.VSS(VSS),.VDD(VDD),.Y(g5021),.A(g943),.B(g4501));
  OR2 OR2_31(.VSS(VSS),.VDD(VDD),.Y(g5036),.A(g4047),.B(g2972));
  OR4 OR4_21(.VSS(VSS),.VDD(VDD),.Y(g5040),.A(g3900),.B(g3895),.C(g3890),.D(g4363));
  OR2 OR2_32(.VSS(VSS),.VDD(VDD),.Y(g5052),.A(g4049),.B(g4054));
  OR4 OR4_22(.VSS(VSS),.VDD(VDD),.Y(g5057),.A(g3939),.B(g3925),.C(g3915),.D(g3907));
  OR2 OR2_33(.VSS(VSS),.VDD(VDD),.Y(g5070),.A(g4052),.B(g4058));
  OR2 OR2_34(.VSS(VSS),.VDD(VDD),.Y(g5138),.A(g4108),.B(g3049));
  OR2 OR2_35(.VSS(VSS),.VDD(VDD),.Y(g5140),.A(g4333),.B(g3509));
  OR2 OR2_36(.VSS(VSS),.VDD(VDD),.Y(g5188),.A(g5008),.B(g4365));
  OR2 OR2_37(.VSS(VSS),.VDD(VDD),.Y(g5193),.A(g5017),.B(g4366));
  OR2 OR2_38(.VSS(VSS),.VDD(VDD),.Y(g5194),.A(g5018),.B(g4367));
  OR2 OR2_39(.VSS(VSS),.VDD(VDD),.Y(g5195),.A(g5019),.B(g4368));
  OR2 OR2_40(.VSS(VSS),.VDD(VDD),.Y(g5196),.A(g5020),.B(g4369));
  OR2 OR2_41(.VSS(VSS),.VDD(VDD),.Y(g5200),.A(g5029),.B(g4375));
  OR2 OR2_42(.VSS(VSS),.VDD(VDD),.Y(g5201),.A(g5030),.B(g4376));
  OR2 OR2_43(.VSS(VSS),.VDD(VDD),.Y(g5202),.A(g5031),.B(g4377));
  OR2 OR2_44(.VSS(VSS),.VDD(VDD),.Y(g5203),.A(g5032),.B(g4378));
  OR2 OR2_45(.VSS(VSS),.VDD(VDD),.Y(g5204),.A(g5033),.B(g4379));
  OR2 OR2_46(.VSS(VSS),.VDD(VDD),.Y(g5205),.A(g5034),.B(g4380));
  OR2 OR2_47(.VSS(VSS),.VDD(VDD),.Y(g5208),.A(g5043),.B(g4383));
  OR2 OR2_48(.VSS(VSS),.VDD(VDD),.Y(g5209),.A(g5044),.B(g4384));
  OR2 OR2_49(.VSS(VSS),.VDD(VDD),.Y(g5210),.A(g5045),.B(g4385));
  OR2 OR2_50(.VSS(VSS),.VDD(VDD),.Y(g5211),.A(g5046),.B(g4386));
  OR2 OR2_51(.VSS(VSS),.VDD(VDD),.Y(g5212),.A(g5047),.B(g4387));
  OR2 OR2_52(.VSS(VSS),.VDD(VDD),.Y(g5213),.A(g5048),.B(g4388));
  OR2 OR2_53(.VSS(VSS),.VDD(VDD),.Y(g5214),.A(g5049),.B(g4389));
  OR2 OR2_54(.VSS(VSS),.VDD(VDD),.Y(g5215),.A(g5050),.B(g4390));
  OR2 OR2_55(.VSS(VSS),.VDD(VDD),.Y(g5216),.A(g5062),.B(g4391));
  OR2 OR2_56(.VSS(VSS),.VDD(VDD),.Y(g5217),.A(g5063),.B(g4392));
  OR2 OR2_57(.VSS(VSS),.VDD(VDD),.Y(g5218),.A(g5064),.B(g4393));
  OR2 OR2_58(.VSS(VSS),.VDD(VDD),.Y(g5219),.A(g5065),.B(g4394));
  OR2 OR2_59(.VSS(VSS),.VDD(VDD),.Y(g5220),.A(g5066),.B(g4395));
  OR2 OR2_60(.VSS(VSS),.VDD(VDD),.Y(g5221),.A(g5067),.B(g4396));
  OR2 OR2_61(.VSS(VSS),.VDD(VDD),.Y(g5222),.A(g5068),.B(g4397));
  OR2 OR2_62(.VSS(VSS),.VDD(VDD),.Y(g5223),.A(g5069),.B(g4398));
  OR2 OR2_63(.VSS(VSS),.VDD(VDD),.Y(g5227),.A(g5077),.B(g4407));
  OR2 OR2_64(.VSS(VSS),.VDD(VDD),.Y(g5228),.A(g5078),.B(g4408));
  OR2 OR2_65(.VSS(VSS),.VDD(VDD),.Y(g5229),.A(g5079),.B(g4409));
  OR2 OR2_66(.VSS(VSS),.VDD(VDD),.Y(g5230),.A(g5080),.B(g4410));
  OR2 OR2_67(.VSS(VSS),.VDD(VDD),.Y(g5231),.A(g5081),.B(g4411));
  OR2 OR2_68(.VSS(VSS),.VDD(VDD),.Y(g5232),.A(g5082),.B(g4412));
  OR2 OR2_69(.VSS(VSS),.VDD(VDD),.Y(g5233),.A(g5089),.B(g4420));
  OR2 OR2_70(.VSS(VSS),.VDD(VDD),.Y(g5234),.A(g5090),.B(g4421));
  OR2 OR2_71(.VSS(VSS),.VDD(VDD),.Y(g5235),.A(g5091),.B(g4422));
  OR2 OR2_72(.VSS(VSS),.VDD(VDD),.Y(g5236),.A(g5092),.B(g4423));
  OR2 OR2_73(.VSS(VSS),.VDD(VDD),.Y(g5237),.A(g5093),.B(g4424));
  OR2 OR2_74(.VSS(VSS),.VDD(VDD),.Y(g5238),.A(g5094),.B(g4425));
  OR2 OR2_75(.VSS(VSS),.VDD(VDD),.Y(g5241),.A(g5104),.B(g4433));
  OR2 OR2_76(.VSS(VSS),.VDD(VDD),.Y(g5242),.A(g5105),.B(g4434));
  OR2 OR2_77(.VSS(VSS),.VDD(VDD),.Y(g5243),.A(g5106),.B(g4435));
  OR2 OR2_78(.VSS(VSS),.VDD(VDD),.Y(g5244),.A(g5107),.B(g4436));
  OR2 OR2_79(.VSS(VSS),.VDD(VDD),.Y(g5245),.A(g5108),.B(g4437));
  OR2 OR2_80(.VSS(VSS),.VDD(VDD),.Y(g5253),.A(g5116),.B(g4451));
  OR2 OR2_81(.VSS(VSS),.VDD(VDD),.Y(g5254),.A(g5117),.B(g4452));
  OR2 OR2_82(.VSS(VSS),.VDD(VDD),.Y(g5255),.A(g5118),.B(g4453));
  OR2 OR2_83(.VSS(VSS),.VDD(VDD),.Y(g5256),.A(g5119),.B(g4454));
  OR2 OR2_84(.VSS(VSS),.VDD(VDD),.Y(g5259),.A(g5122),.B(g4472));
  OR2 OR2_85(.VSS(VSS),.VDD(VDD),.Y(g5260),.A(g5123),.B(g4473));
  OR2 OR2_86(.VSS(VSS),.VDD(VDD),.Y(g5264),.A(g5125),.B(g4490));
  OR2 OR2_87(.VSS(VSS),.VDD(VDD),.Y(g5265),.A(g5126),.B(g4491));
  OR3 OR3_10(.VSS(VSS),.VDD(VDD),.Y(g5317),.A(g4727),.B(g4737),.C(g4735));
  OR2 OR2_88(.VSS(VSS),.VDD(VDD),.Y(g5343),.A(g4690),.B(g2862));
  OR2 OR2_89(.VSS(VSS),.VDD(VDD),.Y(g5345),.A(g4736),.B(g4734));
  OR2 OR2_90(.VSS(VSS),.VDD(VDD),.Y(g5440),.A(g4790),.B(g4786));
  OR2 OR2_91(.VSS(VSS),.VDD(VDD),.Y(g5483),.A(g4740),.B(g4098));
  OR2 OR2_92(.VSS(VSS),.VDD(VDD),.Y(g5511),.A(g4743),.B(g4109));
  OR2 OR2_93(.VSS(VSS),.VDD(VDD),.Y(g5518),.A(g4744),.B(g4118));
  OR2 OR2_94(.VSS(VSS),.VDD(VDD),.Y(g5537),.A(g3617),.B(g4835));
  OR2 OR2_95(.VSS(VSS),.VDD(VDD),.Y(g5545),.A(g3617),.B(g4824));
  OR2 OR2_96(.VSS(VSS),.VDD(VDD),.Y(g5549),.A(g2935),.B(g4712));
  OR2 OR2_97(.VSS(VSS),.VDD(VDD),.Y(g5561),.A(g4168),.B(g4797));
  OR2 OR2_98(.VSS(VSS),.VDD(VDD),.Y(g5566),.A(g3617),.B(g4810));
  OR2 OR2_99(.VSS(VSS),.VDD(VDD),.Y(g5572),.A(g5051),.B(g1236));
  OR2 OR2_100(.VSS(VSS),.VDD(VDD),.Y(g5673),.A(g4823),.B(g4872));
  OR2 OR2_101(.VSS(VSS),.VDD(VDD),.Y(g5698),.A(g5057),.B(g5040));
  OR2 OR2_102(.VSS(VSS),.VDD(VDD),.Y(g5704),.A(g4936),.B(g4334));
  OR2 OR2_103(.VSS(VSS),.VDD(VDD),.Y(g5706),.A(g4955),.B(g4342));
  OR2 OR2_104(.VSS(VSS),.VDD(VDD),.Y(g5707),.A(g4956),.B(g4343));
  OR2 OR2_105(.VSS(VSS),.VDD(VDD),.Y(g5708),.A(g2889),.B(g4699));
  OR2 OR2_106(.VSS(VSS),.VDD(VDD),.Y(g5710),.A(g4958),.B(g4351));
  OR2 OR2_107(.VSS(VSS),.VDD(VDD),.Y(g5711),.A(g4959),.B(g4352));
  OR2 OR2_108(.VSS(VSS),.VDD(VDD),.Y(g5715),.A(g4961),.B(g4355));
  OR2 OR2_109(.VSS(VSS),.VDD(VDD),.Y(g5716),.A(g4962),.B(g4356));
  OR2 OR2_110(.VSS(VSS),.VDD(VDD),.Y(g5722),.A(g5001),.B(g4361));
  OR2 OR2_111(.VSS(VSS),.VDD(VDD),.Y(g5830),.A(g5714),.B(g5142));
  OR2 OR2_112(.VSS(VSS),.VDD(VDD),.Y(g6115),.A(g3617),.B(g5558));
  OR2 OR2_113(.VSS(VSS),.VDD(VDD),.Y(g6116),.A(g5546),.B(g4681));
  OR2 OR2_114(.VSS(VSS),.VDD(VDD),.Y(g6120),.A(g3617),.B(g5555));
  OR2 OR2_115(.VSS(VSS),.VDD(VDD),.Y(g6121),.A(g5425),.B(g4785));
  OR2 OR2_116(.VSS(VSS),.VDD(VDD),.Y(g6123),.A(g3617),.B(g5556));
  OR2 OR2_117(.VSS(VSS),.VDD(VDD),.Y(g6124),.A(g5432),.B(g4789));
  OR2 OR2_118(.VSS(VSS),.VDD(VDD),.Y(g6132),.A(g5436),.B(g4793));
  OR2 OR2_119(.VSS(VSS),.VDD(VDD),.Y(g6138),.A(g5438),.B(g5442));
  OR2 OR2_120(.VSS(VSS),.VDD(VDD),.Y(g6144),.A(g4175),.B(g5458));
  OR2 OR2_121(.VSS(VSS),.VDD(VDD),.Y(g6249),.A(g4066),.B(g5313));
  OR2 OR2_122(.VSS(VSS),.VDD(VDD),.Y(g6262),.A(g4074),.B(g5334));
  OR3 OR3_11(.VSS(VSS),.VDD(VDD),.Y(g6270),.A(g1000),.B(g5335),.C(g1909));
  OR2 OR2_123(.VSS(VSS),.VDD(VDD),.Y(g6436),.A(g6266),.B(g5699));
  OR2 OR2_124(.VSS(VSS),.VDD(VDD),.Y(g6440),.A(g6268),.B(g5700));
  OR2 OR2_125(.VSS(VSS),.VDD(VDD),.Y(g6445),.A(g6105),.B(g6107));
  OR3 OR3_12(.VSS(VSS),.VDD(VDD),.Y(g6457),.A(g6196),.B(g6209),.C(g4937));
  OR4 OR4_23(.VSS(VSS),.VDD(VDD),.Y(g6458),.A(g6184),.B(g6259),.C(g6174),.D(g6214));
  OR3 OR3_13(.VSS(VSS),.VDD(VDD),.Y(I11603),.A(g6193),.B(g6197),.C(g6175));
  OR3 OR3_14(.VSS(VSS),.VDD(VDD),.Y(g6459),.A(g6259),.B(g6185),.C(I11603));
  OR2 OR2_126(.VSS(VSS),.VDD(VDD),.Y(g6470),.A(g5817),.B(g2934));
  OR2 OR2_127(.VSS(VSS),.VDD(VDD),.Y(g6525),.A(g6112),.B(g5547));
  OR2 OR2_128(.VSS(VSS),.VDD(VDD),.Y(g6543),.A(g6125),.B(g1553));
  OR3 OR3_15(.VSS(VSS),.VDD(VDD),.Y(g6565),.A(g2396),.B(g6131),.C(g1603));
  OR2 OR2_129(.VSS(VSS),.VDD(VDD),.Y(g6579),.A(g6098),.B(g1975));
  OR2 OR2_130(.VSS(VSS),.VDD(VDD),.Y(g6580),.A(g6039),.B(g6041));
  OR2 OR2_131(.VSS(VSS),.VDD(VDD),.Y(g6585),.A(g3617),.B(g6119));
  OR2 OR2_132(.VSS(VSS),.VDD(VDD),.Y(g6590),.A(g3617),.B(g6153));
  OR2 OR2_133(.VSS(VSS),.VDD(VDD),.Y(g6600),.A(g5443),.B(g6055));
  OR2 OR2_134(.VSS(VSS),.VDD(VDD),.Y(g6602),.A(g6058),.B(g3092));
  OR2 OR2_135(.VSS(VSS),.VDD(VDD),.Y(g6610),.A(g4180),.B(g6061));
  OR2 OR2_136(.VSS(VSS),.VDD(VDD),.Y(g6673),.A(g4053),.B(g5937));
  OR2 OR2_137(.VSS(VSS),.VDD(VDD),.Y(g6685),.A(g4067),.B(g5969));
  OR2 OR2_138(.VSS(VSS),.VDD(VDD),.Y(g6686),.A(g4068),.B(g5970));
  OR2 OR2_139(.VSS(VSS),.VDD(VDD),.Y(g6688),.A(g6145),.B(g5570));
  OR2 OR2_140(.VSS(VSS),.VDD(VDD),.Y(g6694),.A(g6151),.B(g5573));
  OR2 OR2_141(.VSS(VSS),.VDD(VDD),.Y(g6698),.A(g4073),.B(g6001));
  OR2 OR2_142(.VSS(VSS),.VDD(VDD),.Y(g6699),.A(g6154),.B(g5579));
  OR2 OR2_143(.VSS(VSS),.VDD(VDD),.Y(g6705),.A(g6157),.B(g5583));
  OR2 OR2_144(.VSS(VSS),.VDD(VDD),.Y(g6706),.A(g4077),.B(g6002));
  OR2 OR2_145(.VSS(VSS),.VDD(VDD),.Y(g6707),.A(g6160),.B(g5585));
  OR2 OR2_146(.VSS(VSS),.VDD(VDD),.Y(g6710),.A(g55),.B(g6264));
  OR2 OR2_147(.VSS(VSS),.VDD(VDD),.Y(g6716),.A(g6162),.B(g5588));
  OR2 OR2_148(.VSS(VSS),.VDD(VDD),.Y(g6717),.A(g4082),.B(g6005));
  OR2 OR2_149(.VSS(VSS),.VDD(VDD),.Y(g6718),.A(g4083),.B(g6006));
  OR2 OR2_150(.VSS(VSS),.VDD(VDD),.Y(g6719),.A(g6166),.B(g6171));
  OR2 OR2_151(.VSS(VSS),.VDD(VDD),.Y(g6728),.A(g6168),.B(g5593));
  OR2 OR2_152(.VSS(VSS),.VDD(VDD),.Y(g6734),.A(g6176),.B(g5599));
  OR2 OR2_153(.VSS(VSS),.VDD(VDD),.Y(g6735),.A(g4091),.B(g6013));
  OR2 OR2_154(.VSS(VSS),.VDD(VDD),.Y(g6739),.A(g4099),.B(g6021));
  OR2 OR2_155(.VSS(VSS),.VDD(VDD),.Y(g6740),.A(g4100),.B(g6022));
  OR2 OR2_156(.VSS(VSS),.VDD(VDD),.Y(g6906),.A(g6715),.B(g6726));
  OR2 OR2_157(.VSS(VSS),.VDD(VDD),.Y(g6907),.A(g6727),.B(g6732));
  OR2 OR2_158(.VSS(VSS),.VDD(VDD),.Y(g6912),.A(g4199),.B(g6567));
  OR2 OR2_159(.VSS(VSS),.VDD(VDD),.Y(g6913),.A(g6733),.B(g6738));
  OR2 OR2_160(.VSS(VSS),.VDD(VDD),.Y(g6917),.A(g6743),.B(g6753));
  OR2 OR2_161(.VSS(VSS),.VDD(VDD),.Y(g6919),.A(g6771),.B(g6394));
  OR2 OR2_162(.VSS(VSS),.VDD(VDD),.Y(g6920),.A(g6395),.B(g6399));
  OR2 OR2_163(.VSS(VSS),.VDD(VDD),.Y(g6921),.A(g6396),.B(g6401));
  OR2 OR2_164(.VSS(VSS),.VDD(VDD),.Y(g6924),.A(g6400),.B(g6405));
  OR2 OR2_165(.VSS(VSS),.VDD(VDD),.Y(g6925),.A(g6402),.B(g6407));
  OR2 OR2_166(.VSS(VSS),.VDD(VDD),.Y(g6926),.A(g6406),.B(g6411));
  OR2 OR2_167(.VSS(VSS),.VDD(VDD),.Y(g6927),.A(g6408),.B(g6413));
  OR2 OR2_168(.VSS(VSS),.VDD(VDD),.Y(g6928),.A(g6409),.B(g6415));
  OR2 OR2_169(.VSS(VSS),.VDD(VDD),.Y(g6929),.A(g6412),.B(g6418));
  OR2 OR2_170(.VSS(VSS),.VDD(VDD),.Y(g6930),.A(g6414),.B(g6420));
  OR2 OR2_171(.VSS(VSS),.VDD(VDD),.Y(g6931),.A(g6416),.B(g6421));
  OR2 OR2_172(.VSS(VSS),.VDD(VDD),.Y(g6932),.A(g6417),.B(g6423));
  OR2 OR2_173(.VSS(VSS),.VDD(VDD),.Y(g6933),.A(g6419),.B(g6428));
  OR2 OR2_174(.VSS(VSS),.VDD(VDD),.Y(g6934),.A(g6422),.B(g6430));
  OR2 OR2_175(.VSS(VSS),.VDD(VDD),.Y(g6935),.A(g6429),.B(g6431));
  OR2 OR2_176(.VSS(VSS),.VDD(VDD),.Y(g6952),.A(g6633),.B(g6204));
  OR2 OR2_177(.VSS(VSS),.VDD(VDD),.Y(g6964),.A(g6447),.B(g6448));
  OR2 OR2_178(.VSS(VSS),.VDD(VDD),.Y(g6980),.A(g6745),.B(g6028));
  OR2 OR2_179(.VSS(VSS),.VDD(VDD),.Y(g7016),.A(g6042),.B(g6487));
  OR2 OR2_180(.VSS(VSS),.VDD(VDD),.Y(g7020),.A(g3617),.B(g6578));
  OR2 OR2_181(.VSS(VSS),.VDD(VDD),.Y(g7025),.A(g6541),.B(g3095));
  OR2 OR2_182(.VSS(VSS),.VDD(VDD),.Y(g7026),.A(g4186),.B(g6554));
  OR2 OR2_183(.VSS(VSS),.VDD(VDD),.Y(g7029),.A(g6433),.B(g5765));
  OR2 OR2_184(.VSS(VSS),.VDD(VDD),.Y(g7040),.A(g6439),.B(g5783));
  OR2 OR2_185(.VSS(VSS),.VDD(VDD),.Y(g7062),.A(g4048),.B(g6456));
  OR2 OR2_186(.VSS(VSS),.VDD(VDD),.Y(g7080),.A(g4086),.B(g6462));
  OR2 OR2_187(.VSS(VSS),.VDD(VDD),.Y(g7081),.A(g6172),.B(g6629));
  OR3 OR3_16(.VSS(VSS),.VDD(VDD),.Y(g7083),.A(g5448),.B(g6267),.C(g6710));
  OR2 OR2_188(.VSS(VSS),.VDD(VDD),.Y(g7086),.A(g4101),.B(g6464));
  OR2 OR2_189(.VSS(VSS),.VDD(VDD),.Y(g7088),.A(g6638),.B(g6641));
  OR2 OR2_190(.VSS(VSS),.VDD(VDD),.Y(g7089),.A(g4128),.B(g6474));
  OR2 OR2_191(.VSS(VSS),.VDD(VDD),.Y(g7165),.A(g6434),.B(g6908));
  OR2 OR2_192(.VSS(VSS),.VDD(VDD),.Y(g7166),.A(g6437),.B(g6914));
  OR2 OR2_193(.VSS(VSS),.VDD(VDD),.Y(g7167),.A(g6438),.B(g6915));
  OR2 OR2_194(.VSS(VSS),.VDD(VDD),.Y(g7170),.A(g6916),.B(g6444));
  OR2 OR2_195(.VSS(VSS),.VDD(VDD),.Y(g7191),.A(g7071),.B(g6980));
  OR2 OR2_196(.VSS(VSS),.VDD(VDD),.Y(g7202),.A(g6028),.B(g7071));
  OR2 OR2_197(.VSS(VSS),.VDD(VDD),.Y(g7220),.A(g1304),.B(g7062));
  OR2 OR2_198(.VSS(VSS),.VDD(VDD),.Y(g7222),.A(g6049),.B(g6971));
  OR2 OR2_199(.VSS(VSS),.VDD(VDD),.Y(g7227),.A(g6992),.B(g3128));
  OR2 OR2_200(.VSS(VSS),.VDD(VDD),.Y(g7230),.A(g4190),.B(g6995));
  OR2 OR2_201(.VSS(VSS),.VDD(VDD),.Y(g7248),.A(g7079),.B(g5652));
  OR2 OR2_202(.VSS(VSS),.VDD(VDD),.Y(g7254),.A(g6923),.B(g5298));
  OR3 OR3_17(.VSS(VSS),.VDD(VDD),.Y(I13220),.A(g58),.B(g6258),.C(g5418));
  OR3 OR3_18(.VSS(VSS),.VDD(VDD),.Y(g7258),.A(g7083),.B(g5403),.C(I13220));
  OR2 OR2_203(.VSS(VSS),.VDD(VDD),.Y(g7272),.A(g6182),.B(g7038));
  OR2 OR2_204(.VSS(VSS),.VDD(VDD),.Y(g7337),.A(g7278),.B(g4546));
  OR2 OR2_205(.VSS(VSS),.VDD(VDD),.Y(g7363),.A(g7136),.B(g6903));
  OR2 OR2_206(.VSS(VSS),.VDD(VDD),.Y(g7421),.A(g6745),.B(g7202));
  OR3 OR3_19(.VSS(VSS),.VDD(VDD),.Y(I13553),.A(g1166),.B(g1167),.C(g1170));
  OR3 OR3_20(.VSS(VSS),.VDD(VDD),.Y(g7426),.A(g1173),.B(g7217),.C(I13553));
  OR2 OR2_207(.VSS(VSS),.VDD(VDD),.Y(g7428),.A(g6040),.B(g7175));
  OR2 OR2_208(.VSS(VSS),.VDD(VDD),.Y(g7435),.A(g6052),.B(g7182));
  OR2 OR2_209(.VSS(VSS),.VDD(VDD),.Y(g7436),.A(g7183),.B(g6975));
  OR2 OR2_210(.VSS(VSS),.VDD(VDD),.Y(g7438),.A(g7184),.B(g6978));
  OR2 OR2_211(.VSS(VSS),.VDD(VDD),.Y(g7443),.A(g7192),.B(g3158));
  OR2 OR2_212(.VSS(VSS),.VDD(VDD),.Y(g7445),.A(g4192),.B(g7193));
  OR2 OR2_213(.VSS(VSS),.VDD(VDD),.Y(g7450),.A(g6090),.B(g7195));
  OR2 OR2_214(.VSS(VSS),.VDD(VDD),.Y(g7575),.A(g7323),.B(g7142));
  OR2 OR2_215(.VSS(VSS),.VDD(VDD),.Y(g7682),.A(g6044),.B(g7412));
  OR2 OR2_216(.VSS(VSS),.VDD(VDD),.Y(g7687),.A(g6053),.B(g7416));
  OR2 OR2_217(.VSS(VSS),.VDD(VDD),.Y(g7690),.A(g4181),.B(g7417));
  OR2 OR2_218(.VSS(VSS),.VDD(VDD),.Y(g7697),.A(g7419),.B(g3187));
  OR2 OR2_219(.VSS(VSS),.VDD(VDD),.Y(g7782),.A(g4783),.B(g7598));
  OR2 OR2_220(.VSS(VSS),.VDD(VDD),.Y(g7783),.A(g4787),.B(g7600));
  OR3 OR3_21(.VSS(VSS),.VDD(VDD),.Y(I14219),.A(g979),.B(g7566),.C(g1865));
  OR4 OR4_24(.VSS(VSS),.VDD(VDD),.Y(g7784),.A(g7406),.B(g6664),.C(g3492),.D(I14219));
  OR2 OR2_221(.VSS(VSS),.VDD(VDD),.Y(g7787),.A(g4791),.B(g7602));
  OR2 OR2_222(.VSS(VSS),.VDD(VDD),.Y(g7788),.A(g4794),.B(g7604));
  OR2 OR2_223(.VSS(VSS),.VDD(VDD),.Y(g7791),.A(g4796),.B(g7606));
  OR2 OR2_224(.VSS(VSS),.VDD(VDD),.Y(g7810),.A(g4799),.B(g7609));
  OR2 OR2_225(.VSS(VSS),.VDD(VDD),.Y(g7825),.A(g4801),.B(g7615));
  OR2 OR2_226(.VSS(VSS),.VDD(VDD),.Y(g7826),.A(g4804),.B(g7626));
  OR2 OR2_227(.VSS(VSS),.VDD(VDD),.Y(g7834),.A(g7724),.B(g6762));
  OR3 OR3_22(.VSS(VSS),.VDD(VDD),.Y(I14302),.A(g6664),.B(g3492),.C(g979));
  OR4 OR4_25(.VSS(VSS),.VDD(VDD),.Y(g8009),.A(g3591),.B(g7406),.C(g7566),.D(I14302));
  OR3 OR3_23(.VSS(VSS),.VDD(VDD),.Y(g8082),.A(g7654),.B(g7628),.C(g7611));
  OR3 OR3_24(.VSS(VSS),.VDD(VDD),.Y(I14366),.A(g7566),.B(g1030),.C(g6664));
  OR3 OR3_25(.VSS(VSS),.VDD(VDD),.Y(g8091),.A(g7215),.B(g6452),.C(I14366));
  OR3 OR3_26(.VSS(VSS),.VDD(VDD),.Y(g8128),.A(g7566),.B(g6910),.C(g6452));
  OR2 OR2_228(.VSS(VSS),.VDD(VDD),.Y(g8146),.A(g6045),.B(g7597));
  OR2 OR2_229(.VSS(VSS),.VDD(VDD),.Y(g8154),.A(g6054),.B(g7607));
  OR2 OR2_230(.VSS(VSS),.VDD(VDD),.Y(g8155),.A(g7632),.B(g3219));
  OR4 OR4_26(.VSS(VSS),.VDD(VDD),.Y(g8176),.A(g7566),.B(g1030),.C(g6664),.D(g6452));
  OR4 OR4_27(.VSS(VSS),.VDD(VDD),.Y(I14467),.A(g7993),.B(g7966),.C(g7793),.D(g7811));
  OR4 OR4_28(.VSS(VSS),.VDD(VDD),.Y(I14468),.A(g7937),.B(g7887),.C(g8029),.D(g8018));
  OR4 OR4_29(.VSS(VSS),.VDD(VDD),.Y(I14479),.A(g7993),.B(g7966),.C(g7793),.D(g7811));
  OR4 OR4_30(.VSS(VSS),.VDD(VDD),.Y(I14480),.A(g7937),.B(g7887),.C(g8029),.D(g8018));
  OR4 OR4_31(.VSS(VSS),.VDD(VDD),.Y(I14484),.A(g7993),.B(g7966),.C(g7793),.D(g7811));
  OR4 OR4_32(.VSS(VSS),.VDD(VDD),.Y(I14485),.A(g7937),.B(g7887),.C(g8029),.D(g8018));
  OR4 OR4_33(.VSS(VSS),.VDD(VDD),.Y(I14495),.A(g7993),.B(g7966),.C(g7793),.D(g7811));
  OR4 OR4_34(.VSS(VSS),.VDD(VDD),.Y(I14496),.A(g7937),.B(g7887),.C(g8029),.D(g8018));
  OR2 OR2_231(.VSS(VSS),.VDD(VDD),.Y(g8613),.A(g8082),.B(g7616));
  OR2 OR2_232(.VSS(VSS),.VDD(VDD),.Y(g8634),.A(g6047),.B(g8060));
  OR2 OR2_233(.VSS(VSS),.VDD(VDD),.Y(g8637),.A(g6057),.B(g8071));
  OR4 OR4_35(.VSS(VSS),.VDD(VDD),.Y(I14753),.A(g7993),.B(g7966),.C(g7793),.D(g7811));
  OR4 OR4_36(.VSS(VSS),.VDD(VDD),.Y(I14754),.A(g7937),.B(g7887),.C(g8029),.D(g8018));
  OR4 OR4_37(.VSS(VSS),.VDD(VDD),.Y(I14758),.A(g7993),.B(g7966),.C(g7793),.D(g7811));
  OR4 OR4_38(.VSS(VSS),.VDD(VDD),.Y(I14759),.A(g7937),.B(g7887),.C(g8029),.D(g8018));
  OR4 OR4_39(.VSS(VSS),.VDD(VDD),.Y(I14766),.A(g7993),.B(g7966),.C(g7793),.D(g7811));
  OR4 OR4_40(.VSS(VSS),.VDD(VDD),.Y(I14767),.A(g7937),.B(g7887),.C(g8029),.D(g8018));
  OR4 OR4_41(.VSS(VSS),.VDD(VDD),.Y(I14771),.A(g7993),.B(g7966),.C(g7793),.D(g7811));
  OR4 OR4_42(.VSS(VSS),.VDD(VDD),.Y(I14772),.A(g7937),.B(g7887),.C(g8029),.D(g8018));
  OR3 OR3_27(.VSS(VSS),.VDD(VDD),.Y(I14831),.A(g8483),.B(g8464),.C(g8514));
  OR3 OR3_28(.VSS(VSS),.VDD(VDD),.Y(I14834),.A(g8483),.B(g8464),.C(g8514));
  OR4 OR4_43(.VSS(VSS),.VDD(VDD),.Y(I14932),.A(g8278),.B(g8329),.C(g8461),.D(g8382));
  OR4 OR4_44(.VSS(VSS),.VDD(VDD),.Y(I14933),.A(g8385),.B(g8404),.C(g8441),.D(g8462));
  OR3 OR3_29(.VSS(VSS),.VDD(VDD),.Y(g8758),.A(g8655),.B(I14932),.C(I14933));
  OR4 OR4_45(.VSS(VSS),.VDD(VDD),.Y(I14941),.A(g8275),.B(g8323),.C(g8459),.D(g8380));
  OR4 OR4_46(.VSS(VSS),.VDD(VDD),.Y(I14942),.A(g8439),.B(g8440),.C(g8405),.D(g8460));
  OR3 OR3_30(.VSS(VSS),.VDD(VDD),.Y(g8763),.A(g8232),.B(I14941),.C(I14942));
  OR4 OR4_47(.VSS(VSS),.VDD(VDD),.Y(I14951),.A(g8328),.B(g8316),.C(g8455),.D(g8378));
  OR4 OR4_48(.VSS(VSS),.VDD(VDD),.Y(I14952),.A(g8456),.B(g8513),.C(g8458),.D(g8236));
  OR2 OR2_234(.VSS(VSS),.VDD(VDD),.Y(g8769),.A(I14951),.B(I14952));
  OR4 OR4_49(.VSS(VSS),.VDD(VDD),.Y(I14959),.A(g8322),.B(g8308),.C(g8438),.D(g8612));
  OR4 OR4_50(.VSS(VSS),.VDD(VDD),.Y(I14960),.A(g8621),.B(g8622),.C(g8628),.D(g8230));
  OR2 OR2_235(.VSS(VSS),.VDD(VDD),.Y(g8773),.A(I14959),.B(I14960));
  OR4 OR4_51(.VSS(VSS),.VDD(VDD),.Y(I14969),.A(g8315),.B(g8377),.C(g8359),.D(g8611));
  OR4 OR4_52(.VSS(VSS),.VDD(VDD),.Y(I14970),.A(g8457),.B(g8383),.C(g8626),.D(g8233));
  OR2 OR2_236(.VSS(VSS),.VDD(VDD),.Y(g8777),.A(I14969),.B(I14970));
  OR3 OR3_31(.VSS(VSS),.VDD(VDD),.Y(I14980),.A(g8362),.B(g8403),.C(g8610));
  OR3 OR3_32(.VSS(VSS),.VDD(VDD),.Y(g8782),.A(g8624),.B(g8659),.C(I14980));
  OR3 OR3_33(.VSS(VSS),.VDD(VDD),.Y(I14985),.A(g8341),.B(g8384),.C(g8542));
  OR3 OR3_34(.VSS(VSS),.VDD(VDD),.Y(g8785),.A(g8623),.B(g8656),.C(I14985));
  OR3 OR3_35(.VSS(VSS),.VDD(VDD),.Y(I14990),.A(g8337),.B(g8379),.C(g8543));
  OR3 OR3_36(.VSS(VSS),.VDD(VDD),.Y(g8788),.A(g8620),.B(g8658),.C(I14990));
  OR4 OR4_53(.VSS(VSS),.VDD(VDD),.Y(g8794),.A(g8153),.B(g8074),.C(g8069),.D(g8523));
  OR4 OR4_54(.VSS(VSS),.VDD(VDD),.Y(g8795),.A(g8151),.B(g8077),.C(g8075),.D(g8279));
  OR4 OR4_55(.VSS(VSS),.VDD(VDD),.Y(g8796),.A(g8150),.B(g8078),.C(g8070),.D(g8360));
  OR4 OR4_56(.VSS(VSS),.VDD(VDD),.Y(I15017),.A(g8131),.B(g8111),.C(g8042),.D(g8156));
  OR4 OR4_57(.VSS(VSS),.VDD(VDD),.Y(I15018),.A(g7855),.B(g7838),.C(g7905),.D(g7870));
  OR4 OR4_58(.VSS(VSS),.VDD(VDD),.Y(I15019),.A(g7951),.B(g7920),.C(g7983),.D(g8181));
  OR4 OR4_59(.VSS(VSS),.VDD(VDD),.Y(I15020),.A(g8363),.B(g8342),.C(g8407),.D(g8386));
  OR4 OR4_60(.VSS(VSS),.VDD(VDD),.Y(I15021),.A(I15017),.B(I15018),.C(I15019),.D(I15020));
  OR2 OR2_237(.VSS(VSS),.VDD(VDD),.Y(g8804),.A(g6060),.B(g8609));
  OR4 OR4_61(.VSS(VSS),.VDD(VDD),.Y(I15029),.A(g8131),.B(g8111),.C(g8042),.D(g8156));
  OR4 OR4_62(.VSS(VSS),.VDD(VDD),.Y(I15030),.A(g7855),.B(g7838),.C(g7905),.D(g7870));
  OR4 OR4_63(.VSS(VSS),.VDD(VDD),.Y(I15031),.A(g7951),.B(g7920),.C(g7983),.D(g8181));
  OR4 OR4_64(.VSS(VSS),.VDD(VDD),.Y(I15032),.A(g8363),.B(g8342),.C(g8407),.D(g8386));
  OR4 OR4_65(.VSS(VSS),.VDD(VDD),.Y(I15033),.A(I15029),.B(I15030),.C(I15031),.D(I15032));
  OR4 OR4_66(.VSS(VSS),.VDD(VDD),.Y(I15040),.A(g8131),.B(g8111),.C(g8042),.D(g8156));
  OR4 OR4_67(.VSS(VSS),.VDD(VDD),.Y(I15041),.A(g7855),.B(g7838),.C(g7905),.D(g7870));
  OR4 OR4_68(.VSS(VSS),.VDD(VDD),.Y(I15042),.A(g7951),.B(g7920),.C(g7983),.D(g8181));
  OR4 OR4_69(.VSS(VSS),.VDD(VDD),.Y(I15043),.A(g8363),.B(g8342),.C(g8407),.D(g8386));
  OR4 OR4_70(.VSS(VSS),.VDD(VDD),.Y(I15044),.A(I15040),.B(I15041),.C(I15042),.D(I15043));
  OR4 OR4_71(.VSS(VSS),.VDD(VDD),.Y(I15051),.A(g8131),.B(g8111),.C(g8042),.D(g8156));
  OR4 OR4_72(.VSS(VSS),.VDD(VDD),.Y(I15052),.A(g7855),.B(g7838),.C(g7905),.D(g7870));
  OR4 OR4_73(.VSS(VSS),.VDD(VDD),.Y(I15053),.A(g7951),.B(g7920),.C(g7983),.D(g8181));
  OR4 OR4_74(.VSS(VSS),.VDD(VDD),.Y(I15054),.A(g8363),.B(g8342),.C(g8407),.D(g8386));
  OR4 OR4_75(.VSS(VSS),.VDD(VDD),.Y(I15055),.A(I15051),.B(I15052),.C(I15053),.D(I15054));
  OR4 OR4_76(.VSS(VSS),.VDD(VDD),.Y(I15071),.A(g8131),.B(g8111),.C(g8042),.D(g8156));
  OR4 OR4_77(.VSS(VSS),.VDD(VDD),.Y(I15072),.A(g7855),.B(g7838),.C(g7905),.D(g7870));
  OR4 OR4_78(.VSS(VSS),.VDD(VDD),.Y(I15073),.A(g7951),.B(g7920),.C(g7983),.D(g8181));
  OR4 OR4_79(.VSS(VSS),.VDD(VDD),.Y(I15074),.A(g8363),.B(g8342),.C(g8407),.D(g8386));
  OR4 OR4_80(.VSS(VSS),.VDD(VDD),.Y(I15075),.A(I15071),.B(I15072),.C(I15073),.D(I15074));
  OR4 OR4_81(.VSS(VSS),.VDD(VDD),.Y(I15082),.A(g8131),.B(g8111),.C(g8042),.D(g8156));
  OR4 OR4_82(.VSS(VSS),.VDD(VDD),.Y(I15083),.A(g7855),.B(g7838),.C(g7905),.D(g7870));
  OR4 OR4_83(.VSS(VSS),.VDD(VDD),.Y(I15084),.A(g7951),.B(g7920),.C(g7983),.D(g8181));
  OR4 OR4_84(.VSS(VSS),.VDD(VDD),.Y(I15085),.A(g8363),.B(g8342),.C(g8407),.D(g8386));
  OR4 OR4_85(.VSS(VSS),.VDD(VDD),.Y(I15086),.A(I15082),.B(I15083),.C(I15084),.D(I15085));
  OR4 OR4_86(.VSS(VSS),.VDD(VDD),.Y(I15098),.A(g8131),.B(g8111),.C(g8042),.D(g8156));
  OR4 OR4_87(.VSS(VSS),.VDD(VDD),.Y(I15099),.A(g7855),.B(g7838),.C(g7905),.D(g7870));
  OR4 OR4_88(.VSS(VSS),.VDD(VDD),.Y(I15100),.A(g7951),.B(g7920),.C(g7983),.D(g8181));
  OR4 OR4_89(.VSS(VSS),.VDD(VDD),.Y(I15101),.A(g8363),.B(g8342),.C(g8407),.D(g8386));
  OR4 OR4_90(.VSS(VSS),.VDD(VDD),.Y(I15102),.A(I15098),.B(I15099),.C(I15100),.D(I15101));
  OR4 OR4_91(.VSS(VSS),.VDD(VDD),.Y(I15109),.A(g8131),.B(g8111),.C(g8042),.D(g8156));
  OR4 OR4_92(.VSS(VSS),.VDD(VDD),.Y(I15110),.A(g7855),.B(g7838),.C(g7905),.D(g7870));
  OR4 OR4_93(.VSS(VSS),.VDD(VDD),.Y(I15111),.A(g7951),.B(g7920),.C(g7983),.D(g8181));
  OR4 OR4_94(.VSS(VSS),.VDD(VDD),.Y(I15112),.A(g8363),.B(g8342),.C(g8407),.D(g8386));
  OR4 OR4_95(.VSS(VSS),.VDD(VDD),.Y(I15113),.A(I15109),.B(I15110),.C(I15111),.D(I15112));
  OR2 OR2_238(.VSS(VSS),.VDD(VDD),.Y(g8834),.A(g7096),.B(g8229));
  OR3 OR3_37(.VSS(VSS),.VDD(VDD),.Y(I15147),.A(g8483),.B(g8464),.C(g8514));
  OR3 OR3_38(.VSS(VSS),.VDD(VDD),.Y(I15152),.A(g8483),.B(g8464),.C(g8514));
  OR3 OR3_39(.VSS(VSS),.VDD(VDD),.Y(I15165),.A(g8483),.B(g8464),.C(g8514));
  OR3 OR3_40(.VSS(VSS),.VDD(VDD),.Y(I15169),.A(g8483),.B(g8464),.C(g8514));
  OR3 OR3_41(.VSS(VSS),.VDD(VDD),.Y(I15172),.A(g8483),.B(g8464),.C(g8514));
  OR3 OR3_42(.VSS(VSS),.VDD(VDD),.Y(I15175),.A(g8483),.B(g8464),.C(g8514));
  OR4 OR4_96(.VSS(VSS),.VDD(VDD),.Y(I15228),.A(g8270),.B(g8258),.C(g8281),.D(g8273));
  OR4 OR4_97(.VSS(VSS),.VDD(VDD),.Y(I15229),.A(g8262),.B(g8303),.C(g8268),.D(g8312));
  OR4 OR4_98(.VSS(VSS),.VDD(VDD),.Y(I15230),.A(g8274),.B(g8321),.C(g8298),.D(g8696));
  OR4 OR4_99(.VSS(VSS),.VDD(VDD),.Y(I15231),.A(g8701),.B(g8715),.C(g8730),.D(g8720));
  OR4 OR4_100(.VSS(VSS),.VDD(VDD),.Y(I15232),.A(I15228),.B(I15229),.C(I15230),.D(I15231));
  OR3 OR3_43(.VSS(VSS),.VDD(VDD),.Y(g8884),.A(g8735),.B(g8818),.C(I15232));
  OR4 OR4_101(.VSS(VSS),.VDD(VDD),.Y(I15239),.A(g8264),.B(g8260),.C(g8277),.D(g8301));
  OR4 OR4_102(.VSS(VSS),.VDD(VDD),.Y(I15240),.A(g8259),.B(g8294),.C(g8263),.D(g8305));
  OR4 OR4_103(.VSS(VSS),.VDD(VDD),.Y(I15241),.A(g8269),.B(g8314),.C(g8309),.D(g8695));
  OR4 OR4_104(.VSS(VSS),.VDD(VDD),.Y(I15242),.A(g8697),.B(g8714),.C(g8718),.D(g8719));
  OR4 OR4_105(.VSS(VSS),.VDD(VDD),.Y(I15243),.A(I15239),.B(I15240),.C(I15241),.D(I15242));
  OR3 OR3_44(.VSS(VSS),.VDD(VDD),.Y(g8885),.A(g8723),.B(g8806),.C(I15243));
  OR4 OR4_106(.VSS(VSS),.VDD(VDD),.Y(I15250),.A(g8238),.B(g8265),.C(g8272),.D(g8292));
  OR4 OR4_107(.VSS(VSS),.VDD(VDD),.Y(I15251),.A(g8302),.B(g8288),.C(g8311),.D(g8296));
  OR4 OR4_108(.VSS(VSS),.VDD(VDD),.Y(I15252),.A(g8320),.B(g8307),.C(g8317),.D(g8692));
  OR4 OR4_109(.VSS(VSS),.VDD(VDD),.Y(I15253),.A(g8698),.B(g8711),.C(g8722),.D(g8716));
  OR4 OR4_110(.VSS(VSS),.VDD(VDD),.Y(I15254),.A(I15250),.B(I15251),.C(I15252),.D(I15253));
  OR3 OR3_45(.VSS(VSS),.VDD(VDD),.Y(g8886),.A(g8727),.B(g8812),.C(I15254));
  OR4 OR4_111(.VSS(VSS),.VDD(VDD),.Y(I15261),.A(g8256),.B(g8271),.C(g8267),.D(g8286));
  OR4 OR4_112(.VSS(VSS),.VDD(VDD),.Y(I15262),.A(g8293),.B(g8283),.C(g8304),.D(g8289));
  OR4 OR4_113(.VSS(VSS),.VDD(VDD),.Y(I15263),.A(g8313),.B(g8297),.C(g8310),.D(g8690));
  OR4 OR4_114(.VSS(VSS),.VDD(VDD),.Y(I15264),.A(g8700),.B(g8708),.C(g8726),.D(g8731));
  OR4 OR4_115(.VSS(VSS),.VDD(VDD),.Y(I15265),.A(I15261),.B(I15262),.C(I15263),.D(I15264));
  OR2 OR2_239(.VSS(VSS),.VDD(VDD),.Y(g8887),.A(I15265),.B(g8819));
  OR4 OR4_116(.VSS(VSS),.VDD(VDD),.Y(I15272),.A(g8237),.B(g8300),.C(g8261),.D(g8282));
  OR4 OR4_117(.VSS(VSS),.VDD(VDD),.Y(I15273),.A(g8287),.B(g8334),.C(g8295),.D(g8339));
  OR4 OR4_118(.VSS(VSS),.VDD(VDD),.Y(I15274),.A(g8306),.B(g8361),.C(g8299),.D(g8687));
  OR4 OR4_119(.VSS(VSS),.VDD(VDD),.Y(I15275),.A(g8693),.B(g8703),.C(g8712),.D(g8717));
  OR4 OR4_120(.VSS(VSS),.VDD(VDD),.Y(I15276),.A(I15272),.B(I15273),.C(I15274),.D(I15275));
  OR2 OR2_240(.VSS(VSS),.VDD(VDD),.Y(g8888),.A(I15276),.B(g8807));
  OR4 OR4_121(.VSS(VSS),.VDD(VDD),.Y(I15283),.A(g8291),.B(g8276),.C(g8325),.D(g8330));
  OR4 OR4_122(.VSS(VSS),.VDD(VDD),.Y(I15284),.A(g8335),.B(g8340),.C(g8290),.D(g8691));
  OR3 OR3_46(.VSS(VSS),.VDD(VDD),.Y(I15285),.A(g8709),.B(g8713),.C(g8803));
  OR3 OR3_47(.VSS(VSS),.VDD(VDD),.Y(g8889),.A(I15283),.B(I15284),.C(I15285));
  OR4 OR4_123(.VSS(VSS),.VDD(VDD),.Y(I15290),.A(g8285),.B(g8266),.C(g8318),.D(g8326));
  OR4 OR4_124(.VSS(VSS),.VDD(VDD),.Y(I15291),.A(g8331),.B(g8336),.C(g8338),.D(g8688));
  OR3 OR3_48(.VSS(VSS),.VDD(VDD),.Y(I15292),.A(g8704),.B(g8710),.C(g8805));
  OR3 OR3_49(.VSS(VSS),.VDD(VDD),.Y(g8890),.A(I15290),.B(I15291),.C(I15292));
  OR4 OR4_125(.VSS(VSS),.VDD(VDD),.Y(I15297),.A(g8280),.B(g8257),.C(g8319),.D(g8327));
  OR4 OR4_126(.VSS(VSS),.VDD(VDD),.Y(I15298),.A(g8332),.B(g8333),.C(g8686),.D(g8702));
  OR4 OR4_127(.VSS(VSS),.VDD(VDD),.Y(g8891),.A(g8705),.B(g8811),.C(I15297),.D(I15298));
  OR2 OR2_241(.VSS(VSS),.VDD(VDD),.Y(g8893),.A(g8814),.B(g8643));
  OR2 OR2_242(.VSS(VSS),.VDD(VDD),.Y(g8894),.A(g8817),.B(g8645));
  OR2 OR2_243(.VSS(VSS),.VDD(VDD),.Y(g8895),.A(g8823),.B(g8646));
  OR2 OR2_244(.VSS(VSS),.VDD(VDD),.Y(g8896),.A(g8828),.B(g8648));
  OR2 OR2_245(.VSS(VSS),.VDD(VDD),.Y(g8897),.A(g8833),.B(g8650));
  OR2 OR2_246(.VSS(VSS),.VDD(VDD),.Y(g8899),.A(g8839),.B(g8652));
  OR2 OR2_247(.VSS(VSS),.VDD(VDD),.Y(g8900),.A(g8840),.B(g8653));
  OR2 OR2_248(.VSS(VSS),.VDD(VDD),.Y(g8902),.A(g8844),.B(g8654));
  OR3 OR3_50(.VSS(VSS),.VDD(VDD),.Y(g8904),.A(g8090),.B(g8080),.C(g8706));
  OR3 OR3_51(.VSS(VSS),.VDD(VDD),.Y(g8905),.A(g8089),.B(g8087),.C(g8694));
  OR3 OR3_52(.VSS(VSS),.VDD(VDD),.Y(g8906),.A(g8088),.B(g8062),.C(g8699));
  OR3 OR3_53(.VSS(VSS),.VDD(VDD),.Y(g8907),.A(g8081),.B(g8064),.C(g8707));
  OR3 OR3_54(.VSS(VSS),.VDD(VDD),.Y(g8908),.A(g8079),.B(g8066),.C(g8855));
  OR2 OR2_249(.VSS(VSS),.VDD(VDD),.Y(g8909),.A(g6043),.B(g8764));
  OR3 OR3_55(.VSS(VSS),.VDD(VDD),.Y(I15400),.A(g8736),.B(g8748),.C(g8740));
  OR3 OR3_56(.VSS(VSS),.VDD(VDD),.Y(g8964),.A(g8915),.B(g8863),.C(I15400));
  OR4 OR4_128(.VSS(VSS),.VDD(VDD),.Y(g8965),.A(g8739),.B(g8742),.C(g8914),.D(g8847));
  OR4 OR4_129(.VSS(VSS),.VDD(VDD),.Y(g8966),.A(g8741),.B(g8745),.C(g8912),.D(g8850));
  OR2 OR2_250(.VSS(VSS),.VDD(VDD),.Y(g8979),.A(g8919),.B(g8813));
  OR2 OR2_251(.VSS(VSS),.VDD(VDD),.Y(g8980),.A(g8920),.B(g8815));
  OR2 OR2_252(.VSS(VSS),.VDD(VDD),.Y(g8981),.A(g8921),.B(g8816));
  OR2 OR2_253(.VSS(VSS),.VDD(VDD),.Y(g8982),.A(g8922),.B(g8820));
  OR2 OR2_254(.VSS(VSS),.VDD(VDD),.Y(g8983),.A(g8923),.B(g8821));
  OR2 OR2_255(.VSS(VSS),.VDD(VDD),.Y(g8984),.A(g8924),.B(g8822));
  OR2 OR2_256(.VSS(VSS),.VDD(VDD),.Y(g8985),.A(g8925),.B(g8824));
  OR2 OR2_257(.VSS(VSS),.VDD(VDD),.Y(g8986),.A(g8926),.B(g8825));
  OR2 OR2_258(.VSS(VSS),.VDD(VDD),.Y(g8987),.A(g8927),.B(g8826));
  OR2 OR2_259(.VSS(VSS),.VDD(VDD),.Y(g8988),.A(g8928),.B(g8827));
  OR2 OR2_260(.VSS(VSS),.VDD(VDD),.Y(g8989),.A(g8929),.B(g8829));
  OR2 OR2_261(.VSS(VSS),.VDD(VDD),.Y(g8990),.A(g8930),.B(g8830));
  OR2 OR2_262(.VSS(VSS),.VDD(VDD),.Y(g8991),.A(g8931),.B(g8831));
  OR2 OR2_263(.VSS(VSS),.VDD(VDD),.Y(g8992),.A(g8932),.B(g8832));
  OR2 OR2_264(.VSS(VSS),.VDD(VDD),.Y(g8993),.A(g8933),.B(g8835));
  OR2 OR2_265(.VSS(VSS),.VDD(VDD),.Y(g8994),.A(g8934),.B(g8836));
  OR2 OR2_266(.VSS(VSS),.VDD(VDD),.Y(g8995),.A(g8935),.B(g8837));
  OR2 OR2_267(.VSS(VSS),.VDD(VDD),.Y(g8996),.A(g8936),.B(g8838));
  OR2 OR2_268(.VSS(VSS),.VDD(VDD),.Y(g8997),.A(g8937),.B(g8841));
  OR2 OR2_269(.VSS(VSS),.VDD(VDD),.Y(g8998),.A(g8938),.B(g8842));
  OR2 OR2_270(.VSS(VSS),.VDD(VDD),.Y(g8999),.A(g8939),.B(g8843));
  OR2 OR2_271(.VSS(VSS),.VDD(VDD),.Y(g9000),.A(g8940),.B(g8845));
  OR2 OR2_272(.VSS(VSS),.VDD(VDD),.Y(g9001),.A(g8941),.B(g8846));
  OR2 OR2_273(.VSS(VSS),.VDD(VDD),.Y(g9002),.A(g8942),.B(g8848));
  OR2 OR2_274(.VSS(VSS),.VDD(VDD),.Y(g9003),.A(g8943),.B(g8849));
  OR2 OR2_275(.VSS(VSS),.VDD(VDD),.Y(g9004),.A(g8944),.B(g8851));
  OR2 OR2_276(.VSS(VSS),.VDD(VDD),.Y(g9005),.A(g8945),.B(g8852));
  OR2 OR2_277(.VSS(VSS),.VDD(VDD),.Y(g9006),.A(g8946),.B(g8853));
  OR2 OR2_278(.VSS(VSS),.VDD(VDD),.Y(g9007),.A(g8947),.B(g8854));
  OR2 OR2_279(.VSS(VSS),.VDD(VDD),.Y(g9008),.A(g8948),.B(g8857));
  OR2 OR2_280(.VSS(VSS),.VDD(VDD),.Y(g9009),.A(g8949),.B(g8858));
  OR2 OR2_281(.VSS(VSS),.VDD(VDD),.Y(g9010),.A(g8950),.B(g8860));
  OR2 OR2_282(.VSS(VSS),.VDD(VDD),.Y(g9011),.A(g6046),.B(g8892));
  OR4 OR4_130(.VSS(VSS),.VDD(VDD),.Y(g9046),.A(g8744),.B(g8749),.C(g9016),.D(g8862));
  OR4 OR4_131(.VSS(VSS),.VDD(VDD),.Y(g9049),.A(g8732),.B(g8737),.C(g9015),.D(g8861));
  OR4 OR4_132(.VSS(VSS),.VDD(VDD),.Y(g9052),.A(g8728),.B(g8733),.C(g9014),.D(g8679));
  OR4 OR4_133(.VSS(VSS),.VDD(VDD),.Y(g9054),.A(g8724),.B(g8729),.C(g9013),.D(g8680));
  OR4 OR4_134(.VSS(VSS),.VDD(VDD),.Y(g9055),.A(g8721),.B(g8725),.C(g9012),.D(g8859));
  OR2 OR2_283(.VSS(VSS),.VDD(VDD),.Y(g9122),.A(g8953),.B(g9084));
  OR2 OR2_284(.VSS(VSS),.VDD(VDD),.Y(g9123),.A(g8954),.B(g9037));
  OR2 OR2_285(.VSS(VSS),.VDD(VDD),.Y(g9124),.A(g8876),.B(g9038));
  OR2 OR2_286(.VSS(VSS),.VDD(VDD),.Y(g9135),.A(g8951),.B(g9130));
  OR2 OR2_287(.VSS(VSS),.VDD(VDD),.Y(g9136),.A(g8952),.B(g9131));
  OR2 OR2_288(.VSS(VSS),.VDD(VDD),.Y(g9137),.A(g8877),.B(g9118));
  OR2 OR2_289(.VSS(VSS),.VDD(VDD),.Y(g9138),.A(g8878),.B(g9119));
  OR2 OR2_290(.VSS(VSS),.VDD(VDD),.Y(g9139),.A(g8879),.B(g9120));
  OR2 OR2_291(.VSS(VSS),.VDD(VDD),.Y(g9148),.A(g9143),.B(g9024));
  OR2 OR2_292(.VSS(VSS),.VDD(VDD),.Y(g9151),.A(g9144),.B(g8961));
  OR2 OR2_293(.VSS(VSS),.VDD(VDD),.Y(g9154),.A(g9142),.B(g9021));
  OR2 OR2_294(.VSS(VSS),.VDD(VDD),.Y(g9162),.A(g9158),.B(g9022));
  OR2 OR2_295(.VSS(VSS),.VDD(VDD),.Y(g9165),.A(g9159),.B(g9023));
  OR2 OR2_296(.VSS(VSS),.VDD(VDD),.Y(g9168),.A(g9160),.B(g9025));
  OR2 OR2_297(.VSS(VSS),.VDD(VDD),.Y(g9171),.A(g9146),.B(g8962));
  OR2 OR2_298(.VSS(VSS),.VDD(VDD),.Y(g9174),.A(g9147),.B(g8963));
  OR2 OR2_299(.VSS(VSS),.VDD(VDD),.Y(g9239),.A(g7653),.B(g9226));
  OR2 OR2_300(.VSS(VSS),.VDD(VDD),.Y(g9261),.A(g9238),.B(g6227));
  OR2 OR2_301(.VSS(VSS),.VDD(VDD),.Y(g9264),.A(g9247),.B(g6242));
  OR2 OR2_302(.VSS(VSS),.VDD(VDD),.Y(g9267),.A(g9251),.B(g6225));
  OR2 OR2_303(.VSS(VSS),.VDD(VDD),.Y(g9282),.A(g9270),.B(g6238));
  OR2 OR2_304(.VSS(VSS),.VDD(VDD),.Y(g9285),.A(g9271),.B(g6221));
  OR2 OR2_305(.VSS(VSS),.VDD(VDD),.Y(g9288),.A(g9272),.B(g6235));
  OR2 OR2_306(.VSS(VSS),.VDD(VDD),.Y(g9291),.A(g9273),.B(g6216));
  OR2 OR2_307(.VSS(VSS),.VDD(VDD),.Y(g9294),.A(g9274),.B(g6230));
  OR2 OR2_308(.VSS(VSS),.VDD(VDD),.Y(g9337),.A(g9240),.B(g9327));
  OR2 OR2_309(.VSS(VSS),.VDD(VDD),.Y(g9338),.A(g9258),.B(g9334));
  OR2 OR2_310(.VSS(VSS),.VDD(VDD),.Y(g9339),.A(g9259),.B(g9335));
  OR2 OR2_311(.VSS(VSS),.VDD(VDD),.Y(g9352),.A(g9343),.B(g4526));
  OR2 OR2_312(.VSS(VSS),.VDD(VDD),.Y(g9354),.A(g9275),.B(g9344));
  OR2 OR2_313(.VSS(VSS),.VDD(VDD),.Y(g9355),.A(g9276),.B(g9345));
  OR2 OR2_314(.VSS(VSS),.VDD(VDD),.Y(g9356),.A(g9277),.B(g9346));
  OR2 OR2_315(.VSS(VSS),.VDD(VDD),.Y(g9357),.A(g9278),.B(g9347));
  OR2 OR2_316(.VSS(VSS),.VDD(VDD),.Y(g9358),.A(g9279),.B(g9348));
  OR2 OR2_317(.VSS(VSS),.VDD(VDD),.Y(g9363),.A(g9359),.B(g6210));
  OR2 OR2_318(.VSS(VSS),.VDD(VDD),.Y(g9377),.A(g9371),.B(g6757));
  OR2 OR2_319(.VSS(VSS),.VDD(VDD),.Y(g9387),.A(g9349),.B(g9384));
//
  NAND2 NAND2_0(.VSS(VSS),.VDD(VDD),.Y(I5505),.A(g1532),.B(g1528));
  NAND2 NAND2_1(.VSS(VSS),.VDD(VDD),.Y(I5506),.A(g1532),.B(I5505));
  NAND2 NAND2_2(.VSS(VSS),.VDD(VDD),.Y(I5507),.A(g1528),.B(I5505));
  NAND2 NAND2_3(.VSS(VSS),.VDD(VDD),.Y(g1678),.A(I5506),.B(I5507));
  NAND2 NAND2_4(.VSS(VSS),.VDD(VDD),.Y(I5519),.A(g1087),.B(g1098));
  NAND2 NAND2_5(.VSS(VSS),.VDD(VDD),.Y(I5520),.A(g1087),.B(I5519));
  NAND2 NAND2_6(.VSS(VSS),.VDD(VDD),.Y(I5521),.A(g1098),.B(I5519));
  NAND2 NAND2_7(.VSS(VSS),.VDD(VDD),.Y(g1682),.A(I5520),.B(I5521));
  NAND2 NAND2_8(.VSS(VSS),.VDD(VDD),.Y(I5598),.A(g1481),.B(g1489));
  NAND2 NAND2_9(.VSS(VSS),.VDD(VDD),.Y(I5599),.A(g1481),.B(I5598));
  NAND2 NAND2_10(.VSS(VSS),.VDD(VDD),.Y(I5600),.A(g1489),.B(I5598));
  NAND2 NAND2_11(.VSS(VSS),.VDD(VDD),.Y(g1759),.A(I5599),.B(I5600));
  NAND2 NAND2_12(.VSS(VSS),.VDD(VDD),.Y(I5619),.A(g1092),.B(g1130));
  NAND2 NAND2_13(.VSS(VSS),.VDD(VDD),.Y(I5620),.A(g1092),.B(I5619));
  NAND2 NAND2_14(.VSS(VSS),.VDD(VDD),.Y(I5621),.A(g1130),.B(I5619));
  NAND2 NAND2_15(.VSS(VSS),.VDD(VDD),.Y(g1775),.A(I5620),.B(I5621));
  NAND2 NAND2_16(.VSS(VSS),.VDD(VDD),.Y(I5695),.A(g1513),.B(g1524));
  NAND2 NAND2_17(.VSS(VSS),.VDD(VDD),.Y(I5696),.A(g1513),.B(I5695));
  NAND2 NAND2_18(.VSS(VSS),.VDD(VDD),.Y(I5697),.A(g1524),.B(I5695));
  NAND2 NAND2_19(.VSS(VSS),.VDD(VDD),.Y(g1819),.A(I5696),.B(I5697));
  NAND2 NAND2_20(.VSS(VSS),.VDD(VDD),.Y(g1910),.A(g1435),.B(g1439));
  NAND2 NAND2_21(.VSS(VSS),.VDD(VDD),.Y(g2051),.A(g1444),.B(g1450));
  NAND2 NAND2_22(.VSS(VSS),.VDD(VDD),.Y(I6064),.A(g852),.B(g883));
  NAND2 NAND2_23(.VSS(VSS),.VDD(VDD),.Y(I6065),.A(g852),.B(I6064));
  NAND2 NAND2_24(.VSS(VSS),.VDD(VDD),.Y(I6066),.A(g883),.B(I6064));
  NAND2 NAND2_25(.VSS(VSS),.VDD(VDD),.Y(g2294),.A(I6065),.B(I6066));
  NAND2 NAND2_26(.VSS(VSS),.VDD(VDD),.Y(I6102),.A(g849),.B(g921));
  NAND2 NAND2_27(.VSS(VSS),.VDD(VDD),.Y(I6103),.A(g849),.B(I6102));
  NAND2 NAND2_28(.VSS(VSS),.VDD(VDD),.Y(I6104),.A(g921),.B(I6102));
  NAND2 NAND2_29(.VSS(VSS),.VDD(VDD),.Y(g2315),.A(I6103),.B(I6104));
  NAND2 NAND2_30(.VSS(VSS),.VDD(VDD),.Y(I6133),.A(g846),.B(g916));
  NAND2 NAND2_31(.VSS(VSS),.VDD(VDD),.Y(I6134),.A(g846),.B(I6133));
  NAND2 NAND2_32(.VSS(VSS),.VDD(VDD),.Y(I6135),.A(g916),.B(I6133));
  NAND2 NAND2_33(.VSS(VSS),.VDD(VDD),.Y(g2330),.A(I6134),.B(I6135));
  NAND2 NAND2_34(.VSS(VSS),.VDD(VDD),.Y(g2333),.A(g985),.B(g990));
  NAND2 NAND2_35(.VSS(VSS),.VDD(VDD),.Y(I6170),.A(g843),.B(g911));
  NAND2 NAND2_36(.VSS(VSS),.VDD(VDD),.Y(I6171),.A(g843),.B(I6170));
  NAND2 NAND2_37(.VSS(VSS),.VDD(VDD),.Y(I6172),.A(g911),.B(I6170));
  NAND2 NAND2_38(.VSS(VSS),.VDD(VDD),.Y(g2352),.A(I6171),.B(I6172));
  NAND2 NAND2_39(.VSS(VSS),.VDD(VDD),.Y(I6201),.A(g831),.B(g891));
  NAND2 NAND2_40(.VSS(VSS),.VDD(VDD),.Y(I6202),.A(g831),.B(I6201));
  NAND2 NAND2_41(.VSS(VSS),.VDD(VDD),.Y(I6203),.A(g891),.B(I6201));
  NAND2 NAND2_42(.VSS(VSS),.VDD(VDD),.Y(g2367),.A(I6202),.B(I6203));
  NAND2 NAND2_43(.VSS(VSS),.VDD(VDD),.Y(I6232),.A(g834),.B(g896));
  NAND2 NAND2_44(.VSS(VSS),.VDD(VDD),.Y(I6233),.A(g834),.B(I6232));
  NAND2 NAND2_45(.VSS(VSS),.VDD(VDD),.Y(I6234),.A(g896),.B(I6232));
  NAND2 NAND2_46(.VSS(VSS),.VDD(VDD),.Y(g2378),.A(I6233),.B(I6234));
  NAND2 NAND2_47(.VSS(VSS),.VDD(VDD),.Y(I6257),.A(g837),.B(g901));
  NAND2 NAND2_48(.VSS(VSS),.VDD(VDD),.Y(I6258),.A(g837),.B(I6257));
  NAND2 NAND2_49(.VSS(VSS),.VDD(VDD),.Y(I6259),.A(g901),.B(I6257));
  NAND2 NAND2_50(.VSS(VSS),.VDD(VDD),.Y(g2385),.A(I6258),.B(I6259));
  NAND2 NAND2_51(.VSS(VSS),.VDD(VDD),.Y(I6273),.A(g840),.B(g906));
  NAND2 NAND2_52(.VSS(VSS),.VDD(VDD),.Y(I6274),.A(g840),.B(I6273));
  NAND2 NAND2_53(.VSS(VSS),.VDD(VDD),.Y(I6275),.A(g906),.B(I6273));
  NAND2 NAND2_54(.VSS(VSS),.VDD(VDD),.Y(g2395),.A(I6274),.B(I6275));
  NAND2 NAND2_55(.VSS(VSS),.VDD(VDD),.Y(g2474),.A(g1405),.B(g1412));
  NAND2 NAND2_56(.VSS(VSS),.VDD(VDD),.Y(I6499),.A(g1913),.B(g1537));
  NAND2 NAND2_57(.VSS(VSS),.VDD(VDD),.Y(I6500),.A(g1913),.B(I6499));
  NAND2 NAND2_58(.VSS(VSS),.VDD(VDD),.Y(I6501),.A(g1537),.B(I6499));
  NAND2 NAND2_59(.VSS(VSS),.VDD(VDD),.Y(g2751),.A(I6500),.B(I6501));
  NAND2 NAND2_60(.VSS(VSS),.VDD(VDD),.Y(I6522),.A(g1919),.B(g1102));
  NAND2 NAND2_61(.VSS(VSS),.VDD(VDD),.Y(I6523),.A(g1919),.B(I6522));
  NAND2 NAND2_62(.VSS(VSS),.VDD(VDD),.Y(I6524),.A(g1102),.B(I6522));
  NAND2 NAND2_63(.VSS(VSS),.VDD(VDD),.Y(g2783),.A(I6523),.B(I6524));
  NAND2 NAND2_64(.VSS(VSS),.VDD(VDD),.Y(I6538),.A(g2555),.B(g2557));
  NAND2 NAND2_65(.VSS(VSS),.VDD(VDD),.Y(I6539),.A(g2555),.B(I6538));
  NAND2 NAND2_66(.VSS(VSS),.VDD(VDD),.Y(I6540),.A(g2557),.B(I6538));
  NAND2 NAND2_67(.VSS(VSS),.VDD(VDD),.Y(g2801),.A(I6539),.B(I6540));
  NAND2 NAND2_68(.VSS(VSS),.VDD(VDD),.Y(I6739),.A(g195),.B(g1970));
  NAND2 NAND2_69(.VSS(VSS),.VDD(VDD),.Y(I6740),.A(g195),.B(I6739));
  NAND2 NAND2_70(.VSS(VSS),.VDD(VDD),.Y(I6741),.A(g1970),.B(I6739));
  NAND2 NAND2_71(.VSS(VSS),.VDD(VDD),.Y(g2995),.A(I6740),.B(I6741));
  NAND2 NAND2_72(.VSS(VSS),.VDD(VDD),.Y(I6750),.A(g1733),.B(g1494));
  NAND2 NAND2_73(.VSS(VSS),.VDD(VDD),.Y(I6751),.A(g1733),.B(I6750));
  NAND2 NAND2_74(.VSS(VSS),.VDD(VDD),.Y(I6752),.A(g1494),.B(I6750));
  NAND2 NAND2_75(.VSS(VSS),.VDD(VDD),.Y(g3011),.A(I6751),.B(I6752));
  NAND2 NAND2_76(.VSS(VSS),.VDD(VDD),.Y(I6757),.A(g186),.B(g1983));
  NAND2 NAND2_77(.VSS(VSS),.VDD(VDD),.Y(I6758),.A(g186),.B(I6757));
  NAND2 NAND2_78(.VSS(VSS),.VDD(VDD),.Y(I6759),.A(g1983),.B(I6757));
  NAND2 NAND2_79(.VSS(VSS),.VDD(VDD),.Y(g3012),.A(I6758),.B(I6759));
  NAND2 NAND2_80(.VSS(VSS),.VDD(VDD),.Y(I6774),.A(g2386),.B(g1134));
  NAND2 NAND2_81(.VSS(VSS),.VDD(VDD),.Y(I6775),.A(g2386),.B(I6774));
  NAND2 NAND2_82(.VSS(VSS),.VDD(VDD),.Y(I6776),.A(g1134),.B(I6774));
  NAND2 NAND2_83(.VSS(VSS),.VDD(VDD),.Y(g3028),.A(I6775),.B(I6776));
  NAND2 NAND2_84(.VSS(VSS),.VDD(VDD),.Y(I6813),.A(g210),.B(g2052));
  NAND2 NAND2_85(.VSS(VSS),.VDD(VDD),.Y(I6814),.A(g210),.B(I6813));
  NAND2 NAND2_86(.VSS(VSS),.VDD(VDD),.Y(I6815),.A(g2052),.B(I6813));
  NAND2 NAND2_87(.VSS(VSS),.VDD(VDD),.Y(g3083),.A(I6814),.B(I6815));
  NAND2 NAND2_88(.VSS(VSS),.VDD(VDD),.Y(I6842),.A(g205),.B(g2016));
  NAND2 NAND2_89(.VSS(VSS),.VDD(VDD),.Y(I6843),.A(g205),.B(I6842));
  NAND2 NAND2_90(.VSS(VSS),.VDD(VDD),.Y(I6844),.A(g2016),.B(I6842));
  NAND2 NAND2_91(.VSS(VSS),.VDD(VDD),.Y(g3129),.A(I6843),.B(I6844));
  NAND2 NAND2_92(.VSS(VSS),.VDD(VDD),.Y(I6876),.A(g1967),.B(g1910));
  NAND2 NAND2_93(.VSS(VSS),.VDD(VDD),.Y(I6877),.A(g1967),.B(I6876));
  NAND2 NAND2_94(.VSS(VSS),.VDD(VDD),.Y(I6878),.A(g1910),.B(I6876));
  NAND2 NAND2_95(.VSS(VSS),.VDD(VDD),.Y(g3221),.A(I6877),.B(I6878));
  NAND2 NAND2_96(.VSS(VSS),.VDD(VDD),.Y(g3231),.A(g1889),.B(g1904));
  NAND2 NAND2_97(.VSS(VSS),.VDD(VDD),.Y(g3232),.A(g2298),.B(g2276));
  NAND2 NAND2_98(.VSS(VSS),.VDD(VDD),.Y(I6904),.A(g2105),.B(g1838));
  NAND2 NAND2_99(.VSS(VSS),.VDD(VDD),.Y(I6905),.A(g2105),.B(I6904));
  NAND2 NAND2_100(.VSS(VSS),.VDD(VDD),.Y(I6906),.A(g1838),.B(I6904));
  NAND2 NAND2_101(.VSS(VSS),.VDD(VDD),.Y(g3286),.A(I6905),.B(I6906));
  NAND2 NAND2_102(.VSS(VSS),.VDD(VDD),.Y(I6916),.A(g2360),.B(g1732));
  NAND2 NAND2_103(.VSS(VSS),.VDD(VDD),.Y(I6917),.A(g2360),.B(I6916));
  NAND2 NAND2_104(.VSS(VSS),.VDD(VDD),.Y(I6918),.A(g1732),.B(I6916));
  NAND2 NAND2_105(.VSS(VSS),.VDD(VDD),.Y(g3314),.A(I6917),.B(I6918));
  NAND2 NAND2_106(.VSS(VSS),.VDD(VDD),.Y(I6923),.A(g1728),.B(g33));
  NAND2 NAND2_107(.VSS(VSS),.VDD(VDD),.Y(I6924),.A(g1728),.B(I6923));
  NAND2 NAND2_108(.VSS(VSS),.VDD(VDD),.Y(I6925),.A(g33),.B(I6923));
  NAND2 NAND2_109(.VSS(VSS),.VDD(VDD),.Y(g3315),.A(I6924),.B(I6925));
  NAND2 NAND2_110(.VSS(VSS),.VDD(VDD),.Y(I6939),.A(g2161),.B(g2051));
  NAND2 NAND2_111(.VSS(VSS),.VDD(VDD),.Y(I6940),.A(g2161),.B(I6939));
  NAND2 NAND2_112(.VSS(VSS),.VDD(VDD),.Y(I6941),.A(g2051),.B(I6939));
  NAND2 NAND2_113(.VSS(VSS),.VDD(VDD),.Y(g3358),.A(I6940),.B(I6941));
  NAND2 NAND2_114(.VSS(VSS),.VDD(VDD),.Y(I6996),.A(g2275),.B(g2242));
  NAND2 NAND2_115(.VSS(VSS),.VDD(VDD),.Y(I6997),.A(g2275),.B(I6996));
  NAND2 NAND2_116(.VSS(VSS),.VDD(VDD),.Y(I6998),.A(g2242),.B(I6996));
  NAND2 NAND2_117(.VSS(VSS),.VDD(VDD),.Y(g3518),.A(I6997),.B(I6998));
  NAND2 NAND2_118(.VSS(VSS),.VDD(VDD),.Y(I7009),.A(g2295),.B(g2333));
  NAND2 NAND2_119(.VSS(VSS),.VDD(VDD),.Y(I7010),.A(g2295),.B(I7009));
  NAND2 NAND2_120(.VSS(VSS),.VDD(VDD),.Y(I7011),.A(g2333),.B(I7009));
  NAND2 NAND2_121(.VSS(VSS),.VDD(VDD),.Y(g3525),.A(I7010),.B(I7011));
  NAND2 NAND2_122(.VSS(VSS),.VDD(VDD),.Y(I7068),.A(g1639),.B(g1643));
  NAND2 NAND2_123(.VSS(VSS),.VDD(VDD),.Y(I7069),.A(g1639),.B(I7068));
  NAND2 NAND2_124(.VSS(VSS),.VDD(VDD),.Y(I7070),.A(g1643),.B(I7068));
  NAND2 NAND2_125(.VSS(VSS),.VDD(VDD),.Y(g3602),.A(I7069),.B(I7070));
  NAND2 NAND2_126(.VSS(VSS),.VDD(VDD),.Y(I7085),.A(g1753),.B(g1918));
  NAND2 NAND2_127(.VSS(VSS),.VDD(VDD),.Y(I7086),.A(g1753),.B(I7085));
  NAND2 NAND2_128(.VSS(VSS),.VDD(VDD),.Y(I7087),.A(g1918),.B(I7085));
  NAND2 NAND2_129(.VSS(VSS),.VDD(VDD),.Y(g3613),.A(I7086),.B(I7087));
  NAND2 NAND2_130(.VSS(VSS),.VDD(VDD),.Y(I7138),.A(g2404),.B(g2397));
  NAND2 NAND2_131(.VSS(VSS),.VDD(VDD),.Y(I7139),.A(g2404),.B(I7138));
  NAND2 NAND2_132(.VSS(VSS),.VDD(VDD),.Y(I7140),.A(g2397),.B(I7138));
  NAND2 NAND2_133(.VSS(VSS),.VDD(VDD),.Y(g3656),.A(I7139),.B(I7140));
  NAND2 NAND2_134(.VSS(VSS),.VDD(VDD),.Y(I7148),.A(g799),.B(g1974));
  NAND2 NAND2_135(.VSS(VSS),.VDD(VDD),.Y(I7149),.A(g799),.B(I7148));
  NAND2 NAND2_136(.VSS(VSS),.VDD(VDD),.Y(I7150),.A(g1974),.B(I7148));
  NAND2 NAND2_137(.VSS(VSS),.VDD(VDD),.Y(g3658),.A(I7149),.B(I7150));
  NAND2 NAND2_138(.VSS(VSS),.VDD(VDD),.Y(I7156),.A(g2331),.B(g929));
  NAND2 NAND2_139(.VSS(VSS),.VDD(VDD),.Y(I7157),.A(g2331),.B(I7156));
  NAND2 NAND2_140(.VSS(VSS),.VDD(VDD),.Y(I7158),.A(g929),.B(I7156));
  NAND2 NAND2_141(.VSS(VSS),.VDD(VDD),.Y(g3665),.A(I7157),.B(I7158));
  NAND2 NAND2_142(.VSS(VSS),.VDD(VDD),.Y(I7172),.A(g1739),.B(g2006));
  NAND2 NAND2_143(.VSS(VSS),.VDD(VDD),.Y(I7173),.A(g1739),.B(I7172));
  NAND2 NAND2_144(.VSS(VSS),.VDD(VDD),.Y(I7174),.A(g2006),.B(I7172));
  NAND2 NAND2_145(.VSS(VSS),.VDD(VDD),.Y(g3678),.A(I7173),.B(I7174));
  NAND2 NAND2_146(.VSS(VSS),.VDD(VDD),.Y(I7179),.A(g2351),.B(g795));
  NAND2 NAND2_147(.VSS(VSS),.VDD(VDD),.Y(I7180),.A(g2351),.B(I7179));
  NAND2 NAND2_148(.VSS(VSS),.VDD(VDD),.Y(I7181),.A(g795),.B(I7179));
  NAND2 NAND2_149(.VSS(VSS),.VDD(VDD),.Y(g3679),.A(I7180),.B(I7181));
  NAND2 NAND2_150(.VSS(VSS),.VDD(VDD),.Y(I7186),.A(g2353),.B(g1834));
  NAND2 NAND2_151(.VSS(VSS),.VDD(VDD),.Y(I7187),.A(g2353),.B(I7186));
  NAND2 NAND2_152(.VSS(VSS),.VDD(VDD),.Y(I7188),.A(g1834),.B(I7186));
  NAND2 NAND2_153(.VSS(VSS),.VDD(VDD),.Y(g3680),.A(I7187),.B(I7188));
  NAND2 NAND2_154(.VSS(VSS),.VDD(VDD),.Y(g3681),.A(g866),.B(g2368));
  NAND2 NAND2_155(.VSS(VSS),.VDD(VDD),.Y(g3706),.A(g1556),.B(g2510));
  NAND2 NAND2_156(.VSS(VSS),.VDD(VDD),.Y(I7214),.A(g815),.B(g2091));
  NAND2 NAND2_157(.VSS(VSS),.VDD(VDD),.Y(I7215),.A(g815),.B(I7214));
  NAND2 NAND2_158(.VSS(VSS),.VDD(VDD),.Y(I7216),.A(g2091),.B(I7214));
  NAND2 NAND2_159(.VSS(VSS),.VDD(VDD),.Y(g3722),.A(I7215),.B(I7216));
  NAND2 NAND2_160(.VSS(VSS),.VDD(VDD),.Y(I7239),.A(g1658),.B(g2134));
  NAND2 NAND2_161(.VSS(VSS),.VDD(VDD),.Y(I7240),.A(g1658),.B(I7239));
  NAND2 NAND2_162(.VSS(VSS),.VDD(VDD),.Y(I7241),.A(g2134),.B(I7239));
  NAND2 NAND2_163(.VSS(VSS),.VDD(VDD),.Y(g3767),.A(I7240),.B(I7241));
  NAND2 NAND2_164(.VSS(VSS),.VDD(VDD),.Y(I7268),.A(g2486),.B(g955));
  NAND2 NAND2_165(.VSS(VSS),.VDD(VDD),.Y(I7269),.A(g2486),.B(I7268));
  NAND2 NAND2_166(.VSS(VSS),.VDD(VDD),.Y(I7270),.A(g955),.B(I7268));
  NAND2 NAND2_167(.VSS(VSS),.VDD(VDD),.Y(g3811),.A(I7269),.B(I7270));
  NAND2 NAND2_168(.VSS(VSS),.VDD(VDD),.Y(I7277),.A(g2497),.B(g1898));
  NAND2 NAND2_169(.VSS(VSS),.VDD(VDD),.Y(I7278),.A(g2497),.B(I7277));
  NAND2 NAND2_170(.VSS(VSS),.VDD(VDD),.Y(I7279),.A(g1898),.B(I7277));
  NAND2 NAND2_171(.VSS(VSS),.VDD(VDD),.Y(g3818),.A(I7278),.B(I7279));
  NAND2 NAND2_172(.VSS(VSS),.VDD(VDD),.Y(g3883),.A(g2276),.B(g3188));
  NAND2 NAND2_173(.VSS(VSS),.VDD(VDD),.Y(I7421),.A(g2525),.B(g2703));
  NAND2 NAND2_174(.VSS(VSS),.VDD(VDD),.Y(I7422),.A(g2525),.B(I7421));
  NAND2 NAND2_175(.VSS(VSS),.VDD(VDD),.Y(I7423),.A(g2703),.B(I7421));
  NAND2 NAND2_176(.VSS(VSS),.VDD(VDD),.Y(g3886),.A(I7422),.B(I7423));
  NAND2 NAND2_177(.VSS(VSS),.VDD(VDD),.Y(I7428),.A(g3222),.B(g1541));
  NAND2 NAND2_178(.VSS(VSS),.VDD(VDD),.Y(I7429),.A(g3222),.B(I7428));
  NAND2 NAND2_179(.VSS(VSS),.VDD(VDD),.Y(I7430),.A(g1541),.B(I7428));
  NAND2 NAND2_180(.VSS(VSS),.VDD(VDD),.Y(g3887),.A(I7429),.B(I7430));
  NAND2 NAND2_181(.VSS(VSS),.VDD(VDD),.Y(I7436),.A(g2517),.B(g3822));
  NAND2 NAND2_182(.VSS(VSS),.VDD(VDD),.Y(I7437),.A(g2517),.B(I7436));
  NAND2 NAND2_183(.VSS(VSS),.VDD(VDD),.Y(I7438),.A(g3822),.B(I7436));
  NAND2 NAND2_184(.VSS(VSS),.VDD(VDD),.Y(g3889),.A(I7437),.B(I7438));
  NAND2 NAND2_185(.VSS(VSS),.VDD(VDD),.Y(I7443),.A(g2973),.B(g1701));
  NAND2 NAND2_186(.VSS(VSS),.VDD(VDD),.Y(I7444),.A(g2973),.B(I7443));
  NAND2 NAND2_187(.VSS(VSS),.VDD(VDD),.Y(I7445),.A(g1701),.B(I7443));
  NAND2 NAND2_188(.VSS(VSS),.VDD(VDD),.Y(g3890),.A(I7444),.B(I7445));
  NAND2 NAND2_189(.VSS(VSS),.VDD(VDD),.Y(I7452),.A(g3226),.B(g1106));
  NAND2 NAND2_190(.VSS(VSS),.VDD(VDD),.Y(I7453),.A(g3226),.B(I7452));
  NAND2 NAND2_191(.VSS(VSS),.VDD(VDD),.Y(I7454),.A(g1106),.B(I7452));
  NAND2 NAND2_192(.VSS(VSS),.VDD(VDD),.Y(g3893),.A(I7453),.B(I7454));
  NAND2 NAND2_193(.VSS(VSS),.VDD(VDD),.Y(I7459),.A(g2506),.B(g3815));
  NAND2 NAND2_194(.VSS(VSS),.VDD(VDD),.Y(I7460),.A(g2506),.B(I7459));
  NAND2 NAND2_195(.VSS(VSS),.VDD(VDD),.Y(I7461),.A(g3815),.B(I7459));
  NAND2 NAND2_196(.VSS(VSS),.VDD(VDD),.Y(g3894),.A(I7460),.B(I7461));
  NAND2 NAND2_197(.VSS(VSS),.VDD(VDD),.Y(I7466),.A(g2982),.B(g1704));
  NAND2 NAND2_198(.VSS(VSS),.VDD(VDD),.Y(I7467),.A(g2982),.B(I7466));
  NAND2 NAND2_199(.VSS(VSS),.VDD(VDD),.Y(I7468),.A(g1704),.B(I7466));
  NAND2 NAND2_200(.VSS(VSS),.VDD(VDD),.Y(g3895),.A(I7467),.B(I7468));
  NAND2 NAND2_201(.VSS(VSS),.VDD(VDD),.Y(I7478),.A(g2502),.B(g3808));
  NAND2 NAND2_202(.VSS(VSS),.VDD(VDD),.Y(I7479),.A(g2502),.B(I7478));
  NAND2 NAND2_203(.VSS(VSS),.VDD(VDD),.Y(I7480),.A(g3808),.B(I7478));
  NAND2 NAND2_204(.VSS(VSS),.VDD(VDD),.Y(g3899),.A(I7479),.B(I7480));
  NAND2 NAND2_205(.VSS(VSS),.VDD(VDD),.Y(I7485),.A(g2989),.B(g1708));
  NAND2 NAND2_206(.VSS(VSS),.VDD(VDD),.Y(I7486),.A(g2989),.B(I7485));
  NAND2 NAND2_207(.VSS(VSS),.VDD(VDD),.Y(I7487),.A(g1708),.B(I7485));
  NAND2 NAND2_208(.VSS(VSS),.VDD(VDD),.Y(g3900),.A(I7486),.B(I7487));
  NAND2 NAND2_209(.VSS(VSS),.VDD(VDD),.Y(I7503),.A(g2498),.B(g3802));
  NAND2 NAND2_210(.VSS(VSS),.VDD(VDD),.Y(I7504),.A(g2498),.B(I7503));
  NAND2 NAND2_211(.VSS(VSS),.VDD(VDD),.Y(I7505),.A(g3802),.B(I7503));
  NAND2 NAND2_212(.VSS(VSS),.VDD(VDD),.Y(g3906),.A(I7504),.B(I7505));
  NAND2 NAND2_213(.VSS(VSS),.VDD(VDD),.Y(I7510),.A(g2992),.B(g1711));
  NAND2 NAND2_214(.VSS(VSS),.VDD(VDD),.Y(I7511),.A(g2992),.B(I7510));
  NAND2 NAND2_215(.VSS(VSS),.VDD(VDD),.Y(I7512),.A(g1711),.B(I7510));
  NAND2 NAND2_216(.VSS(VSS),.VDD(VDD),.Y(g3907),.A(I7511),.B(I7512));
  NAND2 NAND2_217(.VSS(VSS),.VDD(VDD),.Y(I7531),.A(g2487),.B(g3787));
  NAND2 NAND2_218(.VSS(VSS),.VDD(VDD),.Y(I7532),.A(g2487),.B(I7531));
  NAND2 NAND2_219(.VSS(VSS),.VDD(VDD),.Y(I7533),.A(g3787),.B(I7531));
  NAND2 NAND2_220(.VSS(VSS),.VDD(VDD),.Y(g3914),.A(I7532),.B(I7533));
  NAND2 NAND2_221(.VSS(VSS),.VDD(VDD),.Y(I7538),.A(g2996),.B(g1715));
  NAND2 NAND2_222(.VSS(VSS),.VDD(VDD),.Y(I7539),.A(g2996),.B(I7538));
  NAND2 NAND2_223(.VSS(VSS),.VDD(VDD),.Y(I7540),.A(g1715),.B(I7538));
  NAND2 NAND2_224(.VSS(VSS),.VDD(VDD),.Y(g3915),.A(I7539),.B(I7540));
  NAND2 NAND2_225(.VSS(VSS),.VDD(VDD),.Y(I7567),.A(g2481),.B(g3780));
  NAND2 NAND2_226(.VSS(VSS),.VDD(VDD),.Y(I7568),.A(g2481),.B(I7567));
  NAND2 NAND2_227(.VSS(VSS),.VDD(VDD),.Y(I7569),.A(g3780),.B(I7567));
  NAND2 NAND2_228(.VSS(VSS),.VDD(VDD),.Y(g3924),.A(I7568),.B(I7569));
  NAND2 NAND2_229(.VSS(VSS),.VDD(VDD),.Y(I7574),.A(g2999),.B(g1718));
  NAND2 NAND2_230(.VSS(VSS),.VDD(VDD),.Y(I7575),.A(g2999),.B(I7574));
  NAND2 NAND2_231(.VSS(VSS),.VDD(VDD),.Y(I7576),.A(g1718),.B(I7574));
  NAND2 NAND2_232(.VSS(VSS),.VDD(VDD),.Y(g3925),.A(I7575),.B(I7576));
  NAND2 NAND2_233(.VSS(VSS),.VDD(VDD),.Y(I7609),.A(g2471),.B(g3771));
  NAND2 NAND2_234(.VSS(VSS),.VDD(VDD),.Y(I7610),.A(g2471),.B(I7609));
  NAND2 NAND2_235(.VSS(VSS),.VDD(VDD),.Y(I7611),.A(g3771),.B(I7609));
  NAND2 NAND2_236(.VSS(VSS),.VDD(VDD),.Y(g3938),.A(I7610),.B(I7611));
  NAND2 NAND2_237(.VSS(VSS),.VDD(VDD),.Y(I7616),.A(g3008),.B(g1721));
  NAND2 NAND2_238(.VSS(VSS),.VDD(VDD),.Y(I7617),.A(g3008),.B(I7616));
  NAND2 NAND2_239(.VSS(VSS),.VDD(VDD),.Y(I7618),.A(g1721),.B(I7616));
  NAND2 NAND2_240(.VSS(VSS),.VDD(VDD),.Y(g3939),.A(I7617),.B(I7618));
  NAND2 NAND2_241(.VSS(VSS),.VDD(VDD),.Y(I7891),.A(g2979),.B(g1499));
  NAND2 NAND2_242(.VSS(VSS),.VDD(VDD),.Y(I7892),.A(g2979),.B(I7891));
  NAND2 NAND2_243(.VSS(VSS),.VDD(VDD),.Y(I7893),.A(g1499),.B(I7891));
  NAND2 NAND2_244(.VSS(VSS),.VDD(VDD),.Y(g4090),.A(I7892),.B(I7893));
  NAND2 NAND2_245(.VSS(VSS),.VDD(VDD),.Y(I7937),.A(g3614),.B(g1138));
  NAND2 NAND2_246(.VSS(VSS),.VDD(VDD),.Y(I7938),.A(g3614),.B(I7937));
  NAND2 NAND2_247(.VSS(VSS),.VDD(VDD),.Y(I7939),.A(g1138),.B(I7937));
  NAND2 NAND2_248(.VSS(VSS),.VDD(VDD),.Y(g4110),.A(I7938),.B(I7939));
  NAND2 NAND2_249(.VSS(VSS),.VDD(VDD),.Y(I8119),.A(g1904),.B(g3220));
  NAND2 NAND2_250(.VSS(VSS),.VDD(VDD),.Y(I8120),.A(g1904),.B(I8119));
  NAND2 NAND2_251(.VSS(VSS),.VDD(VDD),.Y(I8121),.A(g3220),.B(I8119));
  NAND2 NAND2_252(.VSS(VSS),.VDD(VDD),.Y(g4219),.A(I8120),.B(I8121));
  NAND2 NAND2_253(.VSS(VSS),.VDD(VDD),.Y(I8132),.A(g3232),.B(g1646));
  NAND2 NAND2_254(.VSS(VSS),.VDD(VDD),.Y(I8133),.A(g3232),.B(I8132));
  NAND2 NAND2_255(.VSS(VSS),.VDD(VDD),.Y(I8134),.A(g1646),.B(I8132));
  NAND2 NAND2_256(.VSS(VSS),.VDD(VDD),.Y(g4227),.A(I8133),.B(I8134));
  NAND2 NAND2_257(.VSS(VSS),.VDD(VDD),.Y(g4228),.A(g1408),.B(g2665));
  NAND2 NAND2_258(.VSS(VSS),.VDD(VDD),.Y(g4231),.A(g2276),.B(g3258));
  NAND2 NAND2_259(.VSS(VSS),.VDD(VDD),.Y(g4235),.A(g1415),.B(g2668));
  NAND2 NAND2_260(.VSS(VSS),.VDD(VDD),.Y(I8150),.A(g3229),.B(g38));
  NAND2 NAND2_261(.VSS(VSS),.VDD(VDD),.Y(I8151),.A(g3229),.B(I8150));
  NAND2 NAND2_262(.VSS(VSS),.VDD(VDD),.Y(I8152),.A(g38),.B(I8150));
  NAND2 NAND2_263(.VSS(VSS),.VDD(VDD),.Y(g4237),.A(I8151),.B(I8152));
  NAND2 NAND2_264(.VSS(VSS),.VDD(VDD),.Y(I8164),.A(g1943),.B(g3231));
  NAND2 NAND2_265(.VSS(VSS),.VDD(VDD),.Y(I8165),.A(g1943),.B(I8164));
  NAND2 NAND2_266(.VSS(VSS),.VDD(VDD),.Y(I8166),.A(g3231),.B(I8164));
  NAND2 NAND2_267(.VSS(VSS),.VDD(VDD),.Y(g4243),.A(I8165),.B(I8166));
  NAND2 NAND2_268(.VSS(VSS),.VDD(VDD),.Y(g4244),.A(g3549),.B(g3533));
  NAND2 NAND2_269(.VSS(VSS),.VDD(VDD),.Y(g4252),.A(g2276),.B(g3313));
  NAND2 NAND2_270(.VSS(VSS),.VDD(VDD),.Y(g4256),.A(g3233),.B(g1444));
  NAND2 NAND2_271(.VSS(VSS),.VDD(VDD),.Y(g4263),.A(g3260),.B(g1435));
  NAND2 NAND2_272(.VSS(VSS),.VDD(VDD),.Y(I8243),.A(g2011),.B(g3506));
  NAND2 NAND2_273(.VSS(VSS),.VDD(VDD),.Y(I8244),.A(g2011),.B(I8243));
  NAND2 NAND2_274(.VSS(VSS),.VDD(VDD),.Y(I8245),.A(g3506),.B(I8243));
  NAND2 NAND2_275(.VSS(VSS),.VDD(VDD),.Y(g4294),.A(I8244),.B(I8245));
  NAND2 NAND2_276(.VSS(VSS),.VDD(VDD),.Y(I8253),.A(g2454),.B(g3825));
  NAND2 NAND2_277(.VSS(VSS),.VDD(VDD),.Y(I8254),.A(g2454),.B(I8253));
  NAND2 NAND2_278(.VSS(VSS),.VDD(VDD),.Y(I8255),.A(g3825),.B(I8253));
  NAND2 NAND2_279(.VSS(VSS),.VDD(VDD),.Y(g4298),.A(I8254),.B(I8255));
  NAND3 NAND3_0(.VSS(VSS),.VDD(VDD),.Y(g4305),.A(g3712),.B(g3700),.C(g3732));
  NAND3 NAND3_1(.VSS(VSS),.VDD(VDD),.Y(g4309),.A(g3002),.B(g3124),.C(g3659));
  NAND2 NAND2_280(.VSS(VSS),.VDD(VDD),.Y(g4310),.A(g3666),.B(g2460));
  NAND2 NAND2_281(.VSS(VSS),.VDD(VDD),.Y(g4313),.A(g3712),.B(g3700));
  NAND2 NAND2_282(.VSS(VSS),.VDD(VDD),.Y(g4332),.A(g3681),.B(g2368));
  NAND2 NAND2_283(.VSS(VSS),.VDD(VDD),.Y(I8326),.A(g2011),.B(g2721));
  NAND2 NAND2_284(.VSS(VSS),.VDD(VDD),.Y(I8327),.A(g2011),.B(I8326));
  NAND2 NAND2_285(.VSS(VSS),.VDD(VDD),.Y(I8328),.A(g2721),.B(I8326));
  NAND2 NAND2_286(.VSS(VSS),.VDD(VDD),.Y(g4359),.A(I8327),.B(I8328));
  NAND2 NAND2_287(.VSS(VSS),.VDD(VDD),.Y(I8338),.A(g2966),.B(g1698));
  NAND2 NAND2_288(.VSS(VSS),.VDD(VDD),.Y(I8339),.A(g2966),.B(I8338));
  NAND2 NAND2_289(.VSS(VSS),.VDD(VDD),.Y(I8340),.A(g1698),.B(I8338));
  NAND2 NAND2_290(.VSS(VSS),.VDD(VDD),.Y(g4363),.A(I8339),.B(I8340));
  NAND2 NAND2_291(.VSS(VSS),.VDD(VDD),.Y(I8392),.A(g2949),.B(g1925));
  NAND2 NAND2_292(.VSS(VSS),.VDD(VDD),.Y(I8393),.A(g2949),.B(I8392));
  NAND2 NAND2_293(.VSS(VSS),.VDD(VDD),.Y(I8394),.A(g1925),.B(I8392));
  NAND2 NAND2_294(.VSS(VSS),.VDD(VDD),.Y(g4399),.A(I8393),.B(I8394));
  NAND2 NAND2_295(.VSS(VSS),.VDD(VDD),.Y(I8470),.A(g2525),.B(g2821));
  NAND2 NAND2_296(.VSS(VSS),.VDD(VDD),.Y(I8471),.A(g2525),.B(I8470));
  NAND2 NAND2_297(.VSS(VSS),.VDD(VDD),.Y(I8472),.A(g2821),.B(I8470));
  NAND2 NAND2_298(.VSS(VSS),.VDD(VDD),.Y(g4456),.A(I8471),.B(I8472));
  NAND2 NAND2_299(.VSS(VSS),.VDD(VDD),.Y(I8502),.A(g2986),.B(g2038));
  NAND2 NAND2_300(.VSS(VSS),.VDD(VDD),.Y(I8503),.A(g2986),.B(I8502));
  NAND2 NAND2_301(.VSS(VSS),.VDD(VDD),.Y(I8504),.A(g2038),.B(I8502));
  NAND2 NAND2_302(.VSS(VSS),.VDD(VDD),.Y(g4474),.A(I8503),.B(I8504));
  NAND2 NAND2_303(.VSS(VSS),.VDD(VDD),.Y(I8510),.A(g2517),.B(g2807));
  NAND2 NAND2_304(.VSS(VSS),.VDD(VDD),.Y(I8511),.A(g2517),.B(I8510));
  NAND2 NAND2_305(.VSS(VSS),.VDD(VDD),.Y(I8512),.A(g2807),.B(I8510));
  NAND2 NAND2_306(.VSS(VSS),.VDD(VDD),.Y(g4476),.A(I8511),.B(I8512));
  NAND2 NAND2_307(.VSS(VSS),.VDD(VDD),.Y(I8536),.A(g2506),.B(g2798));
  NAND2 NAND2_308(.VSS(VSS),.VDD(VDD),.Y(I8537),.A(g2506),.B(I8536));
  NAND2 NAND2_309(.VSS(VSS),.VDD(VDD),.Y(I8538),.A(g2798),.B(I8536));
  NAND2 NAND2_310(.VSS(VSS),.VDD(VDD),.Y(g4492),.A(I8537),.B(I8538));
  NAND2 NAND2_311(.VSS(VSS),.VDD(VDD),.Y(I8558),.A(g2502),.B(g2790));
  NAND2 NAND2_312(.VSS(VSS),.VDD(VDD),.Y(I8559),.A(g2502),.B(I8558));
  NAND2 NAND2_313(.VSS(VSS),.VDD(VDD),.Y(I8560),.A(g2790),.B(I8558));
  NAND2 NAND2_314(.VSS(VSS),.VDD(VDD),.Y(g4502),.A(I8559),.B(I8560));
  NAND2 NAND2_315(.VSS(VSS),.VDD(VDD),.Y(I8581),.A(g2498),.B(g2777));
  NAND2 NAND2_316(.VSS(VSS),.VDD(VDD),.Y(I8582),.A(g2498),.B(I8581));
  NAND2 NAND2_317(.VSS(VSS),.VDD(VDD),.Y(I8583),.A(g2777),.B(I8581));
  NAND2 NAND2_318(.VSS(VSS),.VDD(VDD),.Y(g4513),.A(I8582),.B(I8583));
  NAND2 NAND2_319(.VSS(VSS),.VDD(VDD),.Y(I8605),.A(g2487),.B(g2764));
  NAND2 NAND2_320(.VSS(VSS),.VDD(VDD),.Y(I8606),.A(g2487),.B(I8605));
  NAND2 NAND2_321(.VSS(VSS),.VDD(VDD),.Y(I8607),.A(g2764),.B(I8605));
  NAND2 NAND2_322(.VSS(VSS),.VDD(VDD),.Y(g4528),.A(I8606),.B(I8607));
  NAND2 NAND2_323(.VSS(VSS),.VDD(VDD),.Y(I8635),.A(g2481),.B(g2743));
  NAND2 NAND2_324(.VSS(VSS),.VDD(VDD),.Y(I8636),.A(g2481),.B(I8635));
  NAND2 NAND2_325(.VSS(VSS),.VDD(VDD),.Y(I8637),.A(g2743),.B(I8635));
  NAND2 NAND2_326(.VSS(VSS),.VDD(VDD),.Y(g4548),.A(I8636),.B(I8637));
  NAND2 NAND2_327(.VSS(VSS),.VDD(VDD),.Y(I8658),.A(g2471),.B(g2724));
  NAND2 NAND2_328(.VSS(VSS),.VDD(VDD),.Y(I8659),.A(g2471),.B(I8658));
  NAND2 NAND2_329(.VSS(VSS),.VDD(VDD),.Y(I8660),.A(g2724),.B(I8658));
  NAND2 NAND2_330(.VSS(VSS),.VDD(VDD),.Y(g4563),.A(I8659),.B(I8660));
  NAND2 NAND2_331(.VSS(VSS),.VDD(VDD),.Y(I8678),.A(g2467),.B(g2706));
  NAND2 NAND2_332(.VSS(VSS),.VDD(VDD),.Y(I8679),.A(g2467),.B(I8678));
  NAND2 NAND2_333(.VSS(VSS),.VDD(VDD),.Y(I8680),.A(g2706),.B(I8678));
  NAND2 NAND2_334(.VSS(VSS),.VDD(VDD),.Y(g4575),.A(I8679),.B(I8680));
  NAND2 NAND2_335(.VSS(VSS),.VDD(VDD),.Y(I8938),.A(g4239),.B(g1545));
  NAND2 NAND2_336(.VSS(VSS),.VDD(VDD),.Y(I8939),.A(g4239),.B(I8938));
  NAND2 NAND2_337(.VSS(VSS),.VDD(VDD),.Y(I8940),.A(g1545),.B(I8938));
  NAND2 NAND2_338(.VSS(VSS),.VDD(VDD),.Y(g4679),.A(I8939),.B(I8940));
  NAND2 NAND2_339(.VSS(VSS),.VDD(VDD),.Y(I8955),.A(g4246),.B(g1110));
  NAND2 NAND2_340(.VSS(VSS),.VDD(VDD),.Y(I8956),.A(g4246),.B(I8955));
  NAND2 NAND2_341(.VSS(VSS),.VDD(VDD),.Y(I8957),.A(g1110),.B(I8955));
  NAND2 NAND2_342(.VSS(VSS),.VDD(VDD),.Y(g4686),.A(I8956),.B(I8957));
  NAND2 NAND2_343(.VSS(VSS),.VDD(VDD),.Y(g4700),.A(g2460),.B(g4271));
  NAND3 NAND3_2(.VSS(VSS),.VDD(VDD),.Y(g4714),.A(g4344),.B(g4335),.C(g4328));
  NAND2 NAND2_344(.VSS(VSS),.VDD(VDD),.Y(I9057),.A(g4059),.B(g1504));
  NAND2 NAND2_345(.VSS(VSS),.VDD(VDD),.Y(I9058),.A(g4059),.B(I9057));
  NAND2 NAND2_346(.VSS(VSS),.VDD(VDD),.Y(I9059),.A(g1504),.B(I9057));
  NAND2 NAND2_347(.VSS(VSS),.VDD(VDD),.Y(g4741),.A(I9058),.B(I9059));
  NAND2 NAND2_348(.VSS(VSS),.VDD(VDD),.Y(I9069),.A(g4400),.B(g1149));
  NAND2 NAND2_349(.VSS(VSS),.VDD(VDD),.Y(I9070),.A(g4400),.B(I9069));
  NAND2 NAND2_350(.VSS(VSS),.VDD(VDD),.Y(I9071),.A(g1149),.B(I9069));
  NAND2 NAND2_351(.VSS(VSS),.VDD(VDD),.Y(g4745),.A(I9070),.B(I9071));
  NAND2 NAND2_352(.VSS(VSS),.VDD(VDD),.Y(I9151),.A(g3883),.B(g1649));
  NAND2 NAND2_353(.VSS(VSS),.VDD(VDD),.Y(I9152),.A(g3883),.B(I9151));
  NAND2 NAND2_354(.VSS(VSS),.VDD(VDD),.Y(I9153),.A(g1649),.B(I9151));
  NAND2 NAND2_355(.VSS(VSS),.VDD(VDD),.Y(g4810),.A(I9152),.B(I9153));
  NAND2 NAND2_356(.VSS(VSS),.VDD(VDD),.Y(I9169),.A(g1935),.B(g4244));
  NAND2 NAND2_357(.VSS(VSS),.VDD(VDD),.Y(I9170),.A(g1935),.B(I9169));
  NAND2 NAND2_358(.VSS(VSS),.VDD(VDD),.Y(I9171),.A(g4244),.B(I9169));
  NAND2 NAND2_359(.VSS(VSS),.VDD(VDD),.Y(g4820),.A(I9170),.B(I9171));
  NAND2 NAND2_360(.VSS(VSS),.VDD(VDD),.Y(g4821),.A(g4220),.B(g3605));
  NAND2 NAND2_361(.VSS(VSS),.VDD(VDD),.Y(I9181),.A(g4231),.B(g2007));
  NAND2 NAND2_362(.VSS(VSS),.VDD(VDD),.Y(I9182),.A(g4231),.B(I9181));
  NAND2 NAND2_363(.VSS(VSS),.VDD(VDD),.Y(I9183),.A(g2007),.B(I9181));
  NAND2 NAND2_364(.VSS(VSS),.VDD(VDD),.Y(g4824),.A(I9182),.B(I9183));
  NAND3 NAND3_3(.VSS(VSS),.VDD(VDD),.Y(g4831),.A(g3635),.B(g3605),.C(g4220));
  NAND2 NAND2_365(.VSS(VSS),.VDD(VDD),.Y(I9194),.A(g4252),.B(g1652));
  NAND2 NAND2_366(.VSS(VSS),.VDD(VDD),.Y(I9195),.A(g4252),.B(I9194));
  NAND2 NAND2_367(.VSS(VSS),.VDD(VDD),.Y(I9196),.A(g1652),.B(I9194));
  NAND2 NAND2_368(.VSS(VSS),.VDD(VDD),.Y(g4835),.A(I9195),.B(I9196));
  NAND2 NAND2_369(.VSS(VSS),.VDD(VDD),.Y(g4836),.A(g4288),.B(g1879));
  NAND2 NAND2_370(.VSS(VSS),.VDD(VDD),.Y(g4839),.A(g1879),.B(g4269));
  NAND2 NAND2_371(.VSS(VSS),.VDD(VDD),.Y(g4869),.A(g4254),.B(g3533));
  NAND4 NAND4_0(.VSS(VSS),.VDD(VDD),.Y(g4871),.A(g3635),.B(g3605),.C(g4220),.D(g3644));
  NAND4 NAND4_1(.VSS(VSS),.VDD(VDD),.Y(g4879),.A(g2595),.B(g2584),.C(g4270),.D(g4281));
  NAND2 NAND2_372(.VSS(VSS),.VDD(VDD),.Y(g4880),.A(g4287),.B(g1879));
  NAND2 NAND2_373(.VSS(VSS),.VDD(VDD),.Y(g4881),.A(g2460),.B(g4315));
  NAND2 NAND2_374(.VSS(VSS),.VDD(VDD),.Y(I9233),.A(g4310),.B(g2180));
  NAND2 NAND2_375(.VSS(VSS),.VDD(VDD),.Y(I9234),.A(g4310),.B(I9233));
  NAND2 NAND2_376(.VSS(VSS),.VDD(VDD),.Y(I9235),.A(g2180),.B(I9233));
  NAND2 NAND2_377(.VSS(VSS),.VDD(VDD),.Y(g4887),.A(I9234),.B(I9235));
  NAND2 NAND2_378(.VSS(VSS),.VDD(VDD),.Y(I9241),.A(g2540),.B(g4305));
  NAND2 NAND2_379(.VSS(VSS),.VDD(VDD),.Y(I9242),.A(g2540),.B(I9241));
  NAND2 NAND2_380(.VSS(VSS),.VDD(VDD),.Y(I9243),.A(g4305),.B(I9241));
  NAND2 NAND2_381(.VSS(VSS),.VDD(VDD),.Y(g4889),.A(I9242),.B(I9243));
  NAND2 NAND2_382(.VSS(VSS),.VDD(VDD),.Y(g4893),.A(g2460),.B(g4312));
  NAND2 NAND2_383(.VSS(VSS),.VDD(VDD),.Y(g4905),.A(g4282),.B(g3533));
  NAND2 NAND2_384(.VSS(VSS),.VDD(VDD),.Y(g4910),.A(g2460),.B(g4314));
  NAND2 NAND2_385(.VSS(VSS),.VDD(VDD),.Y(g4911),.A(g4320),.B(g2044));
  NAND2 NAND2_386(.VSS(VSS),.VDD(VDD),.Y(I9276),.A(g2533),.B(g4313));
  NAND2 NAND2_387(.VSS(VSS),.VDD(VDD),.Y(I9277),.A(g2533),.B(I9276));
  NAND2 NAND2_388(.VSS(VSS),.VDD(VDD),.Y(I9278),.A(g4313),.B(I9276));
  NAND2 NAND2_389(.VSS(VSS),.VDD(VDD),.Y(g4912),.A(I9277),.B(I9278));
  NAND2 NAND2_390(.VSS(VSS),.VDD(VDD),.Y(g4954),.A(g4319),.B(g2460));
  NAND2 NAND2_391(.VSS(VSS),.VDD(VDD),.Y(I9381),.A(g4062),.B(g1908));
  NAND2 NAND2_392(.VSS(VSS),.VDD(VDD),.Y(I9382),.A(g4062),.B(I9381));
  NAND2 NAND2_393(.VSS(VSS),.VDD(VDD),.Y(I9383),.A(g1908),.B(I9381));
  NAND2 NAND2_394(.VSS(VSS),.VDD(VDD),.Y(g5035),.A(I9382),.B(I9383));
  NAND2 NAND2_395(.VSS(VSS),.VDD(VDD),.Y(I9475),.A(g4038),.B(g1942));
  NAND2 NAND2_396(.VSS(VSS),.VDD(VDD),.Y(I9476),.A(g4038),.B(I9475));
  NAND2 NAND2_397(.VSS(VSS),.VDD(VDD),.Y(I9477),.A(g1942),.B(I9475));
  NAND2 NAND2_398(.VSS(VSS),.VDD(VDD),.Y(g5095),.A(I9476),.B(I9477));
  NAND2 NAND2_399(.VSS(VSS),.VDD(VDD),.Y(I9547),.A(g1952),.B(g4307));
  NAND2 NAND2_400(.VSS(VSS),.VDD(VDD),.Y(I9548),.A(g1952),.B(I9547));
  NAND2 NAND2_401(.VSS(VSS),.VDD(VDD),.Y(I9549),.A(g4307),.B(I9547));
  NAND2 NAND2_402(.VSS(VSS),.VDD(VDD),.Y(g5141),.A(I9548),.B(I9549));
  NAND2 NAND2_403(.VSS(VSS),.VDD(VDD),.Y(I9691),.A(g5096),.B(g1037));
  NAND2 NAND2_404(.VSS(VSS),.VDD(VDD),.Y(I9692),.A(g5096),.B(I9691));
  NAND2 NAND2_405(.VSS(VSS),.VDD(VDD),.Y(I9693),.A(g1037),.B(I9691));
  NAND2 NAND2_406(.VSS(VSS),.VDD(VDD),.Y(g5189),.A(I9692),.B(I9693));
  NAND2 NAND2_407(.VSS(VSS),.VDD(VDD),.Y(I9745),.A(g4826),.B(g1549));
  NAND2 NAND2_408(.VSS(VSS),.VDD(VDD),.Y(I9746),.A(g4826),.B(I9745));
  NAND2 NAND2_409(.VSS(VSS),.VDD(VDD),.Y(I9747),.A(g1549),.B(I9745));
  NAND2 NAND2_410(.VSS(VSS),.VDD(VDD),.Y(g5239),.A(I9746),.B(I9747));
  NAND2 NAND2_411(.VSS(VSS),.VDD(VDD),.Y(I9767),.A(g4832),.B(g1114));
  NAND2 NAND2_412(.VSS(VSS),.VDD(VDD),.Y(I9768),.A(g4832),.B(I9767));
  NAND2 NAND2_413(.VSS(VSS),.VDD(VDD),.Y(I9769),.A(g1114),.B(I9767));
  NAND2 NAND2_414(.VSS(VSS),.VDD(VDD),.Y(g5257),.A(I9768),.B(I9769));
  NAND3 NAND3_4(.VSS(VSS),.VDD(VDD),.Y(g5284),.A(g4344),.B(g4335),.C(g4963));
  NAND3 NAND3_5(.VSS(VSS),.VDD(VDD),.Y(g5291),.A(g4344),.B(g5002),.C(g4963));
  NAND3 NAND3_6(.VSS(VSS),.VDD(VDD),.Y(g5305),.A(g5009),.B(g4335),.C(g4328));
  NAND3 NAND3_7(.VSS(VSS),.VDD(VDD),.Y(g5310),.A(g5009),.B(g4335),.C(g4963));
  NAND3 NAND3_8(.VSS(VSS),.VDD(VDD),.Y(g5312),.A(g5009),.B(g5002),.C(g4963));
  NAND2 NAND2_415(.VSS(VSS),.VDD(VDD),.Y(I9826),.A(g4729),.B(g1509));
  NAND2 NAND2_416(.VSS(VSS),.VDD(VDD),.Y(I9827),.A(g4729),.B(I9826));
  NAND2 NAND2_417(.VSS(VSS),.VDD(VDD),.Y(I9828),.A(g1509),.B(I9826));
  NAND2 NAND2_418(.VSS(VSS),.VDD(VDD),.Y(g5363),.A(I9827),.B(I9828));
  NAND2 NAND2_419(.VSS(VSS),.VDD(VDD),.Y(g5512),.A(g1879),.B(g4877));
  NAND2 NAND2_420(.VSS(VSS),.VDD(VDD),.Y(g5538),.A(g5132),.B(g1266));
  NAND2 NAND2_421(.VSS(VSS),.VDD(VDD),.Y(I9946),.A(g2128),.B(g4905));
  NAND2 NAND2_422(.VSS(VSS),.VDD(VDD),.Y(I9947),.A(g2128),.B(I9946));
  NAND2 NAND2_423(.VSS(VSS),.VDD(VDD),.Y(I9948),.A(g4905),.B(I9946));
  NAND2 NAND2_424(.VSS(VSS),.VDD(VDD),.Y(g5539),.A(I9947),.B(I9948));
  NAND2 NAND2_425(.VSS(VSS),.VDD(VDD),.Y(I9953),.A(g2131),.B(g4831));
  NAND2 NAND2_426(.VSS(VSS),.VDD(VDD),.Y(I9954),.A(g2131),.B(I9953));
  NAND2 NAND2_427(.VSS(VSS),.VDD(VDD),.Y(I9955),.A(g4831),.B(I9953));
  NAND2 NAND2_428(.VSS(VSS),.VDD(VDD),.Y(g5540),.A(I9954),.B(I9955));
  NAND2 NAND2_429(.VSS(VSS),.VDD(VDD),.Y(I9963),.A(g1938),.B(g4869));
  NAND2 NAND2_430(.VSS(VSS),.VDD(VDD),.Y(I9964),.A(g1938),.B(I9963));
  NAND2 NAND2_431(.VSS(VSS),.VDD(VDD),.Y(I9965),.A(g4869),.B(I9963));
  NAND2 NAND2_432(.VSS(VSS),.VDD(VDD),.Y(g5546),.A(I9964),.B(I9965));
  NAND2 NAND2_433(.VSS(VSS),.VDD(VDD),.Y(g5550),.A(g1879),.B(g4830));
  NAND2 NAND2_434(.VSS(VSS),.VDD(VDD),.Y(I9978),.A(g4880),.B(g2092));
  NAND2 NAND2_435(.VSS(VSS),.VDD(VDD),.Y(I9979),.A(g4880),.B(I9978));
  NAND2 NAND2_436(.VSS(VSS),.VDD(VDD),.Y(I9980),.A(g2092),.B(I9978));
  NAND2 NAND2_437(.VSS(VSS),.VDD(VDD),.Y(g5555),.A(I9979),.B(I9980));
  NAND2 NAND2_438(.VSS(VSS),.VDD(VDD),.Y(I9985),.A(g4836),.B(g2096));
  NAND2 NAND2_439(.VSS(VSS),.VDD(VDD),.Y(I9986),.A(g4836),.B(I9985));
  NAND2 NAND2_440(.VSS(VSS),.VDD(VDD),.Y(I9987),.A(g2096),.B(I9985));
  NAND2 NAND2_441(.VSS(VSS),.VDD(VDD),.Y(g5556),.A(I9986),.B(I9987));
  NAND2 NAND2_442(.VSS(VSS),.VDD(VDD),.Y(I9992),.A(g2145),.B(g4871));
  NAND2 NAND2_443(.VSS(VSS),.VDD(VDD),.Y(I9993),.A(g2145),.B(I9992));
  NAND2 NAND2_444(.VSS(VSS),.VDD(VDD),.Y(I9994),.A(g4871),.B(I9992));
  NAND2 NAND2_445(.VSS(VSS),.VDD(VDD),.Y(g5557),.A(I9993),.B(I9994));
  NAND2 NAND2_446(.VSS(VSS),.VDD(VDD),.Y(I9999),.A(g4839),.B(g1929));
  NAND2 NAND2_447(.VSS(VSS),.VDD(VDD),.Y(I10000),.A(g4839),.B(I9999));
  NAND2 NAND2_448(.VSS(VSS),.VDD(VDD),.Y(I10001),.A(g1929),.B(I9999));
  NAND2 NAND2_449(.VSS(VSS),.VDD(VDD),.Y(g5558),.A(I10000),.B(I10001));
  NAND2 NAND2_450(.VSS(VSS),.VDD(VDD),.Y(g5559),.A(g5132),.B(g1257));
  NAND2 NAND2_451(.VSS(VSS),.VDD(VDD),.Y(I10009),.A(g1949),.B(g4821));
  NAND2 NAND2_452(.VSS(VSS),.VDD(VDD),.Y(I10010),.A(g1949),.B(I10009));
  NAND2 NAND2_453(.VSS(VSS),.VDD(VDD),.Y(I10011),.A(g4821),.B(I10009));
  NAND2 NAND2_454(.VSS(VSS),.VDD(VDD),.Y(g5562),.A(I10010),.B(I10011));
  NAND2 NAND2_455(.VSS(VSS),.VDD(VDD),.Y(I10017),.A(g4700),.B(g2174));
  NAND2 NAND2_456(.VSS(VSS),.VDD(VDD),.Y(I10018),.A(g4700),.B(I10017));
  NAND2 NAND2_457(.VSS(VSS),.VDD(VDD),.Y(I10019),.A(g2174),.B(I10017));
  NAND2 NAND2_458(.VSS(VSS),.VDD(VDD),.Y(g5564),.A(I10018),.B(I10019));
  NAND2 NAND2_459(.VSS(VSS),.VDD(VDD),.Y(g5565),.A(g2044),.B(g4933));
  NAND2 NAND2_460(.VSS(VSS),.VDD(VDD),.Y(g5567),.A(g1879),.B(g4883));
  NAND3 NAND3_9(.VSS(VSS),.VDD(VDD),.Y(g5568),.A(g2044),.B(g4902),.C(g4320));
  NAND2 NAND2_461(.VSS(VSS),.VDD(VDD),.Y(I10038),.A(g4893),.B(g2202));
  NAND2 NAND2_462(.VSS(VSS),.VDD(VDD),.Y(I10039),.A(g4893),.B(I10038));
  NAND2 NAND2_463(.VSS(VSS),.VDD(VDD),.Y(I10040),.A(g2202),.B(I10038));
  NAND2 NAND2_464(.VSS(VSS),.VDD(VDD),.Y(g5575),.A(I10039),.B(I10040));
  NAND3 NAND3_10(.VSS(VSS),.VDD(VDD),.Y(g5576),.A(g4894),.B(g4888),.C(g4884));
  NAND2 NAND2_465(.VSS(VSS),.VDD(VDD),.Y(I10060),.A(g4910),.B(g2226));
  NAND2 NAND2_466(.VSS(VSS),.VDD(VDD),.Y(I10061),.A(g4910),.B(I10060));
  NAND2 NAND2_467(.VSS(VSS),.VDD(VDD),.Y(I10062),.A(g2226),.B(I10060));
  NAND2 NAND2_468(.VSS(VSS),.VDD(VDD),.Y(g5589),.A(I10061),.B(I10062));
  NAND2 NAND2_469(.VSS(VSS),.VDD(VDD),.Y(g5590),.A(g2044),.B(g4906));
  NAND2 NAND2_470(.VSS(VSS),.VDD(VDD),.Y(I10071),.A(g4954),.B(g2253));
  NAND2 NAND2_471(.VSS(VSS),.VDD(VDD),.Y(I10072),.A(g4954),.B(I10071));
  NAND2 NAND2_472(.VSS(VSS),.VDD(VDD),.Y(I10073),.A(g2253),.B(I10071));
  NAND2 NAND2_473(.VSS(VSS),.VDD(VDD),.Y(g5594),.A(I10072),.B(I10073));
  NAND2 NAND2_474(.VSS(VSS),.VDD(VDD),.Y(I10078),.A(g4911),.B(g2256));
  NAND2 NAND2_475(.VSS(VSS),.VDD(VDD),.Y(I10079),.A(g4911),.B(I10078));
  NAND2 NAND2_476(.VSS(VSS),.VDD(VDD),.Y(I10080),.A(g2256),.B(I10078));
  NAND2 NAND2_477(.VSS(VSS),.VDD(VDD),.Y(g5595),.A(I10079),.B(I10080));
  NAND2 NAND2_478(.VSS(VSS),.VDD(VDD),.Y(I10092),.A(g4881),.B(g2177));
  NAND2 NAND2_479(.VSS(VSS),.VDD(VDD),.Y(I10093),.A(g4881),.B(I10092));
  NAND2 NAND2_480(.VSS(VSS),.VDD(VDD),.Y(I10094),.A(g2177),.B(I10092));
  NAND2 NAND2_481(.VSS(VSS),.VDD(VDD),.Y(g5605),.A(I10093),.B(I10094));
  NAND2 NAND2_482(.VSS(VSS),.VDD(VDD),.Y(g5625),.A(g2044),.B(g4957));
  NAND2 NAND2_483(.VSS(VSS),.VDD(VDD),.Y(g5632),.A(g2276),.B(g4901));
  NAND2 NAND2_484(.VSS(VSS),.VDD(VDD),.Y(g5657),.A(g5021),.B(g4381));
  NAND2 NAND2_485(.VSS(VSS),.VDD(VDD),.Y(I10142),.A(g4707),.B(g1916));
  NAND2 NAND2_486(.VSS(VSS),.VDD(VDD),.Y(I10143),.A(g4707),.B(I10142));
  NAND2 NAND2_487(.VSS(VSS),.VDD(VDD),.Y(I10144),.A(g1916),.B(I10142));
  NAND2 NAND2_488(.VSS(VSS),.VDD(VDD),.Y(g5661),.A(I10143),.B(I10144));
  NAND3 NAND3_11(.VSS(VSS),.VDD(VDD),.Y(g5672),.A(g5056),.B(g5039),.C(g5023));
  NAND2 NAND2_489(.VSS(VSS),.VDD(VDD),.Y(g5681),.A(g5132),.B(g2043));
  NAND2 NAND2_490(.VSS(VSS),.VDD(VDD),.Y(g5686),.A(g5132),.B(g1263));
  NAND2 NAND2_491(.VSS(VSS),.VDD(VDD),.Y(I10196),.A(g4724),.B(g1958));
  NAND2 NAND2_492(.VSS(VSS),.VDD(VDD),.Y(I10197),.A(g4724),.B(I10196));
  NAND2 NAND2_493(.VSS(VSS),.VDD(VDD),.Y(I10198),.A(g1958),.B(I10196));
  NAND2 NAND2_494(.VSS(VSS),.VDD(VDD),.Y(g5689),.A(I10197),.B(I10198));
  NAND2 NAND2_495(.VSS(VSS),.VDD(VDD),.Y(g5697),.A(g2044),.B(g5005));
  NAND2 NAND2_496(.VSS(VSS),.VDD(VDD),.Y(I10223),.A(g2522),.B(g4895));
  NAND2 NAND2_497(.VSS(VSS),.VDD(VDD),.Y(I10224),.A(g2522),.B(I10223));
  NAND2 NAND2_498(.VSS(VSS),.VDD(VDD),.Y(I10225),.A(g4895),.B(I10223));
  NAND2 NAND2_499(.VSS(VSS),.VDD(VDD),.Y(g5712),.A(I10224),.B(I10225));
  NAND2 NAND2_500(.VSS(VSS),.VDD(VDD),.Y(I10298),.A(g5461),.B(g2562));
  NAND2 NAND2_501(.VSS(VSS),.VDD(VDD),.Y(I10299),.A(g5461),.B(I10298));
  NAND2 NAND2_502(.VSS(VSS),.VDD(VDD),.Y(I10300),.A(g2562),.B(I10298));
  NAND2 NAND2_503(.VSS(VSS),.VDD(VDD),.Y(g5747),.A(I10299),.B(I10300));
  NAND2 NAND2_504(.VSS(VSS),.VDD(VDD),.Y(I10305),.A(g5470),.B(g3019));
  NAND2 NAND2_505(.VSS(VSS),.VDD(VDD),.Y(I10306),.A(g5470),.B(I10305));
  NAND2 NAND2_506(.VSS(VSS),.VDD(VDD),.Y(I10307),.A(g3019),.B(I10305));
  NAND2 NAND2_507(.VSS(VSS),.VDD(VDD),.Y(g5748),.A(I10306),.B(I10307));
  NAND2 NAND2_508(.VSS(VSS),.VDD(VDD),.Y(I10313),.A(g5484),.B(g1041));
  NAND2 NAND2_509(.VSS(VSS),.VDD(VDD),.Y(I10314),.A(g5484),.B(I10313));
  NAND2 NAND2_510(.VSS(VSS),.VDD(VDD),.Y(I10315),.A(g1041),.B(I10313));
  NAND2 NAND2_511(.VSS(VSS),.VDD(VDD),.Y(g5750),.A(I10314),.B(I10315));
  NAND2 NAND2_512(.VSS(VSS),.VDD(VDD),.Y(I10320),.A(g5459),.B(g2573));
  NAND2 NAND2_513(.VSS(VSS),.VDD(VDD),.Y(I10321),.A(g5459),.B(I10320));
  NAND2 NAND2_514(.VSS(VSS),.VDD(VDD),.Y(I10322),.A(g2573),.B(I10320));
  NAND2 NAND2_515(.VSS(VSS),.VDD(VDD),.Y(g5751),.A(I10321),.B(I10322));
  NAND2 NAND2_516(.VSS(VSS),.VDD(VDD),.Y(I10327),.A(g5467),.B(g2562));
  NAND2 NAND2_517(.VSS(VSS),.VDD(VDD),.Y(I10328),.A(g5467),.B(I10327));
  NAND2 NAND2_518(.VSS(VSS),.VDD(VDD),.Y(I10329),.A(g2562),.B(I10327));
  NAND2 NAND2_519(.VSS(VSS),.VDD(VDD),.Y(g5752),.A(I10328),.B(I10329));
  NAND2 NAND2_520(.VSS(VSS),.VDD(VDD),.Y(I10334),.A(g5462),.B(g2573));
  NAND2 NAND2_521(.VSS(VSS),.VDD(VDD),.Y(I10335),.A(g5462),.B(I10334));
  NAND2 NAND2_522(.VSS(VSS),.VDD(VDD),.Y(I10336),.A(g2573),.B(I10334));
  NAND2 NAND2_523(.VSS(VSS),.VDD(VDD),.Y(g5753),.A(I10335),.B(I10336));
  NAND2 NAND2_524(.VSS(VSS),.VDD(VDD),.Y(I10359),.A(g5552),.B(g1118));
  NAND2 NAND2_525(.VSS(VSS),.VDD(VDD),.Y(I10360),.A(g5552),.B(I10359));
  NAND2 NAND2_526(.VSS(VSS),.VDD(VDD),.Y(I10361),.A(g1118),.B(I10359));
  NAND2 NAND2_527(.VSS(VSS),.VDD(VDD),.Y(g5762),.A(I10360),.B(I10361));
  NAND2 NAND2_528(.VSS(VSS),.VDD(VDD),.Y(I10625),.A(g5314),.B(g1514));
  NAND2 NAND2_529(.VSS(VSS),.VDD(VDD),.Y(I10626),.A(g5314),.B(I10625));
  NAND2 NAND2_530(.VSS(VSS),.VDD(VDD),.Y(I10627),.A(g1514),.B(I10625));
  NAND2 NAND2_531(.VSS(VSS),.VDD(VDD),.Y(g6023),.A(I10626),.B(I10627));
  NAND2 NAND2_532(.VSS(VSS),.VDD(VDD),.Y(I10743),.A(g5550),.B(g2100));
  NAND2 NAND2_533(.VSS(VSS),.VDD(VDD),.Y(I10744),.A(g5550),.B(I10743));
  NAND2 NAND2_534(.VSS(VSS),.VDD(VDD),.Y(I10745),.A(g2100),.B(I10743));
  NAND2 NAND2_535(.VSS(VSS),.VDD(VDD),.Y(g6119),.A(I10744),.B(I10745));
  NAND2 NAND2_536(.VSS(VSS),.VDD(VDD),.Y(I10789),.A(g5512),.B(g2170));
  NAND2 NAND2_537(.VSS(VSS),.VDD(VDD),.Y(I10790),.A(g5512),.B(I10789));
  NAND2 NAND2_538(.VSS(VSS),.VDD(VDD),.Y(I10791),.A(g2170),.B(I10789));
  NAND2 NAND2_539(.VSS(VSS),.VDD(VDD),.Y(g6142),.A(I10790),.B(I10791));
  NAND2 NAND2_540(.VSS(VSS),.VDD(VDD),.Y(I10818),.A(g5567),.B(g2039));
  NAND2 NAND2_541(.VSS(VSS),.VDD(VDD),.Y(I10819),.A(g5567),.B(I10818));
  NAND2 NAND2_542(.VSS(VSS),.VDD(VDD),.Y(I10820),.A(g2039),.B(I10818));
  NAND2 NAND2_543(.VSS(VSS),.VDD(VDD),.Y(g6153),.A(I10819),.B(I10820));
  NAND4 NAND4_2(.VSS(VSS),.VDD(VDD),.Y(g6158),.A(g3735),.B(g3716),.C(g5633),.D(g3754));
  NAND2 NAND2_544(.VSS(VSS),.VDD(VDD),.Y(I10834),.A(g5514),.B(g2584));
  NAND2 NAND2_545(.VSS(VSS),.VDD(VDD),.Y(I10835),.A(g5514),.B(I10834));
  NAND2 NAND2_546(.VSS(VSS),.VDD(VDD),.Y(I10836),.A(g2584),.B(I10834));
  NAND2 NAND2_547(.VSS(VSS),.VDD(VDD),.Y(g6159),.A(I10835),.B(I10836));
  NAND2 NAND2_548(.VSS(VSS),.VDD(VDD),.Y(g6163),.A(g5633),.B(g3716));
  NAND2 NAND2_549(.VSS(VSS),.VDD(VDD),.Y(I10847),.A(g5490),.B(g2595));
  NAND2 NAND2_550(.VSS(VSS),.VDD(VDD),.Y(I10848),.A(g5490),.B(I10847));
  NAND2 NAND2_551(.VSS(VSS),.VDD(VDD),.Y(I10849),.A(g2595),.B(I10847));
  NAND2 NAND2_552(.VSS(VSS),.VDD(VDD),.Y(g6164),.A(I10848),.B(I10849));
  NAND2 NAND2_553(.VSS(VSS),.VDD(VDD),.Y(I10854),.A(g5521),.B(g2584));
  NAND2 NAND2_554(.VSS(VSS),.VDD(VDD),.Y(I10855),.A(g5521),.B(I10854));
  NAND2 NAND2_555(.VSS(VSS),.VDD(VDD),.Y(I10856),.A(g2584),.B(I10854));
  NAND2 NAND2_556(.VSS(VSS),.VDD(VDD),.Y(g6165),.A(I10855),.B(I10856));
  NAND2 NAND2_557(.VSS(VSS),.VDD(VDD),.Y(I10866),.A(g5480),.B(g2605));
  NAND2 NAND2_558(.VSS(VSS),.VDD(VDD),.Y(I10867),.A(g5480),.B(I10866));
  NAND2 NAND2_559(.VSS(VSS),.VDD(VDD),.Y(I10868),.A(g2605),.B(I10866));
  NAND2 NAND2_560(.VSS(VSS),.VDD(VDD),.Y(g6169),.A(I10867),.B(I10868));
  NAND2 NAND2_561(.VSS(VSS),.VDD(VDD),.Y(I10873),.A(g5516),.B(g2595));
  NAND2 NAND2_562(.VSS(VSS),.VDD(VDD),.Y(I10874),.A(g5516),.B(I10873));
  NAND2 NAND2_563(.VSS(VSS),.VDD(VDD),.Y(I10875),.A(g2595),.B(I10873));
  NAND2 NAND2_564(.VSS(VSS),.VDD(VDD),.Y(g6170),.A(I10874),.B(I10875));
  NAND2 NAND2_565(.VSS(VSS),.VDD(VDD),.Y(I10888),.A(g5590),.B(g2259));
  NAND2 NAND2_566(.VSS(VSS),.VDD(VDD),.Y(I10889),.A(g5590),.B(I10888));
  NAND2 NAND2_567(.VSS(VSS),.VDD(VDD),.Y(I10890),.A(g2259),.B(I10888));
  NAND2 NAND2_568(.VSS(VSS),.VDD(VDD),.Y(g6177),.A(I10889),.B(I10890));
  NAND2 NAND2_569(.VSS(VSS),.VDD(VDD),.Y(g6178),.A(g2205),.B(g5568));
  NAND2 NAND2_570(.VSS(VSS),.VDD(VDD),.Y(I10899),.A(g5520),.B(g2752));
  NAND2 NAND2_571(.VSS(VSS),.VDD(VDD),.Y(I10900),.A(g5520),.B(I10899));
  NAND2 NAND2_572(.VSS(VSS),.VDD(VDD),.Y(I10901),.A(g2752),.B(I10899));
  NAND2 NAND2_573(.VSS(VSS),.VDD(VDD),.Y(g6180),.A(I10900),.B(I10901));
  NAND2 NAND2_574(.VSS(VSS),.VDD(VDD),.Y(I10906),.A(g5492),.B(g2605));
  NAND2 NAND2_575(.VSS(VSS),.VDD(VDD),.Y(I10907),.A(g5492),.B(I10906));
  NAND2 NAND2_576(.VSS(VSS),.VDD(VDD),.Y(I10908),.A(g2605),.B(I10906));
  NAND2 NAND2_577(.VSS(VSS),.VDD(VDD),.Y(g6181),.A(I10907),.B(I10908));
  NAND3 NAND3_12(.VSS(VSS),.VDD(VDD),.Y(g6187),.A(g5633),.B(g3735),.C(g3716));
  NAND2 NAND2_578(.VSS(VSS),.VDD(VDD),.Y(I10923),.A(g5525),.B(g2752));
  NAND2 NAND2_579(.VSS(VSS),.VDD(VDD),.Y(I10924),.A(g5525),.B(I10923));
  NAND2 NAND2_580(.VSS(VSS),.VDD(VDD),.Y(I10925),.A(g2752),.B(I10923));
  NAND2 NAND2_581(.VSS(VSS),.VDD(VDD),.Y(g6188),.A(I10924),.B(I10925));
  NAND2 NAND2_582(.VSS(VSS),.VDD(VDD),.Y(I10952),.A(g5565),.B(g2340));
  NAND2 NAND2_583(.VSS(VSS),.VDD(VDD),.Y(I10953),.A(g5565),.B(I10952));
  NAND2 NAND2_584(.VSS(VSS),.VDD(VDD),.Y(I10954),.A(g2340),.B(I10952));
  NAND2 NAND2_585(.VSS(VSS),.VDD(VDD),.Y(g6203),.A(I10953),.B(I10954));
  NAND2 NAND2_586(.VSS(VSS),.VDD(VDD),.Y(I10980),.A(g5625),.B(g2210));
  NAND2 NAND2_587(.VSS(VSS),.VDD(VDD),.Y(I10981),.A(g5625),.B(I10980));
  NAND2 NAND2_588(.VSS(VSS),.VDD(VDD),.Y(I10982),.A(g2210),.B(I10980));
  NAND2 NAND2_589(.VSS(VSS),.VDD(VDD),.Y(g6215),.A(I10981),.B(I10982));
  NAND2 NAND2_590(.VSS(VSS),.VDD(VDD),.Y(I10991),.A(g5632),.B(g2389));
  NAND2 NAND2_591(.VSS(VSS),.VDD(VDD),.Y(I10992),.A(g5632),.B(I10991));
  NAND2 NAND2_592(.VSS(VSS),.VDD(VDD),.Y(I10993),.A(g2389),.B(I10991));
  NAND2 NAND2_593(.VSS(VSS),.VDD(VDD),.Y(g6218),.A(I10992),.B(I10993));
  NAND2 NAND2_594(.VSS(VSS),.VDD(VDD),.Y(I11078),.A(g5697),.B(g2511));
  NAND2 NAND2_595(.VSS(VSS),.VDD(VDD),.Y(I11079),.A(g5697),.B(I11078));
  NAND2 NAND2_596(.VSS(VSS),.VDD(VDD),.Y(I11080),.A(g2511),.B(I11078));
  NAND2 NAND2_597(.VSS(VSS),.VDD(VDD),.Y(g6265),.A(I11079),.B(I11080));
  NAND2 NAND2_598(.VSS(VSS),.VDD(VDD),.Y(I11094),.A(g5515),.B(g2734));
  NAND2 NAND2_599(.VSS(VSS),.VDD(VDD),.Y(I11095),.A(g5515),.B(I11094));
  NAND2 NAND2_600(.VSS(VSS),.VDD(VDD),.Y(I11096),.A(g2734),.B(I11094));
  NAND2 NAND2_601(.VSS(VSS),.VDD(VDD),.Y(g6273),.A(I11095),.B(I11096));
  NAND2 NAND2_602(.VSS(VSS),.VDD(VDD),.Y(I11101),.A(g5491),.B(g2712));
  NAND2 NAND2_603(.VSS(VSS),.VDD(VDD),.Y(I11102),.A(g5491),.B(I11101));
  NAND2 NAND2_604(.VSS(VSS),.VDD(VDD),.Y(I11103),.A(g2712),.B(I11101));
  NAND2 NAND2_605(.VSS(VSS),.VDD(VDD),.Y(g6274),.A(I11102),.B(I11103));
  NAND2 NAND2_606(.VSS(VSS),.VDD(VDD),.Y(I11108),.A(g5522),.B(g2734));
  NAND2 NAND2_607(.VSS(VSS),.VDD(VDD),.Y(I11109),.A(g5522),.B(I11108));
  NAND2 NAND2_608(.VSS(VSS),.VDD(VDD),.Y(I11110),.A(g2734),.B(I11108));
  NAND2 NAND2_609(.VSS(VSS),.VDD(VDD),.Y(g6275),.A(I11109),.B(I11110));
  NAND2 NAND2_610(.VSS(VSS),.VDD(VDD),.Y(I11115),.A(g5481),.B(g3062));
  NAND2 NAND2_611(.VSS(VSS),.VDD(VDD),.Y(I11116),.A(g5481),.B(I11115));
  NAND2 NAND2_612(.VSS(VSS),.VDD(VDD),.Y(I11117),.A(g3062),.B(I11115));
  NAND2 NAND2_613(.VSS(VSS),.VDD(VDD),.Y(g6276),.A(I11116),.B(I11117));
  NAND2 NAND2_614(.VSS(VSS),.VDD(VDD),.Y(I11122),.A(g5517),.B(g2712));
  NAND2 NAND2_615(.VSS(VSS),.VDD(VDD),.Y(I11123),.A(g5517),.B(I11122));
  NAND2 NAND2_616(.VSS(VSS),.VDD(VDD),.Y(I11124),.A(g2712),.B(I11122));
  NAND2 NAND2_617(.VSS(VSS),.VDD(VDD),.Y(g6277),.A(I11123),.B(I11124));
  NAND2 NAND2_618(.VSS(VSS),.VDD(VDD),.Y(I11135),.A(g5476),.B(g3052));
  NAND2 NAND2_619(.VSS(VSS),.VDD(VDD),.Y(I11136),.A(g5476),.B(I11135));
  NAND2 NAND2_620(.VSS(VSS),.VDD(VDD),.Y(I11137),.A(g3052),.B(I11135));
  NAND2 NAND2_621(.VSS(VSS),.VDD(VDD),.Y(g6280),.A(I11136),.B(I11137));
  NAND2 NAND2_622(.VSS(VSS),.VDD(VDD),.Y(I11142),.A(g5493),.B(g3062));
  NAND2 NAND2_623(.VSS(VSS),.VDD(VDD),.Y(I11143),.A(g5493),.B(I11142));
  NAND2 NAND2_624(.VSS(VSS),.VDD(VDD),.Y(I11144),.A(g3062),.B(I11142));
  NAND2 NAND2_625(.VSS(VSS),.VDD(VDD),.Y(g6281),.A(I11143),.B(I11144));
  NAND2 NAND2_626(.VSS(VSS),.VDD(VDD),.Y(I11149),.A(g5473),.B(g3038));
  NAND2 NAND2_627(.VSS(VSS),.VDD(VDD),.Y(I11150),.A(g5473),.B(I11149));
  NAND2 NAND2_628(.VSS(VSS),.VDD(VDD),.Y(I11151),.A(g3038),.B(I11149));
  NAND2 NAND2_629(.VSS(VSS),.VDD(VDD),.Y(g6282),.A(I11150),.B(I11151));
  NAND2 NAND2_630(.VSS(VSS),.VDD(VDD),.Y(I11156),.A(g5482),.B(g3052));
  NAND2 NAND2_631(.VSS(VSS),.VDD(VDD),.Y(I11157),.A(g5482),.B(I11156));
  NAND2 NAND2_632(.VSS(VSS),.VDD(VDD),.Y(I11158),.A(g3052),.B(I11156));
  NAND2 NAND2_633(.VSS(VSS),.VDD(VDD),.Y(g6283),.A(I11157),.B(I11158));
  NAND2 NAND2_634(.VSS(VSS),.VDD(VDD),.Y(I11163),.A(g5469),.B(g3029));
  NAND2 NAND2_635(.VSS(VSS),.VDD(VDD),.Y(I11164),.A(g5469),.B(I11163));
  NAND2 NAND2_636(.VSS(VSS),.VDD(VDD),.Y(I11165),.A(g3029),.B(I11163));
  NAND2 NAND2_637(.VSS(VSS),.VDD(VDD),.Y(g6284),.A(I11164),.B(I11165));
  NAND2 NAND2_638(.VSS(VSS),.VDD(VDD),.Y(I11170),.A(g5477),.B(g3038));
  NAND2 NAND2_639(.VSS(VSS),.VDD(VDD),.Y(I11171),.A(g5477),.B(I11170));
  NAND2 NAND2_640(.VSS(VSS),.VDD(VDD),.Y(I11172),.A(g3038),.B(I11170));
  NAND2 NAND2_641(.VSS(VSS),.VDD(VDD),.Y(g6285),.A(I11171),.B(I11172));
  NAND2 NAND2_642(.VSS(VSS),.VDD(VDD),.Y(I11177),.A(g5466),.B(g3019));
  NAND2 NAND2_643(.VSS(VSS),.VDD(VDD),.Y(I11178),.A(g5466),.B(I11177));
  NAND2 NAND2_644(.VSS(VSS),.VDD(VDD),.Y(I11179),.A(g3019),.B(I11177));
  NAND2 NAND2_645(.VSS(VSS),.VDD(VDD),.Y(g6286),.A(I11178),.B(I11179));
  NAND2 NAND2_646(.VSS(VSS),.VDD(VDD),.Y(I11184),.A(g5474),.B(g3029));
  NAND2 NAND2_647(.VSS(VSS),.VDD(VDD),.Y(I11185),.A(g5474),.B(I11184));
  NAND2 NAND2_648(.VSS(VSS),.VDD(VDD),.Y(I11186),.A(g3029),.B(I11184));
  NAND2 NAND2_649(.VSS(VSS),.VDD(VDD),.Y(g6287),.A(I11185),.B(I11186));
  NAND2 NAND2_650(.VSS(VSS),.VDD(VDD),.Y(I11549),.A(g5984),.B(g1045));
  NAND2 NAND2_651(.VSS(VSS),.VDD(VDD),.Y(I11550),.A(g5984),.B(I11549));
  NAND2 NAND2_652(.VSS(VSS),.VDD(VDD),.Y(I11551),.A(g1045),.B(I11549));
  NAND2 NAND2_653(.VSS(VSS),.VDD(VDD),.Y(g6424),.A(I11550),.B(I11551));
  NAND2 NAND2_654(.VSS(VSS),.VDD(VDD),.Y(I11574),.A(g5894),.B(g1122));
  NAND2 NAND2_655(.VSS(VSS),.VDD(VDD),.Y(I11575),.A(g5894),.B(I11574));
  NAND2 NAND2_656(.VSS(VSS),.VDD(VDD),.Y(I11576),.A(g1122),.B(I11574));
  NAND2 NAND2_657(.VSS(VSS),.VDD(VDD),.Y(g6435),.A(I11575),.B(I11576));
  NAND2 NAND2_658(.VSS(VSS),.VDD(VDD),.Y(g6463),.A(g5918),.B(g5278));
  NAND2 NAND2_659(.VSS(VSS),.VDD(VDD),.Y(I11614),.A(g6239),.B(g1519));
  NAND2 NAND2_660(.VSS(VSS),.VDD(VDD),.Y(I11615),.A(g6239),.B(I11614));
  NAND2 NAND2_661(.VSS(VSS),.VDD(VDD),.Y(I11616),.A(g1519),.B(I11614));
  NAND2 NAND2_662(.VSS(VSS),.VDD(VDD),.Y(g6466),.A(I11615),.B(I11616));
  NAND2 NAND2_663(.VSS(VSS),.VDD(VDD),.Y(g6467),.A(g5956),.B(g5269));
  NAND2 NAND2_664(.VSS(VSS),.VDD(VDD),.Y(g6469),.A(g5918),.B(g5278));
  NAND2 NAND2_665(.VSS(VSS),.VDD(VDD),.Y(g6472),.A(g5971),.B(g5269));
  NAND2 NAND2_666(.VSS(VSS),.VDD(VDD),.Y(g6473),.A(g5269),.B(g5988));
  NAND2 NAND2_667(.VSS(VSS),.VDD(VDD),.Y(g6476),.A(g5939),.B(g5269));
  NAND2 NAND2_668(.VSS(VSS),.VDD(VDD),.Y(g6477),.A(g5269),.B(g5918));
  NAND2 NAND2_669(.VSS(VSS),.VDD(VDD),.Y(g6482),.A(g5269),.B(g5847));
  NAND2 NAND2_670(.VSS(VSS),.VDD(VDD),.Y(g6497),.A(g5278),.B(g5847));
  NAND2 NAND2_671(.VSS(VSS),.VDD(VDD),.Y(g6503),.A(g5269),.B(g5897));
  NAND2 NAND2_672(.VSS(VSS),.VDD(VDD),.Y(g6504),.A(g5269),.B(g5874));
  NAND2 NAND2_673(.VSS(VSS),.VDD(VDD),.Y(g6510),.A(g5278),.B(g5874));
  NAND2 NAND2_674(.VSS(VSS),.VDD(VDD),.Y(g6516),.A(g5897),.B(g5278));
  NAND2 NAND2_675(.VSS(VSS),.VDD(VDD),.Y(g6559),.A(g5814),.B(g6109));
  NAND2 NAND2_676(.VSS(VSS),.VDD(VDD),.Y(I11750),.A(g6112),.B(g1486));
  NAND2 NAND2_677(.VSS(VSS),.VDD(VDD),.Y(I11751),.A(g6112),.B(I11750));
  NAND2 NAND2_678(.VSS(VSS),.VDD(VDD),.Y(I11752),.A(g1486),.B(I11750));
  NAND2 NAND2_679(.VSS(VSS),.VDD(VDD),.Y(g6570),.A(I11751),.B(I11752));
  NAND2 NAND2_680(.VSS(VSS),.VDD(VDD),.Y(I11757),.A(g1758),.B(g6118));
  NAND2 NAND2_681(.VSS(VSS),.VDD(VDD),.Y(I11758),.A(g1758),.B(I11757));
  NAND2 NAND2_682(.VSS(VSS),.VDD(VDD),.Y(I11759),.A(g6118),.B(I11757));
  NAND2 NAND2_683(.VSS(VSS),.VDD(VDD),.Y(g6571),.A(I11758),.B(I11759));
  NAND2 NAND2_684(.VSS(VSS),.VDD(VDD),.Y(I11841),.A(g2548),.B(g6158));
  NAND2 NAND2_685(.VSS(VSS),.VDD(VDD),.Y(I11842),.A(g2548),.B(I11841));
  NAND2 NAND2_686(.VSS(VSS),.VDD(VDD),.Y(I11843),.A(g6158),.B(I11841));
  NAND2 NAND2_687(.VSS(VSS),.VDD(VDD),.Y(g6615),.A(I11842),.B(I11843));
  NAND2 NAND2_688(.VSS(VSS),.VDD(VDD),.Y(I11873),.A(g2543),.B(g6187));
  NAND2 NAND2_689(.VSS(VSS),.VDD(VDD),.Y(I11874),.A(g2543),.B(I11873));
  NAND2 NAND2_690(.VSS(VSS),.VDD(VDD),.Y(I11875),.A(g6187),.B(I11873));
  NAND2 NAND2_691(.VSS(VSS),.VDD(VDD),.Y(g6627),.A(I11874),.B(I11875));
  NAND2 NAND2_692(.VSS(VSS),.VDD(VDD),.Y(g6680),.A(g5403),.B(g6252));
  NAND2 NAND2_693(.VSS(VSS),.VDD(VDD),.Y(I12015),.A(g5874),.B(g5847));
  NAND2 NAND2_694(.VSS(VSS),.VDD(VDD),.Y(I12016),.A(g5874),.B(I12015));
  NAND2 NAND2_695(.VSS(VSS),.VDD(VDD),.Y(I12017),.A(g5847),.B(I12015));
  NAND2 NAND2_696(.VSS(VSS),.VDD(VDD),.Y(g6695),.A(I12016),.B(I12017));
  NAND2 NAND2_697(.VSS(VSS),.VDD(VDD),.Y(I12031),.A(g5918),.B(g5897));
  NAND2 NAND2_698(.VSS(VSS),.VDD(VDD),.Y(I12032),.A(g5918),.B(I12031));
  NAND2 NAND2_699(.VSS(VSS),.VDD(VDD),.Y(I12033),.A(g5897),.B(I12031));
  NAND2 NAND2_700(.VSS(VSS),.VDD(VDD),.Y(g6701),.A(I12032),.B(I12033));
  NAND2 NAND2_701(.VSS(VSS),.VDD(VDD),.Y(I12051),.A(g5956),.B(g5939));
  NAND2 NAND2_702(.VSS(VSS),.VDD(VDD),.Y(I12052),.A(g5956),.B(I12051));
  NAND2 NAND2_703(.VSS(VSS),.VDD(VDD),.Y(I12053),.A(g5939),.B(I12051));
  NAND2 NAND2_704(.VSS(VSS),.VDD(VDD),.Y(g6709),.A(I12052),.B(I12053));
  NAND2 NAND2_705(.VSS(VSS),.VDD(VDD),.Y(I12078),.A(g5988),.B(g5971));
  NAND2 NAND2_706(.VSS(VSS),.VDD(VDD),.Y(I12079),.A(g5988),.B(I12078));
  NAND2 NAND2_707(.VSS(VSS),.VDD(VDD),.Y(I12080),.A(g5971),.B(I12078));
  NAND2 NAND2_708(.VSS(VSS),.VDD(VDD),.Y(g6722),.A(I12079),.B(I12080));
  NAND2 NAND2_709(.VSS(VSS),.VDD(VDD),.Y(I12179),.A(g1961),.B(g6163));
  NAND2 NAND2_710(.VSS(VSS),.VDD(VDD),.Y(I12180),.A(g1961),.B(I12179));
  NAND2 NAND2_711(.VSS(VSS),.VDD(VDD),.Y(I12181),.A(g6163),.B(I12179));
  NAND2 NAND2_712(.VSS(VSS),.VDD(VDD),.Y(g6770),.A(I12180),.B(I12181));
  NAND2 NAND2_713(.VSS(VSS),.VDD(VDD),.Y(I12550),.A(g6689),.B(g1462));
  NAND2 NAND2_714(.VSS(VSS),.VDD(VDD),.Y(I12551),.A(g6689),.B(I12550));
  NAND2 NAND2_715(.VSS(VSS),.VDD(VDD),.Y(I12552),.A(g1462),.B(I12550));
  NAND2 NAND2_716(.VSS(VSS),.VDD(VDD),.Y(g6893),.A(I12551),.B(I12552));
  NAND2 NAND2_717(.VSS(VSS),.VDD(VDD),.Y(I12575),.A(g6574),.B(g1049));
  NAND2 NAND2_718(.VSS(VSS),.VDD(VDD),.Y(I12576),.A(g6574),.B(I12575));
  NAND2 NAND2_719(.VSS(VSS),.VDD(VDD),.Y(I12577),.A(g1049),.B(I12575));
  NAND2 NAND2_720(.VSS(VSS),.VDD(VDD),.Y(g6902),.A(I12576),.B(I12577));
  NAND2 NAND2_721(.VSS(VSS),.VDD(VDD),.Y(I12596),.A(g6582),.B(g1126));
  NAND2 NAND2_722(.VSS(VSS),.VDD(VDD),.Y(I12597),.A(g6582),.B(I12596));
  NAND2 NAND2_723(.VSS(VSS),.VDD(VDD),.Y(I12598),.A(g1126),.B(I12596));
  NAND2 NAND2_724(.VSS(VSS),.VDD(VDD),.Y(g6911),.A(I12597),.B(I12598));
  NAND2 NAND2_725(.VSS(VSS),.VDD(VDD),.Y(I12832),.A(g6722),.B(g6709));
  NAND2 NAND2_726(.VSS(VSS),.VDD(VDD),.Y(I12833),.A(g6722),.B(I12832));
  NAND2 NAND2_727(.VSS(VSS),.VDD(VDD),.Y(I12834),.A(g6709),.B(I12832));
  NAND2 NAND2_728(.VSS(VSS),.VDD(VDD),.Y(g7065),.A(I12833),.B(I12834));
  NAND2 NAND2_729(.VSS(VSS),.VDD(VDD),.Y(g7069),.A(g5435),.B(g6680));
  NAND2 NAND2_730(.VSS(VSS),.VDD(VDD),.Y(I12852),.A(g6701),.B(g6695));
  NAND2 NAND2_731(.VSS(VSS),.VDD(VDD),.Y(I12853),.A(g6701),.B(I12852));
  NAND2 NAND2_732(.VSS(VSS),.VDD(VDD),.Y(I12854),.A(g6695),.B(I12852));
  NAND2 NAND2_733(.VSS(VSS),.VDD(VDD),.Y(g7082),.A(I12853),.B(I12854));
  NAND2 NAND2_734(.VSS(VSS),.VDD(VDD),.Y(I12869),.A(g2536),.B(g6618));
  NAND2 NAND2_735(.VSS(VSS),.VDD(VDD),.Y(I12870),.A(g2536),.B(I12869));
  NAND2 NAND2_736(.VSS(VSS),.VDD(VDD),.Y(I12871),.A(g6618),.B(I12869));
  NAND2 NAND2_737(.VSS(VSS),.VDD(VDD),.Y(g7093),.A(I12870),.B(I12871));
  NAND2 NAND2_738(.VSS(VSS),.VDD(VDD),.Y(I12951),.A(g7003),.B(g1467));
  NAND2 NAND2_739(.VSS(VSS),.VDD(VDD),.Y(I12952),.A(g7003),.B(I12951));
  NAND2 NAND2_740(.VSS(VSS),.VDD(VDD),.Y(I12953),.A(g1467),.B(I12951));
  NAND2 NAND2_741(.VSS(VSS),.VDD(VDD),.Y(g7121),.A(I12952),.B(I12953));
  NAND2 NAND2_742(.VSS(VSS),.VDD(VDD),.Y(I13002),.A(g7010),.B(g1053));
  NAND2 NAND2_743(.VSS(VSS),.VDD(VDD),.Y(I13003),.A(g7010),.B(I13002));
  NAND2 NAND2_744(.VSS(VSS),.VDD(VDD),.Y(I13004),.A(g1053),.B(I13002));
  NAND2 NAND2_745(.VSS(VSS),.VDD(VDD),.Y(g7140),.A(I13003),.B(I13004));
  NAND2 NAND2_746(.VSS(VSS),.VDD(VDD),.Y(I13016),.A(g6941),.B(g1142));
  NAND2 NAND2_747(.VSS(VSS),.VDD(VDD),.Y(I13017),.A(g6941),.B(I13016));
  NAND2 NAND2_748(.VSS(VSS),.VDD(VDD),.Y(I13018),.A(g1142),.B(I13016));
  NAND2 NAND2_749(.VSS(VSS),.VDD(VDD),.Y(g7144),.A(I13017),.B(I13018));
  NAND4 NAND4_3(.VSS(VSS),.VDD(VDD),.Y(g7234),.A(g3757),.B(g3739),.C(g7050),.D(g3770));
  NAND2 NAND2_750(.VSS(VSS),.VDD(VDD),.Y(g7237),.A(g7050),.B(g3739));
  NAND3 NAND3_13(.VSS(VSS),.VDD(VDD),.Y(g7244),.A(g7050),.B(g3757),.C(g3739));
  NAND2 NAND2_751(.VSS(VSS),.VDD(VDD),.Y(I13213),.A(g7065),.B(g7082));
  NAND2 NAND2_752(.VSS(VSS),.VDD(VDD),.Y(I13214),.A(g7065),.B(I13213));
  NAND2 NAND2_753(.VSS(VSS),.VDD(VDD),.Y(I13215),.A(g7082),.B(I13213));
  NAND2 NAND2_754(.VSS(VSS),.VDD(VDD),.Y(g7257),.A(I13214),.B(I13215));
  NAND2 NAND2_755(.VSS(VSS),.VDD(VDD),.Y(I13376),.A(g7199),.B(g1472));
  NAND2 NAND2_756(.VSS(VSS),.VDD(VDD),.Y(I13377),.A(g7199),.B(I13376));
  NAND2 NAND2_757(.VSS(VSS),.VDD(VDD),.Y(I13378),.A(g1472),.B(I13376));
  NAND2 NAND2_758(.VSS(VSS),.VDD(VDD),.Y(g7316),.A(I13377),.B(I13378));
  NAND2 NAND2_759(.VSS(VSS),.VDD(VDD),.Y(I13395),.A(g7212),.B(g1057));
  NAND2 NAND2_760(.VSS(VSS),.VDD(VDD),.Y(I13396),.A(g7212),.B(I13395));
  NAND2 NAND2_761(.VSS(VSS),.VDD(VDD),.Y(I13397),.A(g1057),.B(I13395));
  NAND2 NAND2_762(.VSS(VSS),.VDD(VDD),.Y(g7325),.A(I13396),.B(I13397));
  NAND2 NAND2_763(.VSS(VSS),.VDD(VDD),.Y(I13587),.A(g2556),.B(g7234));
  NAND2 NAND2_764(.VSS(VSS),.VDD(VDD),.Y(I13588),.A(g2556),.B(I13587));
  NAND2 NAND2_765(.VSS(VSS),.VDD(VDD),.Y(I13589),.A(g7234),.B(I13587));
  NAND2 NAND2_766(.VSS(VSS),.VDD(VDD),.Y(g7444),.A(I13588),.B(I13589));
  NAND2 NAND2_767(.VSS(VSS),.VDD(VDD),.Y(I13598),.A(g2551),.B(g7244));
  NAND2 NAND2_768(.VSS(VSS),.VDD(VDD),.Y(I13599),.A(g2551),.B(I13598));
  NAND2 NAND2_769(.VSS(VSS),.VDD(VDD),.Y(I13600),.A(g7244),.B(I13598));
  NAND2 NAND2_770(.VSS(VSS),.VDD(VDD),.Y(g7447),.A(I13599),.B(I13600));
  NAND2 NAND2_771(.VSS(VSS),.VDD(VDD),.Y(I13638),.A(g7257),.B(g7069));
  NAND2 NAND2_772(.VSS(VSS),.VDD(VDD),.Y(I13639),.A(g7257),.B(I13638));
  NAND2 NAND2_773(.VSS(VSS),.VDD(VDD),.Y(I13640),.A(g7069),.B(I13638));
  NAND2 NAND2_774(.VSS(VSS),.VDD(VDD),.Y(g7480),.A(I13639),.B(I13640));
  NAND2 NAND2_775(.VSS(VSS),.VDD(VDD),.Y(I13685),.A(g1977),.B(g7237));
  NAND2 NAND2_776(.VSS(VSS),.VDD(VDD),.Y(I13686),.A(g1977),.B(I13685));
  NAND2 NAND2_777(.VSS(VSS),.VDD(VDD),.Y(I13687),.A(g7237),.B(I13685));
  NAND2 NAND2_778(.VSS(VSS),.VDD(VDD),.Y(g7503),.A(I13686),.B(I13687));
  NAND2 NAND2_779(.VSS(VSS),.VDD(VDD),.Y(I13785),.A(g7427),.B(g1477));
  NAND2 NAND2_780(.VSS(VSS),.VDD(VDD),.Y(I13786),.A(g7427),.B(I13785));
  NAND2 NAND2_781(.VSS(VSS),.VDD(VDD),.Y(I13787),.A(g1477),.B(I13785));
  NAND2 NAND2_782(.VSS(VSS),.VDD(VDD),.Y(g7535),.A(I13786),.B(I13787));
  NAND2 NAND2_783(.VSS(VSS),.VDD(VDD),.Y(I13800),.A(g7429),.B(g1061));
  NAND2 NAND2_784(.VSS(VSS),.VDD(VDD),.Y(I13801),.A(g7429),.B(I13800));
  NAND2 NAND2_785(.VSS(VSS),.VDD(VDD),.Y(I13802),.A(g1061),.B(I13800));
  NAND2 NAND2_786(.VSS(VSS),.VDD(VDD),.Y(g7540),.A(I13801),.B(I13802));
  NAND2 NAND2_787(.VSS(VSS),.VDD(VDD),.Y(I14244),.A(g7683),.B(g1065));
  NAND2 NAND2_788(.VSS(VSS),.VDD(VDD),.Y(I14245),.A(g7683),.B(I14244));
  NAND2 NAND2_789(.VSS(VSS),.VDD(VDD),.Y(I14246),.A(g1065),.B(I14244));
  NAND2 NAND2_790(.VSS(VSS),.VDD(VDD),.Y(g7828),.A(I14245),.B(I14246));
  NAND2 NAND2_791(.VSS(VSS),.VDD(VDD),.Y(I14472),.A(g8147),.B(g1069));
  NAND2 NAND2_792(.VSS(VSS),.VDD(VDD),.Y(I14473),.A(g8147),.B(I14472));
  NAND2 NAND2_793(.VSS(VSS),.VDD(VDD),.Y(I14474),.A(g1069),.B(I14472));
  NAND2 NAND2_794(.VSS(VSS),.VDD(VDD),.Y(g8231),.A(I14473),.B(I14474));
  NAND2 NAND2_795(.VSS(VSS),.VDD(VDD),.Y(g8239),.A(g8073),.B(g8092));
  NAND2 NAND2_796(.VSS(VSS),.VDD(VDD),.Y(g8627),.A(g6232),.B(g8091));
  NAND2 NAND2_797(.VSS(VSS),.VDD(VDD),.Y(g8633),.A(g8176),.B(g6232));
  NAND2 NAND2_798(.VSS(VSS),.VDD(VDD),.Y(I14837),.A(g8660),.B(g1073));
  NAND2 NAND2_799(.VSS(VSS),.VDD(VDD),.Y(I14838),.A(g8660),.B(I14837));
  NAND2 NAND2_800(.VSS(VSS),.VDD(VDD),.Y(I14839),.A(g1073),.B(I14837));
  NAND2 NAND2_801(.VSS(VSS),.VDD(VDD),.Y(g8681),.A(I14838),.B(I14839));
  NAND2 NAND2_802(.VSS(VSS),.VDD(VDD),.Y(g8798),.A(g6984),.B(g8644));
  NAND2 NAND2_803(.VSS(VSS),.VDD(VDD),.Y(I15817),.A(g9151),.B(g9148));
  NAND2 NAND2_804(.VSS(VSS),.VDD(VDD),.Y(I15818),.A(g9151),.B(I15817));
  NAND2 NAND2_805(.VSS(VSS),.VDD(VDD),.Y(I15819),.A(g9148),.B(I15817));
  NAND2 NAND2_806(.VSS(VSS),.VDD(VDD),.Y(g9179),.A(I15818),.B(I15819));
  NAND2 NAND2_807(.VSS(VSS),.VDD(VDD),.Y(I15848),.A(g9162),.B(g9154));
  NAND2 NAND2_808(.VSS(VSS),.VDD(VDD),.Y(I15849),.A(g9162),.B(I15848));
  NAND2 NAND2_809(.VSS(VSS),.VDD(VDD),.Y(I15850),.A(g9154),.B(I15848));
  NAND2 NAND2_810(.VSS(VSS),.VDD(VDD),.Y(g9190),.A(I15849),.B(I15850));
  NAND2 NAND2_811(.VSS(VSS),.VDD(VDD),.Y(I15855),.A(g9168),.B(g9165));
  NAND2 NAND2_812(.VSS(VSS),.VDD(VDD),.Y(I15856),.A(g9168),.B(I15855));
  NAND2 NAND2_813(.VSS(VSS),.VDD(VDD),.Y(I15857),.A(g9165),.B(I15855));
  NAND2 NAND2_814(.VSS(VSS),.VDD(VDD),.Y(g9191),.A(I15856),.B(I15857));
  NAND2 NAND2_815(.VSS(VSS),.VDD(VDD),.Y(I15862),.A(g9174),.B(g9171));
  NAND2 NAND2_816(.VSS(VSS),.VDD(VDD),.Y(I15863),.A(g9174),.B(I15862));
  NAND2 NAND2_817(.VSS(VSS),.VDD(VDD),.Y(I15864),.A(g9171),.B(I15862));
  NAND2 NAND2_818(.VSS(VSS),.VDD(VDD),.Y(g9192),.A(I15863),.B(I15864));
  NAND2 NAND2_819(.VSS(VSS),.VDD(VDD),.Y(I15880),.A(g9190),.B(g9179));
  NAND2 NAND2_820(.VSS(VSS),.VDD(VDD),.Y(I15881),.A(g9190),.B(I15880));
  NAND2 NAND2_821(.VSS(VSS),.VDD(VDD),.Y(I15882),.A(g9179),.B(I15880));
  NAND2 NAND2_822(.VSS(VSS),.VDD(VDD),.Y(g9202),.A(I15881),.B(I15882));
  NAND2 NAND2_823(.VSS(VSS),.VDD(VDD),.Y(I15887),.A(g9192),.B(g9191));
  NAND2 NAND2_824(.VSS(VSS),.VDD(VDD),.Y(I15888),.A(g9192),.B(I15887));
  NAND2 NAND2_825(.VSS(VSS),.VDD(VDD),.Y(I15889),.A(g9191),.B(I15887));
  NAND2 NAND2_826(.VSS(VSS),.VDD(VDD),.Y(g9203),.A(I15888),.B(I15889));
  NAND2 NAND2_827(.VSS(VSS),.VDD(VDD),.Y(I15897),.A(g9202),.B(g9203));
  NAND2 NAND2_828(.VSS(VSS),.VDD(VDD),.Y(I15898),.A(g9202),.B(I15897));
  NAND2 NAND2_829(.VSS(VSS),.VDD(VDD),.Y(I15899),.A(g9203),.B(I15897));
  NAND2 NAND2_830(.VSS(VSS),.VDD(VDD),.Y(g9205),.A(I15898),.B(I15899));
//
  NOR2 NOR2_0(.VSS(VSS),.VDD(VDD),.Y(g1964),.A(g1428),.B(g1429));
  NOR2 NOR2_1(.VSS(VSS),.VDD(VDD),.Y(g1980),.A(g1430),.B(g1431));
  NOR2 NOR2_2(.VSS(VSS),.VDD(VDD),.Y(g2014),.A(g1421),.B(g1416));
  NOR2 NOR2_3(.VSS(VSS),.VDD(VDD),.Y(g2521),.A(g65),.B(g62));
  NOR3 NOR3_0(.VSS(VSS),.VDD(VDD),.Y(g3225),.A(g1021),.B(g1025),.C(g1889));
  NOR2 NOR2_4(.VSS(VSS),.VDD(VDD),.Y(g3233),.A(g1714),.B(g1459));
  NOR3 NOR3_1(.VSS(VSS),.VDD(VDD),.Y(g3237),.A(g1444),.B(g1838),.C(g1454));
  NOR2 NOR2_5(.VSS(VSS),.VDD(VDD),.Y(g3260),.A(g1728),.B(g2490));
  NOR2 NOR2_6(.VSS(VSS),.VDD(VDD),.Y(g3310),.A(g936),.B(g2557));
  NOR4 NOR4_0(.VSS(VSS),.VDD(VDD),.Y(g3504),.A(g1375),.B(g2229),.C(g2213),.D(g2206));
  NOR2 NOR2_7(.VSS(VSS),.VDD(VDD),.Y(g3505),.A(g2263),.B(g1395));
  NOR4 NOR4_1(.VSS(VSS),.VDD(VDD),.Y(g3515),.A(g1388),.B(g2262),.C(g2230),.D(g2214));
  NOR2 NOR2_8(.VSS(VSS),.VDD(VDD),.Y(g3516),.A(g2282),.B(g1401));
  NOR2 NOR2_9(.VSS(VSS),.VDD(VDD),.Y(g3528),.A(g2343),.B(g1391));
  NOR2 NOR2_10(.VSS(VSS),.VDD(VDD),.Y(g3555),.A(g2359),.B(g1398));
  NOR3 NOR3_2(.VSS(VSS),.VDD(VDD),.Y(g3790),.A(g985),.B(g990),.C(g2295));
  NOR2 NOR2_11(.VSS(VSS),.VDD(VDD),.Y(g3885),.A(g3310),.B(g3466));
  NOR2 NOR2_12(.VSS(VSS),.VDD(VDD),.Y(g4160),.A(g1231),.B(g2834));
  NOR2 NOR2_13(.VSS(VSS),.VDD(VDD),.Y(g4232),.A(g1934),.B(g3591));
  NOR2 NOR2_14(.VSS(VSS),.VDD(VDD),.Y(g4318),.A(g3681),.B(g1590));
  NOR2 NOR2_15(.VSS(VSS),.VDD(VDD),.Y(g4349),.A(g2496),.B(g3310));
  NOR2 NOR2_16(.VSS(VSS),.VDD(VDD),.Y(g4354),.A(g1424),.B(g3541));
  NOR2 NOR2_17(.VSS(VSS),.VDD(VDD),.Y(g4676),.A(g3885),.B(g3094));
  NOR4 NOR4_2(.VSS(VSS),.VDD(VDD),.Y(g4884),.A(g4492),.B(g4476),.C(g4456),.D(g4294));
  NOR4 NOR4_3(.VSS(VSS),.VDD(VDD),.Y(g4888),.A(g4548),.B(g4528),.C(g4513),.D(g4502));
  NOR3 NOR3_3(.VSS(VSS),.VDD(VDD),.Y(g4894),.A(g4298),.B(g4575),.C(g4563));
  NOR4 NOR4_4(.VSS(VSS),.VDD(VDD),.Y(g5023),.A(g3894),.B(g3889),.C(g3886),.D(g4359));
  NOR4 NOR4_5(.VSS(VSS),.VDD(VDD),.Y(g5039),.A(g3924),.B(g3914),.C(g3906),.D(g3899));
  NOR3 NOR3_4(.VSS(VSS),.VDD(VDD),.Y(g5056),.A(g3556),.B(g2872),.C(g3938));
  NOR3 NOR3_5(.VSS(VSS),.VDD(VDD),.Y(g5614),.A(g3002),.B(g1590),.C(g4714));
  NOR2 NOR2_18(.VSS(VSS),.VDD(VDD),.Y(g5615),.A(g4714),.B(g3002));
  NOR2 NOR2_19(.VSS(VSS),.VDD(VDD),.Y(g5772),.A(g5428),.B(g1888));
  NOR2 NOR2_20(.VSS(VSS),.VDD(VDD),.Y(g6174),.A(g1855),.B(g5305));
  NOR2 NOR2_21(.VSS(VSS),.VDD(VDD),.Y(g6184),.A(g875),.B(g5291));
  NOR2 NOR2_22(.VSS(VSS),.VDD(VDD),.Y(g6185),.A(g5305),.B(g1590));
  NOR2 NOR2_23(.VSS(VSS),.VDD(VDD),.Y(g6193),.A(g1926),.B(g5310));
  NOR4 NOR4_6(.VSS(VSS),.VDD(VDD),.Y(g6197),.A(g875),.B(g866),.C(g1590),.D(g5291));
  NOR2 NOR2_24(.VSS(VSS),.VDD(VDD),.Y(g6209),.A(g2332),.B(g5305));
  NOR2 NOR2_25(.VSS(VSS),.VDD(VDD),.Y(g6214),.A(g878),.B(g5284));
  NOR2 NOR2_26(.VSS(VSS),.VDD(VDD),.Y(g6259),.A(g3002),.B(g5312));
  NOR2 NOR2_27(.VSS(VSS),.VDD(VDD),.Y(g6452),.A(g6270),.B(g2245));
  NOR4 NOR4_7(.VSS(VSS),.VDD(VDD),.Y(g6465),.A(g5403),.B(g5802),.C(g5769),.D(g5790));
  NOR3 NOR3_6(.VSS(VSS),.VDD(VDD),.Y(g6489),.A(g5802),.B(g5769),.C(g5790));
  NOR3 NOR3_7(.VSS(VSS),.VDD(VDD),.Y(g6664),.A(g5836),.B(g1901),.C(g1788));
  NOR4 NOR4_8(.VSS(VSS),.VDD(VDD),.Y(g6910),.A(g1011),.B(g1837),.C(g6559),.D(g1008));
  NOR3 NOR3_8(.VSS(VSS),.VDD(VDD),.Y(g7152),.A(g6253),.B(g7083),.C(g5418));
  NOR3 NOR3_9(.VSS(VSS),.VDD(VDD),.Y(g7209),.A(g1789),.B(g146),.C(g6984));
  NOR2 NOR2_28(.VSS(VSS),.VDD(VDD),.Y(g7312),.A(g7178),.B(g6970));
  NOR2 NOR2_29(.VSS(VSS),.VDD(VDD),.Y(g7314),.A(g7180),.B(g6972));
  NOR2 NOR2_30(.VSS(VSS),.VDD(VDD),.Y(g7318),.A(g7185),.B(g6979));
  NOR2 NOR2_31(.VSS(VSS),.VDD(VDD),.Y(g7321),.A(g7187),.B(g6990));
  NOR2 NOR2_32(.VSS(VSS),.VDD(VDD),.Y(g7322),.A(g7188),.B(g6991));
  NOR2 NOR2_33(.VSS(VSS),.VDD(VDD),.Y(g7324),.A(g7189),.B(g6994));
  NOR2 NOR2_34(.VSS(VSS),.VDD(VDD),.Y(g7326),.A(g7194),.B(g6999));
  NOR2 NOR2_35(.VSS(VSS),.VDD(VDD),.Y(g7328),.A(g7196),.B(g7001));
  NOR2 NOR2_36(.VSS(VSS),.VDD(VDD),.Y(g7406),.A(g7191),.B(g1600));
  NOR2 NOR2_37(.VSS(VSS),.VDD(VDD),.Y(g7566),.A(g7421),.B(g1597));
  NOR2 NOR2_38(.VSS(VSS),.VDD(VDD),.Y(g8073),.A(g7658),.B(g7654));
  NOR4 NOR4_9(.VSS(VSS),.VDD(VDD),.Y(g8092),.A(g7634),.B(g7628),.C(g7616),.D(g7611));
  NOR3 NOR3_10(.VSS(VSS),.VDD(VDD),.Y(g8230),.A(g8199),.B(I14467),.C(I14468));
  NOR3 NOR3_11(.VSS(VSS),.VDD(VDD),.Y(g8232),.A(g8199),.B(I14479),.C(I14480));
  NOR3 NOR3_12(.VSS(VSS),.VDD(VDD),.Y(g8233),.A(g8199),.B(I14484),.C(I14485));
  NOR3 NOR3_13(.VSS(VSS),.VDD(VDD),.Y(g8236),.A(g8199),.B(I14495),.C(I14496));
  NOR4 NOR4_10(.VSS(VSS),.VDD(VDD),.Y(g8279),.A(g7658),.B(g7616),.C(g8082),.D(g7634));
  NOR4 NOR4_11(.VSS(VSS),.VDD(VDD),.Y(g8360),.A(g7658),.B(g7616),.C(g8082),.D(g7634));
  NOR4 NOR4_12(.VSS(VSS),.VDD(VDD),.Y(g8523),.A(g7658),.B(g7616),.C(g8082),.D(g7634));
  NOR4 NOR4_13(.VSS(VSS),.VDD(VDD),.Y(g8625),.A(g1000),.B(g6573),.C(g1860),.D(g8009));
  NOR2 NOR2_39(.VSS(VSS),.VDD(VDD),.Y(g8629),.A(g6270),.B(g8009));
  NOR4 NOR4_14(.VSS(VSS),.VDD(VDD),.Y(g8630),.A(g6110),.B(g7784),.C(g3591),.D(g1864));
  NOR2 NOR2_40(.VSS(VSS),.VDD(VDD),.Y(g8635),.A(g1034),.B(g8128));
  NOR4 NOR4_15(.VSS(VSS),.VDD(VDD),.Y(g8641),.A(g6559),.B(g162),.C(g7784),.D(g3591));
  NOR2 NOR2_41(.VSS(VSS),.VDD(VDD),.Y(g8644),.A(g4146),.B(g8128));
  NOR3 NOR3_14(.VSS(VSS),.VDD(VDD),.Y(g8655),.A(g8199),.B(I14753),.C(I14754));
  NOR3 NOR3_15(.VSS(VSS),.VDD(VDD),.Y(g8656),.A(g8199),.B(I14758),.C(I14759));
  NOR3 NOR3_16(.VSS(VSS),.VDD(VDD),.Y(g8658),.A(g8199),.B(I14766),.C(I14767));
  NOR3 NOR3_17(.VSS(VSS),.VDD(VDD),.Y(g8659),.A(g8199),.B(I14771),.C(I14772));
  NOR3 NOR3_18(.VSS(VSS),.VDD(VDD),.Y(g8679),.A(g8493),.B(g8239),.C(I14831));
  NOR3 NOR3_19(.VSS(VSS),.VDD(VDD),.Y(g8680),.A(g8493),.B(g8239),.C(I14834));
  NOR3 NOR3_20(.VSS(VSS),.VDD(VDD),.Y(g8694),.A(g7658),.B(g8613),.C(g7634));
  NOR3 NOR3_21(.VSS(VSS),.VDD(VDD),.Y(g8699),.A(g7658),.B(g8613),.C(g7634));
  NOR3 NOR3_22(.VSS(VSS),.VDD(VDD),.Y(g8706),.A(g7658),.B(g8613),.C(g7634));
  NOR3 NOR3_23(.VSS(VSS),.VDD(VDD),.Y(g8707),.A(g7658),.B(g8613),.C(g7634));
  NOR2 NOR2_42(.VSS(VSS),.VDD(VDD),.Y(g8801),.A(g8635),.B(g3790));
  NOR3 NOR3_24(.VSS(VSS),.VDD(VDD),.Y(g8803),.A(g8443),.B(g8421),.C(I15021));
  NOR3 NOR3_25(.VSS(VSS),.VDD(VDD),.Y(g8805),.A(g8443),.B(g8421),.C(I15033));
  NOR3 NOR3_26(.VSS(VSS),.VDD(VDD),.Y(g8806),.A(g8443),.B(g8421),.C(I15044));
  NOR3 NOR3_27(.VSS(VSS),.VDD(VDD),.Y(g8807),.A(g8443),.B(g8421),.C(I15055));
  NOR3 NOR3_28(.VSS(VSS),.VDD(VDD),.Y(g8811),.A(g8443),.B(g8421),.C(I15075));
  NOR3 NOR3_29(.VSS(VSS),.VDD(VDD),.Y(g8812),.A(g8443),.B(g8421),.C(I15086));
  NOR3 NOR3_30(.VSS(VSS),.VDD(VDD),.Y(g8818),.A(g8443),.B(g8421),.C(I15102));
  NOR3 NOR3_31(.VSS(VSS),.VDD(VDD),.Y(g8819),.A(g8443),.B(g8421),.C(I15113));
  NOR3 NOR3_32(.VSS(VSS),.VDD(VDD),.Y(g8847),.A(g8493),.B(g8239),.C(I15147));
  NOR3 NOR3_33(.VSS(VSS),.VDD(VDD),.Y(g8850),.A(g8493),.B(g8239),.C(I15152));
  NOR3 NOR3_34(.VSS(VSS),.VDD(VDD),.Y(g8855),.A(g7658),.B(g8613),.C(g7634));
  NOR3 NOR3_35(.VSS(VSS),.VDD(VDD),.Y(g8859),.A(g8493),.B(g8239),.C(I15165));
  NOR3 NOR3_36(.VSS(VSS),.VDD(VDD),.Y(g8861),.A(g8493),.B(g8239),.C(I15169));
  NOR3 NOR3_37(.VSS(VSS),.VDD(VDD),.Y(g8862),.A(g8493),.B(g8239),.C(I15172));
  NOR3 NOR3_38(.VSS(VSS),.VDD(VDD),.Y(g8863),.A(g8493),.B(g8239),.C(I15175));

endmodule