module s1423(G727,G701BF,G1,G12,VDD,G7,G0,G2,G14,G16,G13,G4,G6,G5,G3,G11,VSS,G9,G702,CLOCK,G8,G10,G729,G726,G15);
input G7,G14,G13,G5,G3,G11,G1,G12,VDD,G0,G2,G16,G4,G6,VSS,G9,CLOCK,G8,G10,G15;
output G727,G701BF,G702,G729,G726;

  wire G273,G196,G521,G339,G435,G472,G681,G618,G419,G26,G571,G518,G36,G528,G470,G61,G59,G728,G696,G350,G403,G288,G53,G582,G81,G139,G587,G35,G359,G188,G466,G33,G68,G490,G512,G625,G272,G498,G74,G317,G217,G585,G79,G392,G355,G656,G255,G484,G211,G637,G212,G164,G439,G161,G93,G46,G357,G70,G687,G516,G242,G325,I1239,G209,G459,G662,G666,G534,G75,G230,G704,G136,G257,G613,G321,G433,G369,G292,G601,G638,G375,G502,G604,G483,G343,G685,G464,G153,G443,G383,G334,G680,G38,G203,G537,G602,G360,G144,G655,I1,G201,G300,G51,G554,G23,G531,G235,G660,G588,G446,G27,G30,G135,G227,G251,G290,G346,G143,G605,I1245,G387,G441,G452,G128,G49,G244,G52,G269,G547,G178,G428,G563,G326,G494,G386,G208,G123,G394,G241,G57,G333,G458,G550,G539,G510,G154,G460,G598,G90,G39,G640,G214,G191,G545,G595,G294,G373,G659,G578,G644,G440,G491,G306,G649,G195,G486,G482,G331,G377,G425,G710,G259,G708,G92,G171,G220,G83,G603,G551,G236,G505,G89,G673,G467,G129,G388,G457,G268,G519,G311,G40,G718,G612,G586,G462,G199,G32,G529,G579,G310,G575,G165,G329,G583,G137,G302,G378,G705,G270,G677,G473,G608,G180,G499,G474,G485,G181,G297,G100,G356,I1242,G189,G522,I1248,G351,G145,G651,G569,G338,G500,G157,G332,G316,G309,G322,G151,G192,G335,G232,G650,G286,G559,G216,G418,G667,G399,G506,G318,G215,G580,G630,G152,G487,G596,I1227,G308,G376,I1254,I12,G400,G690,G86,G616,G589,G535,G285,G671,I1211,G722,G719,G501,G281,G219,G622,G693,G679,G225,G676,G562,G345,G543,G73,G102,G461,G43,G96,G576,G34,G237,G701,G252,G454,G374,G97,G669,G194,G670,G233,G525,G489,G156,G328BF,G675,G71,G80,G621,G234,G540,G385,G712,G725,G226,G398,G25,G434,G438,G530,G160,G469,G28,G368,G303,G22,G714,G132,G337,G475,G246,G456,G639,G654,G643,G645,G568,G238,G396,G64,G672,G221,G240,G636,G94,G223,G478,G204,G495,G361,G414,G707,G341,G41,G130,G250,G106,I1236,G218,G72,G691,G275,G342,G397,G641,G116,G389,G371,G450,G653,G29,G60,G520,G85,G210,G37,G65,G283,G682,G312,G515,G436,G590,G497,G393,G688,G173,G706,G686,G182,I1203,G426,G176,G597,G54,G88,G508,G362,G111,G614,G406,G332BF,G126,G249,G107,G694,G647,G276,G62,I1251,G553,G683,G271,G158,G390,G567,I1162,G131,G42,G635,G542,G253,G193,G496,G305,G455,G168,G149,G48,G713,G364,G202,G507,G536,G247,G323,G700,G314,G365,G698,G668,G379,G183,G231,G422,G284,G134,G417,G122,G488,G492,G476,G544,G63,G504,G648,G584,G558,G620,G717,G611,G610,G256,G174,G517,G55,G289,G291,G121,G261,G118,G652,G104,G146,G444,G565,G77,G363,G190,G409,G293,G348,G437,G447,G523,G327,G430,G665,G105,G155,G99,G480,G532,G716,G367,G723,G243,G481,G84,G463,G56,G548,G296,G570,G91,G101,G634,G572,G429,G280,G527,G549,G31,G724,G533,G657,G561,G479,G684,G315,G254,G721,G623,G405,G114,G119,G112,G298,G560,G87,G526,G213,G606,G328,G172,G646,G224,G222,G658,G624,G103,G349,G574,G633,G395,G465,G313,G167,G207,G248,G82,G513,G200,G142,I1267,G664,G69,G628,G427,G503,G299,G266,G380,G415,I1260,G262,G471,G556,G493,G170,G477,G692,G423,G370,G169,G468,G179,I1264,G353,G115,G133,G206,G120,G245,G432,G150,G267,G344,G524,I1257,G198,G514,G239,G184,G141,G47,G277,G295,G78,G411,G410,G674,G175,G304,I1230,G594,G631,G445,G564,G420,G566,G600,I1183,G264,G347,G449,I1233,G109,G66,G324,G453,G148,G615,G689,G599,G147,G187,G162,G229,G58,G711,G609,G709,G401,G592,G408,G108,G442,G205,G24,G541,G546,G320,G509,G307,G45,G354,G197,G424,G260,G358,G697,G703,G278,G416,G159,G407,G413,G274,G661,G330,G319,G287,G228,G127,G577,G699,G301,G138,G166,G352,G715,G366,G617,G185,G448,G113,G431,G50,G67,G279,G265,G372,G76,G382,G340,G95,G412,G511,G451,G384,G626,G642,G591,G163,G619,G629,G552,G695,G573,G557,G186,G124,G282,G44,G140,G381,G663,G110,G720,G607,G678,G538,G263,G593,G177,G125,G98,G391,G555,G581,G627,G404,G117,G258,G632,G402,G421,G336;
//# 17 inputs
//# 5 outputs
//# 74 D-type flipflops
//# 167 inverters
//# 490 gates (197 ANDs + 64 NANDs + 137 ORs + 92 NORs)
//
//
//
  MSFF DFF_0(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G22),.DATA(G332BF));
  MSFF DFF_1(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G23),.DATA(G328BF));
  MSFF DFF_2(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G24),.DATA(G109));
  MSFF DFF_3(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G25),.DATA(G113));
  MSFF DFF_4(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G26),.DATA(G118));
  MSFF DFF_5(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G27),.DATA(G125));
  MSFF DFF_6(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G28),.DATA(G129));
  MSFF DFF_7(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G29),.DATA(G140));
  MSFF DFF_8(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G30),.DATA(G144));
  MSFF DFF_9(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G31),.DATA(G149));
  MSFF DFF_10(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G32),.DATA(G154));
  MSFF DFF_11(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G33),.DATA(G159));
  MSFF DFF_12(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G34),.DATA(G166));
  MSFF DFF_13(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G35),.DATA(G175));
  MSFF DFF_14(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G36),.DATA(G189));
  MSFF DFF_15(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G37),.DATA(G193));
  MSFF DFF_16(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G38),.DATA(G198));
  MSFF DFF_17(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G39),.DATA(G208));
  MSFF DFF_18(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G40),.DATA(G214));
  MSFF DFF_19(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G41),.DATA(G218));
  MSFF DFF_20(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G42),.DATA(G237));
  MSFF DFF_21(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G43),.DATA(G242));
  MSFF DFF_22(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G44),.DATA(G247));
  MSFF DFF_23(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G45),.DATA(G252));
  MSFF DFF_24(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G46),.DATA(G260));
  MSFF DFF_25(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G47),.DATA(G303));
  MSFF DFF_26(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G48),.DATA(G309));
  MSFF DFF_27(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G49),.DATA(G315));
  MSFF DFF_28(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G50),.DATA(G321));
  MSFF DFF_29(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G51),.DATA(G360));
  MSFF DFF_30(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G52),.DATA(G365));
  MSFF DFF_31(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G53),.DATA(G373));
  MSFF DFF_32(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G54),.DATA(G379));
  MSFF DFF_33(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G55),.DATA(G384));
  MSFF DFF_34(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G56),.DATA(G392));
  MSFF DFF_35(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G57),.DATA(G397));
  MSFF DFF_36(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G58),.DATA(G405));
  MSFF DFF_37(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G59),.DATA(G408));
  MSFF DFF_38(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G60),.DATA(G416));
  MSFF DFF_39(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G61),.DATA(G424));
  MSFF DFF_40(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G62),.DATA(G427));
  MSFF DFF_41(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G63),.DATA(G438));
  MSFF DFF_42(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G64),.DATA(G441));
  MSFF DFF_43(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G65),.DATA(G447));
  MSFF DFF_44(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G66),.DATA(G451));
  MSFF DFF_45(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G67),.DATA(G459));
  MSFF DFF_46(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G68),.DATA(G464));
  MSFF DFF_47(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G69),.DATA(G469));
  MSFF DFF_48(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G70),.DATA(G477));
  MSFF DFF_49(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G71),.DATA(G494));
  MSFF DFF_50(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G72),.DATA(G498));
  MSFF DFF_51(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G73),.DATA(G503));
  MSFF DFF_52(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G74),.DATA(G526));
  MSFF DFF_53(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G75),.DATA(G531));
  MSFF DFF_54(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G76),.DATA(G536));
  MSFF DFF_55(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G77),.DATA(G541));
  MSFF DFF_56(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G78),.DATA(G548));
  MSFF DFF_57(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G79),.DATA(G565));
  MSFF DFF_58(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G80),.DATA(G569));
  MSFF DFF_59(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G81),.DATA(G573));
  MSFF DFF_60(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G82),.DATA(G577));
  MSFF DFF_61(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G83),.DATA(G590));
  MSFF DFF_62(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G84),.DATA(G608));
  MSFF DFF_63(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G85),.DATA(G613));
  MSFF DFF_64(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G86),.DATA(G657));
  MSFF DFF_65(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G87),.DATA(G663));
  MSFF DFF_66(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G88),.DATA(G669));
  MSFF DFF_67(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G89),.DATA(G675));
  MSFF DFF_68(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G90),.DATA(G682));
  MSFF DFF_69(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G91),.DATA(G687));
  MSFF DFF_70(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G92),.DATA(G693));
  MSFF DFF_71(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G93),.DATA(G705));
  MSFF DFF_72(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G94),.DATA(G707));
  MSFF DFF_73(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G95),.DATA(G713));
//
  NOT NOT1_0(.VSS(VSS),.VDD(VDD),.Y(I1),.A(G332));
  NOT NOT1_1(.VSS(VSS),.VDD(VDD),.Y(G332BF),.A(I1));
  NOT NOT1_2(.VSS(VSS),.VDD(VDD),.Y(I12),.A(G328));
  NOT NOT1_3(.VSS(VSS),.VDD(VDD),.Y(G328BF),.A(I12));
  NOT NOT1_4(.VSS(VSS),.VDD(VDD),.Y(G108),.A(G712));
  NOT NOT1_5(.VSS(VSS),.VDD(VDD),.Y(G111),.A(G24));
  NOT NOT1_6(.VSS(VSS),.VDD(VDD),.Y(G112),.A(G712));
  NOT NOT1_7(.VSS(VSS),.VDD(VDD),.Y(G117),.A(G712));
  NOT NOT1_8(.VSS(VSS),.VDD(VDD),.Y(G124),.A(G712));
  NOT NOT1_9(.VSS(VSS),.VDD(VDD),.Y(G127),.A(G27));
  NOT NOT1_10(.VSS(VSS),.VDD(VDD),.Y(G128),.A(G712));
  NOT NOT1_11(.VSS(VSS),.VDD(VDD),.Y(G139),.A(G712));
  NOT NOT1_12(.VSS(VSS),.VDD(VDD),.Y(G142),.A(G29));
  NOT NOT1_13(.VSS(VSS),.VDD(VDD),.Y(G143),.A(G712));
  NOT NOT1_14(.VSS(VSS),.VDD(VDD),.Y(G148),.A(G712));
  NOT NOT1_15(.VSS(VSS),.VDD(VDD),.Y(G153),.A(G712));
  NOT NOT1_16(.VSS(VSS),.VDD(VDD),.Y(G158),.A(G712));
  NOT NOT1_17(.VSS(VSS),.VDD(VDD),.Y(G165),.A(G712));
  NOT NOT1_18(.VSS(VSS),.VDD(VDD),.Y(G174),.A(G712));
  NOT NOT1_19(.VSS(VSS),.VDD(VDD),.Y(G176),.A(G35));
  NOT NOT1_20(.VSS(VSS),.VDD(VDD),.Y(G178),.A(G34));
  NOT NOT1_21(.VSS(VSS),.VDD(VDD),.Y(G179),.A(G180));
  NOT NOT1_22(.VSS(VSS),.VDD(VDD),.Y(G180),.A(G92));
  NOT NOT1_23(.VSS(VSS),.VDD(VDD),.Y(G188),.A(G712));
  NOT NOT1_24(.VSS(VSS),.VDD(VDD),.Y(G191),.A(G36));
  NOT NOT1_25(.VSS(VSS),.VDD(VDD),.Y(G192),.A(G712));
  NOT NOT1_26(.VSS(VSS),.VDD(VDD),.Y(G197),.A(G712));
  NOT NOT1_27(.VSS(VSS),.VDD(VDD),.Y(G204),.A(G38));
  NOT NOT1_28(.VSS(VSS),.VDD(VDD),.Y(G207),.A(G712));
  NOT NOT1_29(.VSS(VSS),.VDD(VDD),.Y(G210),.A(G39));
  NOT NOT1_30(.VSS(VSS),.VDD(VDD),.Y(G213),.A(G712));
  NOT NOT1_31(.VSS(VSS),.VDD(VDD),.Y(G216),.A(G40));
  NOT NOT1_32(.VSS(VSS),.VDD(VDD),.Y(G217),.A(G712));
  NOT NOT1_33(.VSS(VSS),.VDD(VDD),.Y(G236),.A(G259));
  NOT NOT1_34(.VSS(VSS),.VDD(VDD),.Y(G241),.A(G259));
  NOT NOT1_35(.VSS(VSS),.VDD(VDD),.Y(G246),.A(G259));
  NOT NOT1_36(.VSS(VSS),.VDD(VDD),.Y(G251),.A(G259));
  NOT NOT1_37(.VSS(VSS),.VDD(VDD),.Y(G258),.A(G259));
  NOT NOT1_38(.VSS(VSS),.VDD(VDD),.Y(G296),.A(G297));
  NOT NOT1_39(.VSS(VSS),.VDD(VDD),.Y(G302),.A(G712));
  NOT NOT1_40(.VSS(VSS),.VDD(VDD),.Y(G305),.A(G324));
  NOT NOT1_41(.VSS(VSS),.VDD(VDD),.Y(G308),.A(G712));
  NOT NOT1_42(.VSS(VSS),.VDD(VDD),.Y(G311),.A(G324));
  NOT NOT1_43(.VSS(VSS),.VDD(VDD),.Y(G314),.A(G712));
  NOT NOT1_44(.VSS(VSS),.VDD(VDD),.Y(G317),.A(G324));
  NOT NOT1_45(.VSS(VSS),.VDD(VDD),.Y(G320),.A(G712));
  NOT NOT1_46(.VSS(VSS),.VDD(VDD),.Y(G323),.A(G324));
  NOT NOT1_47(.VSS(VSS),.VDD(VDD),.Y(G336),.A(G355));
  NOT NOT1_48(.VSS(VSS),.VDD(VDD),.Y(G339),.A(G355));
  NOT NOT1_49(.VSS(VSS),.VDD(VDD),.Y(G343),.A(G348));
  NOT NOT1_50(.VSS(VSS),.VDD(VDD),.Y(G347),.A(G348));
  NOT NOT1_51(.VSS(VSS),.VDD(VDD),.Y(G348),.A(G91));
  NOT NOT1_52(.VSS(VSS),.VDD(VDD),.Y(G351),.A(G645));
  NOT NOT1_53(.VSS(VSS),.VDD(VDD),.Y(G354),.A(G355));
  NOT NOT1_54(.VSS(VSS),.VDD(VDD),.Y(G359),.A(G372));
  NOT NOT1_55(.VSS(VSS),.VDD(VDD),.Y(G364),.A(G372));
  NOT NOT1_56(.VSS(VSS),.VDD(VDD),.Y(G371),.A(G372));
  NOT NOT1_57(.VSS(VSS),.VDD(VDD),.Y(G378),.A(G391));
  NOT NOT1_58(.VSS(VSS),.VDD(VDD),.Y(G383),.A(G391));
  NOT NOT1_59(.VSS(VSS),.VDD(VDD),.Y(G390),.A(G391));
  NOT NOT1_60(.VSS(VSS),.VDD(VDD),.Y(G396),.A(G404));
  NOT NOT1_61(.VSS(VSS),.VDD(VDD),.Y(G403),.A(G404));
  NOT NOT1_62(.VSS(VSS),.VDD(VDD),.Y(G407),.A(G712));
  NOT NOT1_63(.VSS(VSS),.VDD(VDD),.Y(G415),.A(G423));
  NOT NOT1_64(.VSS(VSS),.VDD(VDD),.Y(G422),.A(G423));
  NOT NOT1_65(.VSS(VSS),.VDD(VDD),.Y(G426),.A(G712));
  NOT NOT1_66(.VSS(VSS),.VDD(VDD),.Y(G437),.A(G712));
  NOT NOT1_67(.VSS(VSS),.VDD(VDD),.Y(G440),.A(G712));
  NOT NOT1_68(.VSS(VSS),.VDD(VDD),.Y(G445),.A(G65));
  NOT NOT1_69(.VSS(VSS),.VDD(VDD),.Y(G446),.A(G712));
  NOT NOT1_70(.VSS(VSS),.VDD(VDD),.Y(G449),.A(G66));
  NOT NOT1_71(.VSS(VSS),.VDD(VDD),.Y(G450),.A(G712));
  NOT NOT1_72(.VSS(VSS),.VDD(VDD),.Y(G455),.A(G456));
  NOT NOT1_73(.VSS(VSS),.VDD(VDD),.Y(G458),.A(G476));
  NOT NOT1_74(.VSS(VSS),.VDD(VDD),.Y(G463),.A(G476));
  NOT NOT1_75(.VSS(VSS),.VDD(VDD),.Y(G468),.A(G476));
  NOT NOT1_76(.VSS(VSS),.VDD(VDD),.Y(G475),.A(G476));
  NOT NOT1_77(.VSS(VSS),.VDD(VDD),.Y(G486),.A(G712));
  NOT NOT1_78(.VSS(VSS),.VDD(VDD),.Y(G491),.A(G500));
  NOT NOT1_79(.VSS(VSS),.VDD(VDD),.Y(G495),.A(G500));
  NOT NOT1_80(.VSS(VSS),.VDD(VDD),.Y(G499),.A(G500));
  NOT NOT1_81(.VSS(VSS),.VDD(VDD),.Y(G504),.A(G511));
  NOT NOT1_82(.VSS(VSS),.VDD(VDD),.Y(G507),.A(G511));
  NOT NOT1_83(.VSS(VSS),.VDD(VDD),.Y(G510),.A(G511));
  NOT NOT1_84(.VSS(VSS),.VDD(VDD),.Y(G511),.A(G63));
  NOT NOT1_85(.VSS(VSS),.VDD(VDD),.Y(G525),.A(G589));
  NOT NOT1_86(.VSS(VSS),.VDD(VDD),.Y(G530),.A(G589));
  NOT NOT1_87(.VSS(VSS),.VDD(VDD),.Y(G535),.A(G589));
  NOT NOT1_88(.VSS(VSS),.VDD(VDD),.Y(G540),.A(G589));
  NOT NOT1_89(.VSS(VSS),.VDD(VDD),.Y(G547),.A(G589));
  NOT NOT1_90(.VSS(VSS),.VDD(VDD),.Y(G562),.A(G610));
  NOT NOT1_91(.VSS(VSS),.VDD(VDD),.Y(G566),.A(G610));
  NOT NOT1_92(.VSS(VSS),.VDD(VDD),.Y(G570),.A(G610));
  NOT NOT1_93(.VSS(VSS),.VDD(VDD),.Y(G574),.A(G610));
  NOT NOT1_94(.VSS(VSS),.VDD(VDD),.Y(G588),.A(G589));
  NOT NOT1_95(.VSS(VSS),.VDD(VDD),.Y(G595),.A(G593));
  NOT NOT1_96(.VSS(VSS),.VDD(VDD),.Y(G596),.A(G597));
  NOT NOT1_97(.VSS(VSS),.VDD(VDD),.Y(G600),.A(G601));
  NOT NOT1_98(.VSS(VSS),.VDD(VDD),.Y(G605),.A(G610));
  NOT NOT1_99(.VSS(VSS),.VDD(VDD),.Y(G609),.A(G610));
  NOT NOT1_100(.VSS(VSS),.VDD(VDD),.Y(G614),.A(G64));
  NOT NOT1_101(.VSS(VSS),.VDD(VDD),.Y(G615),.A(G616));
  NOT NOT1_102(.VSS(VSS),.VDD(VDD),.Y(G617),.A(G645));
  NOT NOT1_103(.VSS(VSS),.VDD(VDD),.Y(G620),.A(G645));
  NOT NOT1_104(.VSS(VSS),.VDD(VDD),.Y(G623),.A(G645));
  NOT NOT1_105(.VSS(VSS),.VDD(VDD),.Y(G626),.A(G645));
  NOT NOT1_106(.VSS(VSS),.VDD(VDD),.Y(G629),.A(G645));
  NOT NOT1_107(.VSS(VSS),.VDD(VDD),.Y(G632),.A(G645));
  NOT NOT1_108(.VSS(VSS),.VDD(VDD),.Y(G635),.A(G645));
  NOT NOT1_109(.VSS(VSS),.VDD(VDD),.Y(G638),.A(G645));
  NOT NOT1_110(.VSS(VSS),.VDD(VDD),.Y(G641),.A(G645));
  NOT NOT1_111(.VSS(VSS),.VDD(VDD),.Y(G644),.A(G645));
  NOT NOT1_112(.VSS(VSS),.VDD(VDD),.Y(G645),.A(G90));
  NOT NOT1_113(.VSS(VSS),.VDD(VDD),.Y(G656),.A(G712));
  NOT NOT1_114(.VSS(VSS),.VDD(VDD),.Y(G658),.A(G659));
  NOT NOT1_115(.VSS(VSS),.VDD(VDD),.Y(I1162),.A(G13));
  NOT NOT1_116(.VSS(VSS),.VDD(VDD),.Y(G659),.A(I1162));
  NOT NOT1_117(.VSS(VSS),.VDD(VDD),.Y(G661),.A(G94));
  NOT NOT1_118(.VSS(VSS),.VDD(VDD),.Y(G662),.A(G712));
  NOT NOT1_119(.VSS(VSS),.VDD(VDD),.Y(G665),.A(G678));
  NOT NOT1_120(.VSS(VSS),.VDD(VDD),.Y(G668),.A(G712));
  NOT NOT1_121(.VSS(VSS),.VDD(VDD),.Y(G671),.A(G678));
  NOT NOT1_122(.VSS(VSS),.VDD(VDD),.Y(G674),.A(G712));
  NOT NOT1_123(.VSS(VSS),.VDD(VDD),.Y(G677),.A(G678));
  NOT NOT1_124(.VSS(VSS),.VDD(VDD),.Y(I1183),.A(G11));
  NOT NOT1_125(.VSS(VSS),.VDD(VDD),.Y(G678),.A(I1183));
  NOT NOT1_126(.VSS(VSS),.VDD(VDD),.Y(G685),.A(G696));
  NOT NOT1_127(.VSS(VSS),.VDD(VDD),.Y(G689),.A(G696));
  NOT NOT1_128(.VSS(VSS),.VDD(VDD),.Y(G695),.A(G696));
  NOT NOT1_129(.VSS(VSS),.VDD(VDD),.Y(I1203),.A(G10));
  NOT NOT1_130(.VSS(VSS),.VDD(VDD),.Y(G696),.A(I1203));
  NOT NOT1_131(.VSS(VSS),.VDD(VDD),.Y(G701),.A(G15));
  NOT NOT1_132(.VSS(VSS),.VDD(VDD),.Y(I1211),.A(G701));
  NOT NOT1_133(.VSS(VSS),.VDD(VDD),.Y(G701BF),.A(I1211));
  NOT NOT1_134(.VSS(VSS),.VDD(VDD),.Y(G704),.A(G712));
  NOT NOT1_135(.VSS(VSS),.VDD(VDD),.Y(G706),.A(G712));
  NOT NOT1_136(.VSS(VSS),.VDD(VDD),.Y(G711),.A(G712));
  NOT NOT1_137(.VSS(VSS),.VDD(VDD),.Y(G712),.A(G14));
  NOT NOT1_138(.VSS(VSS),.VDD(VDD),.Y(G714),.A(G701));
  NOT NOT1_139(.VSS(VSS),.VDD(VDD),.Y(I1227),.A(G6));
  NOT NOT1_140(.VSS(VSS),.VDD(VDD),.Y(G715),.A(I1227));
  NOT NOT1_141(.VSS(VSS),.VDD(VDD),.Y(I1230),.A(G7));
  NOT NOT1_142(.VSS(VSS),.VDD(VDD),.Y(G716),.A(I1230));
  NOT NOT1_143(.VSS(VSS),.VDD(VDD),.Y(I1233),.A(G8));
  NOT NOT1_144(.VSS(VSS),.VDD(VDD),.Y(G717),.A(I1233));
  NOT NOT1_145(.VSS(VSS),.VDD(VDD),.Y(I1236),.A(G9));
  NOT NOT1_146(.VSS(VSS),.VDD(VDD),.Y(G718),.A(I1236));
  NOT NOT1_147(.VSS(VSS),.VDD(VDD),.Y(I1239),.A(G12));
  NOT NOT1_148(.VSS(VSS),.VDD(VDD),.Y(G719),.A(I1239));
  NOT NOT1_149(.VSS(VSS),.VDD(VDD),.Y(I1242),.A(G0));
  NOT NOT1_150(.VSS(VSS),.VDD(VDD),.Y(G720),.A(I1242));
  NOT NOT1_151(.VSS(VSS),.VDD(VDD),.Y(I1245),.A(G1));
  NOT NOT1_152(.VSS(VSS),.VDD(VDD),.Y(G721),.A(I1245));
  NOT NOT1_153(.VSS(VSS),.VDD(VDD),.Y(I1248),.A(G2));
  NOT NOT1_154(.VSS(VSS),.VDD(VDD),.Y(G722),.A(I1248));
  NOT NOT1_155(.VSS(VSS),.VDD(VDD),.Y(I1251),.A(G3));
  NOT NOT1_156(.VSS(VSS),.VDD(VDD),.Y(G723),.A(I1251));
  NOT NOT1_157(.VSS(VSS),.VDD(VDD),.Y(I1254),.A(G4));
  NOT NOT1_158(.VSS(VSS),.VDD(VDD),.Y(G724),.A(I1254));
  NOT NOT1_159(.VSS(VSS),.VDD(VDD),.Y(I1257),.A(G5));
  NOT NOT1_160(.VSS(VSS),.VDD(VDD),.Y(G725),.A(I1257));
  NOT NOT1_161(.VSS(VSS),.VDD(VDD),.Y(I1260),.A(G93));
  NOT NOT1_162(.VSS(VSS),.VDD(VDD),.Y(G726),.A(I1260));
  NOT NOT1_163(.VSS(VSS),.VDD(VDD),.Y(I1264),.A(G16));
  NOT NOT1_164(.VSS(VSS),.VDD(VDD),.Y(G728),.A(I1264));
  NOT NOT1_165(.VSS(VSS),.VDD(VDD),.Y(I1267),.A(G95));
  NOT NOT1_166(.VSS(VSS),.VDD(VDD),.Y(G729),.A(I1267));
//
  AND2 AND2_0(.VSS(VSS),.VDD(VDD),.Y(G101),.A(G630),.B(G631));
  AND2 AND2_1(.VSS(VSS),.VDD(VDD),.Y(G102),.A(G633),.B(G634));
  AND2 AND2_2(.VSS(VSS),.VDD(VDD),.Y(G103),.A(G636),.B(G637));
  AND2 AND2_3(.VSS(VSS),.VDD(VDD),.Y(G104),.A(G639),.B(G640));
  AND2 AND2_4(.VSS(VSS),.VDD(VDD),.Y(G105),.A(G642),.B(G643));
  AND2 AND2_5(.VSS(VSS),.VDD(VDD),.Y(G109),.A(G106),.B(G108));
  AND2 AND2_6(.VSS(VSS),.VDD(VDD),.Y(G113),.A(G114),.B(G112));
  AND2 AND2_7(.VSS(VSS),.VDD(VDD),.Y(G116),.A(G133),.B(G25));
  AND2 AND2_8(.VSS(VSS),.VDD(VDD),.Y(G118),.A(G119),.B(G117));
  AND2 AND2_9(.VSS(VSS),.VDD(VDD),.Y(G121),.A(G134),.B(G26));
  AND2 AND2_10(.VSS(VSS),.VDD(VDD),.Y(G125),.A(G122),.B(G124));
  AND2 AND2_11(.VSS(VSS),.VDD(VDD),.Y(G129),.A(G130),.B(G128));
  AND2 AND2_12(.VSS(VSS),.VDD(VDD),.Y(G132),.A(G136),.B(G28));
  AND2 AND2_13(.VSS(VSS),.VDD(VDD),.Y(G133),.A(G700),.B(G111));
  AND2 AND2_14(.VSS(VSS),.VDD(VDD),.Y(G134),.A(G133),.B(G25));
  AND2 AND2_15(.VSS(VSS),.VDD(VDD),.Y(G135),.A(G134),.B(G26));
  AND2 AND2_16(.VSS(VSS),.VDD(VDD),.Y(G136),.A(G135),.B(G127));
  AND2 AND2_17(.VSS(VSS),.VDD(VDD),.Y(G140),.A(G137),.B(G139));
  AND2 AND2_18(.VSS(VSS),.VDD(VDD),.Y(G144),.A(G145),.B(G143));
  AND2 AND2_19(.VSS(VSS),.VDD(VDD),.Y(G147),.A(G168),.B(G30));
  AND2 AND2_20(.VSS(VSS),.VDD(VDD),.Y(G149),.A(G150),.B(G148));
  AND2 AND2_21(.VSS(VSS),.VDD(VDD),.Y(G152),.A(G169),.B(G31));
  AND2 AND2_22(.VSS(VSS),.VDD(VDD),.Y(G154),.A(G155),.B(G153));
  AND2 AND2_23(.VSS(VSS),.VDD(VDD),.Y(G157),.A(G170),.B(G32));
  AND2 AND2_24(.VSS(VSS),.VDD(VDD),.Y(G159),.A(G160),.B(G158));
  AND2 AND2_25(.VSS(VSS),.VDD(VDD),.Y(G162),.A(G171),.B(G33));
  AND2 AND2_26(.VSS(VSS),.VDD(VDD),.Y(G166),.A(G163),.B(G165));
  AND2 AND2_27(.VSS(VSS),.VDD(VDD),.Y(G168),.A(G177),.B(G142));
  AND2 AND2_28(.VSS(VSS),.VDD(VDD),.Y(G169),.A(G168),.B(G30));
  AND2 AND2_29(.VSS(VSS),.VDD(VDD),.Y(G170),.A(G169),.B(G31));
  AND2 AND2_30(.VSS(VSS),.VDD(VDD),.Y(G171),.A(G170),.B(G32));
  AND2 AND2_31(.VSS(VSS),.VDD(VDD),.Y(G172),.A(G171),.B(G33));
  AND2 AND2_32(.VSS(VSS),.VDD(VDD),.Y(G173),.A(G172),.B(G34));
  AND2 AND2_33(.VSS(VSS),.VDD(VDD),.Y(G175),.A(G176),.B(G174));
  AND2 AND2_34(.VSS(VSS),.VDD(VDD),.Y(G185),.A(G181),.B(G182));
  AND2 AND2_35(.VSS(VSS),.VDD(VDD),.Y(G189),.A(G186),.B(G188));
  AND2 AND2_36(.VSS(VSS),.VDD(VDD),.Y(G193),.A(G194),.B(G192));
  AND2 AND2_37(.VSS(VSS),.VDD(VDD),.Y(G196),.A(G202),.B(G37));
  AND2 AND2_38(.VSS(VSS),.VDD(VDD),.Y(G198),.A(G199),.B(G197));
  AND2 AND2_39(.VSS(VSS),.VDD(VDD),.Y(G201),.A(G203),.B(G38));
  AND2 AND2_40(.VSS(VSS),.VDD(VDD),.Y(G202),.A(G522),.B(G191));
  AND2 AND2_41(.VSS(VSS),.VDD(VDD),.Y(G203),.A(G202),.B(G37));
  AND2 AND2_42(.VSS(VSS),.VDD(VDD),.Y(G208),.A(G205),.B(G207));
  AND2 AND2_43(.VSS(VSS),.VDD(VDD),.Y(G214),.A(G211),.B(G213));
  AND2 AND2_44(.VSS(VSS),.VDD(VDD),.Y(G218),.A(G219),.B(G217));
  AND2 AND2_45(.VSS(VSS),.VDD(VDD),.Y(G221),.A(G223),.B(G41));
  AND2 AND2_46(.VSS(VSS),.VDD(VDD),.Y(G222),.A(G183),.B(G210));
  AND2 AND2_47(.VSS(VSS),.VDD(VDD),.Y(G223),.A(G222),.B(G216));
  AND2 AND2_48(.VSS(VSS),.VDD(VDD),.Y(G224),.A(G203),.B(G38));
  AND2 AND2_49(.VSS(VSS),.VDD(VDD),.Y(G225),.A(G204),.B(G203));
  AND2 AND2_50(.VSS(VSS),.VDD(VDD),.Y(G226),.A(G136),.B(G28));
  AND2 AND2_51(.VSS(VSS),.VDD(VDD),.Y(G227),.A(G172),.B(G178));
  AND2 AND2_52(.VSS(VSS),.VDD(VDD),.Y(G228),.A(G223),.B(G41));
  AND2 AND2_53(.VSS(VSS),.VDD(VDD),.Y(G229),.A(G432),.B(G62));
  AND2 AND2_54(.VSS(VSS),.VDD(VDD),.Y(G237),.A(G238),.B(G236));
  AND2 AND2_55(.VSS(VSS),.VDD(VDD),.Y(G240),.A(G299),.B(G42));
  AND2 AND2_56(.VSS(VSS),.VDD(VDD),.Y(G242),.A(G243),.B(G241));
  AND2 AND2_57(.VSS(VSS),.VDD(VDD),.Y(G245),.A(G262),.B(G43));
  AND2 AND2_58(.VSS(VSS),.VDD(VDD),.Y(G247),.A(G248),.B(G246));
  AND2 AND2_59(.VSS(VSS),.VDD(VDD),.Y(G250),.A(G263),.B(G44));
  AND2 AND2_60(.VSS(VSS),.VDD(VDD),.Y(G252),.A(G253),.B(G251));
  AND2 AND2_61(.VSS(VSS),.VDD(VDD),.Y(G255),.A(G264),.B(G45));
  AND2 AND2_62(.VSS(VSS),.VDD(VDD),.Y(G259),.A(G624),.B(G625));
  AND2 AND2_63(.VSS(VSS),.VDD(VDD),.Y(G260),.A(G256),.B(G258));
  AND2 AND2_64(.VSS(VSS),.VDD(VDD),.Y(G261),.A(G265),.B(G46));
  AND2 AND2_65(.VSS(VSS),.VDD(VDD),.Y(G262),.A(G299),.B(G42));
  AND2 AND2_66(.VSS(VSS),.VDD(VDD),.Y(G263),.A(G262),.B(G43));
  AND2 AND2_67(.VSS(VSS),.VDD(VDD),.Y(G264),.A(G263),.B(G44));
  AND2 AND2_68(.VSS(VSS),.VDD(VDD),.Y(G265),.A(G264),.B(G45));
  AND2 AND2_69(.VSS(VSS),.VDD(VDD),.Y(G271),.A(G275),.B(G266));
  AND2 AND2_70(.VSS(VSS),.VDD(VDD),.Y(G272),.A(G276),.B(G277));
  AND2 AND2_71(.VSS(VSS),.VDD(VDD),.Y(G273),.A(G278),.B(G279));
  AND2 AND2_72(.VSS(VSS),.VDD(VDD),.Y(G274),.A(G280),.B(G281));
  AND2 AND2_73(.VSS(VSS),.VDD(VDD),.Y(G303),.A(G304),.B(G302));
  AND2 AND2_74(.VSS(VSS),.VDD(VDD),.Y(G304),.A(G306),.B(G307));
  AND2 AND2_75(.VSS(VSS),.VDD(VDD),.Y(G309),.A(G310),.B(G308));
  AND2 AND2_76(.VSS(VSS),.VDD(VDD),.Y(G310),.A(G312),.B(G313));
  AND2 AND2_77(.VSS(VSS),.VDD(VDD),.Y(G315),.A(G316),.B(G314));
  AND2 AND2_78(.VSS(VSS),.VDD(VDD),.Y(G316),.A(G318),.B(G319));
  AND2 AND2_79(.VSS(VSS),.VDD(VDD),.Y(G321),.A(G322),.B(G320));
  AND2 AND2_80(.VSS(VSS),.VDD(VDD),.Y(G322),.A(G325),.B(G326));
  AND2 AND2_81(.VSS(VSS),.VDD(VDD),.Y(G329),.A(G331),.B(G714));
  AND2 AND2_82(.VSS(VSS),.VDD(VDD),.Y(G330),.A(G332),.B(G714));
  AND2 AND2_83(.VSS(VSS),.VDD(VDD),.Y(G335),.A(G337),.B(G338));
  AND2 AND2_84(.VSS(VSS),.VDD(VDD),.Y(G342),.A(G344),.B(G345));
  AND2 AND2_85(.VSS(VSS),.VDD(VDD),.Y(G346),.A(G349),.B(G350));
  AND2 AND2_86(.VSS(VSS),.VDD(VDD),.Y(G358),.A(G523),.B(G53));
  AND2 AND2_87(.VSS(VSS),.VDD(VDD),.Y(G360),.A(G361),.B(G359));
  AND2 AND2_88(.VSS(VSS),.VDD(VDD),.Y(G363),.A(G523),.B(G51));
  AND2 AND2_89(.VSS(VSS),.VDD(VDD),.Y(G365),.A(G366),.B(G364));
  AND2 AND2_90(.VSS(VSS),.VDD(VDD),.Y(G368),.A(G375),.B(G52));
  AND2 AND2_91(.VSS(VSS),.VDD(VDD),.Y(G373),.A(G369),.B(G371));
  AND2 AND2_92(.VSS(VSS),.VDD(VDD),.Y(G374),.A(G376),.B(G53));
  AND2 AND2_93(.VSS(VSS),.VDD(VDD),.Y(G375),.A(G523),.B(G51));
  AND2 AND2_94(.VSS(VSS),.VDD(VDD),.Y(G376),.A(G375),.B(G52));
  AND3 AND3_0(.VSS(VSS),.VDD(VDD),.Y(G377),.A(G183),.B(G54),.C(G56));
  AND2 AND2_95(.VSS(VSS),.VDD(VDD),.Y(G379),.A(G380),.B(G378));
  AND2 AND2_96(.VSS(VSS),.VDD(VDD),.Y(G382),.A(G183),.B(G54));
  AND2 AND2_97(.VSS(VSS),.VDD(VDD),.Y(G384),.A(G385),.B(G383));
  AND2 AND2_98(.VSS(VSS),.VDD(VDD),.Y(G387),.A(G394),.B(G55));
  AND2 AND2_99(.VSS(VSS),.VDD(VDD),.Y(G392),.A(G388),.B(G390));
  AND2 AND2_100(.VSS(VSS),.VDD(VDD),.Y(G393),.A(G395),.B(G56));
  AND2 AND2_101(.VSS(VSS),.VDD(VDD),.Y(G394),.A(G183),.B(G54));
  AND2 AND2_102(.VSS(VSS),.VDD(VDD),.Y(G395),.A(G394),.B(G55));
  AND2 AND2_103(.VSS(VSS),.VDD(VDD),.Y(G397),.A(G398),.B(G396));
  AND2 AND2_104(.VSS(VSS),.VDD(VDD),.Y(G400),.A(G335),.B(G57));
  AND2 AND2_105(.VSS(VSS),.VDD(VDD),.Y(G405),.A(G401),.B(G403));
  AND2 AND2_106(.VSS(VSS),.VDD(VDD),.Y(G406),.A(G412),.B(G58));
  AND2 AND2_107(.VSS(VSS),.VDD(VDD),.Y(G408),.A(G409),.B(G407));
  AND2 AND2_108(.VSS(VSS),.VDD(VDD),.Y(G411),.A(G413),.B(G59));
  AND2 AND2_109(.VSS(VSS),.VDD(VDD),.Y(G412),.A(G335),.B(G57));
  AND2 AND2_110(.VSS(VSS),.VDD(VDD),.Y(G413),.A(G335),.B(G58));
  AND2 AND2_111(.VSS(VSS),.VDD(VDD),.Y(G414),.A(G413),.B(G59));
  AND2 AND2_112(.VSS(VSS),.VDD(VDD),.Y(G416),.A(G417),.B(G415));
  AND2 AND2_113(.VSS(VSS),.VDD(VDD),.Y(G419),.A(G358),.B(G60));
  AND2 AND2_114(.VSS(VSS),.VDD(VDD),.Y(G424),.A(G420),.B(G422));
  AND2 AND2_115(.VSS(VSS),.VDD(VDD),.Y(G425),.A(G431),.B(G61));
  AND2 AND2_116(.VSS(VSS),.VDD(VDD),.Y(G427),.A(G428),.B(G426));
  AND2 AND2_117(.VSS(VSS),.VDD(VDD),.Y(G430),.A(G432),.B(G62));
  AND2 AND2_118(.VSS(VSS),.VDD(VDD),.Y(G431),.A(G358),.B(G60));
  AND2 AND2_119(.VSS(VSS),.VDD(VDD),.Y(G432),.A(G358),.B(G61));
  AND2 AND2_120(.VSS(VSS),.VDD(VDD),.Y(G433),.A(G356),.B(G357));
  AND2 AND2_121(.VSS(VSS),.VDD(VDD),.Y(G435),.A(G340),.B(G341));
  AND2 AND2_122(.VSS(VSS),.VDD(VDD),.Y(G436),.A(G352),.B(G353));
  AND2 AND2_123(.VSS(VSS),.VDD(VDD),.Y(G438),.A(G439),.B(G437));
  AND2 AND2_124(.VSS(VSS),.VDD(VDD),.Y(G441),.A(G442),.B(G440));
  AND2 AND2_125(.VSS(VSS),.VDD(VDD),.Y(G443),.A(G615),.B(G511));
  AND2 AND2_126(.VSS(VSS),.VDD(VDD),.Y(G447),.A(G448),.B(G446));
  AND2 AND2_127(.VSS(VSS),.VDD(VDD),.Y(G451),.A(G452),.B(G450));
  AND2 AND2_128(.VSS(VSS),.VDD(VDD),.Y(G453),.A(G615),.B(G445));
  AND3 AND3_1(.VSS(VSS),.VDD(VDD),.Y(G457),.A(G455),.B(G449),.C(G728));
  AND2 AND2_129(.VSS(VSS),.VDD(VDD),.Y(G459),.A(G460),.B(G458));
  AND2 AND2_130(.VSS(VSS),.VDD(VDD),.Y(G462),.A(G434),.B(G67));
  AND2 AND2_131(.VSS(VSS),.VDD(VDD),.Y(G464),.A(G465),.B(G463));
  AND2 AND2_132(.VSS(VSS),.VDD(VDD),.Y(G467),.A(G479),.B(G68));
  AND2 AND2_133(.VSS(VSS),.VDD(VDD),.Y(G469),.A(G470),.B(G468));
  AND2 AND2_134(.VSS(VSS),.VDD(VDD),.Y(G472),.A(G480),.B(G69));
  AND2 AND2_135(.VSS(VSS),.VDD(VDD),.Y(G477),.A(G473),.B(G475));
  AND2 AND2_136(.VSS(VSS),.VDD(VDD),.Y(G478),.A(G481),.B(G70));
  AND2 AND2_137(.VSS(VSS),.VDD(VDD),.Y(G479),.A(G434),.B(G67));
  AND2 AND2_138(.VSS(VSS),.VDD(VDD),.Y(G480),.A(G479),.B(G68));
  AND2 AND2_139(.VSS(VSS),.VDD(VDD),.Y(G481),.A(G480),.B(G69));
  AND2 AND2_140(.VSS(VSS),.VDD(VDD),.Y(G488),.A(G505),.B(G506));
  AND2 AND2_141(.VSS(VSS),.VDD(VDD),.Y(G489),.A(G508),.B(G509));
  AND2 AND2_142(.VSS(VSS),.VDD(VDD),.Y(G490),.A(G512),.B(G513));
  AND2 AND2_143(.VSS(VSS),.VDD(VDD),.Y(G494),.A(G492),.B(G493));
  AND2 AND2_144(.VSS(VSS),.VDD(VDD),.Y(G498),.A(G496),.B(G497));
  AND2 AND2_145(.VSS(VSS),.VDD(VDD),.Y(G503),.A(G501),.B(G502));
  AND2 AND2_146(.VSS(VSS),.VDD(VDD),.Y(G526),.A(G527),.B(G525));
  AND2 AND2_147(.VSS(VSS),.VDD(VDD),.Y(G529),.A(G604),.B(G74));
  AND2 AND2_148(.VSS(VSS),.VDD(VDD),.Y(G531),.A(G532),.B(G530));
  AND2 AND2_149(.VSS(VSS),.VDD(VDD),.Y(G534),.A(G550),.B(G75));
  AND2 AND2_150(.VSS(VSS),.VDD(VDD),.Y(G536),.A(G537),.B(G535));
  AND2 AND2_151(.VSS(VSS),.VDD(VDD),.Y(G539),.A(G551),.B(G76));
  AND2 AND2_152(.VSS(VSS),.VDD(VDD),.Y(G541),.A(G542),.B(G540));
  AND2 AND2_153(.VSS(VSS),.VDD(VDD),.Y(G544),.A(G552),.B(G77));
  AND2 AND2_154(.VSS(VSS),.VDD(VDD),.Y(G548),.A(G545),.B(G547));
  AND2 AND2_155(.VSS(VSS),.VDD(VDD),.Y(G549),.A(G553),.B(G78));
  AND2 AND2_156(.VSS(VSS),.VDD(VDD),.Y(G550),.A(G604),.B(G74));
  AND2 AND2_157(.VSS(VSS),.VDD(VDD),.Y(G551),.A(G550),.B(G75));
  AND2 AND2_158(.VSS(VSS),.VDD(VDD),.Y(G552),.A(G551),.B(G76));
  AND2 AND2_159(.VSS(VSS),.VDD(VDD),.Y(G553),.A(G552),.B(G77));
  AND2 AND2_160(.VSS(VSS),.VDD(VDD),.Y(G565),.A(G563),.B(G564));
  AND2 AND2_161(.VSS(VSS),.VDD(VDD),.Y(G569),.A(G567),.B(G568));
  AND2 AND2_162(.VSS(VSS),.VDD(VDD),.Y(G573),.A(G571),.B(G572));
  AND2 AND2_163(.VSS(VSS),.VDD(VDD),.Y(G577),.A(G575),.B(G576));
  AND2 AND2_164(.VSS(VSS),.VDD(VDD),.Y(G589),.A(G627),.B(G628));
  AND2 AND2_165(.VSS(VSS),.VDD(VDD),.Y(G590),.A(G591),.B(G588));
  AND2 AND2_166(.VSS(VSS),.VDD(VDD),.Y(G592),.A(G594),.B(G595));
  AND2 AND2_167(.VSS(VSS),.VDD(VDD),.Y(G601),.A(G621),.B(G622));
  AND2 AND2_168(.VSS(VSS),.VDD(VDD),.Y(G604),.A(G433),.B(G524));
  AND2 AND2_169(.VSS(VSS),.VDD(VDD),.Y(G608),.A(G606),.B(G607));
  AND2 AND2_170(.VSS(VSS),.VDD(VDD),.Y(G613),.A(G611),.B(G612));
  AND2 AND2_171(.VSS(VSS),.VDD(VDD),.Y(G648),.A(G646),.B(G647));
  AND2 AND2_172(.VSS(VSS),.VDD(VDD),.Y(G649),.A(G618),.B(G619));
  AND2 AND2_173(.VSS(VSS),.VDD(VDD),.Y(G650),.A(G226),.B(G661));
  AND2 AND2_174(.VSS(VSS),.VDD(VDD),.Y(G651),.A(G227),.B(G87));
  AND2 AND2_175(.VSS(VSS),.VDD(VDD),.Y(G652),.A(G228),.B(G88));
  AND2 AND2_176(.VSS(VSS),.VDD(VDD),.Y(G653),.A(G229),.B(G89));
  AND2 AND2_177(.VSS(VSS),.VDD(VDD),.Y(G654),.A(G90),.B(G476));
  AND2 AND2_178(.VSS(VSS),.VDD(VDD),.Y(G655),.A(G91),.B(G476));
  AND2 AND2_179(.VSS(VSS),.VDD(VDD),.Y(G657),.A(G659),.B(G656));
  AND2 AND2_180(.VSS(VSS),.VDD(VDD),.Y(G663),.A(G664),.B(G662));
  AND2 AND2_181(.VSS(VSS),.VDD(VDD),.Y(G664),.A(G666),.B(G667));
  AND2 AND2_182(.VSS(VSS),.VDD(VDD),.Y(G669),.A(G670),.B(G668));
  AND2 AND2_183(.VSS(VSS),.VDD(VDD),.Y(G670),.A(G672),.B(G673));
  AND2 AND2_184(.VSS(VSS),.VDD(VDD),.Y(G675),.A(G676),.B(G674));
  AND2 AND2_185(.VSS(VSS),.VDD(VDD),.Y(G676),.A(G679),.B(G680));
  AND2 AND2_186(.VSS(VSS),.VDD(VDD),.Y(G683),.A(G684),.B(G685));
  AND2 AND2_187(.VSS(VSS),.VDD(VDD),.Y(G688),.A(G690),.B(G691));
  AND2 AND2_188(.VSS(VSS),.VDD(VDD),.Y(G694),.A(G697),.B(G698));
  AND2 AND2_189(.VSS(VSS),.VDD(VDD),.Y(G702),.A(G703),.B(G645));
  AND2 AND2_190(.VSS(VSS),.VDD(VDD),.Y(G705),.A(G230),.B(G704));
  AND2 AND2_191(.VSS(VSS),.VDD(VDD),.Y(G707),.A(G708),.B(G706));
  AND2 AND2_192(.VSS(VSS),.VDD(VDD),.Y(G709),.A(G678),.B(G89));
  AND2 AND2_193(.VSS(VSS),.VDD(VDD),.Y(G713),.A(G599),.B(G711));
  AND2 AND2_194(.VSS(VSS),.VDD(VDD),.Y(G727),.A(G476),.B(G645));
//
  OR2 OR2_0(.VSS(VSS),.VDD(VDD),.Y(G110),.A(G700),.B(G111));
  OR2 OR2_1(.VSS(VSS),.VDD(VDD),.Y(G126),.A(G135),.B(G127));
  OR2 OR2_2(.VSS(VSS),.VDD(VDD),.Y(G141),.A(G177),.B(G142));
  OR2 OR2_3(.VSS(VSS),.VDD(VDD),.Y(G167),.A(G172),.B(G178));
  OR2 OR2_4(.VSS(VSS),.VDD(VDD),.Y(G177),.A(G180),.B(G226));
  OR2 OR2_5(.VSS(VSS),.VDD(VDD),.Y(G181),.A(G178),.B(G180));
  OR2 OR2_6(.VSS(VSS),.VDD(VDD),.Y(G182),.A(G35),.B(G179));
  OR2 OR2_7(.VSS(VSS),.VDD(VDD),.Y(G183),.A(G180),.B(G227));
  OR2 OR2_8(.VSS(VSS),.VDD(VDD),.Y(G184),.A(G180),.B(G173));
  OR2 OR2_9(.VSS(VSS),.VDD(VDD),.Y(G190),.A(G522),.B(G191));
  OR2 OR2_10(.VSS(VSS),.VDD(VDD),.Y(G209),.A(G183),.B(G210));
  OR2 OR2_11(.VSS(VSS),.VDD(VDD),.Y(G215),.A(G222),.B(G216));
  OR2 OR2_12(.VSS(VSS),.VDD(VDD),.Y(G235),.A(G649),.B(G233));
  OR2 OR2_13(.VSS(VSS),.VDD(VDD),.Y(G275),.A(G101),.B(G42));
  OR2 OR2_14(.VSS(VSS),.VDD(VDD),.Y(G276),.A(G102),.B(G43));
  OR2 OR2_15(.VSS(VSS),.VDD(VDD),.Y(G277),.A(G267),.B(G271));
  OR2 OR2_16(.VSS(VSS),.VDD(VDD),.Y(G278),.A(G103),.B(G44));
  OR2 OR2_17(.VSS(VSS),.VDD(VDD),.Y(G279),.A(G268),.B(G272));
  OR2 OR2_18(.VSS(VSS),.VDD(VDD),.Y(G280),.A(G104),.B(G45));
  OR2 OR2_19(.VSS(VSS),.VDD(VDD),.Y(G281),.A(G269),.B(G273));
  OR2 OR2_20(.VSS(VSS),.VDD(VDD),.Y(G282),.A(G105),.B(G46));
  OR2 OR2_21(.VSS(VSS),.VDD(VDD),.Y(G283),.A(G270),.B(G274));
  OR2 OR2_22(.VSS(VSS),.VDD(VDD),.Y(G291),.A(G42),.B(G101));
  OR2 OR2_23(.VSS(VSS),.VDD(VDD),.Y(G292),.A(G43),.B(G102));
  OR2 OR2_24(.VSS(VSS),.VDD(VDD),.Y(G293),.A(G44),.B(G103));
  OR2 OR2_25(.VSS(VSS),.VDD(VDD),.Y(G294),.A(G45),.B(G104));
  OR2 OR2_26(.VSS(VSS),.VDD(VDD),.Y(G295),.A(G46),.B(G105));
  OR4 OR4_0(.VSS(VSS),.VDD(VDD),.Y(G300),.A(G50),.B(G49),.C(G48),.D(G47));
  OR2 OR2_27(.VSS(VSS),.VDD(VDD),.Y(G306),.A(G47),.B(G324));
  OR2 OR2_28(.VSS(VSS),.VDD(VDD),.Y(G307),.A(G719),.B(G305));
  OR2 OR2_29(.VSS(VSS),.VDD(VDD),.Y(G312),.A(G48),.B(G324));
  OR2 OR2_30(.VSS(VSS),.VDD(VDD),.Y(G313),.A(G47),.B(G311));
  OR2 OR2_31(.VSS(VSS),.VDD(VDD),.Y(G318),.A(G49),.B(G324));
  OR2 OR2_32(.VSS(VSS),.VDD(VDD),.Y(G319),.A(G48),.B(G317));
  OR2 OR2_33(.VSS(VSS),.VDD(VDD),.Y(G324),.A(G377),.B(G348));
  OR2 OR2_34(.VSS(VSS),.VDD(VDD),.Y(G325),.A(G50),.B(G324));
  OR2 OR2_35(.VSS(VSS),.VDD(VDD),.Y(G326),.A(G49),.B(G323));
  OR2 OR2_36(.VSS(VSS),.VDD(VDD),.Y(G333),.A(G300),.B(G714));
  OR2 OR2_37(.VSS(VSS),.VDD(VDD),.Y(G334),.A(G301),.B(G714));
  OR2 OR2_38(.VSS(VSS),.VDD(VDD),.Y(G337),.A(G224),.B(G355));
  OR2 OR2_39(.VSS(VSS),.VDD(VDD),.Y(G338),.A(G183),.B(G336));
  OR2 OR2_40(.VSS(VSS),.VDD(VDD),.Y(G340),.A(G38),.B(G355));
  OR2 OR2_41(.VSS(VSS),.VDD(VDD),.Y(G341),.A(G185),.B(G339));
  OR2 OR2_42(.VSS(VSS),.VDD(VDD),.Y(G344),.A(G229),.B(G348));
  OR2 OR2_43(.VSS(VSS),.VDD(VDD),.Y(G345),.A(G414),.B(G343));
  OR2 OR2_44(.VSS(VSS),.VDD(VDD),.Y(G349),.A(G62),.B(G348));
  OR2 OR2_45(.VSS(VSS),.VDD(VDD),.Y(G350),.A(G59),.B(G347));
  OR2 OR2_46(.VSS(VSS),.VDD(VDD),.Y(G352),.A(G346),.B(G645));
  OR2 OR2_47(.VSS(VSS),.VDD(VDD),.Y(G353),.A(G35),.B(G351));
  OR2 OR2_48(.VSS(VSS),.VDD(VDD),.Y(G355),.A(G457),.B(G645));
  OR2 OR2_49(.VSS(VSS),.VDD(VDD),.Y(G356),.A(G225),.B(G355));
  OR2 OR2_50(.VSS(VSS),.VDD(VDD),.Y(G357),.A(G184),.B(G354));
  OR2 OR2_51(.VSS(VSS),.VDD(VDD),.Y(G372),.A(G712),.B(G358));
  OR2 OR2_52(.VSS(VSS),.VDD(VDD),.Y(G391),.A(G712),.B(G377));
  OR2 OR2_53(.VSS(VSS),.VDD(VDD),.Y(G404),.A(G712),.B(G413));
  OR2 OR2_54(.VSS(VSS),.VDD(VDD),.Y(G423),.A(G712),.B(G432));
  OR2 OR2_55(.VSS(VSS),.VDD(VDD),.Y(G434),.A(G342),.B(G645));
  OR2 OR2_56(.VSS(VSS),.VDD(VDD),.Y(G439),.A(G435),.B(G63));
  OR2 OR2_57(.VSS(VSS),.VDD(VDD),.Y(G448),.A(G615),.B(G65));
  OR2 OR2_58(.VSS(VSS),.VDD(VDD),.Y(G456),.A(G83),.B(G524));
  OR2 OR2_59(.VSS(VSS),.VDD(VDD),.Y(G492),.A(G71),.B(G500));
  OR2 OR2_60(.VSS(VSS),.VDD(VDD),.Y(G493),.A(G488),.B(G491));
  OR2 OR2_61(.VSS(VSS),.VDD(VDD),.Y(G496),.A(G72),.B(G500));
  OR2 OR2_62(.VSS(VSS),.VDD(VDD),.Y(G497),.A(G489),.B(G495));
  OR2 OR2_63(.VSS(VSS),.VDD(VDD),.Y(G500),.A(G654),.B(G712));
  OR2 OR2_64(.VSS(VSS),.VDD(VDD),.Y(G501),.A(G73),.B(G500));
  OR2 OR2_65(.VSS(VSS),.VDD(VDD),.Y(G502),.A(G490),.B(G499));
  OR2 OR2_66(.VSS(VSS),.VDD(VDD),.Y(G505),.A(G723),.B(G511));
  OR2 OR2_67(.VSS(VSS),.VDD(VDD),.Y(G506),.A(G720),.B(G504));
  OR2 OR2_68(.VSS(VSS),.VDD(VDD),.Y(G508),.A(G724),.B(G511));
  OR2 OR2_69(.VSS(VSS),.VDD(VDD),.Y(G509),.A(G721),.B(G507));
  OR2 OR2_70(.VSS(VSS),.VDD(VDD),.Y(G512),.A(G725),.B(G511));
  OR2 OR2_71(.VSS(VSS),.VDD(VDD),.Y(G513),.A(G722),.B(G510));
  OR2 OR2_72(.VSS(VSS),.VDD(VDD),.Y(G518),.A(G71),.B(G67));
  OR2 OR2_73(.VSS(VSS),.VDD(VDD),.Y(G519),.A(G72),.B(G68));
  OR2 OR2_74(.VSS(VSS),.VDD(VDD),.Y(G520),.A(G73),.B(G69));
  OR2 OR2_75(.VSS(VSS),.VDD(VDD),.Y(G521),.A(G487),.B(G70));
  OR2 OR2_76(.VSS(VSS),.VDD(VDD),.Y(G522),.A(G348),.B(G228));
  OR2 OR2_77(.VSS(VSS),.VDD(VDD),.Y(G523),.A(G348),.B(G414));
  OR2 OR2_78(.VSS(VSS),.VDD(VDD),.Y(G524),.A(G554),.B(G555));
  OR2 OR2_79(.VSS(VSS),.VDD(VDD),.Y(G563),.A(G79),.B(G610));
  OR2 OR2_80(.VSS(VSS),.VDD(VDD),.Y(G564),.A(G715),.B(G562));
  OR2 OR2_81(.VSS(VSS),.VDD(VDD),.Y(G567),.A(G80),.B(G610));
  OR2 OR2_82(.VSS(VSS),.VDD(VDD),.Y(G568),.A(G716),.B(G566));
  OR2 OR2_83(.VSS(VSS),.VDD(VDD),.Y(G571),.A(G81),.B(G610));
  OR2 OR2_84(.VSS(VSS),.VDD(VDD),.Y(G572),.A(G717),.B(G570));
  OR2 OR2_85(.VSS(VSS),.VDD(VDD),.Y(G575),.A(G82),.B(G610));
  OR2 OR2_86(.VSS(VSS),.VDD(VDD),.Y(G576),.A(G718),.B(G574));
  OR2 OR2_87(.VSS(VSS),.VDD(VDD),.Y(G583),.A(G79),.B(G74));
  OR2 OR2_88(.VSS(VSS),.VDD(VDD),.Y(G584),.A(G80),.B(G75));
  OR2 OR2_89(.VSS(VSS),.VDD(VDD),.Y(G585),.A(G81),.B(G76));
  OR2 OR2_90(.VSS(VSS),.VDD(VDD),.Y(G586),.A(G82),.B(G77));
  OR2 OR2_91(.VSS(VSS),.VDD(VDD),.Y(G587),.A(G561),.B(G78));
  OR2 OR2_92(.VSS(VSS),.VDD(VDD),.Y(G591),.A(G592),.B(G604));
  OR2 OR2_93(.VSS(VSS),.VDD(VDD),.Y(G594),.A(G83),.B(G593));
  OR2 OR2_94(.VSS(VSS),.VDD(VDD),.Y(G602),.A(G85),.B(G601));
  OR2 OR2_95(.VSS(VSS),.VDD(VDD),.Y(G603),.A(G600),.B(G84));
  OR2 OR2_96(.VSS(VSS),.VDD(VDD),.Y(G606),.A(G84),.B(G610));
  OR2 OR2_97(.VSS(VSS),.VDD(VDD),.Y(G607),.A(G696),.B(G605));
  OR2 OR2_98(.VSS(VSS),.VDD(VDD),.Y(G610),.A(G655),.B(G712));
  OR2 OR2_99(.VSS(VSS),.VDD(VDD),.Y(G611),.A(G85),.B(G610));
  OR2 OR2_100(.VSS(VSS),.VDD(VDD),.Y(G612),.A(G678),.B(G609));
  OR2 OR2_101(.VSS(VSS),.VDD(VDD),.Y(G618),.A(G457),.B(G645));
  OR2 OR2_102(.VSS(VSS),.VDD(VDD),.Y(G619),.A(G715),.B(G617));
  OR2 OR2_103(.VSS(VSS),.VDD(VDD),.Y(G621),.A(G614),.B(G645));
  OR2 OR2_104(.VSS(VSS),.VDD(VDD),.Y(G622),.A(G717),.B(G620));
  OR2 OR2_105(.VSS(VSS),.VDD(VDD),.Y(G624),.A(G476),.B(G645));
  OR2 OR2_106(.VSS(VSS),.VDD(VDD),.Y(G625),.A(G716),.B(G623));
  OR2 OR2_107(.VSS(VSS),.VDD(VDD),.Y(G627),.A(G476),.B(G645));
  OR2 OR2_108(.VSS(VSS),.VDD(VDD),.Y(G628),.A(G718),.B(G626));
  OR2 OR2_109(.VSS(VSS),.VDD(VDD),.Y(G630),.A(G96),.B(G645));
  OR2 OR2_110(.VSS(VSS),.VDD(VDD),.Y(G631),.A(G720),.B(G629));
  OR2 OR2_111(.VSS(VSS),.VDD(VDD),.Y(G633),.A(G97),.B(G645));
  OR2 OR2_112(.VSS(VSS),.VDD(VDD),.Y(G634),.A(G721),.B(G632));
  OR2 OR2_113(.VSS(VSS),.VDD(VDD),.Y(G636),.A(G98),.B(G645));
  OR2 OR2_114(.VSS(VSS),.VDD(VDD),.Y(G637),.A(G722),.B(G635));
  OR2 OR2_115(.VSS(VSS),.VDD(VDD),.Y(G639),.A(G99),.B(G645));
  OR2 OR2_116(.VSS(VSS),.VDD(VDD),.Y(G640),.A(G723),.B(G638));
  OR2 OR2_117(.VSS(VSS),.VDD(VDD),.Y(G642),.A(G100),.B(G645));
  OR2 OR2_118(.VSS(VSS),.VDD(VDD),.Y(G643),.A(G724),.B(G641));
  OR2 OR2_119(.VSS(VSS),.VDD(VDD),.Y(G646),.A(G456),.B(G645));
  OR2 OR2_120(.VSS(VSS),.VDD(VDD),.Y(G647),.A(G725),.B(G644));
  OR2 OR2_121(.VSS(VSS),.VDD(VDD),.Y(G666),.A(G87),.B(G678));
  OR2 OR2_122(.VSS(VSS),.VDD(VDD),.Y(G667),.A(G661),.B(G665));
  OR2 OR2_123(.VSS(VSS),.VDD(VDD),.Y(G672),.A(G88),.B(G678));
  OR2 OR2_124(.VSS(VSS),.VDD(VDD),.Y(G673),.A(G87),.B(G671));
  OR2 OR2_125(.VSS(VSS),.VDD(VDD),.Y(G679),.A(G89),.B(G678));
  OR2 OR2_126(.VSS(VSS),.VDD(VDD),.Y(G680),.A(G88),.B(G677));
  OR2 OR2_127(.VSS(VSS),.VDD(VDD),.Y(G682),.A(G681),.B(G699));
  OR2 OR2_128(.VSS(VSS),.VDD(VDD),.Y(G684),.A(G645),.B(G696));
  OR2 OR2_129(.VSS(VSS),.VDD(VDD),.Y(G687),.A(G686),.B(G699));
  OR2 OR2_130(.VSS(VSS),.VDD(VDD),.Y(G690),.A(G348),.B(G696));
  OR2 OR2_131(.VSS(VSS),.VDD(VDD),.Y(G691),.A(G645),.B(G689));
  OR2 OR2_132(.VSS(VSS),.VDD(VDD),.Y(G693),.A(G692),.B(G699));
  OR2 OR2_133(.VSS(VSS),.VDD(VDD),.Y(G697),.A(G180),.B(G696));
  OR2 OR2_134(.VSS(VSS),.VDD(VDD),.Y(G698),.A(G348),.B(G695));
  OR2 OR2_135(.VSS(VSS),.VDD(VDD),.Y(G699),.A(G658),.B(G712));
//
  NAND2 NAND2_0(.VSS(VSS),.VDD(VDD),.Y(G96),.A(G74),.B(G596));
  NAND2 NAND2_1(.VSS(VSS),.VDD(VDD),.Y(G97),.A(G75),.B(G596));
  NAND2 NAND2_2(.VSS(VSS),.VDD(VDD),.Y(G98),.A(G76),.B(G596));
  NAND2 NAND2_3(.VSS(VSS),.VDD(VDD),.Y(G99),.A(G77),.B(G596));
  NAND2 NAND2_4(.VSS(VSS),.VDD(VDD),.Y(G100),.A(G78),.B(G596));
  NAND2 NAND2_5(.VSS(VSS),.VDD(VDD),.Y(G106),.A(G107),.B(G110));
  NAND2 NAND2_6(.VSS(VSS),.VDD(VDD),.Y(G107),.A(G700),.B(G111));
  NAND2 NAND2_7(.VSS(VSS),.VDD(VDD),.Y(G122),.A(G123),.B(G126));
  NAND2 NAND2_8(.VSS(VSS),.VDD(VDD),.Y(G123),.A(G135),.B(G127));
  NAND2 NAND2_9(.VSS(VSS),.VDD(VDD),.Y(G137),.A(G138),.B(G141));
  NAND2 NAND2_10(.VSS(VSS),.VDD(VDD),.Y(G138),.A(G177),.B(G142));
  NAND2 NAND2_11(.VSS(VSS),.VDD(VDD),.Y(G163),.A(G164),.B(G167));
  NAND2 NAND2_12(.VSS(VSS),.VDD(VDD),.Y(G164),.A(G172),.B(G178));
  NAND2 NAND2_13(.VSS(VSS),.VDD(VDD),.Y(G186),.A(G187),.B(G190));
  NAND2 NAND2_14(.VSS(VSS),.VDD(VDD),.Y(G187),.A(G522),.B(G191));
  NAND2 NAND2_15(.VSS(VSS),.VDD(VDD),.Y(G205),.A(G206),.B(G209));
  NAND2 NAND2_16(.VSS(VSS),.VDD(VDD),.Y(G206),.A(G183),.B(G210));
  NAND2 NAND2_17(.VSS(VSS),.VDD(VDD),.Y(G211),.A(G212),.B(G215));
  NAND2 NAND2_18(.VSS(VSS),.VDD(VDD),.Y(G212),.A(G222),.B(G216));
  NAND2 NAND2_19(.VSS(VSS),.VDD(VDD),.Y(G230),.A(G234),.B(G235));
  NAND2 NAND2_20(.VSS(VSS),.VDD(VDD),.Y(G231),.A(G435),.B(G648));
  NAND3 NAND3_0(.VSS(VSS),.VDD(VDD),.Y(G232),.A(G296),.B(G298),.C(G435));
  NAND3 NAND3_1(.VSS(VSS),.VDD(VDD),.Y(G233),.A(G700),.B(G232),.C(G231));
  NAND2 NAND2_21(.VSS(VSS),.VDD(VDD),.Y(G234),.A(G649),.B(G436));
  NAND2 NAND2_22(.VSS(VSS),.VDD(VDD),.Y(G266),.A(G286),.B(G291));
  NAND2 NAND2_23(.VSS(VSS),.VDD(VDD),.Y(G267),.A(G287),.B(G292));
  NAND2 NAND2_24(.VSS(VSS),.VDD(VDD),.Y(G268),.A(G288),.B(G293));
  NAND2 NAND2_25(.VSS(VSS),.VDD(VDD),.Y(G269),.A(G284),.B(G294));
  NAND2 NAND2_26(.VSS(VSS),.VDD(VDD),.Y(G270),.A(G285),.B(G295));
  NAND2 NAND2_27(.VSS(VSS),.VDD(VDD),.Y(G284),.A(G45),.B(G104));
  NAND2 NAND2_28(.VSS(VSS),.VDD(VDD),.Y(G285),.A(G46),.B(G105));
  NAND2 NAND2_29(.VSS(VSS),.VDD(VDD),.Y(G286),.A(G42),.B(G101));
  NAND2 NAND2_30(.VSS(VSS),.VDD(VDD),.Y(G287),.A(G43),.B(G102));
  NAND2 NAND2_31(.VSS(VSS),.VDD(VDD),.Y(G288),.A(G44),.B(G103));
  NAND2 NAND2_32(.VSS(VSS),.VDD(VDD),.Y(G297),.A(G289),.B(G290));
  NAND2 NAND2_33(.VSS(VSS),.VDD(VDD),.Y(G298),.A(G297),.B(G700));
  NAND4 NAND4_0(.VSS(VSS),.VDD(VDD),.Y(G301),.A(G50),.B(G49),.C(G48),.D(G47));
  NAND2 NAND2_34(.VSS(VSS),.VDD(VDD),.Y(G331),.A(G333),.B(G22));
  NAND2 NAND2_35(.VSS(VSS),.VDD(VDD),.Y(G332),.A(G334),.B(G331));
  NAND2 NAND2_36(.VSS(VSS),.VDD(VDD),.Y(G476),.A(G486),.B(G616));
  NAND2 NAND2_37(.VSS(VSS),.VDD(VDD),.Y(G482),.A(G514),.B(G518));
  NAND2 NAND2_38(.VSS(VSS),.VDD(VDD),.Y(G483),.A(G515),.B(G519));
  NAND2 NAND2_39(.VSS(VSS),.VDD(VDD),.Y(G484),.A(G516),.B(G520));
  NAND2 NAND2_40(.VSS(VSS),.VDD(VDD),.Y(G485),.A(G517),.B(G521));
  NAND2 NAND2_41(.VSS(VSS),.VDD(VDD),.Y(G514),.A(G71),.B(G67));
  NAND2 NAND2_42(.VSS(VSS),.VDD(VDD),.Y(G515),.A(G72),.B(G68));
  NAND2 NAND2_43(.VSS(VSS),.VDD(VDD),.Y(G516),.A(G73),.B(G69));
  NAND2 NAND2_44(.VSS(VSS),.VDD(VDD),.Y(G517),.A(G487),.B(G70));
  NAND3 NAND3_2(.VSS(VSS),.VDD(VDD),.Y(G554),.A(G556),.B(G557),.C(G558));
  NAND2 NAND2_45(.VSS(VSS),.VDD(VDD),.Y(G555),.A(G559),.B(G560));
  NAND2 NAND2_46(.VSS(VSS),.VDD(VDD),.Y(G556),.A(G578),.B(G583));
  NAND2 NAND2_47(.VSS(VSS),.VDD(VDD),.Y(G557),.A(G579),.B(G584));
  NAND2 NAND2_48(.VSS(VSS),.VDD(VDD),.Y(G558),.A(G580),.B(G585));
  NAND2 NAND2_49(.VSS(VSS),.VDD(VDD),.Y(G559),.A(G581),.B(G586));
  NAND2 NAND2_50(.VSS(VSS),.VDD(VDD),.Y(G560),.A(G582),.B(G587));
  NAND2 NAND2_51(.VSS(VSS),.VDD(VDD),.Y(G578),.A(G79),.B(G74));
  NAND2 NAND2_52(.VSS(VSS),.VDD(VDD),.Y(G579),.A(G80),.B(G75));
  NAND2 NAND2_53(.VSS(VSS),.VDD(VDD),.Y(G580),.A(G81),.B(G76));
  NAND2 NAND2_54(.VSS(VSS),.VDD(VDD),.Y(G581),.A(G82),.B(G77));
  NAND2 NAND2_55(.VSS(VSS),.VDD(VDD),.Y(G582),.A(G561),.B(G78));
  NAND2 NAND2_56(.VSS(VSS),.VDD(VDD),.Y(G597),.A(G602),.B(G603));
  NAND2 NAND2_57(.VSS(VSS),.VDD(VDD),.Y(G598),.A(G435),.B(G83));
  NAND4 NAND4_1(.VSS(VSS),.VDD(VDD),.Y(G616),.A(G482),.B(G483),.C(G484),.D(G485));
  NAND2 NAND2_58(.VSS(VSS),.VDD(VDD),.Y(G700),.A(G282),.B(G283));
//
  NOR2 NOR2_0(.VSS(VSS),.VDD(VDD),.Y(G114),.A(G115),.B(G116));
  NOR2 NOR2_1(.VSS(VSS),.VDD(VDD),.Y(G115),.A(G133),.B(G25));
  NOR2 NOR2_2(.VSS(VSS),.VDD(VDD),.Y(G119),.A(G120),.B(G121));
  NOR2 NOR2_3(.VSS(VSS),.VDD(VDD),.Y(G120),.A(G134),.B(G26));
  NOR2 NOR2_4(.VSS(VSS),.VDD(VDD),.Y(G130),.A(G131),.B(G132));
  NOR2 NOR2_5(.VSS(VSS),.VDD(VDD),.Y(G131),.A(G136),.B(G28));
  NOR2 NOR2_6(.VSS(VSS),.VDD(VDD),.Y(G145),.A(G146),.B(G147));
  NOR2 NOR2_7(.VSS(VSS),.VDD(VDD),.Y(G146),.A(G168),.B(G30));
  NOR2 NOR2_8(.VSS(VSS),.VDD(VDD),.Y(G150),.A(G151),.B(G152));
  NOR2 NOR2_9(.VSS(VSS),.VDD(VDD),.Y(G151),.A(G169),.B(G31));
  NOR2 NOR2_10(.VSS(VSS),.VDD(VDD),.Y(G155),.A(G156),.B(G157));
  NOR2 NOR2_11(.VSS(VSS),.VDD(VDD),.Y(G156),.A(G170),.B(G32));
  NOR2 NOR2_12(.VSS(VSS),.VDD(VDD),.Y(G160),.A(G161),.B(G162));
  NOR2 NOR2_13(.VSS(VSS),.VDD(VDD),.Y(G161),.A(G171),.B(G33));
  NOR2 NOR2_14(.VSS(VSS),.VDD(VDD),.Y(G194),.A(G195),.B(G196));
  NOR2 NOR2_15(.VSS(VSS),.VDD(VDD),.Y(G195),.A(G202),.B(G37));
  NOR2 NOR2_16(.VSS(VSS),.VDD(VDD),.Y(G199),.A(G200),.B(G201));
  NOR2 NOR2_17(.VSS(VSS),.VDD(VDD),.Y(G200),.A(G203),.B(G38));
  NOR2 NOR2_18(.VSS(VSS),.VDD(VDD),.Y(G219),.A(G220),.B(G221));
  NOR2 NOR2_19(.VSS(VSS),.VDD(VDD),.Y(G220),.A(G223),.B(G41));
  NOR2 NOR2_20(.VSS(VSS),.VDD(VDD),.Y(G238),.A(G239),.B(G240));
  NOR2 NOR2_21(.VSS(VSS),.VDD(VDD),.Y(G239),.A(G299),.B(G42));
  NOR2 NOR2_22(.VSS(VSS),.VDD(VDD),.Y(G243),.A(G244),.B(G245));
  NOR2 NOR2_23(.VSS(VSS),.VDD(VDD),.Y(G244),.A(G262),.B(G43));
  NOR2 NOR2_24(.VSS(VSS),.VDD(VDD),.Y(G248),.A(G249),.B(G250));
  NOR2 NOR2_25(.VSS(VSS),.VDD(VDD),.Y(G249),.A(G263),.B(G44));
  NOR2 NOR2_26(.VSS(VSS),.VDD(VDD),.Y(G253),.A(G254),.B(G255));
  NOR2 NOR2_27(.VSS(VSS),.VDD(VDD),.Y(G254),.A(G264),.B(G45));
  NOR2 NOR2_28(.VSS(VSS),.VDD(VDD),.Y(G256),.A(G257),.B(G261));
  NOR2 NOR2_29(.VSS(VSS),.VDD(VDD),.Y(G257),.A(G265),.B(G46));
  NOR3 NOR3_0(.VSS(VSS),.VDD(VDD),.Y(G289),.A(G270),.B(G269),.C(G268));
  NOR2 NOR2_30(.VSS(VSS),.VDD(VDD),.Y(G290),.A(G267),.B(G266));
  NOR2 NOR2_31(.VSS(VSS),.VDD(VDD),.Y(G299),.A(G301),.B(G328));
  NOR2 NOR2_32(.VSS(VSS),.VDD(VDD),.Y(G327),.A(G330),.B(G23));
  NOR2 NOR2_33(.VSS(VSS),.VDD(VDD),.Y(G328),.A(G329),.B(G327));
  NOR2 NOR2_34(.VSS(VSS),.VDD(VDD),.Y(G361),.A(G362),.B(G363));
  NOR2 NOR2_35(.VSS(VSS),.VDD(VDD),.Y(G362),.A(G523),.B(G51));
  NOR2 NOR2_36(.VSS(VSS),.VDD(VDD),.Y(G366),.A(G367),.B(G368));
  NOR2 NOR2_37(.VSS(VSS),.VDD(VDD),.Y(G367),.A(G375),.B(G52));
  NOR2 NOR2_38(.VSS(VSS),.VDD(VDD),.Y(G369),.A(G370),.B(G374));
  NOR2 NOR2_39(.VSS(VSS),.VDD(VDD),.Y(G370),.A(G376),.B(G53));
  NOR2 NOR2_40(.VSS(VSS),.VDD(VDD),.Y(G380),.A(G381),.B(G382));
  NOR2 NOR2_41(.VSS(VSS),.VDD(VDD),.Y(G381),.A(G183),.B(G54));
  NOR2 NOR2_42(.VSS(VSS),.VDD(VDD),.Y(G385),.A(G386),.B(G387));
  NOR2 NOR2_43(.VSS(VSS),.VDD(VDD),.Y(G386),.A(G394),.B(G55));
  NOR2 NOR2_44(.VSS(VSS),.VDD(VDD),.Y(G388),.A(G389),.B(G393));
  NOR2 NOR2_45(.VSS(VSS),.VDD(VDD),.Y(G389),.A(G395),.B(G56));
  NOR2 NOR2_46(.VSS(VSS),.VDD(VDD),.Y(G398),.A(G399),.B(G400));
  NOR2 NOR2_47(.VSS(VSS),.VDD(VDD),.Y(G399),.A(G335),.B(G57));
  NOR2 NOR2_48(.VSS(VSS),.VDD(VDD),.Y(G401),.A(G402),.B(G406));
  NOR2 NOR2_49(.VSS(VSS),.VDD(VDD),.Y(G402),.A(G412),.B(G58));
  NOR2 NOR2_50(.VSS(VSS),.VDD(VDD),.Y(G409),.A(G410),.B(G411));
  NOR2 NOR2_51(.VSS(VSS),.VDD(VDD),.Y(G410),.A(G413),.B(G59));
  NOR2 NOR2_52(.VSS(VSS),.VDD(VDD),.Y(G417),.A(G418),.B(G419));
  NOR2 NOR2_53(.VSS(VSS),.VDD(VDD),.Y(G418),.A(G358),.B(G60));
  NOR2 NOR2_54(.VSS(VSS),.VDD(VDD),.Y(G420),.A(G421),.B(G425));
  NOR2 NOR2_55(.VSS(VSS),.VDD(VDD),.Y(G421),.A(G431),.B(G61));
  NOR2 NOR2_56(.VSS(VSS),.VDD(VDD),.Y(G428),.A(G429),.B(G430));
  NOR2 NOR2_57(.VSS(VSS),.VDD(VDD),.Y(G429),.A(G432),.B(G62));
  NOR2 NOR2_58(.VSS(VSS),.VDD(VDD),.Y(G442),.A(G443),.B(G444));
  NOR2 NOR2_59(.VSS(VSS),.VDD(VDD),.Y(G444),.A(G615),.B(G64));
  NOR2 NOR2_60(.VSS(VSS),.VDD(VDD),.Y(G452),.A(G453),.B(G454));
  NOR2 NOR2_61(.VSS(VSS),.VDD(VDD),.Y(G454),.A(G615),.B(G66));
  NOR2 NOR2_62(.VSS(VSS),.VDD(VDD),.Y(G460),.A(G461),.B(G462));
  NOR2 NOR2_63(.VSS(VSS),.VDD(VDD),.Y(G461),.A(G434),.B(G67));
  NOR2 NOR2_64(.VSS(VSS),.VDD(VDD),.Y(G465),.A(G466),.B(G467));
  NOR2 NOR2_65(.VSS(VSS),.VDD(VDD),.Y(G466),.A(G479),.B(G68));
  NOR2 NOR2_66(.VSS(VSS),.VDD(VDD),.Y(G470),.A(G471),.B(G472));
  NOR2 NOR2_67(.VSS(VSS),.VDD(VDD),.Y(G471),.A(G480),.B(G69));
  NOR2 NOR2_68(.VSS(VSS),.VDD(VDD),.Y(G473),.A(G474),.B(G478));
  NOR2 NOR2_69(.VSS(VSS),.VDD(VDD),.Y(G474),.A(G481),.B(G70));
  NOR3 NOR3_1(.VSS(VSS),.VDD(VDD),.Y(G487),.A(G71),.B(G72),.C(G73));
  NOR2 NOR2_70(.VSS(VSS),.VDD(VDD),.Y(G527),.A(G528),.B(G529));
  NOR2 NOR2_71(.VSS(VSS),.VDD(VDD),.Y(G528),.A(G604),.B(G74));
  NOR2 NOR2_72(.VSS(VSS),.VDD(VDD),.Y(G532),.A(G533),.B(G534));
  NOR2 NOR2_73(.VSS(VSS),.VDD(VDD),.Y(G533),.A(G550),.B(G75));
  NOR2 NOR2_74(.VSS(VSS),.VDD(VDD),.Y(G537),.A(G538),.B(G539));
  NOR2 NOR2_75(.VSS(VSS),.VDD(VDD),.Y(G538),.A(G551),.B(G76));
  NOR2 NOR2_76(.VSS(VSS),.VDD(VDD),.Y(G542),.A(G543),.B(G544));
  NOR2 NOR2_77(.VSS(VSS),.VDD(VDD),.Y(G543),.A(G552),.B(G77));
  NOR2 NOR2_78(.VSS(VSS),.VDD(VDD),.Y(G545),.A(G546),.B(G549));
  NOR2 NOR2_79(.VSS(VSS),.VDD(VDD),.Y(G546),.A(G553),.B(G78));
  NOR4 NOR4_0(.VSS(VSS),.VDD(VDD),.Y(G561),.A(G79),.B(G80),.C(G81),.D(G82));
  NOR2 NOR2_80(.VSS(VSS),.VDD(VDD),.Y(G593),.A(G435),.B(G524));
  NOR2 NOR2_81(.VSS(VSS),.VDD(VDD),.Y(G599),.A(G598),.B(G597));
  NOR2 NOR2_82(.VSS(VSS),.VDD(VDD),.Y(G660),.A(G658),.B(G86));
  NOR2 NOR2_83(.VSS(VSS),.VDD(VDD),.Y(G681),.A(G683),.B(G660));
  NOR2 NOR2_84(.VSS(VSS),.VDD(VDD),.Y(G686),.A(G688),.B(G660));
  NOR2 NOR2_85(.VSS(VSS),.VDD(VDD),.Y(G692),.A(G694),.B(G660));
  NOR4 NOR4_1(.VSS(VSS),.VDD(VDD),.Y(G703),.A(G650),.B(G651),.C(G652),.D(G653));
  NOR2 NOR2_86(.VSS(VSS),.VDD(VDD),.Y(G708),.A(G709),.B(G710));
  NOR2 NOR2_87(.VSS(VSS),.VDD(VDD),.Y(G710),.A(G678),.B(G94));

endmodule