module s9234(g6360,g89,g4307,g560,g6282,g4422,g6370,g559,g306,g301,g319,g98,g2584,g6372,g6366,g6362,g558,g102,g5137,g5692,g5469,g4809,g3600,g3222,g564,VDD,g561,g5468,g6374,g107,g6728,g6284,g705,g6368,g563,VSS,g557,g6364,g4321,g310,CLOCK,g314,g562,g94);
input g89,g560,g559,g306,g301,g319,g98,g558,g102,g564,VDD,g561,g107,g705,g563,VSS,g557,g310,CLOCK,g314,g562,g94;
output g6360,g4307,g6282,g4422,g6370,g2584,g6372,g6366,g6362,g5137,g5692,g5469,g4809,g3600,g3222,g5468,g6374,g6728,g6284,g6368,g6364,g4321;

  wire g285,I2464,g6367,g3333,g4181,g1076,g2896,g4129,I3310,g3462,I3596,I6587,g4657,I7007,I7478,g5637,g3964,I2327,g2656,I5195,g2672,I3843,I8872,g5500,g938,g6048,g5444,I2196,g286,I2620,g2883,I2137,g6838,g3353,g4810,g4210,I3890,g6264,g3042,I7541,g3853,g6103,g6114,I8597,g2796,g3744,I5692,g3626,g4407,g4392,I3452,g2809,g4792,g3520,g2604,g6376,g4493,g6070,I3972,I9143,I2890,g5550,g6469,I7209,g2497,g3859,g6704,g5197,I4513,I6473,g606,g1176,g47,g3931,g5121,g3785,I6185,g5448,I5264,I8834,I4273,I7251,I7969,I9059,I3990,g6236,I2442,I2570,I7517,g5135,g3029,I6745,g6889,I3395,g1011,g4126,g6604,g2905,I9052,g2829,I7472,g5024,I6599,g3884,g1829,g5274,g1603,g6537,g4585,g6353,g2056,g2895,g4622,I8854,g3186,I2460,g2768,g1375,g901,g2092,g3880,I5536,g370,I2802,g2172,g3793,I3040,g1902,I5938,I4465,g6799,I5040,I6196,I5457,g84,g74,g1643,g1960,I7640,I8377,g4355,g1576,g3995,g6782,g5164,g4438,g5010,g1756,g4501,I3614,g2701,g6718,g3891,g2887,g2179,g3182,g6697,g2039,g3276,g2903,g6893,g1761,I6359,I8582,g5430,I6078,g4233,g1586,I5910,g791,g5602,g6055,g6342,I8535,g3014,g123,I4252,I8411,g6706,I8860,g5351,I2284,g1256,g2137,I6537,g6455,g695,g6713,I2182,I6812,g5878,I2845,g1037,I5214,g3383,g4370,g5727,g666,g1966,g1416,I8473,g5912,I3215,g5403,g3890,I5360,I2745,g2916,I6661,g122,I8329,g3219,I3047,g6842,I3681,I2306,g4713,I2169,I7035,g4222,g4943,g2330,g3700,g6150,I3251,I2899,g2923,g3761,g3718,g5251,g2080,I1844,I2073,I3717,g6509,I3773,g4424,g3143,g1578,g6254,I5124,I3711,g4767,g6792,I7107,g361,I8690,g4098,I9113,g5952,I5885,g1567,I8857,g5521,g5753,I7119,g6739,g4344,g6348,I7237,g6073,g5236,I5644,g386,g3998,g4360,I7978,I5490,g3953,I2125,g4164,I2293,g3790,g6708,g5598,I5006,I5731,g1088,g6774,g6182,g2747,I2072,g1378,g2650,g2981,g1683,I3127,g2598,I6366,g4428,g3725,g3616,I5766,g3037,g402,I6740,g6489,I8518,g2877,g6517,g6492,g6478,I2204,g2861,g4373,I2296,g965,g3239,g3,I5227,g2576,g111,g2586,I4282,g798,g5672,I8764,g1449,I4809,g6120,g6890,g3028,g45,g2802,I2405,I2491,I8809,g2814,g4517,I8863,g6851,g3668,I2767,g5372,I4243,g4848,g4188,I5454,g4801,I2352,g4017,g1355,g4131,I3028,I3714,I7536,g2734,I5430,g6554,g5451,I8379,I7686,g1852,I2831,g5052,I3155,g804,I3522,I7086,g5491,I2402,I8730,g6837,I4192,g4455,g4706,g654,g3031,g1975,I6289,I7643,g1276,g2738,I8500,I5403,g6682,I6247,g4841,g3778,g2612,g1777,g861,I7372,I2982,g328,g2134,g2867,g5939,I1979,g4114,g932,I5301,g6506,I5640,g1317,g1963,I7698,I8713,I6959,g2256,I5562,g2886,g6938,g5145,g6709,I8211,g3860,g349,g1928,g5310,I4477,g4400,I1847,g4364,g4363,g1620,I3349,g6847,I6448,g3608,I6567,g4707,g1474,g5484,g856,I8335,g4721,g4800,g1762,I6660,g4003,g5493,g5895,g2857,g2582,I3540,g3361,g4662,g4401,I7097,I5300,g6135,I9176,g5169,g2264,g6797,g3287,g3847,g2699,g6910,g3234,g2706,g3448,g4375,g1205,g4840,g3073,g4404,I2760,g2927,g3489,g4580,g4156,g131,g5638,g3354,g3425,g10,g1056,g4673,I2394,g2360,g5358,I9008,g1337,I1970,I3502,g2838,g5395,g3662,g1114,I5187,g3666,g3076,I6081,g4589,I7223,g2860,g5122,I7543,I3635,g2506,g6099,I6573,g2975,g2079,g6824,g5742,g4399,g4492,g6094,g710,g5148,I4312,I1877,I6989,g6653,g288,g4458,I5081,I5484,g2807,g6601,I3989,g926,g3997,g6647,g4362,I2860,g4946,g6508,I5768,g3840,I2343,g6483,I2940,g5429,I5243,I8110,g6473,g207,I2445,g2136,g2029,g4569,g4272,g3365,g3356,g6466,g6272,I5343,g5309,g1946,g6796,g5022,I7245,I1953,g6327,I2014,I5376,g4685,g6565,g4631,I3445,g4112,g3296,g1577,g3835,I4527,g5880,g5439,g5116,g6655,g2081,g1988,g4507,g3135,g3522,g5480,g242,g5872,g6906,g2875,g5331,I8432,g119,g2524,I6012,g4836,g2509,g5900,g3537,g366,g6253,g5364,g1203,g6403,g2864,I3556,g6043,g1665,g3486,g1046,g4719,I8367,g3095,g1315,g2858,g4487,g1978,I2992,g683,I3816,I8638,g1633,g4242,I3953,I3954,g4715,g4756,g4560,g685,I8749,g2675,I2681,I8978,g3123,g5060,I7571,g1110,g2959,I8721,g1054,g6116,I8981,I8806,g5250,g3212,g638,g6134,g3346,I5944,I3840,g6310,g3085,g3935,I2995,I2287,g5470,g5088,I7254,g206,g4433,g5557,g3500,g5225,g1692,g6108,g4168,g3783,g3858,I3569,I2854,I2919,I8659,I4161,g3928,I6630,g2283,g4445,g2995,I3935,g4789,g6520,I5148,g2434,g5497,I7587,g1645,I5307,g3740,g5083,I8727,g4231,g6843,g2870,I5445,g675,g6344,g478,g4403,g5496,I6051,g5697,g2625,I7264,I6308,I6962,g3225,g6056,g1407,g2242,g2904,g5683,g6596,g193,g5467,I9131,g6572,I1862,I6499,g941,I2958,I8891,I4507,g5273,I2724,g6467,g11,I2735,I7555,g3963,g6418,I2883,g5043,I7469,I5933,g6416,g4452,g2177,g4837,I2110,g5751,g4346,g551,g679,g5729,g4950,I5068,g6923,g6786,g1831,g1143,g3457,g4785,g5662,g6518,g5167,g6535,g5077,g152,g38,g3360,I2147,g5180,g2746,g1972,g3317,g6707,g2340,I7295,I4152,g6142,I2753,g4372,I5463,g6877,g3750,I7811,I5448,g1541,g3781,g4434,g1837,g2018,g3797,g3911,g4783,g5231,g6428,g2874,I5496,g680,g4139,g204,I3105,I6783,g3976,g5089,g2792,g1384,g4354,I8346,g5278,g2808,g1646,g6445,g6465,g5323,g6620,g5291,I9137,g5562,g3652,I5736,g1285,I2617,g4292,I6250,g5593,I6789,I6927,I8385,I8626,I7980,g4856,g4702,I5542,g5382,g5569,I6075,I3446,g14,g1345,g6599,g2174,g5996,g6875,g682,g6479,g508,I4166,g6235,g6512,I5252,I8476,I2828,I8635,g3701,g6262,g6612,g4011,I2082,I5879,g5246,I5594,g345,g4613,g4051,g4246,I5094,g6039,g4280,I5394,g6357,g5888,I8195,I2388,g2491,g6600,I4961,g5068,g5154,I3206,g1656,g341,g1847,I5904,g4221,g3869,I3334,g2107,I3509,I2050,I5316,g4626,g5062,I3102,I2361,g4658,g2787,g4393,g6932,I2614,I4964,g5691,g6298,g3512,g69,g5946,g5494,g844,g3053,g6823,g4241,I7596,I7176,g6125,g5087,I3255,g4629,g2789,g3714,I6733,g6715,g5994,g3645,g5433,g3511,I5998,g5217,g4166,I6625,I8984,I8290,g1584,g5660,I8818,I8044,g6676,g3127,g6665,g5157,I5259,g4214,g1305,g6605,g3796,I3590,I3499,I6292,g1918,g5879,g2254,g3848,I6318,g4832,I2476,I7604,g6371,I9005,g1232,g3040,I8189,g5471,I8417,I5577,g4647,I3733,g3765,g6933,g1471,g3117,g2890,g4530,g5902,g5695,I6417,I8359,I5526,I5433,g851,g3641,g6084,g6339,g5475,I7439,g6424,g2996,g6500,g5149,I7193,g2464,g1935,g4229,g6720,I2795,I8541,g2728,I7153,I7522,g4440,I3927,g2095,g6341,g6836,I4327,g3370,g1787,g4448,g686,g5702,g5800,I2925,g1575,I3999,I5568,g6280,I6464,g5601,I8603,g4223,g642,g6585,g6453,g5016,g5808,g5775,g5626,I8255,I3697,g2920,g5066,g4586,g4802,g4515,g3902,g6593,g5587,I9217,g2821,g5685,g5527,I4976,g2781,g5908,g6454,I3115,g2078,g3745,g3622,g6287,g6864,g3349,g6722,I8120,I2330,I3902,I7534,I2716,I7397,g5486,g4659,g4525,g4628,I5857,g3369,g4900,I7608,g4356,g6486,g6631,g4449,g1936,g2865,g4182,g59,g4228,I5890,g4220,g1335,g1556,g2164,I5056,g5992,g2267,g4646,g4352,I5532,g6433,I2143,I1952,I8840,I5228,I9082,g625,g2772,g6438,g4739,g3060,g5226,g3207,g4441,g6498,I6084,g6415,g6159,I8347,I5657,I2700,I2057,g5813,g4224,g4320,g2913,g5951,g3351,g1550,g3690,g3491,g5784,g931,g2997,g1318,g4048,g586,I5002,g5809,g839,g5866,g4865,g6130,g4111,I2301,I5923,g3015,I4133,g2535,I6621,I7583,g4293,g873,g3521,g4526,I9140,I2221,g5941,g2685,g698,I3895,g5025,g4615,g6351,I5385,g6695,g4104,g2117,g2755,g893,I3868,g5723,g5877,I3431,g4838,g5142,g1279,I2044,I8089,I3650,g5316,g4227,I3528,g5048,g114,g6337,g6285,g4461,g1805,g6849,g4342,I8276,I5379,g4854,I5896,g4740,I7077,g2764,I2023,I7231,g2947,g1070,g5377,g6077,g5049,g289,I8758,I4217,I5511,g2004,I2521,I3593,g3079,g3870,g4161,g485,g1772,g1327,g2086,I5359,I2272,g4388,g3328,g3170,g3756,g5406,g2138,g3654,g5477,I6528,I3080,g5234,g5209,g4850,g3593,g3531,g4559,g5350,g1776,I4009,g3183,g6578,g6069,I2485,g1253,g1919,g5363,I3608,g3331,g6892,g6323,g1835,g5069,g5086,I7838,g5953,g574,I5987,I6066,g3315,I6187,g4328,g6768,g4701,I3971,g4639,g3528,g5447,g2765,g4202,g4074,I2367,I2749,I3271,I6324,g6143,g1820,g5544,I5600,g3372,I2544,I3177,g2933,g2346,I3965,g5524,g4178,g2312,I6801,g6176,g2647,I3493,g4494,g1725,I7361,I9134,g1703,g3843,g276,g5922,g1609,g5233,I6546,g2820,I8128,I5537,g357,I8576,g4844,g3669,g5773,g3380,g6119,I9158,I6564,I3611,g5817,I6659,g6128,g5061,g6887,g2924,g2839,g1730,g5328,g3844,g4140,I1924,g5090,g5054,g3973,I4233,g6673,g3653,g3598,I3278,g2085,I6114,g4456,I8674,I5783,g5576,g5541,g4591,g1887,g3697,g6651,g1979,g3302,I3581,g2440,g3660,g1177,I2814,g1842,I3388,g5219,g2782,g3575,g4590,I6437,g3043,g3748,g6712,g5383,g1348,g3688,I9044,g4001,I7528,I7966,g774,g6185,I5743,g3263,I4623,g4793,g2435,g6515,g3378,I6737,g5627,g2113,g4708,I5760,g6762,g5599,I7039,I2358,g3727,g1042,g6212,g5230,g6918,I3874,g2609,g2104,g843,g422,g3914,g784,g4016,g430,I4019,g4353,g1806,g6743,g4052,I5699,g4871,g2044,g4670,g2974,g2171,g5659,I4183,g1341,g6831,g5354,I5612,g4614,I6108,g3109,I7029,I8295,g4609,g709,g1001,I7704,I6087,g6303,g872,g5111,g5269,I5840,g5210,g3171,g2846,I6036,g6614,g4870,g2195,g3459,g3719,I5523,I2574,g3499,g3483,g6534,g6661,g6679,I4198,g6412,I3970,g6648,I2212,g1740,g3228,g6732,I7578,g3329,g6559,g1470,I2970,I2773,g6015,I5793,g6074,g5370,I3212,g6527,g1254,g4250,g5917,g3238,g3904,I4351,I7042,g2585,I2630,g5901,I5556,I7865,g3440,g6193,I9203,I2671,g6652,g2940,g5954,I2033,I5759,I4414,g5190,g4584,I6311,g5456,I7707,g4236,I8716,I5920,I5023,g4603,I3152,I8348,I8127,g1585,g5636,g1997,I3099,g5506,g3967,g1542,g5046,g4368,g2443,g6496,g6555,g4536,g414,I2128,g6929,g3798,I3662,g4683,g5646,g6266,I3894,I5037,I3988,I5481,g5864,g6841,g4128,I6015,I5244,g766,I8665,g5572,g6429,g1699,g4851,I3629,I6570,g6158,g5174,g4936,I7963,I2683,I4291,g3779,I3247,g2575,I3776,g2009,g5680,g4769,g1274,g6553,I3644,g5375,g3301,g3320,g5852,g4777,I2537,I5019,g6909,g1815,g6152,I7829,g1953,I2246,g36,g3284,g4276,I4671,g665,g4775,I3481,g4516,g4610,g668,g6242,I8264,g3810,g6529,g6741,g205,I6343,I3400,I8203,I2887,g3209,g3368,I2417,I2797,g4587,g5095,g4302,g3452,g6336,g6588,g3936,g6902,g2804,g4134,g2885,g3801,g1781,I3428,I8267,I6986,g1998,g6273,g4868,g4712,g3289,g6586,g3872,g1117,g4860,I2785,g1982,I8168,g1038,g6167,g282,g905,g4308,g2512,I6576,I9220,I9098,g3887,I3534,I9085,g3983,g2025,g4385,g6781,g3490,I3767,I3328,I5893,I5774,g6288,I3871,I7358,g6325,I6026,g2780,I8174,I9116,g917,g4032,g4830,I6305,g3465,I8462,g3702,g4568,g5926,g6769,I3109,g2135,I5756,g3857,I3284,g3603,g6736,g3541,g3850,g662,I2581,I4526,g6912,g1415,g4387,g3925,g3940,I9164,g5399,g5163,g4915,g209,g1331,I2973,g5629,g6616,I5418,g3777,I3961,g5349,I2675,I5257,I6474,I2037,g5958,g4127,g667,g3204,I7562,g5085,g3830,g2265,g5248,I6552,I3144,g6730,g2089,g4117,g4132,g3854,g3382,I8040,I5790,g6911,I3179,I2811,I8441,g3955,g6088,I6400,g5449,I6976,g6090,g2841,g2793,g5265,g5590,g6855,g3525,g4623,I2278,I3010,I6410,g5570,g5997,I7239,I7433,g3388,g5681,g3927,g6561,g3559,I3307,g1284,I7146,I8527,g6714,g4561,g6113,I7270,I5649,g894,g2041,g3618,g4524,g3505,g5432,g4490,I3462,g2753,g3723,I2346,g3842,g6657,g6068,g3984,I2228,I5258,g496,I4757,g3968,g3991,I6769,g5425,g6332,g2263,g622,I4437,g4179,g6800,I5907,g4612,g829,g706,g6845,I8567,I3074,I3391,g838,I6612,I3031,g5453,I8662,I2244,g3977,I3575,g4333,g1340,g4050,g6067,I8357,I6139,g1845,I4229,I8261,g1287,g1640,I6001,g5498,g254,g4781,I6666,g6117,g2042,g5178,g1372,g4382,g1661,I3602,I2140,g1950,I2635,g850,I4010,g5947,g4949,I3694,g1695,I3126,I5648,I3361,g6649,I4182,g6345,g3876,g5777,g5144,g1477,I3288,g837,I4003,g4942,g6656,g4158,g1642,g5325,g939,I7230,I2588,g4038,g4866,I6763,g1334,I3399,g6829,I5439,I5271,g6457,g6365,I8243,g1647,I9236,g3952,g4120,I8800,I2172,g248,g2068,I5478,g1563,I3337,g6440,I6759,g6913,g5455,g281,I4547,g5191,I8369,I6923,I8258,I6346,g28,I7805,I2731,I4324,g4405,I5460,g331,g6358,g6425,g3441,g5189,g5152,g4319,g3956,g382,g4446,g6156,g3746,g4234,I4160,g297,I3946,g5295,I5493,g6385,I6444,g1394,g6314,g4171,g6693,g6907,g4654,g2960,I6403,g5821,g3291,I3379,I8994,g3729,g6719,g6450,I7989,g6283,g6640,I2382,g5678,I8081,g6898,g6148,g5938,g4045,g4813,g3224,g3567,g6426,g2308,g4049,g3288,g6411,I3906,g6691,g4700,g406,g1624,I6677,I9110,g6065,I3364,g6936,I6680,g3485,g4447,g291,g3731,g6822,g5415,g2931,g5140,g1755,g5490,g4731,g2276,g4286,g4620,g2066,I7563,I6488,g1797,I2081,g4687,g5679,g2324,g15,g4744,g2433,g4215,g4351,I9038,g1880,g3929,g5454,g4439,g3140,g6507,g2769,g5694,I7808,g5658,I7497,g4192,g5515,g2059,g6319,g4833,g578,I1841,I1986,g5162,I4382,g1710,g1687,I6949,g5919,g1792,g6589,g6525,g5357,I1917,I4903,g3479,g6089,g1588,I3669,I4452,I5647,g6729,g5369,g2827,I6060,I8617,g3332,I2763,g6317,g2986,g2175,g3866,g3878,g949,I7143,g3759,g148,g3424,g4864,g5138,g1636,I4420,I6646,g6669,I3134,I3434,g4133,g5299,I7987,g3232,I7972,g1059,g1540,g6595,g2121,I3090,g5915,g2101,g6407,g3942,g3621,I5746,g2067,I5843,I3235,g5235,g4762,g1914,I9011,g6485,g6582,I7509,I4501,g1560,I2041,g5445,I7481,g6516,g6621,g5200,I5871,g6852,g2671,g4699,g6312,g6903,I4516,g6888,g3961,g6497,g6275,g3766,g3865,g1352,I8349,g1686,g4348,g4621,g2090,g6566,g79,g4057,g4339,I5209,g4806,g2700,g4464,I4919,g5824,g6346,g2806,g2111,g5942,g948,g6767,g5053,g598,g1748,I3638,g6299,I4306,I2185,I2411,g2470,I5091,g2745,g4426,g6087,g6461,I3914,I3659,I5761,g4486,g6141,g4550,g5504,I2004,g3376,g6818,I5030,g5147,g4101,g3259,g3980,g3693,g5559,g4430,g2663,g4152,I6543,g4784,g1048,g4794,g4873,I6028,g2118,I2542,g536,g908,I4294,I8056,g4773,g4914,g3898,I3465,g118,g3630,I7065,g6785,g5812,g5578,g749,I8150,g5705,g3615,g1157,g6583,g6501,g3814,g1685,g6625,g4723,I5337,g3166,g4261,g830,I2376,g5431,g4834,I1947,g3063,I9065,I5603,I2499,g6334,g4396,I2231,g3913,g1690,g4235,g5502,g4816,g3090,g1189,g4007,g6846,I3158,g3846,I2507,g1875,g4277,g4109,g6252,g3451,g4855,I5103,g3300,g5374,I5475,g4437,g1675,g3357,I7475,I3455,g6590,g6295,g6716,g4910,I3086,I8156,g6920,I4297,g516,I6406,g4593,g5172,I7352,g184,I6390,g2353,g1732,I1988,g2315,g2603,g4010,g4500,g6615,g4135,I7051,I8144,I2498,g1808,g6735,g2957,I2943,g5993,g5115,g2036,g1594,g2105,I5825,g3679,I9050,I8202,g6278,g2909,I3268,I3983,g2936,g6417,g2937,g5438,I4492,g1743,g4624,g4967,g6352,I4587,I1938,I1874,g4617,g6502,g3710,I6020,g834,I9182,I8147,I6795,g4146,g5378,g5266,g4130,I2779,I8137,g374,g1659,I8966,g2574,g2962,g2060,g3807,g1,g4760,g6558,g5379,I3623,g1564,g5064,g5770,g6033,g4123,g3820,g2293,g3464,g895,g3379,g2951,g4172,g5367,g5944,g1623,g5428,g2446,I3752,I8693,g1528,g5227,I3053,I2897,g5647,g6721,g6493,g500,g5955,g6361,g6394,I4279,I8093,g5443,I7311,g1985,I4285,I4410,I6315,g5317,I9146,g2580,g6658,g3086,g3158,g6806,g3134,g2709,g3672,g280,g3325,g4173,g3052,g4473,g2835,g2739,g4686,g5899,I5226,g3886,g3921,g4667,g43,I3376,I5106,g1814,g5202,g4718,I4799,g1336,g6315,I2653,g2367,g2156,I2910,g4791,I2986,g4937,g4504,g6147,I7451,g1192,g4124,I3782,I5421,g3297,g3772,I2005,I7692,g6255,g1917,g6737,I1962,g4039,g2643,g3855,I2608,I4347,g3551,g2169,g6244,g3307,g6144,g1289,g2594,g3861,g48,g3502,I4939,g3203,g5605,g5783,g3162,g5063,g4814,g2618,g4206,g5292,g1825,g5435,g6613,g6526,g2688,g677,g3339,I2674,I3025,I2015,g4432,I6792,g5950,g4829,I8591,I4023,g631,g5281,I3488,g6524,g6904,I6195,I6069,g2634,I2768,I4920,g4397,g2170,g6442,I1963,I3587,g4247,g6375,g2760,g2686,g6710,g862,g1419,g6258,g3306,g6567,g1351,g4495,I4480,I5084,g1502,g5474,I8030,I5696,I7484,g2836,I5520,I3830,g1583,g1220,g3074,g4523,g2024,I7098,g2515,g236,g4389,I4159,g2356,g2679,g2108,I7440,g1111,I6972,I5415,g1006,I2788,g6230,I8358,g3167,g6598,g3726,g6194,I3004,g3532,g6107,g1824,I8485,g3324,g3699,I8821,I3037,g5682,I2913,I7349,g5492,g6302,g2163,I3168,g3784,g1118,g1344,I7217,I7170,I6995,g378,I5436,g4443,I8656,g5418,g5376,g2295,g4046,I6895,I8632,g4608,g4080,g5898,g4199,g6556,g3974,I2648,g2159,g6404,g6557,I2473,g6803,g528,g809,g6624,g426,g3144,g3104,g6131,g6545,g5308,g1123,g1782,I4249,I8345,g2381,g1249,g5571,g6373,g943,g5635,I2596,I7466,g4465,g3852,g2485,g2142,I3016,I4593,g4499,I2190,g3832,g64,g6645,I8724,g3957,g2872,g6577,g4599,I7979,g1174,g3334,g4334,I5078,I3496,g4666,g6240,I6495,g6874,g980,g4427,g3118,g4033,I6072,g1649,I4234,g6876,I9233,g5479,g4980,g5327,I1980,I2300,I2199,I6780,g4099,I3298,g1841,g5466,I8943,g5360,g5687,g2327,g3892,I3373,g1570,g6066,g6564,I4681,I5686,I7333,g2457,g3698,g4485,g5568,g4872,g4459,g2538,g5483,g1338,I8183,g6347,g2430,I6352,g1853,g2053,g4322,g3338,I2638,I3811,g2968,g743,g3161,I5197,g1387,g4350,g1593,g3966,I9185,g6901,g1854,g1052,g6243,g6733,g1655,I5514,g4059,g6646,g2868,g5774,g4151,g1481,g672,I8438,I6337,g1573,I7055,I2029,g1119,g3677,I6649,g2914,I4123,I4468,I7167,I4921,I3304,I5535,g4488,g3638,I6531,g492,I5952,g5957,g2,g3667,g3322,g2103,g2712,g2731,g4471,I3331,I6280,g4435,g6879,g910,g3023,I8368,I5831,g5508,g4578,g4565,I4184,g6499,g3057,g1060,g4047,I2370,g6896,g42,I8332,g5688,g4054,g5903,I9057,g4514,I2315,g3223,g4451,g1905,g5538,g2720,g3868,g6304,g1711,I7576,g4022,g6538,g4717,I6579,I4528,g4645,I3189,g2758,g3013,g2640,I6692,I8034,g5616,I5622,g5671,g2894,g1094,g2591,g3246,I8066,g1027,g4436,g5869,g2664,g6106,I3340,g3875,g3237,I1838,g4037,g619,g3841,g692,g2158,g6109,I8136,g1473,g6173,I8444,g2488,g2908,g1101,I6706,g6146,g6488,g3001,I8884,I2663,I6302,I8866,g3816,g4757,g3838,g1660,g6522,g4671,I8002,I8153,g6734,g4116,g398,I1825,g4106,g4270,g4541,g4271,g1716,I5545,g845,g5184,g4693,I6772,I6766,I9128,I7232,g5368,g4243,I8162,g5918,g4198,I6434,g918,g6306,g4849,g4861,g4125,g5143,g6420,I3188,I1961,I8459,I7218,I4471,g2779,I5716,g1838,I2712,I7695,I7527,g1064,g4564,g4187,g6321,g127,g6931,I6420,g5371,g2544,g2361,g2682,g5535,g3933,I5767,I2373,g4842,I2457,g6544,g3180,I7910,g3829,I8888,I7244,g6619,g3558,I7441,I5119,g1789,g5042,g6290,g2316,g6122,g5781,I8414,I8671,g5419,g5533,g4847,g6363,g5300,I9230,g5816,g6343,g1292,g3732,g5179,g3277,I4445,I9092,g4359,g2777,I6296,g4697,I3626,g1742,g6161,g6766,g951,g6825,I6283,g2922,g1793,g5801,g3327,I5293,g5093,g3002,I9024,g6844,g1739,g390,g3094,I6561,g4423,g2958,g1358,g2733,g760,g1644,g6791,I8051,g3377,g714,g5693,I7802,g3864,I2290,g4630,g6698,g1812,g3791,g1678,g2197,g4638,I8107,g5731,g1608,g4607,g5596,g3972,g6687,g5485,g1664,g1339,g6548,g3132,g5860,g5173,g4911,g1638,I2225,g3704,g5260,g3295,g3498,I8229,g4652,g2364,g6748,g6725,g211,g5645,g2357,g2767,g4527,g4636,g4601,I7150,g2347,g5565,g5945,g5956,g33,g1648,I7276,g5935,g4265,g4381,g702,g6793,g4300,g1113,g3636,g4309,g4068,g5099,I5784,g1395,g2098,I2989,I2934,g6549,I7487,g3655,I5382,g3461,g6324,g6584,g3614,I8080,g4020,I8774,g6490,g3774,I7612,g6919,I3050,g6531,I7073,g4416,I2337,I4802,g3742,g2670,I7116,I8117,g6408,g4788,g3762,g3871,g1826,g5119,I6786,g5531,g5434,I6809,g5804,g3970,g2275,g719,g678,g4668,I2159,I2776,g3453,g5352,I4510,g6229,I8538,g3597,g696,g4894,g3526,g3941,g5625,I4371,g857,I3883,I8135,g1514,g4928,I5207,I8916,g1222,I3022,g6083,I8843,I2479,g582,g1039,g1422,g3350,I5451,I4498,g2119,g687,g5373,I6942,g5356,I2334,I6382,g5791,I8171,g3620,g3128,g6239,g5501,g6,g5067,g6610,I1865,g4736,g3226,g2788,g4732,g6798,I8681,g5861,g4522,g6279,g5532,g3752,g927,g3788,g6307,g2795,g6772,I7556,g2955,g2323,I6231,I2022,g1770,I3934,g6573,I8946,g3373,g940,g2818,g2921,g3932,g3689,g6308,I4941,I1942,g3631,I8647,g5110,g6104,I4040,I7593,I7432,g3906,g6513,I6425,g2891,I7817,g6777,g1681,I8273,g3136,g5019,g5097,I2870,g3075,g4843,I8961,I3411,I2108,I5865,I5728,I4276,I6143,I8875,g5442,I7679,g2944,I5851,g6915,I4646,g5623,g835,I8509,g3538,g2882,g1436,I7799,g6536,g3482,I8687,g4532,g135,g6749,g6530,I6452,g5536,I3222,g6093,g1332,g4041,g4141,I2658,I3190,g5924,I3584,I2526,g1549,g3108,I3408,I8456,g676,I8831,g6817,g4618,g6401,g909,I2154,g5921,I5837,I1951,g1925,I7999,g2902,g3305,g6354,g6406,g5925,g6166,g5699,g2889,g6179,g4289,g2587,I3422,g6289,g4463,I7164,g3768,g3364,I5233,g4036,g2551,g4371,I8710,g4644,I3749,g2770,g1108,g6297,I5406,I8684,g5361,g5664,g1819,g4655,g5911,I3370,I3441,I4486,g3601,g5509,g6257,I2021,g3934,g4340,g2157,g5380,g4948,I2949,g1322,g2667,g3685,g1783,I5217,g5534,g2941,g6281,g5212,g4831,I4246,I2162,g3181,g1320,g410,g3336,g5353,g3619,g3665,I8594,g3352,I2566,I2207,g1791,g3437,g4103,g3678,g5499,g3724,g928,g1460,I8395,g3374,g2722,g1729,I4334,g4641,I2688,I3886,I2552,g1821,g6035,I8837,I5157,g6129,g326,g6082,g6820,g6770,g1257,I5529,g3771,I7990,g37,g1484,I4303,g1333,g5092,I4459,g4651,g5673,g6247,g4512,g5741,g179,g3926,g5923,g4798,I2074,g2845,g2084,g3316,g4323,g3155,g6905,g2035,g3458,g3041,I8005,I8387,g208,g1543,g1161,g5530,I7988,I6485,I6689,g594,g6643,I8958,g4177,I8165,I9119,g3321,g2007,I1996,g4347,g4205,g6916,g4827,g5446,g1726,g5385,g6790,g1858,g2950,g3982,g1861,g5420,I8103,g3996,I1971,g5663,g613,g4149,I1987,I2508,g1884,I4546,g3546,g5241,g1589,g996,g689,I4210,g1498,I6750,I8828,g5684,g2778,g3337,g2893,g697,g5886,g6160,g3770,I4264,g1759,g453,g5503,I9058,g6504,g2166,g3659,g6878,g6726,g1628,g4602,g6301,g3899,I1932,I2857,g1175,g3612,g1991,g465,g1063,g2419,g1790,I7267,I7261,g3540,I6355,I5615,g6519,g5311,g684,I5400,I4455,g2588,I9104,I3740,I1880,g4625,I2604,g4180,g6170,g3644,g1954,I7224,g2416,g1267,g1823,g4040,I9173,I2047,g4252,g5603,g5424,I3641,I2109,g1631,g3456,I3316,g3527,g3280,I5391,g946,g3684,g283,g1894,I7852,g41,I2842,g3480,g2062,g3133,g4267,g6133,g4669,I4678,g5136,g6895,I6701,g1283,g6826,g5481,g5597,I4008,g6313,I8515,g898,I2935,g4741,I8650,g4410,g4425,g1922,I5469,g5091,g6105,g6747,g2518,g5518,I7549,g3216,I4309,g4508,g6359,g688,g6052,I3083,I9031,g4121,I4031,g4391,g2554,I7835,I5637,I2593,g3363,g5082,g1030,g6400,g6286,I2682,g394,g855,g3978,g4862,g4230,g4534,g2906,g5045,g5407,I9002,g4170,g6338,g4677,g4378,g2800,g3519,g3229,g6608,I9208,I8226,g6773,g279,g5314,g5160,g3275,g3657,I5991,g590,g6914,g6611,I6048,g3240,g4619,g6271,g6439,g3187,g900,I7091,g5553,g1138,I2933,g1733,g2692,g4248,g1857,I3425,I9152,I7550,I5223,g3775,I4354,g6414,g3330,g4771,I7548,I4331,g4694,I1958,g6833,g2339,I6672,I3848,g4770,I5302,I9028,g1546,g5648,I4391,I5977,g6634,g4845,g2866,g5245,g6778,I8126,g6188,g4941,g3910,g1294,g3617,g545,g3536,g2803,g5787,g5728,g1499,g6246,I3665,g4144,g1109,g5255,g6724,g6431,g6484,I7045,I2218,g3611,g6309,g2759,g3463,g2088,g2268,I5862,g1116,g4358,g4863,g3739,g4653,g6260,I7210,g6248,g2336,I5169,g6934,I7535,g1833,g5242,g520,g3862,g1319,g3083,I5723,g2956,g290,I3746,g6505,g5563,g6145,I7463,I3979,g6617,g2660,I5777,I4545,g5218,g3282,I4777,g5355,g4035,g5473,g913,I8488,g5177,g5863,g6886,g3851,g2873,g650,I8761,g3312,g3633,g3658,g5326,g3154,I8778,I3791,g3084,g4632,I7336,g4839,g6305,I4050,g6607,I4474,g4807,I8450,g6684,g1671,g3780,g5910,g4642,I9051,g669,g4797,I8232,g5579,g1754,g2599,g5555,g6576,g4376,g4903,g1491,g2850,I5502,g4727,g6683,I3225,g6044,g6924,g23,g6514,I2873,I7161,I3875,g5633,g5948,g610,g4511,g3863,g3836,I6175,I4444,g1878,g166,g922,g2106,g4491,g3196,g353,g5495,g4119,g6935,I5591,I7971,I3779,I8629,g3335,g197,g6265,g5240,g6468,I5739,g6448,g4285,I2215,g4563,I8282,g3233,g3656,g6165,g3535,I5324,g1899,I5929,g3355,I7683,g6080,g3683,g4377,g3632,g1363,g3874,g5318,g2953,I3059,I8429,g5582,g6795,I3044,g1898,g1233,g4472,I2707,I6057,I9125,g6397,g4528,g1084,I2318,I5702,g5214,I2061,g1219,g6705,I7569,g6118,I8447,I2961,g2776,I7061,g1044,g6939,g461,g6245,g4634,I3125,g6602,g3477,g6702,I6867,I2703,g1934,g5228,g128,I3833,g5013,g5151,g5854,g5937,g4597,g2945,I3294,I3698,g694,g2727,g4562,g4160,g6828,I4446,g4826,I6946,g3625,I5720,g628,g5478,I8913,g3877,I5659,g4600,I2578,I2805,I5182,g2010,g3122,g5118,g3113,g754,I3281,g5176,I6118,I6105,g6075,g4869,g6540,g6481,g4730,g6449,g4812,g1734,g6474,g4266,I7246,g2394,I1927,g6036,I3093,g4705,I5308,g5905,I7514,g1273,g1411,g2397,g5124,I6111,g3604,g4703,g5778,g39,I3804,g6511,g1535,g6696,g1650,I8220,I5427,g4238,g293,g1329,g6430,g5423,g3235,g4190,g4633,g3834,g6163,g3342,g1587,g1255,I6392,I6549,g4616,g1702,g2120,g1533,I2998,g2602,I3367,g2099,g5552,g5165,g2541,g5256,g4582,g1771,I9035,g6320,I8588,g1518,I6555,g3985,g1417,g4237,g5201,g3150,g2214,I2738,g1637,I2696,g5402,I2808,I2060,g6269,I2420,I5269,g3907,g937,g1749,g5546,g3960,I3699,g2954,I7104,I3785,g6014,g3901,I8246,I8997,I4270,I2324,I3915,I7906,g2565,g18,g2856,g4468,g3999,g5512,I4433,g5543,I3398,g6427,g1947,I8435,I2424,g6294,I8210,I4504,g2721,g2659,g277,g4720,g3230,I6937,g1293,g5892,I8512,I3741,g4804,g4345,g3682,I4212,g1480,g4367,g3664,I4189,I3325,g1688,g3067,g5098,I8342,g6925,g3831,g6091,g6882,g4637,g6154,I8074,g6092,g2862,g3789,g4929,g2834,g6422,g4374,g4774,I2867,g5436,g1459,g3258,g2695,g4191,I4340,g4107,I8779,g1832,g6330,g2155,g2213,I8300,g1250,I3056,I3258,I3505,g6787,g4044,g4592,g6816,g3145,I2796,I8061,g3421,g3012,g336,g2644,g6622,g6758,g5050,I8079,g2555,g3481,g3241,I8506,g3176,g6606,g4531,I5868,g5304,g5440,I8180,g4824,g6523,g6686,g6688,g6121,g3323,g1682,g3371,g715,g4143,I3516,I6269,g3049,g5381,g1784,g5168,I4240,g4549,I5309,g6296,g6034,g1055,g4497,I7434,g1741,g1911,g2410,I3198,I3301,g2294,I9064,g6854,g6318,I5027,g5621,g4606,I8177,g3484,I3726,g4656,I3232,g5577,g2976,I2907,g1834,g2912,I4288,I2839,g2350,I6874,g3799,g5012,g1735,g1654,I9101,g2160,I4986,I8497,I5848,g3767,I8940,g4460,I5109,g5714,I2193,g4759,g1142,I3355,g46,I3313,g6711,g1295,I3385,I3739,g2243,I8702,I6023,g3304,g5139,g4588,I6470,I3034,g5153,g170,g1513,I8356,g1391,g889,g4105,I2399,g1890,g3466,g4014,g5600,g5873,g2744,g6853,g2628,I2240,g6873,I3755,g5296,g332,g6835,g5545,g3517,I3563,g3293,g3557,g6543,I5424,I4205,g5237,g6821,I5409,g3642,I7490,I6952,g4660,I2449,I4743,g663,g5198,g5051,I5926,g5488,I8249,g729,g2505,g6692,g1047,I2721,g1325,g3802,I2782,I4267,g3281,I3855,g139,g3691,g5604,I6102,g3114,g1879,g6268,g5752,g4380,I3471,g5540,g2390,g4938,g5890,I2627,g2296,g5362,g2473,I5630,g6794,g4442,g5458,I3062,g4110,g3366,g4394,I5705,g1402,g3345,g4567,g4299,I2946,I6090,g5185,g1846,g4113,g2525,g2871,g6694,g3278,g6291,g3093,I6096,g6521,g6100,I3413,g2740,g6079,g5074,I2234,g2307,I8521,g2691,I4940,g5277,I3826,g4680,g3236,I3274,g3384,I8878,g5441,g3885,g6127,I7970,g6801,g6812,I4203,g5011,g567,g6563,g6189,g5615,g1940,I3770,I8118,g5411,g6689,I8752,g4819,I5249,g4349,g6900,g4115,g5183,g6830,g1706,g4004,g5141,g1075,I9041,g2001,g449,g1891,I3019,I4176,g5797,g3763,g4209,g3292,I6685,I2623,I2864,g2863,g6700,g6880,g899,g5875,g1503,g5505,I8641,g3627,g5539,g4043,g6580,g1193,g6541,I5059,I6534,I6963,g6487,I7564,g3912,I3761,g1773,g5330,g1326,g4357,I3620,I7342,I7190,g157,I9227,g3533,g4457,g5410,g6750,g2461,I7494,g434,g2378,g2043,g6784,g5188,g4176,I7197,g6703,g3749,I8491,g5437,g2484,g1290,g6192,g5014,I1969,g4145,g6292,I6186,g2794,I6744,g3157,g4815,g6740,I1850,g1908,g6263,g4811,g1674,I3543,I3170,I8524,I2964,g1291,I3513,g1689,g2897,g5472,g1221,g2754,g736,g1112,g6443,I3007,g3649,g2967,g1160,g3358,I2741,g5670,g5216,g2026,g4147,g4184,g3449,g5158,g3813,g5329,g6085,g4648,I2825,g3247,g5893,g6937,g6928,g5720,g4853,g6560,g5161,g2437,I7577,g4947,g2961,g5573,I8812,I9179,g5634,g3896,I2756,I9107,g964,g5665,g3100,I5050,I3858,g4761,g3539,I2391,g2819,I2090,g1418,g2752,I9077,g3589,g2178,g6591,g1830,g4823,I6194,g865,g5398,I3893,g6494,g4213,g4768,g6819,g2998,g6231,g3703,g4453,g4296,I2929,g5897,I4151,g4244,g3613,I3864,g1366,g4232,g5392,g5113,g3686,g437,g1204,g4520,g6409,g6930,I8564,I3599,I2728,g821,g6322,g1156,I3800,I6099,g4262,g4186,g5182,g6123,I4495,I4534,g24,g5117,g5620,g6249,I5116,g2837,I2067,g1931,g2757,g5023,g5112,g6157,g1450,g3776,I6414,g4150,g2241,g2973,g929,g489,g6788,I2791,I4784,g602,g1115,g4058,I8370,g6827,g4529,g4154,g6809,g2215,g5776,g897,g327,I4402,I3836,g5391,I7313,g7,g3147,I2385,g2805,g4245,g6528,I6798,g4454,I7814,g6164,g2687,g4933,I7689,I2601,I4255,g6140,I4424,g6251,I6027,g3806,g5726,g6745,g5556,g854,g6623,I9021,g1461,g2932,I4343,g3173,g3599,g2568,I7521,g4053,g4042,g1043,g3564,g5414,g945,g4021,I2955,I6391,I5196,I6507,g1666,I4366,I3605,I2340,g3819,g4877,I3723,g4808,I8975,g4402,g3845,g4640,g6233,I8972,I8119,g3208,g2230,g6261,g6637,g1813,g2212,g6434,g6574,g4766,I4791,g3671,g4799,g4513,g4162,I1868,g6413,g486,g3146,I3071,I8223,g3319,g6040,g1760,g6789,I6054,g3903,g2716,g2422,I8129,I4706,g1937,I6819,g1555,I4537,g3629,g3986,I8555,g6891,I4223,g5649,I2979,g3251,I9167,g2284,g3172,g5564,I9161,I6441,g5114,I2165,I4752,g3897,I8620,I3933,g3800,g1769,g3303,g2949,g6660,g5264,g6495,I8420,g2333,g1672,g5487,g3922,I3169,g1764,g1627,g1282,g2653,g985,g2405,I2692,g5853,g5192,g3764,g3367,g2790,g4674,g2391,g4314,I7701,g6333,g6594,I2309,g6256,g4273,g1534,I9095,I6430,g1410,g6738,g699,I2312,I5333,g1696,I6558,g6437,g212,g4153,g6410,g230,I3632,g1994,I8668,g6162,g693,g4704,g5181,I5618,g143,g6441,I8600,g5883,I8907,g5940,g4611,I5948,g2110,g2678,g4691,g5489,g4635,g3340,I2091,g6078,g4450,g6754,g5632,g3124,g2306,I4258,I2355,g6587,g3022,g4583,g6211,I3352,I5782,I8201,g1263,I5352,g5450,I5351,g6451,g3283,g2467,g5711,g5175,g4643,g5701,g5159,g6927,g2719,I9122,g3792,g1316,g4253,g4627,I7856,I8910,g3673,I4783,I2848,I7542,I6607,g4828,g2031,g6447,g3663,g4779,g3979,g5884,g2173,I6170,g5307,g5698,I3322,I9074,I8309,I8585,I8881,g1581,I3797,g5171,I5548,g418,g853,g1763,g1529,I7113,g4533,g2631,I5499,g6575,I1856,g4225,g3199,g1558,I2179,I7339,g5782,g6644,I6377,g3308,g1328,I4362,I8494,I7557,g1106,g3286,g6883,g6293,g3873,I2275,g5788,g4722,g6571,I8897,g1680,g6329,g4684,g3815,g4444,g6110,g3530,g5507,I2414,I8815,I4226,g4726,g2087,g2194,I5708,g5187,I7871,g3755,g691,I5876,g2791,I2122,g5857,g5150,I2131,g3311,g441,g2311,g5936,g6062,g5059,g19,g5270,g1775,g2460,g2550,g3883,I3202,g2637,g4169,g5537,I6093,g6238,I5517,g5359,g3518,I3546,g2743,I6723,g3646,g6132,I7529,I2134,g6402,I4429,g5668,g6270,g2343,I5658,I7208,g5386,g3019,I4235,g6723,I4688,I7501,I6321,g287,I3847,g6482,g4155,I3909,g2756,I4318,g2096,I8082,g5084,g3905,g1731,g3787,I2321,g3751,I2364,g532,g639,g25,g5696,g2291,I3691,g2705,g6326,g3959,g3030,I8279,g3743,I2497,I4173,g4758,I8186,I2506,g4581,g5213,g6436,g3375,I5597,g4503,g1519,g3381,g1286,I4667,I7859,g6316,g866,g4219,I5609,I3553,I7404,I1835,g6098,g1673,g4661,I5388,I2821,g4786,g2766,I3550,I5071,g3195,I6362,g5581,I7520,g32,I3537,g3054,I7646,g2100,I1853,g2577,I2349,g2032,g5876,g3602,g2109,g3200,g4489,I7173,g878,g3341,g896,I3823,I6004,g6060,g5995,I7187,g2853,I7960,g5170,g6731,g6701,g5674,I6756,g6884,I8138,g6503,g3889,g1807,g4165,I8573,I7346,g4429,I4398,g5862,I2453,g681,I6349,g2826,g4772,g2935,g5740,g6832,g1552,g1381,g1190,I8696,g5583,g4803,I8531,g5156,g5094,g2481,g3545,I1832,g3271,g1582,I3525,I7355,I3819,g5780,I5674,g5666,g4688,g858,g3387,I7796,g3343,g4240,I8678,I5750,g1679,g6432,g2145,I6327,g6086,g5015,g6155,g3747,I7892,g5224,I3678,I4762,I2877,g6834,g950,g3192,I2893,I5508,g3089,I6008,g278,g218,I6500,g6885,g5622,I7506,I8503,I8360,g2494,I8991,I4315,g210,g1539,g5889,g3628,I6177,g6232,I2916,g3670,g3939,g3839,g5885,I3672,I3952,g5387,I3161,g4874,I3140,g6452,g29,g4361,I5328,g3989,g1236,g6331,g5708,g5874,g971,g4537,g3651,I1859,g4535,g3016,g6542,g2097,I8386,g6081,g2748,g445,I3653,g3634,g1017,g2008,g3285,I6063,I7012,g1557,I5713,g4137,g5220,g4251,I8470,g1691,g6628,g4092,g4932,g1574,I3531,g2292,g5580,g554,g4714,I3096,g4598,g4765,I2150,g3007,I8767,g1330,g541,g5452,g2783,g3534,I6132,g4369,I3478,g1426,g5348,I4211,g3680,I7981,g1324,g3882,g1720,g5920,g3681,g3110,I6340,I3419,g3988,g3893,g5975,g3299,I7258,g5017,I8070,g1321,g4716,g3279,g1641,I7069,g2615,g3687,I4483,g4780,g5232,I3447,g6405,I8869,I6456,I5292,I2880,g571,I8240,I2611,g2409,I8113,g3034,g5575,g2102,g1957,g6569,I7216,g1369,g4167,g1943,I3148,g1788,g6369,g3648,g3757,g1849,g6097,g5676,g5818,I6126,I3065,g4822,g4787,g2040,I4170,g5215,g6124,g3529,g6897,g4390,I3456,I6956,g3833,g5193,I3729,g2915,I6033,I5208,I5633,g1684,I8159,g6783,I2528,g1288,I2904,g4825,I7312,I2428,g2030,g2876,g1897,g6102,g117,I3942,I3474,g1053,I8570,I5753,g1724,g1045,g2317,g3741,g548,g512,g1551,g6727,I4489,I8423,g921,I1935,g1323,g4835,g4566,g1504,I3861,g4579,g3888,g3803,g3310,I4684,I3788,g4015,I4519,g3298,g6101,g2622,I2053,g2928,g3705,g3478,I7002,g5044,I4935,g1721,g2892,g2154,g3930,I8270,I3656,I3675,I4664,I7570,g2842,g5482,g4672,g6670,g6802,g337,I5242,g2828,g6234,g5120,g22,g3544,I4782,g3096,g2698,g2253,g3692,g6597,g6894,g4521,I5854,g4904,g6311,g6552,g947,I4441,g847,I5466,I2299,I3412,I3001,g4122,I3758,g4148,g3064,g5047,g846,g3046,g6771,g54,g3971,g6076,g2061,I8426,g6444,g2266,g5794,I5294,I6039,g4510,I1995,g1714,g3571,I8548,I2527,g5700,g2817,g260,I5053,I6182,g6267,g6922,g5560,g1423,I5472,g5891,I3244,I4261,g6153,I8745,I8453,g3867,g2608,g3455,g44,g2244,g4239,g6335,g2822,g4431,I2175,g2231,g3900,g3103,g3318,g2713,I3319,g1270,I4195,I9047,I7637,I4794,g5730,g815,g849,I8653,I6525,g4502,I3617,g3487,g3694,I6992,I8803,g5618,I8699,g2934,g2869,g4301,I2379,I3457,I5442,g2413,I8196,g1206,I3261,I6885,g6941,g4142,g2449,g4545,I1978,I5153,g269,g3099,I2080,I6045,I5606,g6539,g6940,I5505,g3647,I5654,g4386,g3661,g2196,I8579,g4000,g1715,g1639,g4544,g1774,g5865,g4857,g6340,g2830,g1173,g3359,I7110,g3879,g6926,g3730,g6259,g6047,g4398,g3488,g4805,g4867,I9066,g658,I2062,g3326,g5566,g3242,g2581,g266,g3504,g4852,I3572,I5397,g3460,g6562,I8773,g1612,I5188,g6840,g2232,I7081,g292,g5619,g3454,I8544,I2922,I8285,g6839,g49,I3343,g4136,I5177,I3346,g2370,I3808,g6654,I8235,g1822,I8378,g2583,g5324,I6635,g3434,g2907,g2946,I6582,g5584,g716,I5270,g4379,g3954,g457,I7600,g3856,I3485,g5247,g4698,g6032,g6423,I5189,g175,g5249,g6328,g6568,I2115,g3177,g5457,I3468,I6933,g5065,g2849,I6775,I2245,g1398,g3191,g4596,I2013,I8376,I8217,I4204,g5628,g5558,I2408,g3070,g3605,g3782,I8552,g5211,g161,I5320,I6753,I2643,g4745,g6744,g6581,g3635,g4790,g5630,I8394,I6176,g4679,g2801,I5626,g3962,g1209,I6334,I7284,g1359,I1871,g2726,g1122,g3965,g5018,I8393,g1883,g1848,g1439,I3736,g5551,I6386,g5904,g6435,I4522,g6419,g338,g4284,I6816,g4163,g2091,g3082,g2112,I7832,g1653,g4509,g3992,I8209,g5779,g2859,I7634,I6371,g2619,g3849,g6456,I3684,g5909,g2408,I9014,I6615,g5624,g2771,g6699,g2320,I3705,g4218,I6540,g4183,g842,I5204,I5882,I3068,g4159,I8969,g6717,g5229,I3382,g6480,g6603,g2919,g4993,g616,I8479,g5894,g634,g4086,I8027,g4194,g5186,I5668,I6397,I6964,I2543,g2125,g4384,g3760,I2003,g1836,I4321,g4692,g4577,g3503,g4776,g2888,g5916,g5887,g6061,g3923,g5549,g40,I5551,g4764,I6501,g2436,I4980,g944,I2237,I3240,g3758,g1107,g4859,g6659,I3578,g6137,g5717,g6446,I3560,g323,g5123,g3294,g3637,I8482,g3650,g6237,I5487,g4100,g524,g5476,g4118,g4034,I2952,g5315,g5617,I8755,I3291,g6685,g4281,g836,g6510,g3773,g4343,I8988,I8623,g3190,g6274,I5412,g2813,g5896,g4193,g6921,g848,g923,g284,I9170,g4858,g2176,g3609,I2766,g4782,I6253,g6250,g3728,g4406,g3227,g5677,I4462,g4496,I7225,g5194,g4735,g2234,g5943,I2668,g4138,g4185,I3846,g646,g3975,g1738,I3764,I7099,g1747,I8614,g1191,g1559,I2967,g6690,g4778,g4763,g1246,I3112,g3733,g3215,g3881,g5465,I3178,g6848,g4518,g6095,I6697,g5199,g5146,g3231,I4300,I1994,I5899,I3647,g6277,g4846,g6126,g930,g6908,I6930,I4220,g3290,g5675,g6532,I4066,I2817,g3344,g3828,g6881,g6057,I3358,g2884,I8252,I8467,g5166,g3969,g5949,I3687,g4002,g6115,g6533,g1472,g6096,I8644,g224,I4150,I3519,g5567,g1595,I9149,I5033,I2898,g942,g6570,g6241,g5661,g5574,g6300,g6149,g3450,g4249,I7590,I8894,g4383,g1632,g2952,g6151,g6650,g2948,g664,g2966,I7996,g2245,g3643,I8707,I7058,g4102,g3924,g3510,g1036,g2607,g2073,g852,g5542,g2255,g6051,g3837,g4752,g2732,I3923,g6850,g3309,I4358,g6421,g2233,g6746,I8194,g4711,g2015,I6475,I5913,I4059,g2831,g4195,g2165,I3794,I3876,I2676,g3554,I4337,I2584,g6917,I3720,g4189,g6742,I3916,g4519,g5096,g6609,g1969,g3981,g1811,I2269,g3267,g3987,g2021,g6592,g4341,I6918,g6899,g2840,g1802,g5561,g5303,I6743,I4955,g4462,g3362,g3958,I3405,g3610,g4678,g3156,I6299,g3433,I9155,I2281,I5065,g690,g504,g6579,g471,g4108,g3769,I3013,I3708,I8208,g6276,g1275,I6330,I6042,g5805,I4821,I6244,g5667,g6491,g2252,g4157,g188,I5043,g5686,g4498,g6618,g4226,I3137,g5384,I7238,g6136,g5554,g3821,g4395,I7318,I3077,g3990,g5669,g952,I4375,g5155,g3709,I2119,g1670,I2089,g3501,I5236,g4753,g5261,I2835,g5631,g1049,g3786,g5388;
//# 19 inputs
//# 22 outputs
//# 228 D-type flipflops
//# 3570 inverters
//# 2027 gates (955 ANDs + 528 NANDs + 431 ORs + 113 NORs)
//
//
//
  MSFF DFF_0(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g46),.DATA(g4109));
  MSFF DFF_1(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g45),.DATA(g4108));
  MSFF DFF_2(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g44),.DATA(g4107));
  MSFF DFF_3(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g42),.DATA(g4106));
  MSFF DFF_4(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g40),.DATA(g4105));
  MSFF DFF_5(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g39),.DATA(g4103));
  MSFF DFF_6(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g38),.DATA(g4102));
  MSFF DFF_7(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g37),.DATA(g4101));
  MSFF DFF_8(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g36),.DATA(g4100));
  MSFF DFF_9(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g32),.DATA(g4099));
  MSFF DFF_10(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g28),.DATA(g6727));
  MSFF DFF_11(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g24),.DATA(g6726));
  MSFF DFF_12(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g18),.DATA(g6725));
  MSFF DFF_13(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g14),.DATA(g6724));
  MSFF DFF_14(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g10),.DATA(g6723));
  MSFF DFF_15(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g6),.DATA(g6722));
  MSFF DFF_16(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2),.DATA(g6721));
  MSFF DFF_17(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1),.DATA(g6720));
  MSFF DFF_18(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g48),.DATA(g6729));
  MSFF DFF_19(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g47),.DATA(g4112));
  MSFF DFF_20(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g41),.DATA(g4110));
  MSFF DFF_21(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g22),.DATA(g4104));
  MSFF DFF_22(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g23),.DATA(g4098));
  MSFF DFF_23(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g284),.DATA(g3224));
  MSFF DFF_24(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g285),.DATA(g3225));
  MSFF DFF_25(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g286),.DATA(g3226));
  MSFF DFF_26(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g287),.DATA(g3227));
  MSFF DFF_27(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g288),.DATA(g3228));
  MSFF DFF_28(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g289),.DATA(g3229));
  MSFF DFF_29(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g290),.DATA(g3230));
  MSFF DFF_30(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g291),.DATA(g3231));
  MSFF DFF_31(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g292),.DATA(g3232));
  MSFF DFF_32(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g338),.DATA(g5475));
  MSFF DFF_33(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g341),.DATA(g5476));
  MSFF DFF_34(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g345),.DATA(g5477));
  MSFF DFF_35(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g349),.DATA(g5478));
  MSFF DFF_36(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g353),.DATA(g5479));
  MSFF DFF_37(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g357),.DATA(g5480));
  MSFF DFF_38(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g361),.DATA(g6582));
  MSFF DFF_39(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g49),.DATA(g6583));
  MSFF DFF_40(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g54),.DATA(g6584));
  MSFF DFF_41(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g59),.DATA(g6585));
  MSFF DFF_42(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g64),.DATA(g6586));
  MSFF DFF_43(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g69),.DATA(g6587));
  MSFF DFF_44(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g74),.DATA(g6588));
  MSFF DFF_45(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g79),.DATA(g6589));
  MSFF DFF_46(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g84),.DATA(g6590));
  MSFF DFF_47(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g366),.DATA(g6278));
  MSFF DFF_48(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g370),.DATA(g5693));
  MSFF DFF_49(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g374),.DATA(g5694));
  MSFF DFF_50(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g378),.DATA(g5695));
  MSFF DFF_51(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g382),.DATA(g5696));
  MSFF DFF_52(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g386),.DATA(g5697));
  MSFF DFF_53(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g390),.DATA(g5698));
  MSFF DFF_54(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g394),.DATA(g5699));
  MSFF DFF_55(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g398),.DATA(g5700));
  MSFF DFF_56(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g326),.DATA(g4840));
  MSFF DFF_57(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g327),.DATA(g4117));
  MSFF DFF_58(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g328),.DATA(g4118));
  MSFF DFF_59(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g331),.DATA(g4119));
  MSFF DFF_60(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g323),.DATA(g4120));
  MSFF DFF_61(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g332),.DATA(g6823));
  MSFF DFF_62(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g336),.DATA(g6925));
  MSFF DFF_63(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g337),.DATA(g2585));
  MSFF DFF_64(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g128),.DATA(g5138));
  MSFF DFF_65(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g131),.DATA(g5139));
  MSFF DFF_66(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g135),.DATA(g5140));
  MSFF DFF_67(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g139),.DATA(g5141));
  MSFF DFF_68(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g143),.DATA(g6401));
  MSFF DFF_69(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g152),.DATA(g6402));
  MSFF DFF_70(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g161),.DATA(g6403));
  MSFF DFF_71(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g170),.DATA(g6404));
  MSFF DFF_72(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g179),.DATA(g6405));
  MSFF DFF_73(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g188),.DATA(g6406));
  MSFF DFF_74(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g148),.DATA(g5874));
  MSFF DFF_75(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g157),.DATA(g5470));
  MSFF DFF_76(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g166),.DATA(g5471));
  MSFF DFF_77(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g175),.DATA(g5472));
  MSFF DFF_78(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g184),.DATA(g5473));
  MSFF DFF_79(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g193),.DATA(g5474));
  MSFF DFF_80(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g117),.DATA(g4839));
  MSFF DFF_81(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g118),.DATA(g4113));
  MSFF DFF_82(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g119),.DATA(g4114));
  MSFF DFF_83(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g122),.DATA(g4115));
  MSFF DFF_84(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g114),.DATA(g4116));
  MSFF DFF_85(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g123),.DATA(g6940));
  MSFF DFF_86(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g111),.DATA(g6277));
  MSFF DFF_87(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g127),.DATA(g6941));
  MSFF DFF_88(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g276),.DATA(g5877));
  MSFF DFF_89(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g277),.DATA(g6104));
  MSFF DFF_90(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g278),.DATA(g6105));
  MSFF DFF_91(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g279),.DATA(g6106));
  MSFF DFF_92(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g280),.DATA(g5878));
  MSFF DFF_93(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g281),.DATA(g6107));
  MSFF DFF_94(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g282),.DATA(g6841));
  MSFF DFF_95(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g283),.DATA(g6842));
  MSFF DFF_96(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g204),.DATA(g5875));
  MSFF DFF_97(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g205),.DATA(g6100));
  MSFF DFF_98(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g206),.DATA(g6101));
  MSFF DFF_99(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g207),.DATA(g6102));
  MSFF DFF_100(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g208),.DATA(g5876));
  MSFF DFF_101(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g209),.DATA(g6103));
  MSFF DFF_102(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g210),.DATA(g6839));
  MSFF DFF_103(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g211),.DATA(g6840));
  MSFF DFF_104(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g212),.DATA(g3233));
  MSFF DFF_105(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g218),.DATA(g3234));
  MSFF DFF_106(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g224),.DATA(g3235));
  MSFF DFF_107(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g230),.DATA(g3236));
  MSFF DFF_108(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g236),.DATA(g3237));
  MSFF DFF_109(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g242),.DATA(g3238));
  MSFF DFF_110(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g248),.DATA(g3239));
  MSFF DFF_111(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g254),.DATA(g3240));
  MSFF DFF_112(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g260),.DATA(g3241));
  MSFF DFF_113(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g567),.DATA(g4121));
  MSFF DFF_114(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g598),.DATA(g4122));
  MSFF DFF_115(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g634),.DATA(g4424));
  MSFF DFF_116(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g642),.DATA(g4658));
  MSFF DFF_117(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g606),.DATA(g4857));
  MSFF DFF_118(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g646),.DATA(g5148));
  MSFF DFF_119(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g650),.DATA(g5329));
  MSFF DFF_120(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g654),.DATA(g5490));
  MSFF DFF_121(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g571),.DATA(g5580));
  MSFF DFF_122(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g578),.DATA(g6592));
  MSFF DFF_123(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g582),.DATA(g6593));
  MSFF DFF_124(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g586),.DATA(g6594));
  MSFF DFF_125(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g574),.DATA(g6591));
  MSFF DFF_126(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g590),.DATA(g6595));
  MSFF DFF_127(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g594),.DATA(g6596));
  MSFF DFF_128(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g602),.DATA(g4123));
  MSFF DFF_129(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g610),.DATA(g4124));
  MSFF DFF_130(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g613),.DATA(g4423));
  MSFF DFF_131(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g616),.DATA(g4657));
  MSFF DFF_132(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g619),.DATA(g4858));
  MSFF DFF_133(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g622),.DATA(g5147));
  MSFF DFF_134(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g625),.DATA(g5328));
  MSFF DFF_135(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g628),.DATA(g5489));
  MSFF DFF_136(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g631),.DATA(g5581));
  MSFF DFF_137(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g43),.DATA(g6407));
  MSFF DFF_138(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g266),.DATA(g4659));
  MSFF DFF_139(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g658),.DATA(g4425));
  MSFF DFF_140(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g667),.DATA(g4127));
  MSFF DFF_141(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g666),.DATA(g4128));
  MSFF DFF_142(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g662),.DATA(g1831));
  MSFF DFF_143(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g663),.DATA(g4125));
  MSFF DFF_144(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g664),.DATA(g1288));
  MSFF DFF_145(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g471),.DATA(g1291));
  MSFF DFF_146(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g665),.DATA(g4126));
  MSFF DFF_147(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g478),.DATA(g1292));
  MSFF DFF_148(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g638),.DATA(g1289));
  MSFF DFF_149(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g639),.DATA(g1290));
  MSFF DFF_150(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g699),.DATA(g4426));
  MSFF DFF_151(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g702),.DATA(g1293));
  MSFF DFF_152(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g675),.DATA(g1294));
  MSFF DFF_153(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g669),.DATA(g5582));
  MSFF DFF_154(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g676),.DATA(g5330));
  MSFF DFF_155(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g672),.DATA(g5491));
  MSFF DFF_156(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3),.DATA(g6597));
  MSFF DFF_157(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g7),.DATA(g6598));
  MSFF DFF_158(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g11),.DATA(g6599));
  MSFF DFF_159(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g15),.DATA(g6602));
  MSFF DFF_160(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g19),.DATA(g6600));
  MSFF DFF_161(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g25),.DATA(g6601));
  MSFF DFF_162(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g29),.DATA(g6853));
  MSFF DFF_163(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g33),.DATA(g6854));
  MSFF DFF_164(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g690),.DATA(g4142));
  MSFF DFF_165(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g691),.DATA(g4143));
  MSFF DFF_166(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g692),.DATA(g4144));
  MSFF DFF_167(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g693),.DATA(g4145));
  MSFF DFF_168(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g694),.DATA(g4146));
  MSFF DFF_169(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g695),.DATA(g4147));
  MSFF DFF_170(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g696),.DATA(g4148));
  MSFF DFF_171(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g697),.DATA(g4149));
  MSFF DFF_172(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g677),.DATA(g4129));
  MSFF DFF_173(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g678),.DATA(g4130));
  MSFF DFF_174(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g679),.DATA(g4131));
  MSFF DFF_175(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g680),.DATA(g4132));
  MSFF DFF_176(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g681),.DATA(g4133));
  MSFF DFF_177(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g682),.DATA(g4134));
  MSFF DFF_178(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g683),.DATA(g4135));
  MSFF DFF_179(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g684),.DATA(g4136));
  MSFF DFF_180(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g685),.DATA(g4137));
  MSFF DFF_181(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g686),.DATA(g4138));
  MSFF DFF_182(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g687),.DATA(g4139));
  MSFF DFF_183(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g688),.DATA(g4140));
  MSFF DFF_184(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g689),.DATA(g4141));
  MSFF DFF_185(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g698),.DATA(g4150));
  MSFF DFF_186(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g668),.DATA(g6800));
  MSFF DFF_187(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g485),.DATA(g6801));
  MSFF DFF_188(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g402),.DATA(g4849));
  MSFF DFF_189(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g406),.DATA(g4850));
  MSFF DFF_190(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g410),.DATA(g4851));
  MSFF DFF_191(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g414),.DATA(g4852));
  MSFF DFF_192(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g418),.DATA(g4853));
  MSFF DFF_193(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g422),.DATA(g4854));
  MSFF DFF_194(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g426),.DATA(g4855));
  MSFF DFF_195(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g430),.DATA(g4856));
  MSFF DFF_196(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g461),.DATA(g4841));
  MSFF DFF_197(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g457),.DATA(g4842));
  MSFF DFF_198(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g453),.DATA(g4843));
  MSFF DFF_199(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g449),.DATA(g4844));
  MSFF DFF_200(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g445),.DATA(g4845));
  MSFF DFF_201(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g441),.DATA(g4846));
  MSFF DFF_202(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g437),.DATA(g4847));
  MSFF DFF_203(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g434),.DATA(g4848));
  MSFF DFF_204(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g545),.DATA(g6824));
  MSFF DFF_205(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g548),.DATA(g6825));
  MSFF DFF_206(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g551),.DATA(g6826));
  MSFF DFF_207(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g554),.DATA(g6827));
  MSFF DFF_208(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g197),.DATA(g6509));
  MSFF DFF_209(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g269),.DATA(g6510));
  MSFF DFF_210(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g293),.DATA(g6511));
  MSFF DFF_211(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g297),.DATA(g6512));
  MSFF DFF_212(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g500),.DATA(g6497));
  MSFF DFF_213(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g504),.DATA(g6498));
  MSFF DFF_214(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g508),.DATA(g6499));
  MSFF DFF_215(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g512),.DATA(g6500));
  MSFF DFF_216(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g516),.DATA(g6501));
  MSFF DFF_217(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g520),.DATA(g6502));
  MSFF DFF_218(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g524),.DATA(g6503));
  MSFF DFF_219(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g528),.DATA(g6504));
  MSFF DFF_220(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g532),.DATA(g6508));
  MSFF DFF_221(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g465),.DATA(g6507));
  MSFF DFF_222(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g536),.DATA(g6506));
  MSFF DFF_223(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g541),.DATA(g6505));
  MSFF DFF_224(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g486),.DATA(g2586));
  MSFF DFF_225(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g489),.DATA(g2587));
  MSFF DFF_226(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g496),.DATA(g6745));
  MSFF DFF_227(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g492),.DATA(g6744));
//
  NOT NOT1_0(.VSS(VSS),.VDD(VDD),.Y(I1825),.A(g361));
  NOT NOT1_1(.VSS(VSS),.VDD(VDD),.Y(g706),.A(I1825));
  NOT NOT1_2(.VSS(VSS),.VDD(VDD),.Y(g709),.A(g114));
  NOT NOT1_3(.VSS(VSS),.VDD(VDD),.Y(g710),.A(g128));
  NOT NOT1_4(.VSS(VSS),.VDD(VDD),.Y(g714),.A(g131));
  NOT NOT1_5(.VSS(VSS),.VDD(VDD),.Y(g715),.A(g135));
  NOT NOT1_6(.VSS(VSS),.VDD(VDD),.Y(I1832),.A(g143));
  NOT NOT1_7(.VSS(VSS),.VDD(VDD),.Y(g716),.A(I1832));
  NOT NOT1_8(.VSS(VSS),.VDD(VDD),.Y(I1835),.A(g205));
  NOT NOT1_9(.VSS(VSS),.VDD(VDD),.Y(g719),.A(I1835));
  NOT NOT1_10(.VSS(VSS),.VDD(VDD),.Y(I1838),.A(g206));
  NOT NOT1_11(.VSS(VSS),.VDD(VDD),.Y(g729),.A(I1838));
  NOT NOT1_12(.VSS(VSS),.VDD(VDD),.Y(I1841),.A(g207));
  NOT NOT1_13(.VSS(VSS),.VDD(VDD),.Y(g736),.A(I1841));
  NOT NOT1_14(.VSS(VSS),.VDD(VDD),.Y(I1844),.A(g208));
  NOT NOT1_15(.VSS(VSS),.VDD(VDD),.Y(g743),.A(I1844));
  NOT NOT1_16(.VSS(VSS),.VDD(VDD),.Y(I1847),.A(g209));
  NOT NOT1_17(.VSS(VSS),.VDD(VDD),.Y(g749),.A(I1847));
  NOT NOT1_18(.VSS(VSS),.VDD(VDD),.Y(I1850),.A(g210));
  NOT NOT1_19(.VSS(VSS),.VDD(VDD),.Y(g754),.A(I1850));
  NOT NOT1_20(.VSS(VSS),.VDD(VDD),.Y(I1853),.A(g211));
  NOT NOT1_21(.VSS(VSS),.VDD(VDD),.Y(g760),.A(I1853));
  NOT NOT1_22(.VSS(VSS),.VDD(VDD),.Y(I1856),.A(g204));
  NOT NOT1_23(.VSS(VSS),.VDD(VDD),.Y(g766),.A(I1856));
  NOT NOT1_24(.VSS(VSS),.VDD(VDD),.Y(I1859),.A(g277));
  NOT NOT1_25(.VSS(VSS),.VDD(VDD),.Y(g774),.A(I1859));
  NOT NOT1_26(.VSS(VSS),.VDD(VDD),.Y(I1862),.A(g278));
  NOT NOT1_27(.VSS(VSS),.VDD(VDD),.Y(g784),.A(I1862));
  NOT NOT1_28(.VSS(VSS),.VDD(VDD),.Y(I1865),.A(g279));
  NOT NOT1_29(.VSS(VSS),.VDD(VDD),.Y(g791),.A(I1865));
  NOT NOT1_30(.VSS(VSS),.VDD(VDD),.Y(I1868),.A(g280));
  NOT NOT1_31(.VSS(VSS),.VDD(VDD),.Y(g798),.A(I1868));
  NOT NOT1_32(.VSS(VSS),.VDD(VDD),.Y(I1871),.A(g281));
  NOT NOT1_33(.VSS(VSS),.VDD(VDD),.Y(g804),.A(I1871));
  NOT NOT1_34(.VSS(VSS),.VDD(VDD),.Y(I1874),.A(g282));
  NOT NOT1_35(.VSS(VSS),.VDD(VDD),.Y(g809),.A(I1874));
  NOT NOT1_36(.VSS(VSS),.VDD(VDD),.Y(I1877),.A(g283));
  NOT NOT1_37(.VSS(VSS),.VDD(VDD),.Y(g815),.A(I1877));
  NOT NOT1_38(.VSS(VSS),.VDD(VDD),.Y(I1880),.A(g276));
  NOT NOT1_39(.VSS(VSS),.VDD(VDD),.Y(g821),.A(I1880));
  NOT NOT1_40(.VSS(VSS),.VDD(VDD),.Y(g829),.A(g323));
  NOT NOT1_41(.VSS(VSS),.VDD(VDD),.Y(g830),.A(g338));
  NOT NOT1_42(.VSS(VSS),.VDD(VDD),.Y(g834),.A(g341));
  NOT NOT1_43(.VSS(VSS),.VDD(VDD),.Y(g835),.A(g345));
  NOT NOT1_44(.VSS(VSS),.VDD(VDD),.Y(g836),.A(g349));
  NOT NOT1_45(.VSS(VSS),.VDD(VDD),.Y(g837),.A(g353));
  NOT NOT1_46(.VSS(VSS),.VDD(VDD),.Y(g838),.A(g564));
  NOT NOT1_47(.VSS(VSS),.VDD(VDD),.Y(g839),.A(g567));
  NOT NOT1_48(.VSS(VSS),.VDD(VDD),.Y(g842),.A(g571));
  NOT NOT1_49(.VSS(VSS),.VDD(VDD),.Y(g843),.A(g574));
  NOT NOT1_50(.VSS(VSS),.VDD(VDD),.Y(g844),.A(g578));
  NOT NOT1_51(.VSS(VSS),.VDD(VDD),.Y(g845),.A(g582));
  NOT NOT1_52(.VSS(VSS),.VDD(VDD),.Y(g846),.A(g586));
  NOT NOT1_53(.VSS(VSS),.VDD(VDD),.Y(g847),.A(g590));
  NOT NOT1_54(.VSS(VSS),.VDD(VDD),.Y(g848),.A(g594));
  NOT NOT1_55(.VSS(VSS),.VDD(VDD),.Y(g849),.A(g598));
  NOT NOT1_56(.VSS(VSS),.VDD(VDD),.Y(g850),.A(g602));
  NOT NOT1_57(.VSS(VSS),.VDD(VDD),.Y(g851),.A(g606));
  NOT NOT1_58(.VSS(VSS),.VDD(VDD),.Y(g852),.A(g634));
  NOT NOT1_59(.VSS(VSS),.VDD(VDD),.Y(g853),.A(g642));
  NOT NOT1_60(.VSS(VSS),.VDD(VDD),.Y(g854),.A(g646));
  NOT NOT1_61(.VSS(VSS),.VDD(VDD),.Y(g855),.A(g650));
  NOT NOT1_62(.VSS(VSS),.VDD(VDD),.Y(g856),.A(g654));
  NOT NOT1_63(.VSS(VSS),.VDD(VDD),.Y(g857),.A(g170));
  NOT NOT1_64(.VSS(VSS),.VDD(VDD),.Y(g858),.A(g301));
  NOT NOT1_65(.VSS(VSS),.VDD(VDD),.Y(g861),.A(g179));
  NOT NOT1_66(.VSS(VSS),.VDD(VDD),.Y(g862),.A(g319));
  NOT NOT1_67(.VSS(VSS),.VDD(VDD),.Y(g865),.A(g188));
  NOT NOT1_68(.VSS(VSS),.VDD(VDD),.Y(g866),.A(g314));
  NOT NOT1_69(.VSS(VSS),.VDD(VDD),.Y(g872),.A(g143));
  NOT NOT1_70(.VSS(VSS),.VDD(VDD),.Y(g873),.A(g306));
  NOT NOT1_71(.VSS(VSS),.VDD(VDD),.Y(g878),.A(g639));
  NOT NOT1_72(.VSS(VSS),.VDD(VDD),.Y(g889),.A(g310));
  NOT NOT1_73(.VSS(VSS),.VDD(VDD),.Y(g893),.A(g23));
  NOT NOT1_74(.VSS(VSS),.VDD(VDD),.Y(I1917),.A(g48));
  NOT NOT1_75(.VSS(VSS),.VDD(VDD),.Y(g894),.A(I1917));
  NOT NOT1_76(.VSS(VSS),.VDD(VDD),.Y(g895),.A(g139));
  NOT NOT1_77(.VSS(VSS),.VDD(VDD),.Y(g896),.A(g22));
  NOT NOT1_78(.VSS(VSS),.VDD(VDD),.Y(g897),.A(g41));
  NOT NOT1_79(.VSS(VSS),.VDD(VDD),.Y(g898),.A(g47));
  NOT NOT1_80(.VSS(VSS),.VDD(VDD),.Y(I1924),.A(g663));
  NOT NOT1_81(.VSS(VSS),.VDD(VDD),.Y(g899),.A(I1924));
  NOT NOT1_82(.VSS(VSS),.VDD(VDD),.Y(I1927),.A(g665));
  NOT NOT1_83(.VSS(VSS),.VDD(VDD),.Y(g900),.A(I1927));
  NOT NOT1_84(.VSS(VSS),.VDD(VDD),.Y(I1932),.A(g667));
  NOT NOT1_85(.VSS(VSS),.VDD(VDD),.Y(g908),.A(I1932));
  NOT NOT1_86(.VSS(VSS),.VDD(VDD),.Y(I1935),.A(g666));
  NOT NOT1_87(.VSS(VSS),.VDD(VDD),.Y(g909),.A(I1935));
  NOT NOT1_88(.VSS(VSS),.VDD(VDD),.Y(I1938),.A(g332));
  NOT NOT1_89(.VSS(VSS),.VDD(VDD),.Y(g910),.A(I1938));
  NOT NOT1_90(.VSS(VSS),.VDD(VDD),.Y(g913),.A(g658));
  NOT NOT1_91(.VSS(VSS),.VDD(VDD),.Y(I1942),.A(g664));
  NOT NOT1_92(.VSS(VSS),.VDD(VDD),.Y(g917),.A(I1942));
  NOT NOT1_93(.VSS(VSS),.VDD(VDD),.Y(g921),.A(g111));
  NOT NOT1_94(.VSS(VSS),.VDD(VDD),.Y(I1947),.A(g699));
  NOT NOT1_95(.VSS(VSS),.VDD(VDD),.Y(g922),.A(I1947));
  NOT NOT1_96(.VSS(VSS),.VDD(VDD),.Y(g923),.A(g332));
  NOT NOT1_97(.VSS(VSS),.VDD(VDD),.Y(I1958),.A(g702));
  NOT NOT1_98(.VSS(VSS),.VDD(VDD),.Y(g927),.A(I1958));
  NOT NOT1_99(.VSS(VSS),.VDD(VDD),.Y(g929),.A(g49));
  NOT NOT1_100(.VSS(VSS),.VDD(VDD),.Y(g931),.A(g54));
  NOT NOT1_101(.VSS(VSS),.VDD(VDD),.Y(g932),.A(g337));
  NOT NOT1_102(.VSS(VSS),.VDD(VDD),.Y(g938),.A(g59));
  NOT NOT1_103(.VSS(VSS),.VDD(VDD),.Y(g940),.A(g64));
  NOT NOT1_104(.VSS(VSS),.VDD(VDD),.Y(g942),.A(g69));
  NOT NOT1_105(.VSS(VSS),.VDD(VDD),.Y(g943),.A(g496));
  NOT NOT1_106(.VSS(VSS),.VDD(VDD),.Y(g945),.A(g536));
  NOT NOT1_107(.VSS(VSS),.VDD(VDD),.Y(g946),.A(g361));
  NOT NOT1_108(.VSS(VSS),.VDD(VDD),.Y(g947),.A(g74));
  NOT NOT1_109(.VSS(VSS),.VDD(VDD),.Y(g949),.A(g79));
  NOT NOT1_110(.VSS(VSS),.VDD(VDD),.Y(g951),.A(g84));
  NOT NOT1_111(.VSS(VSS),.VDD(VDD),.Y(I2029),.A(g677));
  NOT NOT1_112(.VSS(VSS),.VDD(VDD),.Y(g952),.A(I2029));
  NOT NOT1_113(.VSS(VSS),.VDD(VDD),.Y(g964),.A(g357));
  NOT NOT1_114(.VSS(VSS),.VDD(VDD),.Y(I2033),.A(g678));
  NOT NOT1_115(.VSS(VSS),.VDD(VDD),.Y(g965),.A(I2033));
  NOT NOT1_116(.VSS(VSS),.VDD(VDD),.Y(g971),.A(g658));
  NOT NOT1_117(.VSS(VSS),.VDD(VDD),.Y(I2037),.A(g679));
  NOT NOT1_118(.VSS(VSS),.VDD(VDD),.Y(g980),.A(I2037));
  NOT NOT1_119(.VSS(VSS),.VDD(VDD),.Y(g985),.A(g638));
  NOT NOT1_120(.VSS(VSS),.VDD(VDD),.Y(I2041),.A(g680));
  NOT NOT1_121(.VSS(VSS),.VDD(VDD),.Y(g996),.A(I2041));
  NOT NOT1_122(.VSS(VSS),.VDD(VDD),.Y(I2044),.A(g681));
  NOT NOT1_123(.VSS(VSS),.VDD(VDD),.Y(g1001),.A(I2044));
  NOT NOT1_124(.VSS(VSS),.VDD(VDD),.Y(I2047),.A(g682));
  NOT NOT1_125(.VSS(VSS),.VDD(VDD),.Y(g1006),.A(I2047));
  NOT NOT1_126(.VSS(VSS),.VDD(VDD),.Y(I2050),.A(g683));
  NOT NOT1_127(.VSS(VSS),.VDD(VDD),.Y(g1011),.A(I2050));
  NOT NOT1_128(.VSS(VSS),.VDD(VDD),.Y(I2053),.A(g684));
  NOT NOT1_129(.VSS(VSS),.VDD(VDD),.Y(g1017),.A(I2053));
  NOT NOT1_130(.VSS(VSS),.VDD(VDD),.Y(I2057),.A(g685));
  NOT NOT1_131(.VSS(VSS),.VDD(VDD),.Y(g1030),.A(I2057));
  NOT NOT1_132(.VSS(VSS),.VDD(VDD),.Y(I2067),.A(g686));
  NOT NOT1_133(.VSS(VSS),.VDD(VDD),.Y(g1037),.A(I2067));
  NOT NOT1_134(.VSS(VSS),.VDD(VDD),.Y(g1038),.A(g127));
  NOT NOT1_135(.VSS(VSS),.VDD(VDD),.Y(g1039),.A(g662));
  NOT NOT1_136(.VSS(VSS),.VDD(VDD),.Y(g1043),.A(g486));
  NOT NOT1_137(.VSS(VSS),.VDD(VDD),.Y(g1045),.A(g699));
  NOT NOT1_138(.VSS(VSS),.VDD(VDD),.Y(g1046),.A(g489));
  NOT NOT1_139(.VSS(VSS),.VDD(VDD),.Y(g1048),.A(g492));
  NOT NOT1_140(.VSS(VSS),.VDD(VDD),.Y(g1049),.A(g266));
  NOT NOT1_141(.VSS(VSS),.VDD(VDD),.Y(g1052),.A(g668));
  NOT NOT1_142(.VSS(VSS),.VDD(VDD),.Y(g1053),.A(g197));
  NOT NOT1_143(.VSS(VSS),.VDD(VDD),.Y(g1054),.A(g485));
  NOT NOT1_144(.VSS(VSS),.VDD(VDD),.Y(g1055),.A(g269));
  NOT NOT1_145(.VSS(VSS),.VDD(VDD),.Y(g1056),.A(g89));
  NOT NOT1_146(.VSS(VSS),.VDD(VDD),.Y(g1059),.A(g702));
  NOT NOT1_147(.VSS(VSS),.VDD(VDD),.Y(g1060),.A(g107));
  NOT NOT1_148(.VSS(VSS),.VDD(VDD),.Y(g1063),.A(g675));
  NOT NOT1_149(.VSS(VSS),.VDD(VDD),.Y(g1064),.A(g102));
  NOT NOT1_150(.VSS(VSS),.VDD(VDD),.Y(g1070),.A(g94));
  NOT NOT1_151(.VSS(VSS),.VDD(VDD),.Y(I2115),.A(g687));
  NOT NOT1_152(.VSS(VSS),.VDD(VDD),.Y(g1076),.A(I2115));
  NOT NOT1_153(.VSS(VSS),.VDD(VDD),.Y(g1084),.A(g98));
  NOT NOT1_154(.VSS(VSS),.VDD(VDD),.Y(I2119),.A(g688));
  NOT NOT1_155(.VSS(VSS),.VDD(VDD),.Y(g1088),.A(I2119));
  NOT NOT1_156(.VSS(VSS),.VDD(VDD),.Y(I2122),.A(g689));
  NOT NOT1_157(.VSS(VSS),.VDD(VDD),.Y(g1094),.A(I2122));
  NOT NOT1_158(.VSS(VSS),.VDD(VDD),.Y(I2125),.A(g698));
  NOT NOT1_159(.VSS(VSS),.VDD(VDD),.Y(g1101),.A(I2125));
  NOT NOT1_160(.VSS(VSS),.VDD(VDD),.Y(I2128),.A(g18));
  NOT NOT1_161(.VSS(VSS),.VDD(VDD),.Y(g1106),.A(I2128));
  NOT NOT1_162(.VSS(VSS),.VDD(VDD),.Y(I2131),.A(g24));
  NOT NOT1_163(.VSS(VSS),.VDD(VDD),.Y(g1107),.A(I2131));
  NOT NOT1_164(.VSS(VSS),.VDD(VDD),.Y(I2134),.A(g705));
  NOT NOT1_165(.VSS(VSS),.VDD(VDD),.Y(g1108),.A(I2134));
  NOT NOT1_166(.VSS(VSS),.VDD(VDD),.Y(I2137),.A(g1));
  NOT NOT1_167(.VSS(VSS),.VDD(VDD),.Y(g1109),.A(I2137));
  NOT NOT1_168(.VSS(VSS),.VDD(VDD),.Y(I2140),.A(g28));
  NOT NOT1_169(.VSS(VSS),.VDD(VDD),.Y(g1110),.A(I2140));
  NOT NOT1_170(.VSS(VSS),.VDD(VDD),.Y(I2143),.A(g2));
  NOT NOT1_171(.VSS(VSS),.VDD(VDD),.Y(g1111),.A(I2143));
  NOT NOT1_172(.VSS(VSS),.VDD(VDD),.Y(g1112),.A(g336));
  NOT NOT1_173(.VSS(VSS),.VDD(VDD),.Y(I2147),.A(g6));
  NOT NOT1_174(.VSS(VSS),.VDD(VDD),.Y(g1113),.A(I2147));
  NOT NOT1_175(.VSS(VSS),.VDD(VDD),.Y(I2150),.A(g10));
  NOT NOT1_176(.VSS(VSS),.VDD(VDD),.Y(g1114),.A(I2150));
  NOT NOT1_177(.VSS(VSS),.VDD(VDD),.Y(g1115),.A(g40));
  NOT NOT1_178(.VSS(VSS),.VDD(VDD),.Y(I2154),.A(g14));
  NOT NOT1_179(.VSS(VSS),.VDD(VDD),.Y(g1116),.A(I2154));
  NOT NOT1_180(.VSS(VSS),.VDD(VDD),.Y(g1117),.A(g32));
  NOT NOT1_181(.VSS(VSS),.VDD(VDD),.Y(g1118),.A(g36));
  NOT NOT1_182(.VSS(VSS),.VDD(VDD),.Y(I2159),.A(g465));
  NOT NOT1_183(.VSS(VSS),.VDD(VDD),.Y(g1119),.A(I2159));
  NOT NOT1_184(.VSS(VSS),.VDD(VDD),.Y(I2162),.A(g197));
  NOT NOT1_185(.VSS(VSS),.VDD(VDD),.Y(g1122),.A(I2162));
  NOT NOT1_186(.VSS(VSS),.VDD(VDD),.Y(I2165),.A(g690));
  NOT NOT1_187(.VSS(VSS),.VDD(VDD),.Y(g1123),.A(I2165));
  NOT NOT1_188(.VSS(VSS),.VDD(VDD),.Y(I2169),.A(g269));
  NOT NOT1_189(.VSS(VSS),.VDD(VDD),.Y(g1142),.A(I2169));
  NOT NOT1_190(.VSS(VSS),.VDD(VDD),.Y(I2172),.A(g691));
  NOT NOT1_191(.VSS(VSS),.VDD(VDD),.Y(g1143),.A(I2172));
  NOT NOT1_192(.VSS(VSS),.VDD(VDD),.Y(I2175),.A(g25));
  NOT NOT1_193(.VSS(VSS),.VDD(VDD),.Y(g1156),.A(I2175));
  NOT NOT1_194(.VSS(VSS),.VDD(VDD),.Y(I2179),.A(g293));
  NOT NOT1_195(.VSS(VSS),.VDD(VDD),.Y(g1160),.A(I2179));
  NOT NOT1_196(.VSS(VSS),.VDD(VDD),.Y(I2182),.A(g692));
  NOT NOT1_197(.VSS(VSS),.VDD(VDD),.Y(g1161),.A(I2182));
  NOT NOT1_198(.VSS(VSS),.VDD(VDD),.Y(I2185),.A(g29));
  NOT NOT1_199(.VSS(VSS),.VDD(VDD),.Y(g1173),.A(I2185));
  NOT NOT1_200(.VSS(VSS),.VDD(VDD),.Y(g1174),.A(g37));
  NOT NOT1_201(.VSS(VSS),.VDD(VDD),.Y(g1175),.A(g42));
  NOT NOT1_202(.VSS(VSS),.VDD(VDD),.Y(I2190),.A(g297));
  NOT NOT1_203(.VSS(VSS),.VDD(VDD),.Y(g1176),.A(I2190));
  NOT NOT1_204(.VSS(VSS),.VDD(VDD),.Y(I2193),.A(g693));
  NOT NOT1_205(.VSS(VSS),.VDD(VDD),.Y(g1177),.A(I2193));
  NOT NOT1_206(.VSS(VSS),.VDD(VDD),.Y(I2196),.A(g3));
  NOT NOT1_207(.VSS(VSS),.VDD(VDD),.Y(g1189),.A(I2196));
  NOT NOT1_208(.VSS(VSS),.VDD(VDD),.Y(I2199),.A(g33));
  NOT NOT1_209(.VSS(VSS),.VDD(VDD),.Y(g1190),.A(I2199));
  NOT NOT1_210(.VSS(VSS),.VDD(VDD),.Y(g1191),.A(g38));
  NOT NOT1_211(.VSS(VSS),.VDD(VDD),.Y(g1192),.A(g44));
  NOT NOT1_212(.VSS(VSS),.VDD(VDD),.Y(I2204),.A(g694));
  NOT NOT1_213(.VSS(VSS),.VDD(VDD),.Y(g1193),.A(I2204));
  NOT NOT1_214(.VSS(VSS),.VDD(VDD),.Y(I2207),.A(g7));
  NOT NOT1_215(.VSS(VSS),.VDD(VDD),.Y(g1203),.A(I2207));
  NOT NOT1_216(.VSS(VSS),.VDD(VDD),.Y(g1204),.A(g39));
  NOT NOT1_217(.VSS(VSS),.VDD(VDD),.Y(g1205),.A(g45));
  NOT NOT1_218(.VSS(VSS),.VDD(VDD),.Y(I2212),.A(g123));
  NOT NOT1_219(.VSS(VSS),.VDD(VDD),.Y(g1206),.A(I2212));
  NOT NOT1_220(.VSS(VSS),.VDD(VDD),.Y(I2215),.A(g695));
  NOT NOT1_221(.VSS(VSS),.VDD(VDD),.Y(g1209),.A(I2215));
  NOT NOT1_222(.VSS(VSS),.VDD(VDD),.Y(I2218),.A(g11));
  NOT NOT1_223(.VSS(VSS),.VDD(VDD),.Y(g1219),.A(I2218));
  NOT NOT1_224(.VSS(VSS),.VDD(VDD),.Y(I2221),.A(g43));
  NOT NOT1_225(.VSS(VSS),.VDD(VDD),.Y(g1220),.A(I2221));
  NOT NOT1_226(.VSS(VSS),.VDD(VDD),.Y(g1221),.A(g46));
  NOT NOT1_227(.VSS(VSS),.VDD(VDD),.Y(I2225),.A(g696));
  NOT NOT1_228(.VSS(VSS),.VDD(VDD),.Y(g1222),.A(I2225));
  NOT NOT1_229(.VSS(VSS),.VDD(VDD),.Y(I2228),.A(g15));
  NOT NOT1_230(.VSS(VSS),.VDD(VDD),.Y(g1232),.A(I2228));
  NOT NOT1_231(.VSS(VSS),.VDD(VDD),.Y(I2231),.A(g465));
  NOT NOT1_232(.VSS(VSS),.VDD(VDD),.Y(g1233),.A(I2231));
  NOT NOT1_233(.VSS(VSS),.VDD(VDD),.Y(I2234),.A(g697));
  NOT NOT1_234(.VSS(VSS),.VDD(VDD),.Y(g1236),.A(I2234));
  NOT NOT1_235(.VSS(VSS),.VDD(VDD),.Y(I2237),.A(g465));
  NOT NOT1_236(.VSS(VSS),.VDD(VDD),.Y(g1246),.A(I2237));
  NOT NOT1_237(.VSS(VSS),.VDD(VDD),.Y(I2240),.A(g19));
  NOT NOT1_238(.VSS(VSS),.VDD(VDD),.Y(g1249),.A(I2240));
  NOT NOT1_239(.VSS(VSS),.VDD(VDD),.Y(g1250),.A(g123));
  NOT NOT1_240(.VSS(VSS),.VDD(VDD),.Y(g1254),.A(g152));
  NOT NOT1_241(.VSS(VSS),.VDD(VDD),.Y(g1255),.A(g161));
  NOT NOT1_242(.VSS(VSS),.VDD(VDD),.Y(g1256),.A(g838));
  NOT NOT1_243(.VSS(VSS),.VDD(VDD),.Y(g1257),.A(g845));
  NOT NOT1_244(.VSS(VSS),.VDD(VDD),.Y(g1263),.A(g846));
  NOT NOT1_245(.VSS(VSS),.VDD(VDD),.Y(g1267),.A(g843));
  NOT NOT1_246(.VSS(VSS),.VDD(VDD),.Y(g1270),.A(g844));
  NOT NOT1_247(.VSS(VSS),.VDD(VDD),.Y(g1273),.A(g839));
  NOT NOT1_248(.VSS(VSS),.VDD(VDD),.Y(g1274),.A(g856));
  NOT NOT1_249(.VSS(VSS),.VDD(VDD),.Y(g1275),.A(g842));
  NOT NOT1_250(.VSS(VSS),.VDD(VDD),.Y(g1276),.A(g847));
  NOT NOT1_251(.VSS(VSS),.VDD(VDD),.Y(g1279),.A(g848));
  NOT NOT1_252(.VSS(VSS),.VDD(VDD),.Y(g1282),.A(g849));
  NOT NOT1_253(.VSS(VSS),.VDD(VDD),.Y(g1283),.A(g853));
  NOT NOT1_254(.VSS(VSS),.VDD(VDD),.Y(g1284),.A(g851));
  NOT NOT1_255(.VSS(VSS),.VDD(VDD),.Y(g1285),.A(g852));
  NOT NOT1_256(.VSS(VSS),.VDD(VDD),.Y(g1286),.A(g854));
  NOT NOT1_257(.VSS(VSS),.VDD(VDD),.Y(g1287),.A(g855));
  NOT NOT1_258(.VSS(VSS),.VDD(VDD),.Y(I2269),.A(g899));
  NOT NOT1_259(.VSS(VSS),.VDD(VDD),.Y(g1288),.A(I2269));
  NOT NOT1_260(.VSS(VSS),.VDD(VDD),.Y(I2272),.A(g908));
  NOT NOT1_261(.VSS(VSS),.VDD(VDD),.Y(g1289),.A(I2272));
  NOT NOT1_262(.VSS(VSS),.VDD(VDD),.Y(I2275),.A(g909));
  NOT NOT1_263(.VSS(VSS),.VDD(VDD),.Y(g1290),.A(I2275));
  NOT NOT1_264(.VSS(VSS),.VDD(VDD),.Y(I2278),.A(g917));
  NOT NOT1_265(.VSS(VSS),.VDD(VDD),.Y(g1291),.A(I2278));
  NOT NOT1_266(.VSS(VSS),.VDD(VDD),.Y(I2281),.A(g900));
  NOT NOT1_267(.VSS(VSS),.VDD(VDD),.Y(g1292),.A(I2281));
  NOT NOT1_268(.VSS(VSS),.VDD(VDD),.Y(I2284),.A(g922));
  NOT NOT1_269(.VSS(VSS),.VDD(VDD),.Y(g1293),.A(I2284));
  NOT NOT1_270(.VSS(VSS),.VDD(VDD),.Y(I2287),.A(g927));
  NOT NOT1_271(.VSS(VSS),.VDD(VDD),.Y(g1294),.A(I2287));
  NOT NOT1_272(.VSS(VSS),.VDD(VDD),.Y(I2290),.A(g971));
  NOT NOT1_273(.VSS(VSS),.VDD(VDD),.Y(g1295),.A(I2290));
  NOT NOT1_274(.VSS(VSS),.VDD(VDD),.Y(I2293),.A(g971));
  NOT NOT1_275(.VSS(VSS),.VDD(VDD),.Y(g1305),.A(I2293));
  NOT NOT1_276(.VSS(VSS),.VDD(VDD),.Y(I2296),.A(g893));
  NOT NOT1_277(.VSS(VSS),.VDD(VDD),.Y(g1315),.A(I2296));
  NOT NOT1_278(.VSS(VSS),.VDD(VDD),.Y(I2306),.A(g896));
  NOT NOT1_279(.VSS(VSS),.VDD(VDD),.Y(g1317),.A(I2306));
  NOT NOT1_280(.VSS(VSS),.VDD(VDD),.Y(I2309),.A(g1236));
  NOT NOT1_281(.VSS(VSS),.VDD(VDD),.Y(g1318),.A(I2309));
  NOT NOT1_282(.VSS(VSS),.VDD(VDD),.Y(I2312),.A(g897));
  NOT NOT1_283(.VSS(VSS),.VDD(VDD),.Y(g1319),.A(I2312));
  NOT NOT1_284(.VSS(VSS),.VDD(VDD),.Y(I2315),.A(g1222));
  NOT NOT1_285(.VSS(VSS),.VDD(VDD),.Y(g1320),.A(I2315));
  NOT NOT1_286(.VSS(VSS),.VDD(VDD),.Y(I2318),.A(g1236));
  NOT NOT1_287(.VSS(VSS),.VDD(VDD),.Y(g1321),.A(I2318));
  NOT NOT1_288(.VSS(VSS),.VDD(VDD),.Y(I2321),.A(g898));
  NOT NOT1_289(.VSS(VSS),.VDD(VDD),.Y(g1322),.A(I2321));
  NOT NOT1_290(.VSS(VSS),.VDD(VDD),.Y(I2324),.A(g1209));
  NOT NOT1_291(.VSS(VSS),.VDD(VDD),.Y(g1323),.A(I2324));
  NOT NOT1_292(.VSS(VSS),.VDD(VDD),.Y(I2327),.A(g1222));
  NOT NOT1_293(.VSS(VSS),.VDD(VDD),.Y(g1324),.A(I2327));
  NOT NOT1_294(.VSS(VSS),.VDD(VDD),.Y(I2330),.A(g1122));
  NOT NOT1_295(.VSS(VSS),.VDD(VDD),.Y(g1325),.A(I2330));
  NOT NOT1_296(.VSS(VSS),.VDD(VDD),.Y(g1326),.A(g894));
  NOT NOT1_297(.VSS(VSS),.VDD(VDD),.Y(I2334),.A(g1193));
  NOT NOT1_298(.VSS(VSS),.VDD(VDD),.Y(g1327),.A(I2334));
  NOT NOT1_299(.VSS(VSS),.VDD(VDD),.Y(I2337),.A(g1209));
  NOT NOT1_300(.VSS(VSS),.VDD(VDD),.Y(g1328),.A(I2337));
  NOT NOT1_301(.VSS(VSS),.VDD(VDD),.Y(I2340),.A(g1142));
  NOT NOT1_302(.VSS(VSS),.VDD(VDD),.Y(g1329),.A(I2340));
  NOT NOT1_303(.VSS(VSS),.VDD(VDD),.Y(I2343),.A(g1177));
  NOT NOT1_304(.VSS(VSS),.VDD(VDD),.Y(g1330),.A(I2343));
  NOT NOT1_305(.VSS(VSS),.VDD(VDD),.Y(I2346),.A(g1193));
  NOT NOT1_306(.VSS(VSS),.VDD(VDD),.Y(g1331),.A(I2346));
  NOT NOT1_307(.VSS(VSS),.VDD(VDD),.Y(I2349),.A(g1160));
  NOT NOT1_308(.VSS(VSS),.VDD(VDD),.Y(g1332),.A(I2349));
  NOT NOT1_309(.VSS(VSS),.VDD(VDD),.Y(I2352),.A(g1161));
  NOT NOT1_310(.VSS(VSS),.VDD(VDD),.Y(g1333),.A(I2352));
  NOT NOT1_311(.VSS(VSS),.VDD(VDD),.Y(I2355),.A(g1177));
  NOT NOT1_312(.VSS(VSS),.VDD(VDD),.Y(g1334),.A(I2355));
  NOT NOT1_313(.VSS(VSS),.VDD(VDD),.Y(I2358),.A(g1176));
  NOT NOT1_314(.VSS(VSS),.VDD(VDD),.Y(g1335),.A(I2358));
  NOT NOT1_315(.VSS(VSS),.VDD(VDD),.Y(I2361),.A(g1075));
  NOT NOT1_316(.VSS(VSS),.VDD(VDD),.Y(g1336),.A(I2361));
  NOT NOT1_317(.VSS(VSS),.VDD(VDD),.Y(I2364),.A(g1143));
  NOT NOT1_318(.VSS(VSS),.VDD(VDD),.Y(g1337),.A(I2364));
  NOT NOT1_319(.VSS(VSS),.VDD(VDD),.Y(I2367),.A(g1161));
  NOT NOT1_320(.VSS(VSS),.VDD(VDD),.Y(g1338),.A(I2367));
  NOT NOT1_321(.VSS(VSS),.VDD(VDD),.Y(I2370),.A(g1123));
  NOT NOT1_322(.VSS(VSS),.VDD(VDD),.Y(g1339),.A(I2370));
  NOT NOT1_323(.VSS(VSS),.VDD(VDD),.Y(I2373),.A(g1143));
  NOT NOT1_324(.VSS(VSS),.VDD(VDD),.Y(g1340),.A(I2373));
  NOT NOT1_325(.VSS(VSS),.VDD(VDD),.Y(I2376),.A(g729));
  NOT NOT1_326(.VSS(VSS),.VDD(VDD),.Y(g1341),.A(I2376));
  NOT NOT1_327(.VSS(VSS),.VDD(VDD),.Y(I2379),.A(g1123));
  NOT NOT1_328(.VSS(VSS),.VDD(VDD),.Y(g1344),.A(I2379));
  NOT NOT1_329(.VSS(VSS),.VDD(VDD),.Y(I2382),.A(g719));
  NOT NOT1_330(.VSS(VSS),.VDD(VDD),.Y(g1345),.A(I2382));
  NOT NOT1_331(.VSS(VSS),.VDD(VDD),.Y(I2385),.A(g784));
  NOT NOT1_332(.VSS(VSS),.VDD(VDD),.Y(g1348),.A(I2385));
  NOT NOT1_333(.VSS(VSS),.VDD(VDD),.Y(I2388),.A(g878));
  NOT NOT1_334(.VSS(VSS),.VDD(VDD),.Y(g1351),.A(I2388));
  NOT NOT1_335(.VSS(VSS),.VDD(VDD),.Y(I2391),.A(g774));
  NOT NOT1_336(.VSS(VSS),.VDD(VDD),.Y(g1352),.A(I2391));
  NOT NOT1_337(.VSS(VSS),.VDD(VDD),.Y(I2394),.A(g719));
  NOT NOT1_338(.VSS(VSS),.VDD(VDD),.Y(g1355),.A(I2394));
  NOT NOT1_339(.VSS(VSS),.VDD(VDD),.Y(g1358),.A(g1119));
  NOT NOT1_340(.VSS(VSS),.VDD(VDD),.Y(I2399),.A(g729));
  NOT NOT1_341(.VSS(VSS),.VDD(VDD),.Y(g1363),.A(I2399));
  NOT NOT1_342(.VSS(VSS),.VDD(VDD),.Y(I2402),.A(g774));
  NOT NOT1_343(.VSS(VSS),.VDD(VDD),.Y(g1366),.A(I2402));
  NOT NOT1_344(.VSS(VSS),.VDD(VDD),.Y(I2405),.A(g1112));
  NOT NOT1_345(.VSS(VSS),.VDD(VDD),.Y(g1369),.A(I2405));
  NOT NOT1_346(.VSS(VSS),.VDD(VDD),.Y(I2408),.A(g719));
  NOT NOT1_347(.VSS(VSS),.VDD(VDD),.Y(g1372),.A(I2408));
  NOT NOT1_348(.VSS(VSS),.VDD(VDD),.Y(I2411),.A(g736));
  NOT NOT1_349(.VSS(VSS),.VDD(VDD),.Y(g1375),.A(I2411));
  NOT NOT1_350(.VSS(VSS),.VDD(VDD),.Y(I2414),.A(g784));
  NOT NOT1_351(.VSS(VSS),.VDD(VDD),.Y(g1378),.A(I2414));
  NOT NOT1_352(.VSS(VSS),.VDD(VDD),.Y(I2417),.A(g774));
  NOT NOT1_353(.VSS(VSS),.VDD(VDD),.Y(g1381),.A(I2417));
  NOT NOT1_354(.VSS(VSS),.VDD(VDD),.Y(I2420),.A(g791));
  NOT NOT1_355(.VSS(VSS),.VDD(VDD),.Y(g1384),.A(I2420));
  NOT NOT1_356(.VSS(VSS),.VDD(VDD),.Y(I2424),.A(g719));
  NOT NOT1_357(.VSS(VSS),.VDD(VDD),.Y(g1391),.A(I2424));
  NOT NOT1_358(.VSS(VSS),.VDD(VDD),.Y(g1394),.A(g1206));
  NOT NOT1_359(.VSS(VSS),.VDD(VDD),.Y(I2428),.A(g774));
  NOT NOT1_360(.VSS(VSS),.VDD(VDD),.Y(g1395),.A(I2428));
  NOT NOT1_361(.VSS(VSS),.VDD(VDD),.Y(g1410),.A(g1233));
  NOT NOT1_362(.VSS(VSS),.VDD(VDD),.Y(g1415),.A(g1246));
  NOT NOT1_363(.VSS(VSS),.VDD(VDD),.Y(I2442),.A(g872));
  NOT NOT1_364(.VSS(VSS),.VDD(VDD),.Y(g1423),.A(I2442));
  NOT NOT1_365(.VSS(VSS),.VDD(VDD),.Y(I2445),.A(g971));
  NOT NOT1_366(.VSS(VSS),.VDD(VDD),.Y(g1426),.A(I2445));
  NOT NOT1_367(.VSS(VSS),.VDD(VDD),.Y(I2449),.A(g971));
  NOT NOT1_368(.VSS(VSS),.VDD(VDD),.Y(g1439),.A(I2449));
  NOT NOT1_369(.VSS(VSS),.VDD(VDD),.Y(I2453),.A(g952));
  NOT NOT1_370(.VSS(VSS),.VDD(VDD),.Y(g1450),.A(I2453));
  NOT NOT1_371(.VSS(VSS),.VDD(VDD),.Y(I2457),.A(g1253));
  NOT NOT1_372(.VSS(VSS),.VDD(VDD),.Y(g1460),.A(I2457));
  NOT NOT1_373(.VSS(VSS),.VDD(VDD),.Y(I2460),.A(g952));
  NOT NOT1_374(.VSS(VSS),.VDD(VDD),.Y(g1461),.A(I2460));
  NOT NOT1_375(.VSS(VSS),.VDD(VDD),.Y(I2464),.A(g850));
  NOT NOT1_376(.VSS(VSS),.VDD(VDD),.Y(g1471),.A(I2464));
  NOT NOT1_377(.VSS(VSS),.VDD(VDD),.Y(g1472),.A(g952));
  NOT NOT1_378(.VSS(VSS),.VDD(VDD),.Y(g1477),.A(g952));
  NOT NOT1_379(.VSS(VSS),.VDD(VDD),.Y(g1480),.A(g985));
  NOT NOT1_380(.VSS(VSS),.VDD(VDD),.Y(I2473),.A(g971));
  NOT NOT1_381(.VSS(VSS),.VDD(VDD),.Y(g1484),.A(I2473));
  NOT NOT1_382(.VSS(VSS),.VDD(VDD),.Y(I2476),.A(g971));
  NOT NOT1_383(.VSS(VSS),.VDD(VDD),.Y(g1491),.A(I2476));
  NOT NOT1_384(.VSS(VSS),.VDD(VDD),.Y(I2479),.A(g1049));
  NOT NOT1_385(.VSS(VSS),.VDD(VDD),.Y(g1498),.A(I2479));
  NOT NOT1_386(.VSS(VSS),.VDD(VDD),.Y(g1502),.A(g709));
  NOT NOT1_387(.VSS(VSS),.VDD(VDD),.Y(g1503),.A(g878));
  NOT NOT1_388(.VSS(VSS),.VDD(VDD),.Y(I2485),.A(g766));
  NOT NOT1_389(.VSS(VSS),.VDD(VDD),.Y(g1504),.A(I2485));
  NOT NOT1_390(.VSS(VSS),.VDD(VDD),.Y(g1513),.A(g878));
  NOT NOT1_391(.VSS(VSS),.VDD(VDD),.Y(I2491),.A(g821));
  NOT NOT1_392(.VSS(VSS),.VDD(VDD),.Y(g1519),.A(I2491));
  NOT NOT1_393(.VSS(VSS),.VDD(VDD),.Y(g1528),.A(g878));
  NOT NOT1_394(.VSS(VSS),.VDD(VDD),.Y(g1529),.A(g1076));
  NOT NOT1_395(.VSS(VSS),.VDD(VDD),.Y(g1533),.A(g878));
  NOT NOT1_396(.VSS(VSS),.VDD(VDD),.Y(g1535),.A(g1088));
  NOT NOT1_397(.VSS(VSS),.VDD(VDD),.Y(g1539),.A(g878));
  NOT NOT1_398(.VSS(VSS),.VDD(VDD),.Y(g1541),.A(g1094));
  NOT NOT1_399(.VSS(VSS),.VDD(VDD),.Y(g1542),.A(g878));
  NOT NOT1_400(.VSS(VSS),.VDD(VDD),.Y(g1543),.A(g1006));
  NOT NOT1_401(.VSS(VSS),.VDD(VDD),.Y(g1546),.A(g1101));
  NOT NOT1_402(.VSS(VSS),.VDD(VDD),.Y(g1549),.A(g878));
  NOT NOT1_403(.VSS(VSS),.VDD(VDD),.Y(g1550),.A(g996));
  NOT NOT1_404(.VSS(VSS),.VDD(VDD),.Y(g1551),.A(g1011));
  NOT NOT1_405(.VSS(VSS),.VDD(VDD),.Y(g1552),.A(g1030));
  NOT NOT1_406(.VSS(VSS),.VDD(VDD),.Y(I2521),.A(g1063));
  NOT NOT1_407(.VSS(VSS),.VDD(VDD),.Y(g1555),.A(I2521));
  NOT NOT1_408(.VSS(VSS),.VDD(VDD),.Y(g1556),.A(g878));
  NOT NOT1_409(.VSS(VSS),.VDD(VDD),.Y(g1557),.A(g1017));
  NOT NOT1_410(.VSS(VSS),.VDD(VDD),.Y(g1559),.A(g965));
  NOT NOT1_411(.VSS(VSS),.VDD(VDD),.Y(g1563),.A(g1006));
  NOT NOT1_412(.VSS(VSS),.VDD(VDD),.Y(g1564),.A(g1030));
  NOT NOT1_413(.VSS(VSS),.VDD(VDD),.Y(I2537),.A(g971));
  NOT NOT1_414(.VSS(VSS),.VDD(VDD),.Y(g1567),.A(I2537));
  NOT NOT1_415(.VSS(VSS),.VDD(VDD),.Y(g1577),.A(g1001));
  NOT NOT1_416(.VSS(VSS),.VDD(VDD),.Y(I2552),.A(g971));
  NOT NOT1_417(.VSS(VSS),.VDD(VDD),.Y(g1578),.A(I2552));
  NOT NOT1_418(.VSS(VSS),.VDD(VDD),.Y(g1581),.A(g910));
  NOT NOT1_419(.VSS(VSS),.VDD(VDD),.Y(g1583),.A(g1001));
  NOT NOT1_420(.VSS(VSS),.VDD(VDD),.Y(g1584),.A(g743));
  NOT NOT1_421(.VSS(VSS),.VDD(VDD),.Y(g1586),.A(g1052));
  NOT NOT1_422(.VSS(VSS),.VDD(VDD),.Y(g1587),.A(g1123));
  NOT NOT1_423(.VSS(VSS),.VDD(VDD),.Y(g1588),.A(g798));
  NOT NOT1_424(.VSS(VSS),.VDD(VDD),.Y(g1593),.A(g1054));
  NOT NOT1_425(.VSS(VSS),.VDD(VDD),.Y(g1594),.A(g1143));
  NOT NOT1_426(.VSS(VSS),.VDD(VDD),.Y(I2570),.A(g1222));
  NOT NOT1_427(.VSS(VSS),.VDD(VDD),.Y(g1608),.A(I2570));
  NOT NOT1_428(.VSS(VSS),.VDD(VDD),.Y(I2578),.A(g1209));
  NOT NOT1_429(.VSS(VSS),.VDD(VDD),.Y(g1623),.A(I2578));
  NOT NOT1_430(.VSS(VSS),.VDD(VDD),.Y(I2581),.A(g946));
  NOT NOT1_431(.VSS(VSS),.VDD(VDD),.Y(g1624),.A(I2581));
  NOT NOT1_432(.VSS(VSS),.VDD(VDD),.Y(I2584),.A(g839));
  NOT NOT1_433(.VSS(VSS),.VDD(VDD),.Y(g1627),.A(I2584));
  NOT NOT1_434(.VSS(VSS),.VDD(VDD),.Y(I2588),.A(g1193));
  NOT NOT1_435(.VSS(VSS),.VDD(VDD),.Y(g1631),.A(I2588));
  NOT NOT1_436(.VSS(VSS),.VDD(VDD),.Y(g1632),.A(g760));
  NOT NOT1_437(.VSS(VSS),.VDD(VDD),.Y(I2593),.A(g1177));
  NOT NOT1_438(.VSS(VSS),.VDD(VDD),.Y(g1636),.A(I2593));
  NOT NOT1_439(.VSS(VSS),.VDD(VDD),.Y(I2596),.A(g985));
  NOT NOT1_440(.VSS(VSS),.VDD(VDD),.Y(g1637),.A(I2596));
  NOT NOT1_441(.VSS(VSS),.VDD(VDD),.Y(g1638),.A(g754));
  NOT NOT1_442(.VSS(VSS),.VDD(VDD),.Y(g1639),.A(g815));
  NOT NOT1_443(.VSS(VSS),.VDD(VDD),.Y(I2601),.A(g1161));
  NOT NOT1_444(.VSS(VSS),.VDD(VDD),.Y(g1640),.A(I2601));
  NOT NOT1_445(.VSS(VSS),.VDD(VDD),.Y(I2604),.A(g1222));
  NOT NOT1_446(.VSS(VSS),.VDD(VDD),.Y(g1641),.A(I2604));
  NOT NOT1_447(.VSS(VSS),.VDD(VDD),.Y(g1642),.A(g809));
  NOT NOT1_448(.VSS(VSS),.VDD(VDD),.Y(I2608),.A(g1143));
  NOT NOT1_449(.VSS(VSS),.VDD(VDD),.Y(g1643),.A(I2608));
  NOT NOT1_450(.VSS(VSS),.VDD(VDD),.Y(I2611),.A(g1209));
  NOT NOT1_451(.VSS(VSS),.VDD(VDD),.Y(g1644),.A(I2611));
  NOT NOT1_452(.VSS(VSS),.VDD(VDD),.Y(I2614),.A(g1123));
  NOT NOT1_453(.VSS(VSS),.VDD(VDD),.Y(g1645),.A(I2614));
  NOT NOT1_454(.VSS(VSS),.VDD(VDD),.Y(I2617),.A(g1193));
  NOT NOT1_455(.VSS(VSS),.VDD(VDD),.Y(g1646),.A(I2617));
  NOT NOT1_456(.VSS(VSS),.VDD(VDD),.Y(I2620),.A(g1177));
  NOT NOT1_457(.VSS(VSS),.VDD(VDD),.Y(g1647),.A(I2620));
  NOT NOT1_458(.VSS(VSS),.VDD(VDD),.Y(I2623),.A(g1161));
  NOT NOT1_459(.VSS(VSS),.VDD(VDD),.Y(g1648),.A(I2623));
  NOT NOT1_460(.VSS(VSS),.VDD(VDD),.Y(g1649),.A(g985));
  NOT NOT1_461(.VSS(VSS),.VDD(VDD),.Y(I2627),.A(g1053));
  NOT NOT1_462(.VSS(VSS),.VDD(VDD),.Y(g1650),.A(I2627));
  NOT NOT1_463(.VSS(VSS),.VDD(VDD),.Y(I2630),.A(g1143));
  NOT NOT1_464(.VSS(VSS),.VDD(VDD),.Y(g1653),.A(I2630));
  NOT NOT1_465(.VSS(VSS),.VDD(VDD),.Y(g1654),.A(g878));
  NOT NOT1_466(.VSS(VSS),.VDD(VDD),.Y(g1655),.A(g985));
  NOT NOT1_467(.VSS(VSS),.VDD(VDD),.Y(I2635),.A(g1055));
  NOT NOT1_468(.VSS(VSS),.VDD(VDD),.Y(g1656),.A(I2635));
  NOT NOT1_469(.VSS(VSS),.VDD(VDD),.Y(I2638),.A(g1123));
  NOT NOT1_470(.VSS(VSS),.VDD(VDD),.Y(g1659),.A(I2638));
  NOT NOT1_471(.VSS(VSS),.VDD(VDD),.Y(g1660),.A(g985));
  NOT NOT1_472(.VSS(VSS),.VDD(VDD),.Y(g1661),.A(g1076));
  NOT NOT1_473(.VSS(VSS),.VDD(VDD),.Y(I2643),.A(g965));
  NOT NOT1_474(.VSS(VSS),.VDD(VDD),.Y(g1664),.A(I2643));
  NOT NOT1_475(.VSS(VSS),.VDD(VDD),.Y(g1665),.A(g985));
  NOT NOT1_476(.VSS(VSS),.VDD(VDD),.Y(g1666),.A(g1088));
  NOT NOT1_477(.VSS(VSS),.VDD(VDD),.Y(I2648),.A(g980));
  NOT NOT1_478(.VSS(VSS),.VDD(VDD),.Y(g1670),.A(I2648));
  NOT NOT1_479(.VSS(VSS),.VDD(VDD),.Y(g1671),.A(g985));
  NOT NOT1_480(.VSS(VSS),.VDD(VDD),.Y(g1672),.A(g1094));
  NOT NOT1_481(.VSS(VSS),.VDD(VDD),.Y(I2653),.A(g996));
  NOT NOT1_482(.VSS(VSS),.VDD(VDD),.Y(g1673),.A(I2653));
  NOT NOT1_483(.VSS(VSS),.VDD(VDD),.Y(g1674),.A(g985));
  NOT NOT1_484(.VSS(VSS),.VDD(VDD),.Y(g1675),.A(g1101));
  NOT NOT1_485(.VSS(VSS),.VDD(VDD),.Y(I2658),.A(g1001));
  NOT NOT1_486(.VSS(VSS),.VDD(VDD),.Y(g1678),.A(I2658));
  NOT NOT1_487(.VSS(VSS),.VDD(VDD),.Y(g1679),.A(g985));
  NOT NOT1_488(.VSS(VSS),.VDD(VDD),.Y(g1680),.A(g1011));
  NOT NOT1_489(.VSS(VSS),.VDD(VDD),.Y(I2663),.A(g1006));
  NOT NOT1_490(.VSS(VSS),.VDD(VDD),.Y(g1681),.A(I2663));
  NOT NOT1_491(.VSS(VSS),.VDD(VDD),.Y(g1682),.A(g829));
  NOT NOT1_492(.VSS(VSS),.VDD(VDD),.Y(g1683),.A(g1017));
  NOT NOT1_493(.VSS(VSS),.VDD(VDD),.Y(I2668),.A(g1011));
  NOT NOT1_494(.VSS(VSS),.VDD(VDD),.Y(g1684),.A(I2668));
  NOT NOT1_495(.VSS(VSS),.VDD(VDD),.Y(I2671),.A(g1017));
  NOT NOT1_496(.VSS(VSS),.VDD(VDD),.Y(g1685),.A(I2671));
  NOT NOT1_497(.VSS(VSS),.VDD(VDD),.Y(I2688),.A(g1030));
  NOT NOT1_498(.VSS(VSS),.VDD(VDD),.Y(g1688),.A(I2688));
  NOT NOT1_499(.VSS(VSS),.VDD(VDD),.Y(I2692),.A(g1037));
  NOT NOT1_500(.VSS(VSS),.VDD(VDD),.Y(g1690),.A(I2692));
  NOT NOT1_501(.VSS(VSS),.VDD(VDD),.Y(I2696),.A(g1156));
  NOT NOT1_502(.VSS(VSS),.VDD(VDD),.Y(g1692),.A(I2696));
  NOT NOT1_503(.VSS(VSS),.VDD(VDD),.Y(g1695),.A(g1106));
  NOT NOT1_504(.VSS(VSS),.VDD(VDD),.Y(I2700),.A(g1173));
  NOT NOT1_505(.VSS(VSS),.VDD(VDD),.Y(g1696),.A(I2700));
  NOT NOT1_506(.VSS(VSS),.VDD(VDD),.Y(I2703),.A(g1189));
  NOT NOT1_507(.VSS(VSS),.VDD(VDD),.Y(g1699),.A(I2703));
  NOT NOT1_508(.VSS(VSS),.VDD(VDD),.Y(g1702),.A(g1107));
  NOT NOT1_509(.VSS(VSS),.VDD(VDD),.Y(I2707),.A(g1190));
  NOT NOT1_510(.VSS(VSS),.VDD(VDD),.Y(g1703),.A(I2707));
  NOT NOT1_511(.VSS(VSS),.VDD(VDD),.Y(g1710),.A(g1109));
  NOT NOT1_512(.VSS(VSS),.VDD(VDD),.Y(I2712),.A(g1203));
  NOT NOT1_513(.VSS(VSS),.VDD(VDD),.Y(g1711),.A(I2712));
  NOT NOT1_514(.VSS(VSS),.VDD(VDD),.Y(g1714),.A(g1110));
  NOT NOT1_515(.VSS(VSS),.VDD(VDD),.Y(I2716),.A(g1115));
  NOT NOT1_516(.VSS(VSS),.VDD(VDD),.Y(g1715),.A(I2716));
  NOT NOT1_517(.VSS(VSS),.VDD(VDD),.Y(g1720),.A(g1111));
  NOT NOT1_518(.VSS(VSS),.VDD(VDD),.Y(I2721),.A(g1219));
  NOT NOT1_519(.VSS(VSS),.VDD(VDD),.Y(g1721),.A(I2721));
  NOT NOT1_520(.VSS(VSS),.VDD(VDD),.Y(I2724),.A(g1220));
  NOT NOT1_521(.VSS(VSS),.VDD(VDD),.Y(g1724),.A(I2724));
  NOT NOT1_522(.VSS(VSS),.VDD(VDD),.Y(g1725),.A(g1113));
  NOT NOT1_523(.VSS(VSS),.VDD(VDD),.Y(I2728),.A(g1232));
  NOT NOT1_524(.VSS(VSS),.VDD(VDD),.Y(g1726),.A(I2728));
  NOT NOT1_525(.VSS(VSS),.VDD(VDD),.Y(I2731),.A(g1117));
  NOT NOT1_526(.VSS(VSS),.VDD(VDD),.Y(g1729),.A(I2731));
  NOT NOT1_527(.VSS(VSS),.VDD(VDD),.Y(g1730),.A(g1114));
  NOT NOT1_528(.VSS(VSS),.VDD(VDD),.Y(I2735),.A(g1118));
  NOT NOT1_529(.VSS(VSS),.VDD(VDD),.Y(g1731),.A(I2735));
  NOT NOT1_530(.VSS(VSS),.VDD(VDD),.Y(I2738),.A(g1236));
  NOT NOT1_531(.VSS(VSS),.VDD(VDD),.Y(g1732),.A(I2738));
  NOT NOT1_532(.VSS(VSS),.VDD(VDD),.Y(I2741),.A(g1222));
  NOT NOT1_533(.VSS(VSS),.VDD(VDD),.Y(g1733),.A(I2741));
  NOT NOT1_534(.VSS(VSS),.VDD(VDD),.Y(g1734),.A(g952));
  NOT NOT1_535(.VSS(VSS),.VDD(VDD),.Y(I2745),.A(g1249));
  NOT NOT1_536(.VSS(VSS),.VDD(VDD),.Y(g1735),.A(I2745));
  NOT NOT1_537(.VSS(VSS),.VDD(VDD),.Y(g1738),.A(g1108));
  NOT NOT1_538(.VSS(VSS),.VDD(VDD),.Y(I2749),.A(g1209));
  NOT NOT1_539(.VSS(VSS),.VDD(VDD),.Y(g1739),.A(I2749));
  NOT NOT1_540(.VSS(VSS),.VDD(VDD),.Y(g1740),.A(g1116));
  NOT NOT1_541(.VSS(VSS),.VDD(VDD),.Y(I2753),.A(g1174));
  NOT NOT1_542(.VSS(VSS),.VDD(VDD),.Y(g1741),.A(I2753));
  NOT NOT1_543(.VSS(VSS),.VDD(VDD),.Y(I2756),.A(g1175));
  NOT NOT1_544(.VSS(VSS),.VDD(VDD),.Y(g1742),.A(I2756));
  NOT NOT1_545(.VSS(VSS),.VDD(VDD),.Y(I2760),.A(g1193));
  NOT NOT1_546(.VSS(VSS),.VDD(VDD),.Y(g1747),.A(I2760));
  NOT NOT1_547(.VSS(VSS),.VDD(VDD),.Y(I2763),.A(g1236));
  NOT NOT1_548(.VSS(VSS),.VDD(VDD),.Y(g1748),.A(I2763));
  NOT NOT1_549(.VSS(VSS),.VDD(VDD),.Y(I2773),.A(g1191));
  NOT NOT1_550(.VSS(VSS),.VDD(VDD),.Y(g1754),.A(I2773));
  NOT NOT1_551(.VSS(VSS),.VDD(VDD),.Y(I2776),.A(g1192));
  NOT NOT1_552(.VSS(VSS),.VDD(VDD),.Y(g1755),.A(I2776));
  NOT NOT1_553(.VSS(VSS),.VDD(VDD),.Y(I2779),.A(g1038));
  NOT NOT1_554(.VSS(VSS),.VDD(VDD),.Y(g1756),.A(I2779));
  NOT NOT1_555(.VSS(VSS),.VDD(VDD),.Y(I2782),.A(g1177));
  NOT NOT1_556(.VSS(VSS),.VDD(VDD),.Y(g1759),.A(I2782));
  NOT NOT1_557(.VSS(VSS),.VDD(VDD),.Y(I2785),.A(g1222));
  NOT NOT1_558(.VSS(VSS),.VDD(VDD),.Y(g1760),.A(I2785));
  NOT NOT1_559(.VSS(VSS),.VDD(VDD),.Y(I2788),.A(g1236));
  NOT NOT1_560(.VSS(VSS),.VDD(VDD),.Y(g1761),.A(I2788));
  NOT NOT1_561(.VSS(VSS),.VDD(VDD),.Y(I2791),.A(g1236));
  NOT NOT1_562(.VSS(VSS),.VDD(VDD),.Y(g1762),.A(I2791));
  NOT NOT1_563(.VSS(VSS),.VDD(VDD),.Y(I2802),.A(g1204));
  NOT NOT1_564(.VSS(VSS),.VDD(VDD),.Y(g1769),.A(I2802));
  NOT NOT1_565(.VSS(VSS),.VDD(VDD),.Y(I2805),.A(g1205));
  NOT NOT1_566(.VSS(VSS),.VDD(VDD),.Y(g1770),.A(I2805));
  NOT NOT1_567(.VSS(VSS),.VDD(VDD),.Y(I2808),.A(g1161));
  NOT NOT1_568(.VSS(VSS),.VDD(VDD),.Y(g1771),.A(I2808));
  NOT NOT1_569(.VSS(VSS),.VDD(VDD),.Y(I2811),.A(g1209));
  NOT NOT1_570(.VSS(VSS),.VDD(VDD),.Y(g1772),.A(I2811));
  NOT NOT1_571(.VSS(VSS),.VDD(VDD),.Y(I2814),.A(g1222));
  NOT NOT1_572(.VSS(VSS),.VDD(VDD),.Y(g1773),.A(I2814));
  NOT NOT1_573(.VSS(VSS),.VDD(VDD),.Y(I2817),.A(g1222));
  NOT NOT1_574(.VSS(VSS),.VDD(VDD),.Y(g1774),.A(I2817));
  NOT NOT1_575(.VSS(VSS),.VDD(VDD),.Y(g1775),.A(g952));
  NOT NOT1_576(.VSS(VSS),.VDD(VDD),.Y(I2821),.A(g1221));
  NOT NOT1_577(.VSS(VSS),.VDD(VDD),.Y(g1776),.A(I2821));
  NOT NOT1_578(.VSS(VSS),.VDD(VDD),.Y(I2825),.A(g1143));
  NOT NOT1_579(.VSS(VSS),.VDD(VDD),.Y(g1781),.A(I2825));
  NOT NOT1_580(.VSS(VSS),.VDD(VDD),.Y(I2828),.A(g1193));
  NOT NOT1_581(.VSS(VSS),.VDD(VDD),.Y(g1782),.A(I2828));
  NOT NOT1_582(.VSS(VSS),.VDD(VDD),.Y(I2831),.A(g1209));
  NOT NOT1_583(.VSS(VSS),.VDD(VDD),.Y(g1783),.A(I2831));
  NOT NOT1_584(.VSS(VSS),.VDD(VDD),.Y(I2835),.A(g1209));
  NOT NOT1_585(.VSS(VSS),.VDD(VDD),.Y(g1787),.A(I2835));
  NOT NOT1_586(.VSS(VSS),.VDD(VDD),.Y(g1788),.A(g985));
  NOT NOT1_587(.VSS(VSS),.VDD(VDD),.Y(I2839),.A(g1123));
  NOT NOT1_588(.VSS(VSS),.VDD(VDD),.Y(g1789),.A(I2839));
  NOT NOT1_589(.VSS(VSS),.VDD(VDD),.Y(I2842),.A(g1177));
  NOT NOT1_590(.VSS(VSS),.VDD(VDD),.Y(g1790),.A(I2842));
  NOT NOT1_591(.VSS(VSS),.VDD(VDD),.Y(I2845),.A(g1193));
  NOT NOT1_592(.VSS(VSS),.VDD(VDD),.Y(g1791),.A(I2845));
  NOT NOT1_593(.VSS(VSS),.VDD(VDD),.Y(I2848),.A(g1193));
  NOT NOT1_594(.VSS(VSS),.VDD(VDD),.Y(g1792),.A(I2848));
  NOT NOT1_595(.VSS(VSS),.VDD(VDD),.Y(I2854),.A(g1236));
  NOT NOT1_596(.VSS(VSS),.VDD(VDD),.Y(g1805),.A(I2854));
  NOT NOT1_597(.VSS(VSS),.VDD(VDD),.Y(I2857),.A(g1161));
  NOT NOT1_598(.VSS(VSS),.VDD(VDD),.Y(g1806),.A(I2857));
  NOT NOT1_599(.VSS(VSS),.VDD(VDD),.Y(I2860),.A(g1177));
  NOT NOT1_600(.VSS(VSS),.VDD(VDD),.Y(g1807),.A(I2860));
  NOT NOT1_601(.VSS(VSS),.VDD(VDD),.Y(I2864),.A(g1177));
  NOT NOT1_602(.VSS(VSS),.VDD(VDD),.Y(g1811),.A(I2864));
  NOT NOT1_603(.VSS(VSS),.VDD(VDD),.Y(I2867),.A(g1143));
  NOT NOT1_604(.VSS(VSS),.VDD(VDD),.Y(g1812),.A(I2867));
  NOT NOT1_605(.VSS(VSS),.VDD(VDD),.Y(I2870),.A(g1161));
  NOT NOT1_606(.VSS(VSS),.VDD(VDD),.Y(g1813),.A(I2870));
  NOT NOT1_607(.VSS(VSS),.VDD(VDD),.Y(I2873),.A(g1161));
  NOT NOT1_608(.VSS(VSS),.VDD(VDD),.Y(g1814),.A(I2873));
  NOT NOT1_609(.VSS(VSS),.VDD(VDD),.Y(I2877),.A(g1123));
  NOT NOT1_610(.VSS(VSS),.VDD(VDD),.Y(g1819),.A(I2877));
  NOT NOT1_611(.VSS(VSS),.VDD(VDD),.Y(I2880),.A(g1143));
  NOT NOT1_612(.VSS(VSS),.VDD(VDD),.Y(g1820),.A(I2880));
  NOT NOT1_613(.VSS(VSS),.VDD(VDD),.Y(I2883),.A(g1143));
  NOT NOT1_614(.VSS(VSS),.VDD(VDD),.Y(g1821),.A(I2883));
  NOT NOT1_615(.VSS(VSS),.VDD(VDD),.Y(I2887),.A(g1123));
  NOT NOT1_616(.VSS(VSS),.VDD(VDD),.Y(g1823),.A(I2887));
  NOT NOT1_617(.VSS(VSS),.VDD(VDD),.Y(I2890),.A(g1123));
  NOT NOT1_618(.VSS(VSS),.VDD(VDD),.Y(g1824),.A(I2890));
  NOT NOT1_619(.VSS(VSS),.VDD(VDD),.Y(I2893),.A(g1236));
  NOT NOT1_620(.VSS(VSS),.VDD(VDD),.Y(g1825),.A(I2893));
  NOT NOT1_621(.VSS(VSS),.VDD(VDD),.Y(I2904),.A(g1256));
  NOT NOT1_622(.VSS(VSS),.VDD(VDD),.Y(g1830),.A(I2904));
  NOT NOT1_623(.VSS(VSS),.VDD(VDD),.Y(I2907),.A(g1498));
  NOT NOT1_624(.VSS(VSS),.VDD(VDD),.Y(g1831),.A(I2907));
  NOT NOT1_625(.VSS(VSS),.VDD(VDD),.Y(I2910),.A(g1645));
  NOT NOT1_626(.VSS(VSS),.VDD(VDD),.Y(g1832),.A(I2910));
  NOT NOT1_627(.VSS(VSS),.VDD(VDD),.Y(I2913),.A(g1792));
  NOT NOT1_628(.VSS(VSS),.VDD(VDD),.Y(g1833),.A(I2913));
  NOT NOT1_629(.VSS(VSS),.VDD(VDD),.Y(I2916),.A(g1643));
  NOT NOT1_630(.VSS(VSS),.VDD(VDD),.Y(g1834),.A(I2916));
  NOT NOT1_631(.VSS(VSS),.VDD(VDD),.Y(I2919),.A(g1787));
  NOT NOT1_632(.VSS(VSS),.VDD(VDD),.Y(g1835),.A(I2919));
  NOT NOT1_633(.VSS(VSS),.VDD(VDD),.Y(I2922),.A(g1774));
  NOT NOT1_634(.VSS(VSS),.VDD(VDD),.Y(g1836),.A(I2922));
  NOT NOT1_635(.VSS(VSS),.VDD(VDD),.Y(I2925),.A(g1762));
  NOT NOT1_636(.VSS(VSS),.VDD(VDD),.Y(g1837),.A(I2925));
  NOT NOT1_637(.VSS(VSS),.VDD(VDD),.Y(g1838),.A(g1595));
  NOT NOT1_638(.VSS(VSS),.VDD(VDD),.Y(I2929),.A(g1659));
  NOT NOT1_639(.VSS(VSS),.VDD(VDD),.Y(g1841),.A(I2929));
  NOT NOT1_640(.VSS(VSS),.VDD(VDD),.Y(g1842),.A(g1612));
  NOT NOT1_641(.VSS(VSS),.VDD(VDD),.Y(I2940),.A(g1653));
  NOT NOT1_642(.VSS(VSS),.VDD(VDD),.Y(g1846),.A(I2940));
  NOT NOT1_643(.VSS(VSS),.VDD(VDD),.Y(I2943),.A(g1715));
  NOT NOT1_644(.VSS(VSS),.VDD(VDD),.Y(g1847),.A(I2943));
  NOT NOT1_645(.VSS(VSS),.VDD(VDD),.Y(I2946),.A(g1587));
  NOT NOT1_646(.VSS(VSS),.VDD(VDD),.Y(g1848),.A(I2946));
  NOT NOT1_647(.VSS(VSS),.VDD(VDD),.Y(I2949),.A(g1263));
  NOT NOT1_648(.VSS(VSS),.VDD(VDD),.Y(g1849),.A(I2949));
  NOT NOT1_649(.VSS(VSS),.VDD(VDD),.Y(I2952),.A(g1594));
  NOT NOT1_650(.VSS(VSS),.VDD(VDD),.Y(g1852),.A(I2952));
  NOT NOT1_651(.VSS(VSS),.VDD(VDD),.Y(I2955),.A(g1729));
  NOT NOT1_652(.VSS(VSS),.VDD(VDD),.Y(g1853),.A(I2955));
  NOT NOT1_653(.VSS(VSS),.VDD(VDD),.Y(I2958),.A(g1257));
  NOT NOT1_654(.VSS(VSS),.VDD(VDD),.Y(g1854),.A(I2958));
  NOT NOT1_655(.VSS(VSS),.VDD(VDD),.Y(I2961),.A(g1731));
  NOT NOT1_656(.VSS(VSS),.VDD(VDD),.Y(g1857),.A(I2961));
  NOT NOT1_657(.VSS(VSS),.VDD(VDD),.Y(I2964),.A(g1257));
  NOT NOT1_658(.VSS(VSS),.VDD(VDD),.Y(g1858),.A(I2964));
  NOT NOT1_659(.VSS(VSS),.VDD(VDD),.Y(I2967),.A(g1682));
  NOT NOT1_660(.VSS(VSS),.VDD(VDD),.Y(g1861),.A(I2967));
  NOT NOT1_661(.VSS(VSS),.VDD(VDD),.Y(I2970),.A(g1504));
  NOT NOT1_662(.VSS(VSS),.VDD(VDD),.Y(g1875),.A(I2970));
  NOT NOT1_663(.VSS(VSS),.VDD(VDD),.Y(I2973),.A(g1687));
  NOT NOT1_664(.VSS(VSS),.VDD(VDD),.Y(g1878),.A(I2973));
  NOT NOT1_665(.VSS(VSS),.VDD(VDD),.Y(g1880),.A(g1603));
  NOT NOT1_666(.VSS(VSS),.VDD(VDD),.Y(g1883),.A(g1797));
  NOT NOT1_667(.VSS(VSS),.VDD(VDD),.Y(I2979),.A(g1263));
  NOT NOT1_668(.VSS(VSS),.VDD(VDD),.Y(g1884),.A(I2979));
  NOT NOT1_669(.VSS(VSS),.VDD(VDD),.Y(I2982),.A(g1426));
  NOT NOT1_670(.VSS(VSS),.VDD(VDD),.Y(g1887),.A(I2982));
  NOT NOT1_671(.VSS(VSS),.VDD(VDD),.Y(g1890),.A(g1359));
  NOT NOT1_672(.VSS(VSS),.VDD(VDD),.Y(I2986),.A(g1504));
  NOT NOT1_673(.VSS(VSS),.VDD(VDD),.Y(g1891),.A(I2986));
  NOT NOT1_674(.VSS(VSS),.VDD(VDD),.Y(I2989),.A(g1519));
  NOT NOT1_675(.VSS(VSS),.VDD(VDD),.Y(g1894),.A(I2989));
  NOT NOT1_676(.VSS(VSS),.VDD(VDD),.Y(I2992),.A(g1741));
  NOT NOT1_677(.VSS(VSS),.VDD(VDD),.Y(g1897),.A(I2992));
  NOT NOT1_678(.VSS(VSS),.VDD(VDD),.Y(I2995),.A(g1742));
  NOT NOT1_679(.VSS(VSS),.VDD(VDD),.Y(g1898),.A(I2995));
  NOT NOT1_680(.VSS(VSS),.VDD(VDD),.Y(I2998),.A(g1257));
  NOT NOT1_681(.VSS(VSS),.VDD(VDD),.Y(g1899),.A(I2998));
  NOT NOT1_682(.VSS(VSS),.VDD(VDD),.Y(I3001),.A(g1267));
  NOT NOT1_683(.VSS(VSS),.VDD(VDD),.Y(g1902),.A(I3001));
  NOT NOT1_684(.VSS(VSS),.VDD(VDD),.Y(I3004),.A(g1426));
  NOT NOT1_685(.VSS(VSS),.VDD(VDD),.Y(g1905),.A(I3004));
  NOT NOT1_686(.VSS(VSS),.VDD(VDD),.Y(I3007),.A(g1439));
  NOT NOT1_687(.VSS(VSS),.VDD(VDD),.Y(g1908),.A(I3007));
  NOT NOT1_688(.VSS(VSS),.VDD(VDD),.Y(I3010),.A(g1504));
  NOT NOT1_689(.VSS(VSS),.VDD(VDD),.Y(g1911),.A(I3010));
  NOT NOT1_690(.VSS(VSS),.VDD(VDD),.Y(I3013),.A(g1519));
  NOT NOT1_691(.VSS(VSS),.VDD(VDD),.Y(g1914),.A(I3013));
  NOT NOT1_692(.VSS(VSS),.VDD(VDD),.Y(I3016),.A(g1754));
  NOT NOT1_693(.VSS(VSS),.VDD(VDD),.Y(g1917),.A(I3016));
  NOT NOT1_694(.VSS(VSS),.VDD(VDD),.Y(I3019),.A(g1755));
  NOT NOT1_695(.VSS(VSS),.VDD(VDD),.Y(g1918),.A(I3019));
  NOT NOT1_696(.VSS(VSS),.VDD(VDD),.Y(I3022),.A(g1426));
  NOT NOT1_697(.VSS(VSS),.VDD(VDD),.Y(g1919),.A(I3022));
  NOT NOT1_698(.VSS(VSS),.VDD(VDD),.Y(I3025),.A(g1439));
  NOT NOT1_699(.VSS(VSS),.VDD(VDD),.Y(g1922),.A(I3025));
  NOT NOT1_700(.VSS(VSS),.VDD(VDD),.Y(I3028),.A(g1504));
  NOT NOT1_701(.VSS(VSS),.VDD(VDD),.Y(g1925),.A(I3028));
  NOT NOT1_702(.VSS(VSS),.VDD(VDD),.Y(I3031),.A(g1504));
  NOT NOT1_703(.VSS(VSS),.VDD(VDD),.Y(g1928),.A(I3031));
  NOT NOT1_704(.VSS(VSS),.VDD(VDD),.Y(I3034),.A(g1519));
  NOT NOT1_705(.VSS(VSS),.VDD(VDD),.Y(g1931),.A(I3034));
  NOT NOT1_706(.VSS(VSS),.VDD(VDD),.Y(I3037),.A(g1769));
  NOT NOT1_707(.VSS(VSS),.VDD(VDD),.Y(g1934),.A(I3037));
  NOT NOT1_708(.VSS(VSS),.VDD(VDD),.Y(I3040),.A(g1770));
  NOT NOT1_709(.VSS(VSS),.VDD(VDD),.Y(g1935),.A(I3040));
  NOT NOT1_710(.VSS(VSS),.VDD(VDD),.Y(g1936),.A(g1756));
  NOT NOT1_711(.VSS(VSS),.VDD(VDD),.Y(I3044),.A(g1257));
  NOT NOT1_712(.VSS(VSS),.VDD(VDD),.Y(g1937),.A(I3044));
  NOT NOT1_713(.VSS(VSS),.VDD(VDD),.Y(I3047),.A(g1426));
  NOT NOT1_714(.VSS(VSS),.VDD(VDD),.Y(g1940),.A(I3047));
  NOT NOT1_715(.VSS(VSS),.VDD(VDD),.Y(I3050),.A(g1439));
  NOT NOT1_716(.VSS(VSS),.VDD(VDD),.Y(g1943),.A(I3050));
  NOT NOT1_717(.VSS(VSS),.VDD(VDD),.Y(I3053),.A(g1407));
  NOT NOT1_718(.VSS(VSS),.VDD(VDD),.Y(g1946),.A(I3053));
  NOT NOT1_719(.VSS(VSS),.VDD(VDD),.Y(I3056),.A(g1519));
  NOT NOT1_720(.VSS(VSS),.VDD(VDD),.Y(g1947),.A(I3056));
  NOT NOT1_721(.VSS(VSS),.VDD(VDD),.Y(I3059),.A(g1519));
  NOT NOT1_722(.VSS(VSS),.VDD(VDD),.Y(g1950),.A(I3059));
  NOT NOT1_723(.VSS(VSS),.VDD(VDD),.Y(I3062),.A(g1776));
  NOT NOT1_724(.VSS(VSS),.VDD(VDD),.Y(g1953),.A(I3062));
  NOT NOT1_725(.VSS(VSS),.VDD(VDD),.Y(I3065),.A(g1426));
  NOT NOT1_726(.VSS(VSS),.VDD(VDD),.Y(g1954),.A(I3065));
  NOT NOT1_727(.VSS(VSS),.VDD(VDD),.Y(I3068),.A(g1439));
  NOT NOT1_728(.VSS(VSS),.VDD(VDD),.Y(g1957),.A(I3068));
  NOT NOT1_729(.VSS(VSS),.VDD(VDD),.Y(I3071),.A(g1504));
  NOT NOT1_730(.VSS(VSS),.VDD(VDD),.Y(g1960),.A(I3071));
  NOT NOT1_731(.VSS(VSS),.VDD(VDD),.Y(I3074),.A(g1426));
  NOT NOT1_732(.VSS(VSS),.VDD(VDD),.Y(g1963),.A(I3074));
  NOT NOT1_733(.VSS(VSS),.VDD(VDD),.Y(I3077),.A(g1439));
  NOT NOT1_734(.VSS(VSS),.VDD(VDD),.Y(g1966),.A(I3077));
  NOT NOT1_735(.VSS(VSS),.VDD(VDD),.Y(I3080),.A(g1519));
  NOT NOT1_736(.VSS(VSS),.VDD(VDD),.Y(g1969),.A(I3080));
  NOT NOT1_737(.VSS(VSS),.VDD(VDD),.Y(I3083),.A(g1426));
  NOT NOT1_738(.VSS(VSS),.VDD(VDD),.Y(g1972),.A(I3083));
  NOT NOT1_739(.VSS(VSS),.VDD(VDD),.Y(I3086),.A(g1439));
  NOT NOT1_740(.VSS(VSS),.VDD(VDD),.Y(g1975),.A(I3086));
  NOT NOT1_741(.VSS(VSS),.VDD(VDD),.Y(g1978),.A(g1387));
  NOT NOT1_742(.VSS(VSS),.VDD(VDD),.Y(I3090),.A(g1504));
  NOT NOT1_743(.VSS(VSS),.VDD(VDD),.Y(g1979),.A(I3090));
  NOT NOT1_744(.VSS(VSS),.VDD(VDD),.Y(I3093),.A(g1426));
  NOT NOT1_745(.VSS(VSS),.VDD(VDD),.Y(g1982),.A(I3093));
  NOT NOT1_746(.VSS(VSS),.VDD(VDD),.Y(I3096),.A(g1439));
  NOT NOT1_747(.VSS(VSS),.VDD(VDD),.Y(g1985),.A(I3096));
  NOT NOT1_748(.VSS(VSS),.VDD(VDD),.Y(I3099),.A(g1519));
  NOT NOT1_749(.VSS(VSS),.VDD(VDD),.Y(g1988),.A(I3099));
  NOT NOT1_750(.VSS(VSS),.VDD(VDD),.Y(I3102),.A(g1426));
  NOT NOT1_751(.VSS(VSS),.VDD(VDD),.Y(g1991),.A(I3102));
  NOT NOT1_752(.VSS(VSS),.VDD(VDD),.Y(I3105),.A(g1439));
  NOT NOT1_753(.VSS(VSS),.VDD(VDD),.Y(g1994),.A(I3105));
  NOT NOT1_754(.VSS(VSS),.VDD(VDD),.Y(g1997),.A(g1398));
  NOT NOT1_755(.VSS(VSS),.VDD(VDD),.Y(I3109),.A(g1504));
  NOT NOT1_756(.VSS(VSS),.VDD(VDD),.Y(g1998),.A(I3109));
  NOT NOT1_757(.VSS(VSS),.VDD(VDD),.Y(I3112),.A(g1439));
  NOT NOT1_758(.VSS(VSS),.VDD(VDD),.Y(g2001),.A(I3112));
  NOT NOT1_759(.VSS(VSS),.VDD(VDD),.Y(I3115),.A(g1519));
  NOT NOT1_760(.VSS(VSS),.VDD(VDD),.Y(g2004),.A(I3115));
  NOT NOT1_761(.VSS(VSS),.VDD(VDD),.Y(g2007),.A(g1411));
  NOT NOT1_762(.VSS(VSS),.VDD(VDD),.Y(g2025),.A(g1276));
  NOT NOT1_763(.VSS(VSS),.VDD(VDD),.Y(I3134),.A(g1336));
  NOT NOT1_764(.VSS(VSS),.VDD(VDD),.Y(g2029),.A(I3134));
  NOT NOT1_765(.VSS(VSS),.VDD(VDD),.Y(I3137),.A(g1315));
  NOT NOT1_766(.VSS(VSS),.VDD(VDD),.Y(g2030),.A(I3137));
  NOT NOT1_767(.VSS(VSS),.VDD(VDD),.Y(I3140),.A(g1317));
  NOT NOT1_768(.VSS(VSS),.VDD(VDD),.Y(g2031),.A(I3140));
  NOT NOT1_769(.VSS(VSS),.VDD(VDD),.Y(g2032),.A(g1749));
  NOT NOT1_770(.VSS(VSS),.VDD(VDD),.Y(I3144),.A(g1319));
  NOT NOT1_771(.VSS(VSS),.VDD(VDD),.Y(g2035),.A(I3144));
  NOT NOT1_772(.VSS(VSS),.VDD(VDD),.Y(g2036),.A(g1764));
  NOT NOT1_773(.VSS(VSS),.VDD(VDD),.Y(I3148),.A(g1595));
  NOT NOT1_774(.VSS(VSS),.VDD(VDD),.Y(g2039),.A(I3148));
  NOT NOT1_775(.VSS(VSS),.VDD(VDD),.Y(g2040),.A(g1738));
  NOT NOT1_776(.VSS(VSS),.VDD(VDD),.Y(I3152),.A(g1322));
  NOT NOT1_777(.VSS(VSS),.VDD(VDD),.Y(g2041),.A(I3152));
  NOT NOT1_778(.VSS(VSS),.VDD(VDD),.Y(I3155),.A(g1612));
  NOT NOT1_779(.VSS(VSS),.VDD(VDD),.Y(g2042),.A(I3155));
  NOT NOT1_780(.VSS(VSS),.VDD(VDD),.Y(I3158),.A(g1829));
  NOT NOT1_781(.VSS(VSS),.VDD(VDD),.Y(g2043),.A(I3158));
  NOT NOT1_782(.VSS(VSS),.VDD(VDD),.Y(I3161),.A(g1270));
  NOT NOT1_783(.VSS(VSS),.VDD(VDD),.Y(g2044),.A(I3161));
  NOT NOT1_784(.VSS(VSS),.VDD(VDD),.Y(g2059),.A(g1402));
  NOT NOT1_785(.VSS(VSS),.VDD(VDD),.Y(g2060),.A(g1369));
  NOT NOT1_786(.VSS(VSS),.VDD(VDD),.Y(g2066),.A(g1341));
  NOT NOT1_787(.VSS(VSS),.VDD(VDD),.Y(g2078),.A(g1345));
  NOT NOT1_788(.VSS(VSS),.VDD(VDD),.Y(g2079),.A(g1348));
  NOT NOT1_789(.VSS(VSS),.VDD(VDD),.Y(I3198),.A(g1819));
  NOT NOT1_790(.VSS(VSS),.VDD(VDD),.Y(g2086),.A(I3198));
  NOT NOT1_791(.VSS(VSS),.VDD(VDD),.Y(g2087),.A(g1352));
  NOT NOT1_792(.VSS(VSS),.VDD(VDD),.Y(I3202),.A(g1812));
  NOT NOT1_793(.VSS(VSS),.VDD(VDD),.Y(g2088),.A(I3202));
  NOT NOT1_794(.VSS(VSS),.VDD(VDD),.Y(I3206),.A(g1823));
  NOT NOT1_795(.VSS(VSS),.VDD(VDD),.Y(g2090),.A(I3206));
  NOT NOT1_796(.VSS(VSS),.VDD(VDD),.Y(g2091),.A(g1355));
  NOT NOT1_797(.VSS(VSS),.VDD(VDD),.Y(I3212),.A(g1806));
  NOT NOT1_798(.VSS(VSS),.VDD(VDD),.Y(g2096),.A(I3212));
  NOT NOT1_799(.VSS(VSS),.VDD(VDD),.Y(I3215),.A(g1820));
  NOT NOT1_800(.VSS(VSS),.VDD(VDD),.Y(g2097),.A(I3215));
  NOT NOT1_801(.VSS(VSS),.VDD(VDD),.Y(g2098),.A(g1363));
  NOT NOT1_802(.VSS(VSS),.VDD(VDD),.Y(g2099),.A(g1366));
  NOT NOT1_803(.VSS(VSS),.VDD(VDD),.Y(I3222),.A(g1790));
  NOT NOT1_804(.VSS(VSS),.VDD(VDD),.Y(g2102),.A(I3222));
  NOT NOT1_805(.VSS(VSS),.VDD(VDD),.Y(I3225),.A(g1813));
  NOT NOT1_806(.VSS(VSS),.VDD(VDD),.Y(g2103),.A(I3225));
  NOT NOT1_807(.VSS(VSS),.VDD(VDD),.Y(g2104),.A(g1372));
  NOT NOT1_808(.VSS(VSS),.VDD(VDD),.Y(g2105),.A(g1375));
  NOT NOT1_809(.VSS(VSS),.VDD(VDD),.Y(g2106),.A(g1378));
  NOT NOT1_810(.VSS(VSS),.VDD(VDD),.Y(I3232),.A(g1782));
  NOT NOT1_811(.VSS(VSS),.VDD(VDD),.Y(g2108),.A(I3232));
  NOT NOT1_812(.VSS(VSS),.VDD(VDD),.Y(I3235),.A(g1807));
  NOT NOT1_813(.VSS(VSS),.VDD(VDD),.Y(g2109),.A(I3235));
  NOT NOT1_814(.VSS(VSS),.VDD(VDD),.Y(g2110),.A(g1381));
  NOT NOT1_815(.VSS(VSS),.VDD(VDD),.Y(g2111),.A(g1384));
  NOT NOT1_816(.VSS(VSS),.VDD(VDD),.Y(I3240),.A(g1460));
  NOT NOT1_817(.VSS(VSS),.VDD(VDD),.Y(g2112),.A(I3240));
  NOT NOT1_818(.VSS(VSS),.VDD(VDD),.Y(I3244),.A(g1772));
  NOT NOT1_819(.VSS(VSS),.VDD(VDD),.Y(g2117),.A(I3244));
  NOT NOT1_820(.VSS(VSS),.VDD(VDD),.Y(I3247),.A(g1791));
  NOT NOT1_821(.VSS(VSS),.VDD(VDD),.Y(g2118),.A(I3247));
  NOT NOT1_822(.VSS(VSS),.VDD(VDD),.Y(g2119),.A(g1391));
  NOT NOT1_823(.VSS(VSS),.VDD(VDD),.Y(I3251),.A(g1471));
  NOT NOT1_824(.VSS(VSS),.VDD(VDD),.Y(g2120),.A(I3251));
  NOT NOT1_825(.VSS(VSS),.VDD(VDD),.Y(I3255),.A(g1650));
  NOT NOT1_826(.VSS(VSS),.VDD(VDD),.Y(g2125),.A(I3255));
  NOT NOT1_827(.VSS(VSS),.VDD(VDD),.Y(I3258),.A(g1760));
  NOT NOT1_828(.VSS(VSS),.VDD(VDD),.Y(g2134),.A(I3258));
  NOT NOT1_829(.VSS(VSS),.VDD(VDD),.Y(I3261),.A(g1783));
  NOT NOT1_830(.VSS(VSS),.VDD(VDD),.Y(g2135),.A(I3261));
  NOT NOT1_831(.VSS(VSS),.VDD(VDD),.Y(g2136),.A(g1395));
  NOT NOT1_832(.VSS(VSS),.VDD(VDD),.Y(I3268),.A(g1656));
  NOT NOT1_833(.VSS(VSS),.VDD(VDD),.Y(g2145),.A(I3268));
  NOT NOT1_834(.VSS(VSS),.VDD(VDD),.Y(I3271),.A(g1748));
  NOT NOT1_835(.VSS(VSS),.VDD(VDD),.Y(g2154),.A(I3271));
  NOT NOT1_836(.VSS(VSS),.VDD(VDD),.Y(I3274),.A(g1773));
  NOT NOT1_837(.VSS(VSS),.VDD(VDD),.Y(g2155),.A(I3274));
  NOT NOT1_838(.VSS(VSS),.VDD(VDD),.Y(I3278),.A(g1695));
  NOT NOT1_839(.VSS(VSS),.VDD(VDD),.Y(g2157),.A(I3278));
  NOT NOT1_840(.VSS(VSS),.VDD(VDD),.Y(I3281),.A(g1761));
  NOT NOT1_841(.VSS(VSS),.VDD(VDD),.Y(g2158),.A(I3281));
  NOT NOT1_842(.VSS(VSS),.VDD(VDD),.Y(I3284),.A(g1702));
  NOT NOT1_843(.VSS(VSS),.VDD(VDD),.Y(g2159),.A(I3284));
  NOT NOT1_844(.VSS(VSS),.VDD(VDD),.Y(I3288),.A(g1710));
  NOT NOT1_845(.VSS(VSS),.VDD(VDD),.Y(g2163),.A(I3288));
  NOT NOT1_846(.VSS(VSS),.VDD(VDD),.Y(I3291),.A(g1714));
  NOT NOT1_847(.VSS(VSS),.VDD(VDD),.Y(g2164),.A(I3291));
  NOT NOT1_848(.VSS(VSS),.VDD(VDD),.Y(I3294),.A(g1720));
  NOT NOT1_849(.VSS(VSS),.VDD(VDD),.Y(g2165),.A(I3294));
  NOT NOT1_850(.VSS(VSS),.VDD(VDD),.Y(I3298),.A(g1725));
  NOT NOT1_851(.VSS(VSS),.VDD(VDD),.Y(g2169),.A(I3298));
  NOT NOT1_852(.VSS(VSS),.VDD(VDD),.Y(I3301),.A(g1730));
  NOT NOT1_853(.VSS(VSS),.VDD(VDD),.Y(g2170),.A(I3301));
  NOT NOT1_854(.VSS(VSS),.VDD(VDD),.Y(I3304),.A(g1740));
  NOT NOT1_855(.VSS(VSS),.VDD(VDD),.Y(g2171),.A(I3304));
  NOT NOT1_856(.VSS(VSS),.VDD(VDD),.Y(I3307),.A(g1339));
  NOT NOT1_857(.VSS(VSS),.VDD(VDD),.Y(g2172),.A(I3307));
  NOT NOT1_858(.VSS(VSS),.VDD(VDD),.Y(I3310),.A(g1640));
  NOT NOT1_859(.VSS(VSS),.VDD(VDD),.Y(g2173),.A(I3310));
  NOT NOT1_860(.VSS(VSS),.VDD(VDD),.Y(I3313),.A(g1337));
  NOT NOT1_861(.VSS(VSS),.VDD(VDD),.Y(g2174),.A(I3313));
  NOT NOT1_862(.VSS(VSS),.VDD(VDD),.Y(I3316),.A(g1344));
  NOT NOT1_863(.VSS(VSS),.VDD(VDD),.Y(g2175),.A(I3316));
  NOT NOT1_864(.VSS(VSS),.VDD(VDD),.Y(I3319),.A(g1636));
  NOT NOT1_865(.VSS(VSS),.VDD(VDD),.Y(g2176),.A(I3319));
  NOT NOT1_866(.VSS(VSS),.VDD(VDD),.Y(I3322),.A(g1333));
  NOT NOT1_867(.VSS(VSS),.VDD(VDD),.Y(g2177),.A(I3322));
  NOT NOT1_868(.VSS(VSS),.VDD(VDD),.Y(I3325),.A(g1340));
  NOT NOT1_869(.VSS(VSS),.VDD(VDD),.Y(g2178),.A(I3325));
  NOT NOT1_870(.VSS(VSS),.VDD(VDD),.Y(I3328),.A(g1273));
  NOT NOT1_871(.VSS(VSS),.VDD(VDD),.Y(g2179),.A(I3328));
  NOT NOT1_872(.VSS(VSS),.VDD(VDD),.Y(I3331),.A(g1631));
  NOT NOT1_873(.VSS(VSS),.VDD(VDD),.Y(g2194),.A(I3331));
  NOT NOT1_874(.VSS(VSS),.VDD(VDD),.Y(I3334),.A(g1330));
  NOT NOT1_875(.VSS(VSS),.VDD(VDD),.Y(g2195),.A(I3334));
  NOT NOT1_876(.VSS(VSS),.VDD(VDD),.Y(I3337),.A(g1338));
  NOT NOT1_877(.VSS(VSS),.VDD(VDD),.Y(g2196),.A(I3337));
  NOT NOT1_878(.VSS(VSS),.VDD(VDD),.Y(I3340),.A(g1282));
  NOT NOT1_879(.VSS(VSS),.VDD(VDD),.Y(g2197),.A(I3340));
  NOT NOT1_880(.VSS(VSS),.VDD(VDD),.Y(I3343),.A(g1623));
  NOT NOT1_881(.VSS(VSS),.VDD(VDD),.Y(g2212),.A(I3343));
  NOT NOT1_882(.VSS(VSS),.VDD(VDD),.Y(I3346),.A(g1327));
  NOT NOT1_883(.VSS(VSS),.VDD(VDD),.Y(g2213),.A(I3346));
  NOT NOT1_884(.VSS(VSS),.VDD(VDD),.Y(I3349),.A(g1334));
  NOT NOT1_885(.VSS(VSS),.VDD(VDD),.Y(g2214),.A(I3349));
  NOT NOT1_886(.VSS(VSS),.VDD(VDD),.Y(I3352),.A(g1285));
  NOT NOT1_887(.VSS(VSS),.VDD(VDD),.Y(g2215),.A(I3352));
  NOT NOT1_888(.VSS(VSS),.VDD(VDD),.Y(I3355),.A(g1608));
  NOT NOT1_889(.VSS(VSS),.VDD(VDD),.Y(g2230),.A(I3355));
  NOT NOT1_890(.VSS(VSS),.VDD(VDD),.Y(I3358),.A(g1323));
  NOT NOT1_891(.VSS(VSS),.VDD(VDD),.Y(g2231),.A(I3358));
  NOT NOT1_892(.VSS(VSS),.VDD(VDD),.Y(I3361),.A(g1331));
  NOT NOT1_893(.VSS(VSS),.VDD(VDD),.Y(g2232),.A(I3361));
  NOT NOT1_894(.VSS(VSS),.VDD(VDD),.Y(I3364),.A(g1648));
  NOT NOT1_895(.VSS(VSS),.VDD(VDD),.Y(g2233),.A(I3364));
  NOT NOT1_896(.VSS(VSS),.VDD(VDD),.Y(I3367),.A(g1283));
  NOT NOT1_897(.VSS(VSS),.VDD(VDD),.Y(g2234),.A(I3367));
  NOT NOT1_898(.VSS(VSS),.VDD(VDD),.Y(I3370),.A(g1805));
  NOT NOT1_899(.VSS(VSS),.VDD(VDD),.Y(g2241),.A(I3370));
  NOT NOT1_900(.VSS(VSS),.VDD(VDD),.Y(I3373),.A(g1320));
  NOT NOT1_901(.VSS(VSS),.VDD(VDD),.Y(g2242),.A(I3373));
  NOT NOT1_902(.VSS(VSS),.VDD(VDD),.Y(I3376),.A(g1328));
  NOT NOT1_903(.VSS(VSS),.VDD(VDD),.Y(g2243),.A(I3376));
  NOT NOT1_904(.VSS(VSS),.VDD(VDD),.Y(I3379),.A(g1647));
  NOT NOT1_905(.VSS(VSS),.VDD(VDD),.Y(g2244),.A(I3379));
  NOT NOT1_906(.VSS(VSS),.VDD(VDD),.Y(I3382),.A(g1284));
  NOT NOT1_907(.VSS(VSS),.VDD(VDD),.Y(g2245),.A(I3382));
  NOT NOT1_908(.VSS(VSS),.VDD(VDD),.Y(I3385),.A(g1318));
  NOT NOT1_909(.VSS(VSS),.VDD(VDD),.Y(g2252),.A(I3385));
  NOT NOT1_910(.VSS(VSS),.VDD(VDD),.Y(I3388),.A(g1324));
  NOT NOT1_911(.VSS(VSS),.VDD(VDD),.Y(g2253),.A(I3388));
  NOT NOT1_912(.VSS(VSS),.VDD(VDD),.Y(I3391),.A(g1646));
  NOT NOT1_913(.VSS(VSS),.VDD(VDD),.Y(g2254),.A(I3391));
  NOT NOT1_914(.VSS(VSS),.VDD(VDD),.Y(I3395),.A(g1286));
  NOT NOT1_915(.VSS(VSS),.VDD(VDD),.Y(g2256),.A(I3395));
  NOT NOT1_916(.VSS(VSS),.VDD(VDD),.Y(I3405),.A(g1321));
  NOT NOT1_917(.VSS(VSS),.VDD(VDD),.Y(g2264),.A(I3405));
  NOT NOT1_918(.VSS(VSS),.VDD(VDD),.Y(I3408),.A(g1644));
  NOT NOT1_919(.VSS(VSS),.VDD(VDD),.Y(g2265),.A(I3408));
  NOT NOT1_920(.VSS(VSS),.VDD(VDD),.Y(I3419),.A(g1287));
  NOT NOT1_921(.VSS(VSS),.VDD(VDD),.Y(g2268),.A(I3419));
  NOT NOT1_922(.VSS(VSS),.VDD(VDD),.Y(I3422),.A(g1641));
  NOT NOT1_923(.VSS(VSS),.VDD(VDD),.Y(g2275),.A(I3422));
  NOT NOT1_924(.VSS(VSS),.VDD(VDD),.Y(I3425),.A(g1274));
  NOT NOT1_925(.VSS(VSS),.VDD(VDD),.Y(g2276),.A(I3425));
  NOT NOT1_926(.VSS(VSS),.VDD(VDD),.Y(I3428),.A(g1825));
  NOT NOT1_927(.VSS(VSS),.VDD(VDD),.Y(g2283),.A(I3428));
  NOT NOT1_928(.VSS(VSS),.VDD(VDD),.Y(I3431),.A(g1275));
  NOT NOT1_929(.VSS(VSS),.VDD(VDD),.Y(g2284),.A(I3431));
  NOT NOT1_930(.VSS(VSS),.VDD(VDD),.Y(I3434),.A(g1627));
  NOT NOT1_931(.VSS(VSS),.VDD(VDD),.Y(g2291),.A(I3434));
  NOT NOT1_932(.VSS(VSS),.VDD(VDD),.Y(g2293),.A(g1567));
  NOT NOT1_933(.VSS(VSS),.VDD(VDD),.Y(g2295),.A(g1578));
  NOT NOT1_934(.VSS(VSS),.VDD(VDD),.Y(I3441),.A(g1502));
  NOT NOT1_935(.VSS(VSS),.VDD(VDD),.Y(g2296),.A(I3441));
  NOT NOT1_936(.VSS(VSS),.VDD(VDD),.Y(g2306),.A(g1743));
  NOT NOT1_937(.VSS(VSS),.VDD(VDD),.Y(I3452),.A(g1450));
  NOT NOT1_938(.VSS(VSS),.VDD(VDD),.Y(g2308),.A(I3452));
  NOT NOT1_939(.VSS(VSS),.VDD(VDD),.Y(I3462),.A(g1450));
  NOT NOT1_940(.VSS(VSS),.VDD(VDD),.Y(g2312),.A(I3462));
  NOT NOT1_941(.VSS(VSS),.VDD(VDD),.Y(I3465),.A(g1724));
  NOT NOT1_942(.VSS(VSS),.VDD(VDD),.Y(g2315),.A(I3465));
  NOT NOT1_943(.VSS(VSS),.VDD(VDD),.Y(I3468),.A(g1802));
  NOT NOT1_944(.VSS(VSS),.VDD(VDD),.Y(g2316),.A(I3468));
  NOT NOT1_945(.VSS(VSS),.VDD(VDD),.Y(I3471),.A(g1450));
  NOT NOT1_946(.VSS(VSS),.VDD(VDD),.Y(g2317),.A(I3471));
  NOT NOT1_947(.VSS(VSS),.VDD(VDD),.Y(I3474),.A(g1450));
  NOT NOT1_948(.VSS(VSS),.VDD(VDD),.Y(g2320),.A(I3474));
  NOT NOT1_949(.VSS(VSS),.VDD(VDD),.Y(I3478),.A(g1450));
  NOT NOT1_950(.VSS(VSS),.VDD(VDD),.Y(g2324),.A(I3478));
  NOT NOT1_951(.VSS(VSS),.VDD(VDD),.Y(I3481),.A(g1461));
  NOT NOT1_952(.VSS(VSS),.VDD(VDD),.Y(g2327),.A(I3481));
  NOT NOT1_953(.VSS(VSS),.VDD(VDD),.Y(g2330),.A(g1777));
  NOT NOT1_954(.VSS(VSS),.VDD(VDD),.Y(I3485),.A(g1450));
  NOT NOT1_955(.VSS(VSS),.VDD(VDD),.Y(g2333),.A(I3485));
  NOT NOT1_956(.VSS(VSS),.VDD(VDD),.Y(I3488),.A(g1295));
  NOT NOT1_957(.VSS(VSS),.VDD(VDD),.Y(g2336),.A(I3488));
  NOT NOT1_958(.VSS(VSS),.VDD(VDD),.Y(I3493),.A(g1461));
  NOT NOT1_959(.VSS(VSS),.VDD(VDD),.Y(g2343),.A(I3493));
  NOT NOT1_960(.VSS(VSS),.VDD(VDD),.Y(I3496),.A(g1326));
  NOT NOT1_961(.VSS(VSS),.VDD(VDD),.Y(g2346),.A(I3496));
  NOT NOT1_962(.VSS(VSS),.VDD(VDD),.Y(I3499),.A(g1450));
  NOT NOT1_963(.VSS(VSS),.VDD(VDD),.Y(g2347),.A(I3499));
  NOT NOT1_964(.VSS(VSS),.VDD(VDD),.Y(I3502),.A(g1295));
  NOT NOT1_965(.VSS(VSS),.VDD(VDD),.Y(g2350),.A(I3502));
  NOT NOT1_966(.VSS(VSS),.VDD(VDD),.Y(I3505),.A(g1305));
  NOT NOT1_967(.VSS(VSS),.VDD(VDD),.Y(g2353),.A(I3505));
  NOT NOT1_968(.VSS(VSS),.VDD(VDD),.Y(I3509),.A(g1461));
  NOT NOT1_969(.VSS(VSS),.VDD(VDD),.Y(g2357),.A(I3509));
  NOT NOT1_970(.VSS(VSS),.VDD(VDD),.Y(g2360),.A(g1793));
  NOT NOT1_971(.VSS(VSS),.VDD(VDD),.Y(I3513),.A(g1450));
  NOT NOT1_972(.VSS(VSS),.VDD(VDD),.Y(g2361),.A(I3513));
  NOT NOT1_973(.VSS(VSS),.VDD(VDD),.Y(I3516),.A(g1295));
  NOT NOT1_974(.VSS(VSS),.VDD(VDD),.Y(g2364),.A(I3516));
  NOT NOT1_975(.VSS(VSS),.VDD(VDD),.Y(I3519),.A(g1305));
  NOT NOT1_976(.VSS(VSS),.VDD(VDD),.Y(g2367),.A(I3519));
  NOT NOT1_977(.VSS(VSS),.VDD(VDD),.Y(I3522),.A(g1664));
  NOT NOT1_978(.VSS(VSS),.VDD(VDD),.Y(g2370),.A(I3522));
  NOT NOT1_979(.VSS(VSS),.VDD(VDD),.Y(I3525),.A(g1461));
  NOT NOT1_980(.VSS(VSS),.VDD(VDD),.Y(g2378),.A(I3525));
  NOT NOT1_981(.VSS(VSS),.VDD(VDD),.Y(I3528),.A(g1422));
  NOT NOT1_982(.VSS(VSS),.VDD(VDD),.Y(g2381),.A(I3528));
  NOT NOT1_983(.VSS(VSS),.VDD(VDD),.Y(I3531),.A(g1593));
  NOT NOT1_984(.VSS(VSS),.VDD(VDD),.Y(g2390),.A(I3531));
  NOT NOT1_985(.VSS(VSS),.VDD(VDD),.Y(I3534),.A(g1295));
  NOT NOT1_986(.VSS(VSS),.VDD(VDD),.Y(g2391),.A(I3534));
  NOT NOT1_987(.VSS(VSS),.VDD(VDD),.Y(I3537),.A(g1305));
  NOT NOT1_988(.VSS(VSS),.VDD(VDD),.Y(g2394),.A(I3537));
  NOT NOT1_989(.VSS(VSS),.VDD(VDD),.Y(I3540),.A(g1670));
  NOT NOT1_990(.VSS(VSS),.VDD(VDD),.Y(g2397),.A(I3540));
  NOT NOT1_991(.VSS(VSS),.VDD(VDD),.Y(I3543),.A(g1461));
  NOT NOT1_992(.VSS(VSS),.VDD(VDD),.Y(g2405),.A(I3543));
  NOT NOT1_993(.VSS(VSS),.VDD(VDD),.Y(I3546),.A(g1586));
  NOT NOT1_994(.VSS(VSS),.VDD(VDD),.Y(g2408),.A(I3546));
  NOT NOT1_995(.VSS(VSS),.VDD(VDD),.Y(g2409),.A(g1815));
  NOT NOT1_996(.VSS(VSS),.VDD(VDD),.Y(I3550),.A(g1295));
  NOT NOT1_997(.VSS(VSS),.VDD(VDD),.Y(g2410),.A(I3550));
  NOT NOT1_998(.VSS(VSS),.VDD(VDD),.Y(I3553),.A(g1305));
  NOT NOT1_999(.VSS(VSS),.VDD(VDD),.Y(g2413),.A(I3553));
  NOT NOT1_1000(.VSS(VSS),.VDD(VDD),.Y(I3556),.A(g1484));
  NOT NOT1_1001(.VSS(VSS),.VDD(VDD),.Y(g2416),.A(I3556));
  NOT NOT1_1002(.VSS(VSS),.VDD(VDD),.Y(I3560),.A(g1673));
  NOT NOT1_1003(.VSS(VSS),.VDD(VDD),.Y(g2422),.A(I3560));
  NOT NOT1_1004(.VSS(VSS),.VDD(VDD),.Y(I3563),.A(g1461));
  NOT NOT1_1005(.VSS(VSS),.VDD(VDD),.Y(g2430),.A(I3563));
  NOT NOT1_1006(.VSS(VSS),.VDD(VDD),.Y(I3569),.A(g1789));
  NOT NOT1_1007(.VSS(VSS),.VDD(VDD),.Y(g2436),.A(I3569));
  NOT NOT1_1008(.VSS(VSS),.VDD(VDD),.Y(I3572),.A(g1295));
  NOT NOT1_1009(.VSS(VSS),.VDD(VDD),.Y(g2437),.A(I3572));
  NOT NOT1_1010(.VSS(VSS),.VDD(VDD),.Y(I3575),.A(g1305));
  NOT NOT1_1011(.VSS(VSS),.VDD(VDD),.Y(g2440),.A(I3575));
  NOT NOT1_1012(.VSS(VSS),.VDD(VDD),.Y(I3578),.A(g1484));
  NOT NOT1_1013(.VSS(VSS),.VDD(VDD),.Y(g2443),.A(I3578));
  NOT NOT1_1014(.VSS(VSS),.VDD(VDD),.Y(I3581),.A(g1491));
  NOT NOT1_1015(.VSS(VSS),.VDD(VDD),.Y(g2446),.A(I3581));
  NOT NOT1_1016(.VSS(VSS),.VDD(VDD),.Y(I3584),.A(g1678));
  NOT NOT1_1017(.VSS(VSS),.VDD(VDD),.Y(g2449),.A(I3584));
  NOT NOT1_1018(.VSS(VSS),.VDD(VDD),.Y(I3587),.A(g1461));
  NOT NOT1_1019(.VSS(VSS),.VDD(VDD),.Y(g2457),.A(I3587));
  NOT NOT1_1020(.VSS(VSS),.VDD(VDD),.Y(I3590),.A(g1781));
  NOT NOT1_1021(.VSS(VSS),.VDD(VDD),.Y(g2460),.A(I3590));
  NOT NOT1_1022(.VSS(VSS),.VDD(VDD),.Y(I3593),.A(g1295));
  NOT NOT1_1023(.VSS(VSS),.VDD(VDD),.Y(g2461),.A(I3593));
  NOT NOT1_1024(.VSS(VSS),.VDD(VDD),.Y(I3596),.A(g1305));
  NOT NOT1_1025(.VSS(VSS),.VDD(VDD),.Y(g2464),.A(I3596));
  NOT NOT1_1026(.VSS(VSS),.VDD(VDD),.Y(I3599),.A(g1484));
  NOT NOT1_1027(.VSS(VSS),.VDD(VDD),.Y(g2467),.A(I3599));
  NOT NOT1_1028(.VSS(VSS),.VDD(VDD),.Y(I3602),.A(g1491));
  NOT NOT1_1029(.VSS(VSS),.VDD(VDD),.Y(g2470),.A(I3602));
  NOT NOT1_1030(.VSS(VSS),.VDD(VDD),.Y(I3605),.A(g1681));
  NOT NOT1_1031(.VSS(VSS),.VDD(VDD),.Y(g2473),.A(I3605));
  NOT NOT1_1032(.VSS(VSS),.VDD(VDD),.Y(I3608),.A(g1461));
  NOT NOT1_1033(.VSS(VSS),.VDD(VDD),.Y(g2481),.A(I3608));
  NOT NOT1_1034(.VSS(VSS),.VDD(VDD),.Y(I3611),.A(g1771));
  NOT NOT1_1035(.VSS(VSS),.VDD(VDD),.Y(g2484),.A(I3611));
  NOT NOT1_1036(.VSS(VSS),.VDD(VDD),.Y(I3614),.A(g1295));
  NOT NOT1_1037(.VSS(VSS),.VDD(VDD),.Y(g2485),.A(I3614));
  NOT NOT1_1038(.VSS(VSS),.VDD(VDD),.Y(I3617),.A(g1305));
  NOT NOT1_1039(.VSS(VSS),.VDD(VDD),.Y(g2488),.A(I3617));
  NOT NOT1_1040(.VSS(VSS),.VDD(VDD),.Y(I3620),.A(g1484));
  NOT NOT1_1041(.VSS(VSS),.VDD(VDD),.Y(g2491),.A(I3620));
  NOT NOT1_1042(.VSS(VSS),.VDD(VDD),.Y(I3623),.A(g1491));
  NOT NOT1_1043(.VSS(VSS),.VDD(VDD),.Y(g2494),.A(I3623));
  NOT NOT1_1044(.VSS(VSS),.VDD(VDD),.Y(I3626),.A(g1684));
  NOT NOT1_1045(.VSS(VSS),.VDD(VDD),.Y(g2497),.A(I3626));
  NOT NOT1_1046(.VSS(VSS),.VDD(VDD),.Y(I3629),.A(g1759));
  NOT NOT1_1047(.VSS(VSS),.VDD(VDD),.Y(g2505),.A(I3629));
  NOT NOT1_1048(.VSS(VSS),.VDD(VDD),.Y(I3632),.A(g1295));
  NOT NOT1_1049(.VSS(VSS),.VDD(VDD),.Y(g2506),.A(I3632));
  NOT NOT1_1050(.VSS(VSS),.VDD(VDD),.Y(I3635),.A(g1305));
  NOT NOT1_1051(.VSS(VSS),.VDD(VDD),.Y(g2509),.A(I3635));
  NOT NOT1_1052(.VSS(VSS),.VDD(VDD),.Y(I3638),.A(g1484));
  NOT NOT1_1053(.VSS(VSS),.VDD(VDD),.Y(g2512),.A(I3638));
  NOT NOT1_1054(.VSS(VSS),.VDD(VDD),.Y(I3641),.A(g1491));
  NOT NOT1_1055(.VSS(VSS),.VDD(VDD),.Y(g2515),.A(I3641));
  NOT NOT1_1056(.VSS(VSS),.VDD(VDD),.Y(I3644),.A(g1685));
  NOT NOT1_1057(.VSS(VSS),.VDD(VDD),.Y(g2518),.A(I3644));
  NOT NOT1_1058(.VSS(VSS),.VDD(VDD),.Y(I3647),.A(g1747));
  NOT NOT1_1059(.VSS(VSS),.VDD(VDD),.Y(g2524),.A(I3647));
  NOT NOT1_1060(.VSS(VSS),.VDD(VDD),.Y(I3650),.A(g1650));
  NOT NOT1_1061(.VSS(VSS),.VDD(VDD),.Y(g2525),.A(I3650));
  NOT NOT1_1062(.VSS(VSS),.VDD(VDD),.Y(I3653),.A(g1305));
  NOT NOT1_1063(.VSS(VSS),.VDD(VDD),.Y(g2535),.A(I3653));
  NOT NOT1_1064(.VSS(VSS),.VDD(VDD),.Y(I3656),.A(g1484));
  NOT NOT1_1065(.VSS(VSS),.VDD(VDD),.Y(g2538),.A(I3656));
  NOT NOT1_1066(.VSS(VSS),.VDD(VDD),.Y(I3659),.A(g1491));
  NOT NOT1_1067(.VSS(VSS),.VDD(VDD),.Y(g2541),.A(I3659));
  NOT NOT1_1068(.VSS(VSS),.VDD(VDD),.Y(I3662),.A(g1688));
  NOT NOT1_1069(.VSS(VSS),.VDD(VDD),.Y(g2544),.A(I3662));
  NOT NOT1_1070(.VSS(VSS),.VDD(VDD),.Y(I3665),.A(g1824));
  NOT NOT1_1071(.VSS(VSS),.VDD(VDD),.Y(g2550),.A(I3665));
  NOT NOT1_1072(.VSS(VSS),.VDD(VDD),.Y(I3669),.A(g1739));
  NOT NOT1_1073(.VSS(VSS),.VDD(VDD),.Y(g2554),.A(I3669));
  NOT NOT1_1074(.VSS(VSS),.VDD(VDD),.Y(I3672),.A(g1656));
  NOT NOT1_1075(.VSS(VSS),.VDD(VDD),.Y(g2555),.A(I3672));
  NOT NOT1_1076(.VSS(VSS),.VDD(VDD),.Y(I3675),.A(g1491));
  NOT NOT1_1077(.VSS(VSS),.VDD(VDD),.Y(g2565),.A(I3675));
  NOT NOT1_1078(.VSS(VSS),.VDD(VDD),.Y(I3678),.A(g1690));
  NOT NOT1_1079(.VSS(VSS),.VDD(VDD),.Y(g2568),.A(I3678));
  NOT NOT1_1080(.VSS(VSS),.VDD(VDD),.Y(I3681),.A(g1821));
  NOT NOT1_1081(.VSS(VSS),.VDD(VDD),.Y(g2574),.A(I3681));
  NOT NOT1_1082(.VSS(VSS),.VDD(VDD),.Y(I3684),.A(g1733));
  NOT NOT1_1083(.VSS(VSS),.VDD(VDD),.Y(g2575),.A(I3684));
  NOT NOT1_1084(.VSS(VSS),.VDD(VDD),.Y(I3687),.A(g1814));
  NOT NOT1_1085(.VSS(VSS),.VDD(VDD),.Y(g2576),.A(I3687));
  NOT NOT1_1086(.VSS(VSS),.VDD(VDD),.Y(I3691),.A(g1732));
  NOT NOT1_1087(.VSS(VSS),.VDD(VDD),.Y(g2580),.A(I3691));
  NOT NOT1_1088(.VSS(VSS),.VDD(VDD),.Y(I3694),.A(g1811));
  NOT NOT1_1089(.VSS(VSS),.VDD(VDD),.Y(g2581),.A(I3694));
  NOT NOT1_1090(.VSS(VSS),.VDD(VDD),.Y(g2583),.A(g1830));
  NOT NOT1_1091(.VSS(VSS),.VDD(VDD),.Y(I3705),.A(g2316));
  NOT NOT1_1092(.VSS(VSS),.VDD(VDD),.Y(g2584),.A(I3705));
  NOT NOT1_1093(.VSS(VSS),.VDD(VDD),.Y(I3708),.A(g1946));
  NOT NOT1_1094(.VSS(VSS),.VDD(VDD),.Y(g2585),.A(I3708));
  NOT NOT1_1095(.VSS(VSS),.VDD(VDD),.Y(I3711),.A(g1848));
  NOT NOT1_1096(.VSS(VSS),.VDD(VDD),.Y(g2586),.A(I3711));
  NOT NOT1_1097(.VSS(VSS),.VDD(VDD),.Y(I3714),.A(g1852));
  NOT NOT1_1098(.VSS(VSS),.VDD(VDD),.Y(g2587),.A(I3714));
  NOT NOT1_1099(.VSS(VSS),.VDD(VDD),.Y(I3717),.A(g2154));
  NOT NOT1_1100(.VSS(VSS),.VDD(VDD),.Y(g2588),.A(I3717));
  NOT NOT1_1101(.VSS(VSS),.VDD(VDD),.Y(I3720),.A(g2155));
  NOT NOT1_1102(.VSS(VSS),.VDD(VDD),.Y(g2591),.A(I3720));
  NOT NOT1_1103(.VSS(VSS),.VDD(VDD),.Y(I3723),.A(g2158));
  NOT NOT1_1104(.VSS(VSS),.VDD(VDD),.Y(g2594),.A(I3723));
  NOT NOT1_1105(.VSS(VSS),.VDD(VDD),.Y(I3726),.A(g2030));
  NOT NOT1_1106(.VSS(VSS),.VDD(VDD),.Y(g2598),.A(I3726));
  NOT NOT1_1107(.VSS(VSS),.VDD(VDD),.Y(I3729),.A(g2436));
  NOT NOT1_1108(.VSS(VSS),.VDD(VDD),.Y(g2599),.A(I3729));
  NOT NOT1_1109(.VSS(VSS),.VDD(VDD),.Y(g2602),.A(g2061));
  NOT NOT1_1110(.VSS(VSS),.VDD(VDD),.Y(I3733),.A(g2031));
  NOT NOT1_1111(.VSS(VSS),.VDD(VDD),.Y(g2603),.A(I3733));
  NOT NOT1_1112(.VSS(VSS),.VDD(VDD),.Y(I3736),.A(g2460));
  NOT NOT1_1113(.VSS(VSS),.VDD(VDD),.Y(g2604),.A(I3736));
  NOT NOT1_1114(.VSS(VSS),.VDD(VDD),.Y(I3746),.A(g2035));
  NOT NOT1_1115(.VSS(VSS),.VDD(VDD),.Y(g2608),.A(I3746));
  NOT NOT1_1116(.VSS(VSS),.VDD(VDD),.Y(I3749),.A(g2484));
  NOT NOT1_1117(.VSS(VSS),.VDD(VDD),.Y(g2609),.A(I3749));
  NOT NOT1_1118(.VSS(VSS),.VDD(VDD),.Y(I3752),.A(g2044));
  NOT NOT1_1119(.VSS(VSS),.VDD(VDD),.Y(g2612),.A(I3752));
  NOT NOT1_1120(.VSS(VSS),.VDD(VDD),.Y(I3755),.A(g2125));
  NOT NOT1_1121(.VSS(VSS),.VDD(VDD),.Y(g2615),.A(I3755));
  NOT NOT1_1122(.VSS(VSS),.VDD(VDD),.Y(I3758),.A(g2041));
  NOT NOT1_1123(.VSS(VSS),.VDD(VDD),.Y(g2618),.A(I3758));
  NOT NOT1_1124(.VSS(VSS),.VDD(VDD),.Y(I3761),.A(g2505));
  NOT NOT1_1125(.VSS(VSS),.VDD(VDD),.Y(g2619),.A(I3761));
  NOT NOT1_1126(.VSS(VSS),.VDD(VDD),.Y(I3764),.A(g2044));
  NOT NOT1_1127(.VSS(VSS),.VDD(VDD),.Y(g2622),.A(I3764));
  NOT NOT1_1128(.VSS(VSS),.VDD(VDD),.Y(I3767),.A(g2125));
  NOT NOT1_1129(.VSS(VSS),.VDD(VDD),.Y(g2625),.A(I3767));
  NOT NOT1_1130(.VSS(VSS),.VDD(VDD),.Y(I3770),.A(g2145));
  NOT NOT1_1131(.VSS(VSS),.VDD(VDD),.Y(g2628),.A(I3770));
  NOT NOT1_1132(.VSS(VSS),.VDD(VDD),.Y(I3773),.A(g2524));
  NOT NOT1_1133(.VSS(VSS),.VDD(VDD),.Y(g2631),.A(I3773));
  NOT NOT1_1134(.VSS(VSS),.VDD(VDD),.Y(I3776),.A(g2044));
  NOT NOT1_1135(.VSS(VSS),.VDD(VDD),.Y(g2634),.A(I3776));
  NOT NOT1_1136(.VSS(VSS),.VDD(VDD),.Y(I3779),.A(g2125));
  NOT NOT1_1137(.VSS(VSS),.VDD(VDD),.Y(g2637),.A(I3779));
  NOT NOT1_1138(.VSS(VSS),.VDD(VDD),.Y(I3782),.A(g2145));
  NOT NOT1_1139(.VSS(VSS),.VDD(VDD),.Y(g2640),.A(I3782));
  NOT NOT1_1140(.VSS(VSS),.VDD(VDD),.Y(I3785),.A(g2346));
  NOT NOT1_1141(.VSS(VSS),.VDD(VDD),.Y(g2643),.A(I3785));
  NOT NOT1_1142(.VSS(VSS),.VDD(VDD),.Y(I3788),.A(g2554));
  NOT NOT1_1143(.VSS(VSS),.VDD(VDD),.Y(g2644),.A(I3788));
  NOT NOT1_1144(.VSS(VSS),.VDD(VDD),.Y(I3791),.A(g2044));
  NOT NOT1_1145(.VSS(VSS),.VDD(VDD),.Y(g2647),.A(I3791));
  NOT NOT1_1146(.VSS(VSS),.VDD(VDD),.Y(I3794),.A(g2044));
  NOT NOT1_1147(.VSS(VSS),.VDD(VDD),.Y(g2650),.A(I3794));
  NOT NOT1_1148(.VSS(VSS),.VDD(VDD),.Y(I3797),.A(g2125));
  NOT NOT1_1149(.VSS(VSS),.VDD(VDD),.Y(g2653),.A(I3797));
  NOT NOT1_1150(.VSS(VSS),.VDD(VDD),.Y(I3800),.A(g2145));
  NOT NOT1_1151(.VSS(VSS),.VDD(VDD),.Y(g2656),.A(I3800));
  NOT NOT1_1152(.VSS(VSS),.VDD(VDD),.Y(I3804),.A(g2575));
  NOT NOT1_1153(.VSS(VSS),.VDD(VDD),.Y(g2660),.A(I3804));
  NOT NOT1_1154(.VSS(VSS),.VDD(VDD),.Y(g2663),.A(g2308));
  NOT NOT1_1155(.VSS(VSS),.VDD(VDD),.Y(I3808),.A(g2125));
  NOT NOT1_1156(.VSS(VSS),.VDD(VDD),.Y(g2664),.A(I3808));
  NOT NOT1_1157(.VSS(VSS),.VDD(VDD),.Y(I3811),.A(g2145));
  NOT NOT1_1158(.VSS(VSS),.VDD(VDD),.Y(g2667),.A(I3811));
  NOT NOT1_1159(.VSS(VSS),.VDD(VDD),.Y(I3816),.A(g2580));
  NOT NOT1_1160(.VSS(VSS),.VDD(VDD),.Y(g2672),.A(I3816));
  NOT NOT1_1161(.VSS(VSS),.VDD(VDD),.Y(I3819),.A(g2044));
  NOT NOT1_1162(.VSS(VSS),.VDD(VDD),.Y(g2675),.A(I3819));
  NOT NOT1_1163(.VSS(VSS),.VDD(VDD),.Y(g2678),.A(g2312));
  NOT NOT1_1164(.VSS(VSS),.VDD(VDD),.Y(I3823),.A(g2125));
  NOT NOT1_1165(.VSS(VSS),.VDD(VDD),.Y(g2679),.A(I3823));
  NOT NOT1_1166(.VSS(VSS),.VDD(VDD),.Y(I3826),.A(g2145));
  NOT NOT1_1167(.VSS(VSS),.VDD(VDD),.Y(g2682),.A(I3826));
  NOT NOT1_1168(.VSS(VSS),.VDD(VDD),.Y(I3830),.A(g2179));
  NOT NOT1_1169(.VSS(VSS),.VDD(VDD),.Y(g2686),.A(I3830));
  NOT NOT1_1170(.VSS(VSS),.VDD(VDD),.Y(I3833),.A(g2266));
  NOT NOT1_1171(.VSS(VSS),.VDD(VDD),.Y(g2687),.A(I3833));
  NOT NOT1_1172(.VSS(VSS),.VDD(VDD),.Y(I3836),.A(g1832));
  NOT NOT1_1173(.VSS(VSS),.VDD(VDD),.Y(g2688),.A(I3836));
  NOT NOT1_1174(.VSS(VSS),.VDD(VDD),.Y(g2691),.A(g2317));
  NOT NOT1_1175(.VSS(VSS),.VDD(VDD),.Y(I3840),.A(g2125));
  NOT NOT1_1176(.VSS(VSS),.VDD(VDD),.Y(g2692),.A(I3840));
  NOT NOT1_1177(.VSS(VSS),.VDD(VDD),.Y(I3843),.A(g2145));
  NOT NOT1_1178(.VSS(VSS),.VDD(VDD),.Y(g2695),.A(I3843));
  NOT NOT1_1179(.VSS(VSS),.VDD(VDD),.Y(I3855),.A(g2550));
  NOT NOT1_1180(.VSS(VSS),.VDD(VDD),.Y(g2701),.A(I3855));
  NOT NOT1_1181(.VSS(VSS),.VDD(VDD),.Y(I3858),.A(g2197));
  NOT NOT1_1182(.VSS(VSS),.VDD(VDD),.Y(g2705),.A(I3858));
  NOT NOT1_1183(.VSS(VSS),.VDD(VDD),.Y(I3861),.A(g1834));
  NOT NOT1_1184(.VSS(VSS),.VDD(VDD),.Y(g2706),.A(I3861));
  NOT NOT1_1185(.VSS(VSS),.VDD(VDD),.Y(I3864),.A(g2044));
  NOT NOT1_1186(.VSS(VSS),.VDD(VDD),.Y(g2709),.A(I3864));
  NOT NOT1_1187(.VSS(VSS),.VDD(VDD),.Y(g2712),.A(g2320));
  NOT NOT1_1188(.VSS(VSS),.VDD(VDD),.Y(I3868),.A(g2125));
  NOT NOT1_1189(.VSS(VSS),.VDD(VDD),.Y(g2713),.A(I3868));
  NOT NOT1_1190(.VSS(VSS),.VDD(VDD),.Y(I3871),.A(g2145));
  NOT NOT1_1191(.VSS(VSS),.VDD(VDD),.Y(g2716),.A(I3871));
  NOT NOT1_1192(.VSS(VSS),.VDD(VDD),.Y(I3883),.A(g2574));
  NOT NOT1_1193(.VSS(VSS),.VDD(VDD),.Y(g2722),.A(I3883));
  NOT NOT1_1194(.VSS(VSS),.VDD(VDD),.Y(I3886),.A(g2215));
  NOT NOT1_1195(.VSS(VSS),.VDD(VDD),.Y(g2726),.A(I3886));
  NOT NOT1_1196(.VSS(VSS),.VDD(VDD),.Y(g2727),.A(g2324));
  NOT NOT1_1197(.VSS(VSS),.VDD(VDD),.Y(I3890),.A(g2145));
  NOT NOT1_1198(.VSS(VSS),.VDD(VDD),.Y(g2728),.A(I3890));
  NOT NOT1_1199(.VSS(VSS),.VDD(VDD),.Y(I3902),.A(g2576));
  NOT NOT1_1200(.VSS(VSS),.VDD(VDD),.Y(g2734),.A(I3902));
  NOT NOT1_1201(.VSS(VSS),.VDD(VDD),.Y(g2738),.A(g2327));
  NOT NOT1_1202(.VSS(VSS),.VDD(VDD),.Y(I3906),.A(g2234));
  NOT NOT1_1203(.VSS(VSS),.VDD(VDD),.Y(g2739),.A(I3906));
  NOT NOT1_1204(.VSS(VSS),.VDD(VDD),.Y(I3909),.A(g2044));
  NOT NOT1_1205(.VSS(VSS),.VDD(VDD),.Y(g2740),.A(I3909));
  NOT NOT1_1206(.VSS(VSS),.VDD(VDD),.Y(g2743),.A(g2333));
  NOT NOT1_1207(.VSS(VSS),.VDD(VDD),.Y(g2744),.A(g2336));
  NOT NOT1_1208(.VSS(VSS),.VDD(VDD),.Y(I3923),.A(g2581));
  NOT NOT1_1209(.VSS(VSS),.VDD(VDD),.Y(g2748),.A(I3923));
  NOT NOT1_1210(.VSS(VSS),.VDD(VDD),.Y(g2752),.A(g2343));
  NOT NOT1_1211(.VSS(VSS),.VDD(VDD),.Y(I3927),.A(g2245));
  NOT NOT1_1212(.VSS(VSS),.VDD(VDD),.Y(g2753),.A(I3927));
  NOT NOT1_1213(.VSS(VSS),.VDD(VDD),.Y(g2754),.A(g2347));
  NOT NOT1_1214(.VSS(VSS),.VDD(VDD),.Y(g2755),.A(g2350));
  NOT NOT1_1215(.VSS(VSS),.VDD(VDD),.Y(g2756),.A(g2353));
  NOT NOT1_1216(.VSS(VSS),.VDD(VDD),.Y(I3942),.A(g1833));
  NOT NOT1_1217(.VSS(VSS),.VDD(VDD),.Y(g2760),.A(I3942));
  NOT NOT1_1218(.VSS(VSS),.VDD(VDD),.Y(g2764),.A(g2357));
  NOT NOT1_1219(.VSS(VSS),.VDD(VDD),.Y(I3946),.A(g2256));
  NOT NOT1_1220(.VSS(VSS),.VDD(VDD),.Y(g2765),.A(I3946));
  NOT NOT1_1221(.VSS(VSS),.VDD(VDD),.Y(g2766),.A(g2361));
  NOT NOT1_1222(.VSS(VSS),.VDD(VDD),.Y(g2767),.A(g2364));
  NOT NOT1_1223(.VSS(VSS),.VDD(VDD),.Y(g2768),.A(g2367));
  NOT NOT1_1224(.VSS(VSS),.VDD(VDD),.Y(I3961),.A(g1835));
  NOT NOT1_1225(.VSS(VSS),.VDD(VDD),.Y(g2772),.A(I3961));
  NOT NOT1_1226(.VSS(VSS),.VDD(VDD),.Y(g2776),.A(g2378));
  NOT NOT1_1227(.VSS(VSS),.VDD(VDD),.Y(I3965),.A(g2268));
  NOT NOT1_1228(.VSS(VSS),.VDD(VDD),.Y(g2777),.A(I3965));
  NOT NOT1_1229(.VSS(VSS),.VDD(VDD),.Y(g2778),.A(g2391));
  NOT NOT1_1230(.VSS(VSS),.VDD(VDD),.Y(g2779),.A(g2394));
  NOT NOT1_1231(.VSS(VSS),.VDD(VDD),.Y(I3979),.A(g1836));
  NOT NOT1_1232(.VSS(VSS),.VDD(VDD),.Y(g2783),.A(I3979));
  NOT NOT1_1233(.VSS(VSS),.VDD(VDD),.Y(g2787),.A(g2405));
  NOT NOT1_1234(.VSS(VSS),.VDD(VDD),.Y(I3983),.A(g2276));
  NOT NOT1_1235(.VSS(VSS),.VDD(VDD),.Y(g2788),.A(I3983));
  NOT NOT1_1236(.VSS(VSS),.VDD(VDD),.Y(g2789),.A(g2410));
  NOT NOT1_1237(.VSS(VSS),.VDD(VDD),.Y(g2790),.A(g2413));
  NOT NOT1_1238(.VSS(VSS),.VDD(VDD),.Y(g2792),.A(g2416));
  NOT NOT1_1239(.VSS(VSS),.VDD(VDD),.Y(I3999),.A(g1837));
  NOT NOT1_1240(.VSS(VSS),.VDD(VDD),.Y(g2796),.A(I3999));
  NOT NOT1_1241(.VSS(VSS),.VDD(VDD),.Y(g2800),.A(g2430));
  NOT NOT1_1242(.VSS(VSS),.VDD(VDD),.Y(I4003),.A(g2284));
  NOT NOT1_1243(.VSS(VSS),.VDD(VDD),.Y(g2801),.A(I4003));
  NOT NOT1_1244(.VSS(VSS),.VDD(VDD),.Y(g2802),.A(g2437));
  NOT NOT1_1245(.VSS(VSS),.VDD(VDD),.Y(g2803),.A(g2440));
  NOT NOT1_1246(.VSS(VSS),.VDD(VDD),.Y(g2805),.A(g2443));
  NOT NOT1_1247(.VSS(VSS),.VDD(VDD),.Y(g2806),.A(g2446));
  NOT NOT1_1248(.VSS(VSS),.VDD(VDD),.Y(I4019),.A(g1841));
  NOT NOT1_1249(.VSS(VSS),.VDD(VDD),.Y(g2809),.A(I4019));
  NOT NOT1_1250(.VSS(VSS),.VDD(VDD),.Y(g2813),.A(g2457));
  NOT NOT1_1251(.VSS(VSS),.VDD(VDD),.Y(I4023),.A(g2315));
  NOT NOT1_1252(.VSS(VSS),.VDD(VDD),.Y(g2814),.A(I4023));
  NOT NOT1_1253(.VSS(VSS),.VDD(VDD),.Y(g2817),.A(g2461));
  NOT NOT1_1254(.VSS(VSS),.VDD(VDD),.Y(g2818),.A(g2464));
  NOT NOT1_1255(.VSS(VSS),.VDD(VDD),.Y(g2819),.A(g2467));
  NOT NOT1_1256(.VSS(VSS),.VDD(VDD),.Y(g2820),.A(g2470));
  NOT NOT1_1257(.VSS(VSS),.VDD(VDD),.Y(I4031),.A(g1846));
  NOT NOT1_1258(.VSS(VSS),.VDD(VDD),.Y(g2822),.A(I4031));
  NOT NOT1_1259(.VSS(VSS),.VDD(VDD),.Y(g2826),.A(g2481));
  NOT NOT1_1260(.VSS(VSS),.VDD(VDD),.Y(g2827),.A(g2485));
  NOT NOT1_1261(.VSS(VSS),.VDD(VDD),.Y(g2828),.A(g2488));
  NOT NOT1_1262(.VSS(VSS),.VDD(VDD),.Y(g2829),.A(g2491));
  NOT NOT1_1263(.VSS(VSS),.VDD(VDD),.Y(g2830),.A(g2494));
  NOT NOT1_1264(.VSS(VSS),.VDD(VDD),.Y(g2835),.A(g2506));
  NOT NOT1_1265(.VSS(VSS),.VDD(VDD),.Y(g2836),.A(g2509));
  NOT NOT1_1266(.VSS(VSS),.VDD(VDD),.Y(g2837),.A(g2512));
  NOT NOT1_1267(.VSS(VSS),.VDD(VDD),.Y(g2838),.A(g2515));
  NOT NOT1_1268(.VSS(VSS),.VDD(VDD),.Y(g2839),.A(g2535));
  NOT NOT1_1269(.VSS(VSS),.VDD(VDD),.Y(g2840),.A(g2538));
  NOT NOT1_1270(.VSS(VSS),.VDD(VDD),.Y(g2841),.A(g2541));
  NOT NOT1_1271(.VSS(VSS),.VDD(VDD),.Y(I4050),.A(g2059));
  NOT NOT1_1272(.VSS(VSS),.VDD(VDD),.Y(g2842),.A(I4050));
  NOT NOT1_1273(.VSS(VSS),.VDD(VDD),.Y(g2845),.A(g2565));
  NOT NOT1_1274(.VSS(VSS),.VDD(VDD),.Y(g2849),.A(g2577));
  NOT NOT1_1275(.VSS(VSS),.VDD(VDD),.Y(g2856),.A(g2010));
  NOT NOT1_1276(.VSS(VSS),.VDD(VDD),.Y(I4059),.A(g1878));
  NOT NOT1_1277(.VSS(VSS),.VDD(VDD),.Y(g2857),.A(I4059));
  NOT NOT1_1278(.VSS(VSS),.VDD(VDD),.Y(I4066),.A(g2582));
  NOT NOT1_1279(.VSS(VSS),.VDD(VDD),.Y(g2862),.A(I4066));
  NOT NOT1_1280(.VSS(VSS),.VDD(VDD),.Y(g2863),.A(g2296));
  NOT NOT1_1281(.VSS(VSS),.VDD(VDD),.Y(g2864),.A(g1887));
  NOT NOT1_1282(.VSS(VSS),.VDD(VDD),.Y(g2865),.A(g2296));
  NOT NOT1_1283(.VSS(VSS),.VDD(VDD),.Y(g2866),.A(g1905));
  NOT NOT1_1284(.VSS(VSS),.VDD(VDD),.Y(g2867),.A(g1908));
  NOT NOT1_1285(.VSS(VSS),.VDD(VDD),.Y(g2869),.A(g2433));
  NOT NOT1_1286(.VSS(VSS),.VDD(VDD),.Y(g2870),.A(g2296));
  NOT NOT1_1287(.VSS(VSS),.VDD(VDD),.Y(g2871),.A(g1919));
  NOT NOT1_1288(.VSS(VSS),.VDD(VDD),.Y(g2872),.A(g1922));
  NOT NOT1_1289(.VSS(VSS),.VDD(VDD),.Y(g2874),.A(g1849));
  NOT NOT1_1290(.VSS(VSS),.VDD(VDD),.Y(g2875),.A(g1940));
  NOT NOT1_1291(.VSS(VSS),.VDD(VDD),.Y(g2876),.A(g1943));
  NOT NOT1_1292(.VSS(VSS),.VDD(VDD),.Y(g2877),.A(g2434));
  NOT NOT1_1293(.VSS(VSS),.VDD(VDD),.Y(g2882),.A(g1854));
  NOT NOT1_1294(.VSS(VSS),.VDD(VDD),.Y(g2883),.A(g1954));
  NOT NOT1_1295(.VSS(VSS),.VDD(VDD),.Y(g2884),.A(g1957));
  NOT NOT1_1296(.VSS(VSS),.VDD(VDD),.Y(g2885),.A(g1963));
  NOT NOT1_1297(.VSS(VSS),.VDD(VDD),.Y(g2886),.A(g1966));
  NOT NOT1_1298(.VSS(VSS),.VDD(VDD),.Y(g2887),.A(g1858));
  NOT NOT1_1299(.VSS(VSS),.VDD(VDD),.Y(g2888),.A(g1972));
  NOT NOT1_1300(.VSS(VSS),.VDD(VDD),.Y(g2889),.A(g1975));
  NOT NOT1_1301(.VSS(VSS),.VDD(VDD),.Y(g2890),.A(g1875));
  NOT NOT1_1302(.VSS(VSS),.VDD(VDD),.Y(g2891),.A(g1884));
  NOT NOT1_1303(.VSS(VSS),.VDD(VDD),.Y(g2892),.A(g1982));
  NOT NOT1_1304(.VSS(VSS),.VDD(VDD),.Y(g2893),.A(g1985));
  NOT NOT1_1305(.VSS(VSS),.VDD(VDD),.Y(g2894),.A(g1891));
  NOT NOT1_1306(.VSS(VSS),.VDD(VDD),.Y(g2895),.A(g1894));
  NOT NOT1_1307(.VSS(VSS),.VDD(VDD),.Y(g2902),.A(g1899));
  NOT NOT1_1308(.VSS(VSS),.VDD(VDD),.Y(g2903),.A(g1902));
  NOT NOT1_1309(.VSS(VSS),.VDD(VDD),.Y(g2904),.A(g1991));
  NOT NOT1_1310(.VSS(VSS),.VDD(VDD),.Y(g2905),.A(g1994));
  NOT NOT1_1311(.VSS(VSS),.VDD(VDD),.Y(g2906),.A(g1911));
  NOT NOT1_1312(.VSS(VSS),.VDD(VDD),.Y(g2907),.A(g1914));
  NOT NOT1_1313(.VSS(VSS),.VDD(VDD),.Y(g2912),.A(g2001));
  NOT NOT1_1314(.VSS(VSS),.VDD(VDD),.Y(g2913),.A(g1925));
  NOT NOT1_1315(.VSS(VSS),.VDD(VDD),.Y(g2914),.A(g1928));
  NOT NOT1_1316(.VSS(VSS),.VDD(VDD),.Y(g2915),.A(g1931));
  NOT NOT1_1317(.VSS(VSS),.VDD(VDD),.Y(g2919),.A(g1937));
  NOT NOT1_1318(.VSS(VSS),.VDD(VDD),.Y(g2920),.A(g1947));
  NOT NOT1_1319(.VSS(VSS),.VDD(VDD),.Y(g2921),.A(g1950));
  NOT NOT1_1320(.VSS(VSS),.VDD(VDD),.Y(g2922),.A(g1960));
  NOT NOT1_1321(.VSS(VSS),.VDD(VDD),.Y(g2923),.A(g1969));
  NOT NOT1_1322(.VSS(VSS),.VDD(VDD),.Y(g2927),.A(g1979));
  NOT NOT1_1323(.VSS(VSS),.VDD(VDD),.Y(g2931),.A(g1988));
  NOT NOT1_1324(.VSS(VSS),.VDD(VDD),.Y(g2932),.A(g1998));
  NOT NOT1_1325(.VSS(VSS),.VDD(VDD),.Y(I4123),.A(g2043));
  NOT NOT1_1326(.VSS(VSS),.VDD(VDD),.Y(g2933),.A(I4123));
  NOT NOT1_1327(.VSS(VSS),.VDD(VDD),.Y(g2934),.A(g2004));
  NOT NOT1_1328(.VSS(VSS),.VDD(VDD),.Y(g2936),.A(g2026));
  NOT NOT1_1329(.VSS(VSS),.VDD(VDD),.Y(I4133),.A(g2040));
  NOT NOT1_1330(.VSS(VSS),.VDD(VDD),.Y(g2945),.A(I4133));
  NOT NOT1_1331(.VSS(VSS),.VDD(VDD),.Y(g2946),.A(g2296));
  NOT NOT1_1332(.VSS(VSS),.VDD(VDD),.Y(g2952),.A(g2381));
  NOT NOT1_1333(.VSS(VSS),.VDD(VDD),.Y(g2954),.A(g2381));
  NOT NOT1_1334(.VSS(VSS),.VDD(VDD),.Y(g2956),.A(g1861));
  NOT NOT1_1335(.VSS(VSS),.VDD(VDD),.Y(g2957),.A(g1861));
  NOT NOT1_1336(.VSS(VSS),.VDD(VDD),.Y(g2958),.A(g1861));
  NOT NOT1_1337(.VSS(VSS),.VDD(VDD),.Y(g2959),.A(g1861));
  NOT NOT1_1338(.VSS(VSS),.VDD(VDD),.Y(g2961),.A(g1861));
  NOT NOT1_1339(.VSS(VSS),.VDD(VDD),.Y(g2962),.A(g2008));
  NOT NOT1_1340(.VSS(VSS),.VDD(VDD),.Y(I4166),.A(g2390));
  NOT NOT1_1341(.VSS(VSS),.VDD(VDD),.Y(g2967),.A(I4166));
  NOT NOT1_1342(.VSS(VSS),.VDD(VDD),.Y(g2968),.A(g2179));
  NOT NOT1_1343(.VSS(VSS),.VDD(VDD),.Y(I4170),.A(g2157));
  NOT NOT1_1344(.VSS(VSS),.VDD(VDD),.Y(g2973),.A(I4170));
  NOT NOT1_1345(.VSS(VSS),.VDD(VDD),.Y(I4173),.A(g2408));
  NOT NOT1_1346(.VSS(VSS),.VDD(VDD),.Y(g2974),.A(I4173));
  NOT NOT1_1347(.VSS(VSS),.VDD(VDD),.Y(I4176),.A(g2268));
  NOT NOT1_1348(.VSS(VSS),.VDD(VDD),.Y(g2975),.A(I4176));
  NOT NOT1_1349(.VSS(VSS),.VDD(VDD),.Y(g2976),.A(g2197));
  NOT NOT1_1350(.VSS(VSS),.VDD(VDD),.Y(g2981),.A(g2179));
  NOT NOT1_1351(.VSS(VSS),.VDD(VDD),.Y(g2986),.A(g2010));
  NOT NOT1_1352(.VSS(VSS),.VDD(VDD),.Y(I4189),.A(g2159));
  NOT NOT1_1353(.VSS(VSS),.VDD(VDD),.Y(g2996),.A(I4189));
  NOT NOT1_1354(.VSS(VSS),.VDD(VDD),.Y(I4192),.A(g1847));
  NOT NOT1_1355(.VSS(VSS),.VDD(VDD),.Y(g2997),.A(I4192));
  NOT NOT1_1356(.VSS(VSS),.VDD(VDD),.Y(I4195),.A(g2173));
  NOT NOT1_1357(.VSS(VSS),.VDD(VDD),.Y(g2998),.A(I4195));
  NOT NOT1_1358(.VSS(VSS),.VDD(VDD),.Y(I4198),.A(g2276));
  NOT NOT1_1359(.VSS(VSS),.VDD(VDD),.Y(g3001),.A(I4198));
  NOT NOT1_1360(.VSS(VSS),.VDD(VDD),.Y(g3002),.A(g2215));
  NOT NOT1_1361(.VSS(VSS),.VDD(VDD),.Y(g3007),.A(g2197));
  NOT NOT1_1362(.VSS(VSS),.VDD(VDD),.Y(I4217),.A(g2163));
  NOT NOT1_1363(.VSS(VSS),.VDD(VDD),.Y(g3014),.A(I4217));
  NOT NOT1_1364(.VSS(VSS),.VDD(VDD),.Y(I4220),.A(g2164));
  NOT NOT1_1365(.VSS(VSS),.VDD(VDD),.Y(g3015),.A(I4220));
  NOT NOT1_1366(.VSS(VSS),.VDD(VDD),.Y(I4223),.A(g2176));
  NOT NOT1_1367(.VSS(VSS),.VDD(VDD),.Y(g3016),.A(I4223));
  NOT NOT1_1368(.VSS(VSS),.VDD(VDD),.Y(I4226),.A(g2525));
  NOT NOT1_1369(.VSS(VSS),.VDD(VDD),.Y(g3019),.A(I4226));
  NOT NOT1_1370(.VSS(VSS),.VDD(VDD),.Y(I4229),.A(g2284));
  NOT NOT1_1371(.VSS(VSS),.VDD(VDD),.Y(g3022),.A(I4229));
  NOT NOT1_1372(.VSS(VSS),.VDD(VDD),.Y(g3023),.A(g2215));
  NOT NOT1_1373(.VSS(VSS),.VDD(VDD),.Y(I4240),.A(g2165));
  NOT NOT1_1374(.VSS(VSS),.VDD(VDD),.Y(g3029),.A(I4240));
  NOT NOT1_1375(.VSS(VSS),.VDD(VDD),.Y(I4243),.A(g1853));
  NOT NOT1_1376(.VSS(VSS),.VDD(VDD),.Y(g3030),.A(I4243));
  NOT NOT1_1377(.VSS(VSS),.VDD(VDD),.Y(I4246),.A(g2194));
  NOT NOT1_1378(.VSS(VSS),.VDD(VDD),.Y(g3031),.A(I4246));
  NOT NOT1_1379(.VSS(VSS),.VDD(VDD),.Y(I4249),.A(g2525));
  NOT NOT1_1380(.VSS(VSS),.VDD(VDD),.Y(g3034),.A(I4249));
  NOT NOT1_1381(.VSS(VSS),.VDD(VDD),.Y(I4252),.A(g2555));
  NOT NOT1_1382(.VSS(VSS),.VDD(VDD),.Y(g3037),.A(I4252));
  NOT NOT1_1383(.VSS(VSS),.VDD(VDD),.Y(I4255),.A(g2179));
  NOT NOT1_1384(.VSS(VSS),.VDD(VDD),.Y(g3040),.A(I4255));
  NOT NOT1_1385(.VSS(VSS),.VDD(VDD),.Y(I4258),.A(g2169));
  NOT NOT1_1386(.VSS(VSS),.VDD(VDD),.Y(g3041),.A(I4258));
  NOT NOT1_1387(.VSS(VSS),.VDD(VDD),.Y(I4261),.A(g1857));
  NOT NOT1_1388(.VSS(VSS),.VDD(VDD),.Y(g3042),.A(I4261));
  NOT NOT1_1389(.VSS(VSS),.VDD(VDD),.Y(I4264),.A(g2212));
  NOT NOT1_1390(.VSS(VSS),.VDD(VDD),.Y(g3043),.A(I4264));
  NOT NOT1_1391(.VSS(VSS),.VDD(VDD),.Y(I4267),.A(g2525));
  NOT NOT1_1392(.VSS(VSS),.VDD(VDD),.Y(g3046),.A(I4267));
  NOT NOT1_1393(.VSS(VSS),.VDD(VDD),.Y(I4270),.A(g2555));
  NOT NOT1_1394(.VSS(VSS),.VDD(VDD),.Y(g3049),.A(I4270));
  NOT NOT1_1395(.VSS(VSS),.VDD(VDD),.Y(I4273),.A(g2197));
  NOT NOT1_1396(.VSS(VSS),.VDD(VDD),.Y(g3052),.A(I4273));
  NOT NOT1_1397(.VSS(VSS),.VDD(VDD),.Y(I4276),.A(g2170));
  NOT NOT1_1398(.VSS(VSS),.VDD(VDD),.Y(g3053),.A(I4276));
  NOT NOT1_1399(.VSS(VSS),.VDD(VDD),.Y(I4279),.A(g2230));
  NOT NOT1_1400(.VSS(VSS),.VDD(VDD),.Y(g3054),.A(I4279));
  NOT NOT1_1401(.VSS(VSS),.VDD(VDD),.Y(I4282),.A(g2525));
  NOT NOT1_1402(.VSS(VSS),.VDD(VDD),.Y(g3057),.A(I4282));
  NOT NOT1_1403(.VSS(VSS),.VDD(VDD),.Y(I4285),.A(g2555));
  NOT NOT1_1404(.VSS(VSS),.VDD(VDD),.Y(g3060),.A(I4285));
  NOT NOT1_1405(.VSS(VSS),.VDD(VDD),.Y(I4288),.A(g2215));
  NOT NOT1_1406(.VSS(VSS),.VDD(VDD),.Y(g3063),.A(I4288));
  NOT NOT1_1407(.VSS(VSS),.VDD(VDD),.Y(I4291),.A(g2241));
  NOT NOT1_1408(.VSS(VSS),.VDD(VDD),.Y(g3064),.A(I4291));
  NOT NOT1_1409(.VSS(VSS),.VDD(VDD),.Y(I4294),.A(g2525));
  NOT NOT1_1410(.VSS(VSS),.VDD(VDD),.Y(g3067),.A(I4294));
  NOT NOT1_1411(.VSS(VSS),.VDD(VDD),.Y(I4297),.A(g2555));
  NOT NOT1_1412(.VSS(VSS),.VDD(VDD),.Y(g3070),.A(I4297));
  NOT NOT1_1413(.VSS(VSS),.VDD(VDD),.Y(I4300),.A(g2234));
  NOT NOT1_1414(.VSS(VSS),.VDD(VDD),.Y(g3073),.A(I4300));
  NOT NOT1_1415(.VSS(VSS),.VDD(VDD),.Y(I4303),.A(g1897));
  NOT NOT1_1416(.VSS(VSS),.VDD(VDD),.Y(g3074),.A(I4303));
  NOT NOT1_1417(.VSS(VSS),.VDD(VDD),.Y(I4306),.A(g1898));
  NOT NOT1_1418(.VSS(VSS),.VDD(VDD),.Y(g3075),.A(I4306));
  NOT NOT1_1419(.VSS(VSS),.VDD(VDD),.Y(I4309),.A(g2525));
  NOT NOT1_1420(.VSS(VSS),.VDD(VDD),.Y(g3076),.A(I4309));
  NOT NOT1_1421(.VSS(VSS),.VDD(VDD),.Y(I4312),.A(g2555));
  NOT NOT1_1422(.VSS(VSS),.VDD(VDD),.Y(g3079),.A(I4312));
  NOT NOT1_1423(.VSS(VSS),.VDD(VDD),.Y(I4315),.A(g2245));
  NOT NOT1_1424(.VSS(VSS),.VDD(VDD),.Y(g3082),.A(I4315));
  NOT NOT1_1425(.VSS(VSS),.VDD(VDD),.Y(I4318),.A(g2171));
  NOT NOT1_1426(.VSS(VSS),.VDD(VDD),.Y(g3083),.A(I4318));
  NOT NOT1_1427(.VSS(VSS),.VDD(VDD),.Y(I4321),.A(g1917));
  NOT NOT1_1428(.VSS(VSS),.VDD(VDD),.Y(g3084),.A(I4321));
  NOT NOT1_1429(.VSS(VSS),.VDD(VDD),.Y(I4324),.A(g1918));
  NOT NOT1_1430(.VSS(VSS),.VDD(VDD),.Y(g3085),.A(I4324));
  NOT NOT1_1431(.VSS(VSS),.VDD(VDD),.Y(I4327),.A(g2525));
  NOT NOT1_1432(.VSS(VSS),.VDD(VDD),.Y(g3086),.A(I4327));
  NOT NOT1_1433(.VSS(VSS),.VDD(VDD),.Y(I4331),.A(g2555));
  NOT NOT1_1434(.VSS(VSS),.VDD(VDD),.Y(g3090),.A(I4331));
  NOT NOT1_1435(.VSS(VSS),.VDD(VDD),.Y(I4334),.A(g2256));
  NOT NOT1_1436(.VSS(VSS),.VDD(VDD),.Y(g3093),.A(I4334));
  NOT NOT1_1437(.VSS(VSS),.VDD(VDD),.Y(I4337),.A(g1934));
  NOT NOT1_1438(.VSS(VSS),.VDD(VDD),.Y(g3094),.A(I4337));
  NOT NOT1_1439(.VSS(VSS),.VDD(VDD),.Y(I4340),.A(g1935));
  NOT NOT1_1440(.VSS(VSS),.VDD(VDD),.Y(g3095),.A(I4340));
  NOT NOT1_1441(.VSS(VSS),.VDD(VDD),.Y(I4343),.A(g2525));
  NOT NOT1_1442(.VSS(VSS),.VDD(VDD),.Y(g3096),.A(I4343));
  NOT NOT1_1443(.VSS(VSS),.VDD(VDD),.Y(I4347),.A(g2555));
  NOT NOT1_1444(.VSS(VSS),.VDD(VDD),.Y(g3100),.A(I4347));
  NOT NOT1_1445(.VSS(VSS),.VDD(VDD),.Y(I4351),.A(g2233));
  NOT NOT1_1446(.VSS(VSS),.VDD(VDD),.Y(g3104),.A(I4351));
  NOT NOT1_1447(.VSS(VSS),.VDD(VDD),.Y(I4354),.A(g1953));
  NOT NOT1_1448(.VSS(VSS),.VDD(VDD),.Y(g3108),.A(I4354));
  NOT NOT1_1449(.VSS(VSS),.VDD(VDD),.Y(I4358),.A(g2525));
  NOT NOT1_1450(.VSS(VSS),.VDD(VDD),.Y(g3110),.A(I4358));
  NOT NOT1_1451(.VSS(VSS),.VDD(VDD),.Y(I4362),.A(g2555));
  NOT NOT1_1452(.VSS(VSS),.VDD(VDD),.Y(g3114),.A(I4362));
  NOT NOT1_1453(.VSS(VSS),.VDD(VDD),.Y(I4366),.A(g2244));
  NOT NOT1_1454(.VSS(VSS),.VDD(VDD),.Y(g3118),.A(I4366));
  NOT NOT1_1455(.VSS(VSS),.VDD(VDD),.Y(I4371),.A(g2555));
  NOT NOT1_1456(.VSS(VSS),.VDD(VDD),.Y(g3124),.A(I4371));
  NOT NOT1_1457(.VSS(VSS),.VDD(VDD),.Y(I4375),.A(g2254));
  NOT NOT1_1458(.VSS(VSS),.VDD(VDD),.Y(g3128),.A(I4375));
  NOT NOT1_1459(.VSS(VSS),.VDD(VDD),.Y(I4382),.A(g2265));
  NOT NOT1_1460(.VSS(VSS),.VDD(VDD),.Y(g3136),.A(I4382));
  NOT NOT1_1461(.VSS(VSS),.VDD(VDD),.Y(I4391),.A(g2275));
  NOT NOT1_1462(.VSS(VSS),.VDD(VDD),.Y(g3150),.A(I4391));
  NOT NOT1_1463(.VSS(VSS),.VDD(VDD),.Y(I4398),.A(g2086));
  NOT NOT1_1464(.VSS(VSS),.VDD(VDD),.Y(g3158),.A(I4398));
  NOT NOT1_1465(.VSS(VSS),.VDD(VDD),.Y(I4402),.A(g2283));
  NOT NOT1_1466(.VSS(VSS),.VDD(VDD),.Y(g3162),.A(I4402));
  NOT NOT1_1467(.VSS(VSS),.VDD(VDD),.Y(I4410),.A(g2088));
  NOT NOT1_1468(.VSS(VSS),.VDD(VDD),.Y(g3173),.A(I4410));
  NOT NOT1_1469(.VSS(VSS),.VDD(VDD),.Y(I4414),.A(g2090));
  NOT NOT1_1470(.VSS(VSS),.VDD(VDD),.Y(g3177),.A(I4414));
  NOT NOT1_1471(.VSS(VSS),.VDD(VDD),.Y(I4420),.A(g2096));
  NOT NOT1_1472(.VSS(VSS),.VDD(VDD),.Y(g3183),.A(I4420));
  NOT NOT1_1473(.VSS(VSS),.VDD(VDD),.Y(I4424),.A(g2097));
  NOT NOT1_1474(.VSS(VSS),.VDD(VDD),.Y(g3187),.A(I4424));
  NOT NOT1_1475(.VSS(VSS),.VDD(VDD),.Y(I4429),.A(g2102));
  NOT NOT1_1476(.VSS(VSS),.VDD(VDD),.Y(g3192),.A(I4429));
  NOT NOT1_1477(.VSS(VSS),.VDD(VDD),.Y(I4433),.A(g2103));
  NOT NOT1_1478(.VSS(VSS),.VDD(VDD),.Y(g3196),.A(I4433));
  NOT NOT1_1479(.VSS(VSS),.VDD(VDD),.Y(g3199),.A(g1861));
  NOT NOT1_1480(.VSS(VSS),.VDD(VDD),.Y(I4437),.A(g2108));
  NOT NOT1_1481(.VSS(VSS),.VDD(VDD),.Y(g3200),.A(I4437));
  NOT NOT1_1482(.VSS(VSS),.VDD(VDD),.Y(I4441),.A(g2109));
  NOT NOT1_1483(.VSS(VSS),.VDD(VDD),.Y(g3204),.A(I4441));
  NOT NOT1_1484(.VSS(VSS),.VDD(VDD),.Y(I4452),.A(g2117));
  NOT NOT1_1485(.VSS(VSS),.VDD(VDD),.Y(g3209),.A(I4452));
  NOT NOT1_1486(.VSS(VSS),.VDD(VDD),.Y(I4455),.A(g2118));
  NOT NOT1_1487(.VSS(VSS),.VDD(VDD),.Y(g3212),.A(I4455));
  NOT NOT1_1488(.VSS(VSS),.VDD(VDD),.Y(I4459),.A(g2134));
  NOT NOT1_1489(.VSS(VSS),.VDD(VDD),.Y(g3216),.A(I4459));
  NOT NOT1_1490(.VSS(VSS),.VDD(VDD),.Y(I4462),.A(g2135));
  NOT NOT1_1491(.VSS(VSS),.VDD(VDD),.Y(g3219),.A(I4462));
  NOT NOT1_1492(.VSS(VSS),.VDD(VDD),.Y(I4465),.A(g2945));
  NOT NOT1_1493(.VSS(VSS),.VDD(VDD),.Y(g3222),.A(I4465));
  NOT NOT1_1494(.VSS(VSS),.VDD(VDD),.Y(I4468),.A(g2583));
  NOT NOT1_1495(.VSS(VSS),.VDD(VDD),.Y(g3223),.A(I4468));
  NOT NOT1_1496(.VSS(VSS),.VDD(VDD),.Y(I4471),.A(g3040));
  NOT NOT1_1497(.VSS(VSS),.VDD(VDD),.Y(g3224),.A(I4471));
  NOT NOT1_1498(.VSS(VSS),.VDD(VDD),.Y(I4474),.A(g3052));
  NOT NOT1_1499(.VSS(VSS),.VDD(VDD),.Y(g3225),.A(I4474));
  NOT NOT1_1500(.VSS(VSS),.VDD(VDD),.Y(I4477),.A(g3063));
  NOT NOT1_1501(.VSS(VSS),.VDD(VDD),.Y(g3226),.A(I4477));
  NOT NOT1_1502(.VSS(VSS),.VDD(VDD),.Y(I4480),.A(g3073));
  NOT NOT1_1503(.VSS(VSS),.VDD(VDD),.Y(g3227),.A(I4480));
  NOT NOT1_1504(.VSS(VSS),.VDD(VDD),.Y(I4483),.A(g3082));
  NOT NOT1_1505(.VSS(VSS),.VDD(VDD),.Y(g3228),.A(I4483));
  NOT NOT1_1506(.VSS(VSS),.VDD(VDD),.Y(I4486),.A(g3093));
  NOT NOT1_1507(.VSS(VSS),.VDD(VDD),.Y(g3229),.A(I4486));
  NOT NOT1_1508(.VSS(VSS),.VDD(VDD),.Y(I4489),.A(g2975));
  NOT NOT1_1509(.VSS(VSS),.VDD(VDD),.Y(g3230),.A(I4489));
  NOT NOT1_1510(.VSS(VSS),.VDD(VDD),.Y(I4492),.A(g3001));
  NOT NOT1_1511(.VSS(VSS),.VDD(VDD),.Y(g3231),.A(I4492));
  NOT NOT1_1512(.VSS(VSS),.VDD(VDD),.Y(I4495),.A(g3022));
  NOT NOT1_1513(.VSS(VSS),.VDD(VDD),.Y(g3232),.A(I4495));
  NOT NOT1_1514(.VSS(VSS),.VDD(VDD),.Y(I4498),.A(g2686));
  NOT NOT1_1515(.VSS(VSS),.VDD(VDD),.Y(g3233),.A(I4498));
  NOT NOT1_1516(.VSS(VSS),.VDD(VDD),.Y(I4501),.A(g2705));
  NOT NOT1_1517(.VSS(VSS),.VDD(VDD),.Y(g3234),.A(I4501));
  NOT NOT1_1518(.VSS(VSS),.VDD(VDD),.Y(I4504),.A(g2726));
  NOT NOT1_1519(.VSS(VSS),.VDD(VDD),.Y(g3235),.A(I4504));
  NOT NOT1_1520(.VSS(VSS),.VDD(VDD),.Y(I4507),.A(g2739));
  NOT NOT1_1521(.VSS(VSS),.VDD(VDD),.Y(g3236),.A(I4507));
  NOT NOT1_1522(.VSS(VSS),.VDD(VDD),.Y(I4510),.A(g2753));
  NOT NOT1_1523(.VSS(VSS),.VDD(VDD),.Y(g3237),.A(I4510));
  NOT NOT1_1524(.VSS(VSS),.VDD(VDD),.Y(I4513),.A(g2765));
  NOT NOT1_1525(.VSS(VSS),.VDD(VDD),.Y(g3238),.A(I4513));
  NOT NOT1_1526(.VSS(VSS),.VDD(VDD),.Y(I4516),.A(g2777));
  NOT NOT1_1527(.VSS(VSS),.VDD(VDD),.Y(g3239),.A(I4516));
  NOT NOT1_1528(.VSS(VSS),.VDD(VDD),.Y(I4519),.A(g2788));
  NOT NOT1_1529(.VSS(VSS),.VDD(VDD),.Y(g3240),.A(I4519));
  NOT NOT1_1530(.VSS(VSS),.VDD(VDD),.Y(I4522),.A(g2801));
  NOT NOT1_1531(.VSS(VSS),.VDD(VDD),.Y(g3241),.A(I4522));
  NOT NOT1_1532(.VSS(VSS),.VDD(VDD),.Y(g3242),.A(g3083));
  NOT NOT1_1533(.VSS(VSS),.VDD(VDD),.Y(g3247),.A(g2973));
  NOT NOT1_1534(.VSS(VSS),.VDD(VDD),.Y(I4534),.A(g2858));
  NOT NOT1_1535(.VSS(VSS),.VDD(VDD),.Y(g3251),.A(I4534));
  NOT NOT1_1536(.VSS(VSS),.VDD(VDD),.Y(I4537),.A(g2877));
  NOT NOT1_1537(.VSS(VSS),.VDD(VDD),.Y(g3258),.A(I4537));
  NOT NOT1_1538(.VSS(VSS),.VDD(VDD),.Y(g3259),.A(g2996));
  NOT NOT1_1539(.VSS(VSS),.VDD(VDD),.Y(g3263),.A(g3015));
  NOT NOT1_1540(.VSS(VSS),.VDD(VDD),.Y(g3267),.A(g3030));
  NOT NOT1_1541(.VSS(VSS),.VDD(VDD),.Y(g3271),.A(g3042));
  NOT NOT1_1542(.VSS(VSS),.VDD(VDD),.Y(g3284),.A(g3019));
  NOT NOT1_1543(.VSS(VSS),.VDD(VDD),.Y(g3289),.A(g3034));
  NOT NOT1_1544(.VSS(VSS),.VDD(VDD),.Y(g3291),.A(g3037));
  NOT NOT1_1545(.VSS(VSS),.VDD(VDD),.Y(g3297),.A(g3046));
  NOT NOT1_1546(.VSS(VSS),.VDD(VDD),.Y(g3299),.A(g3049));
  NOT NOT1_1547(.VSS(VSS),.VDD(VDD),.Y(g3306),.A(g3057));
  NOT NOT1_1548(.VSS(VSS),.VDD(VDD),.Y(g3308),.A(g3060));
  NOT NOT1_1549(.VSS(VSS),.VDD(VDD),.Y(I4587),.A(g2962));
  NOT NOT1_1550(.VSS(VSS),.VDD(VDD),.Y(g3312),.A(I4587));
  NOT NOT1_1551(.VSS(VSS),.VDD(VDD),.Y(I4593),.A(g2966));
  NOT NOT1_1552(.VSS(VSS),.VDD(VDD),.Y(g3318),.A(I4593));
  NOT NOT1_1553(.VSS(VSS),.VDD(VDD),.Y(g3320),.A(g3067));
  NOT NOT1_1554(.VSS(VSS),.VDD(VDD),.Y(g3322),.A(g3070));
  NOT NOT1_1555(.VSS(VSS),.VDD(VDD),.Y(g3331),.A(g3076));
  NOT NOT1_1556(.VSS(VSS),.VDD(VDD),.Y(g3332),.A(g3079));
  NOT NOT1_1557(.VSS(VSS),.VDD(VDD),.Y(g3342),.A(g3086));
  NOT NOT1_1558(.VSS(VSS),.VDD(VDD),.Y(g3343),.A(g3090));
  NOT NOT1_1559(.VSS(VSS),.VDD(VDD),.Y(I4623),.A(g2962));
  NOT NOT1_1560(.VSS(VSS),.VDD(VDD),.Y(g3346),.A(I4623));
  NOT NOT1_1561(.VSS(VSS),.VDD(VDD),.Y(g3354),.A(g3096));
  NOT NOT1_1562(.VSS(VSS),.VDD(VDD),.Y(g3355),.A(g3100));
  NOT NOT1_1563(.VSS(VSS),.VDD(VDD),.Y(g3363),.A(g3110));
  NOT NOT1_1564(.VSS(VSS),.VDD(VDD),.Y(g3364),.A(g3114));
  NOT NOT1_1565(.VSS(VSS),.VDD(VDD),.Y(I4646),.A(g2602));
  NOT NOT1_1566(.VSS(VSS),.VDD(VDD),.Y(g3369),.A(I4646));
  NOT NOT1_1567(.VSS(VSS),.VDD(VDD),.Y(g3370),.A(g3124));
  NOT NOT1_1568(.VSS(VSS),.VDD(VDD),.Y(g3380),.A(g2831));
  NOT NOT1_1569(.VSS(VSS),.VDD(VDD),.Y(g3384),.A(g2834));
  NOT NOT1_1570(.VSS(VSS),.VDD(VDD),.Y(I4664),.A(g2924));
  NOT NOT1_1571(.VSS(VSS),.VDD(VDD),.Y(g3387),.A(I4664));
  NOT NOT1_1572(.VSS(VSS),.VDD(VDD),.Y(I4667),.A(g2908));
  NOT NOT1_1573(.VSS(VSS),.VDD(VDD),.Y(g3388),.A(I4667));
  NOT NOT1_1574(.VSS(VSS),.VDD(VDD),.Y(I4671),.A(g2928));
  NOT NOT1_1575(.VSS(VSS),.VDD(VDD),.Y(g3424),.A(I4671));
  NOT NOT1_1576(.VSS(VSS),.VDD(VDD),.Y(I4678),.A(g2670));
  NOT NOT1_1577(.VSS(VSS),.VDD(VDD),.Y(g3440),.A(I4678));
  NOT NOT1_1578(.VSS(VSS),.VDD(VDD),.Y(I4681),.A(g2947));
  NOT NOT1_1579(.VSS(VSS),.VDD(VDD),.Y(g3441),.A(I4681));
  NOT NOT1_1580(.VSS(VSS),.VDD(VDD),.Y(I4684),.A(g2687));
  NOT NOT1_1581(.VSS(VSS),.VDD(VDD),.Y(g3448),.A(I4684));
  NOT NOT1_1582(.VSS(VSS),.VDD(VDD),.Y(I4688),.A(g3207));
  NOT NOT1_1583(.VSS(VSS),.VDD(VDD),.Y(g3450),.A(I4688));
  NOT NOT1_1584(.VSS(VSS),.VDD(VDD),.Y(g3451),.A(g2615));
  NOT NOT1_1585(.VSS(VSS),.VDD(VDD),.Y(g3452),.A(g2625));
  NOT NOT1_1586(.VSS(VSS),.VDD(VDD),.Y(g3453),.A(g2628));
  NOT NOT1_1587(.VSS(VSS),.VDD(VDD),.Y(g3455),.A(g2637));
  NOT NOT1_1588(.VSS(VSS),.VDD(VDD),.Y(g3456),.A(g2640));
  NOT NOT1_1589(.VSS(VSS),.VDD(VDD),.Y(g3457),.A(g2653));
  NOT NOT1_1590(.VSS(VSS),.VDD(VDD),.Y(g3458),.A(g2656));
  NOT NOT1_1591(.VSS(VSS),.VDD(VDD),.Y(g3459),.A(g2664));
  NOT NOT1_1592(.VSS(VSS),.VDD(VDD),.Y(g3460),.A(g2667));
  NOT NOT1_1593(.VSS(VSS),.VDD(VDD),.Y(g3461),.A(g2986));
  NOT NOT1_1594(.VSS(VSS),.VDD(VDD),.Y(g3462),.A(g2679));
  NOT NOT1_1595(.VSS(VSS),.VDD(VDD),.Y(g3463),.A(g2682));
  NOT NOT1_1596(.VSS(VSS),.VDD(VDD),.Y(g3465),.A(g2986));
  NOT NOT1_1597(.VSS(VSS),.VDD(VDD),.Y(I4706),.A(g2877));
  NOT NOT1_1598(.VSS(VSS),.VDD(VDD),.Y(g3466),.A(I4706));
  NOT NOT1_1599(.VSS(VSS),.VDD(VDD),.Y(g3477),.A(g2692));
  NOT NOT1_1600(.VSS(VSS),.VDD(VDD),.Y(g3478),.A(g2695));
  NOT NOT1_1601(.VSS(VSS),.VDD(VDD),.Y(g3480),.A(g2986));
  NOT NOT1_1602(.VSS(VSS),.VDD(VDD),.Y(g3481),.A(g2612));
  NOT NOT1_1603(.VSS(VSS),.VDD(VDD),.Y(g3482),.A(g2713));
  NOT NOT1_1604(.VSS(VSS),.VDD(VDD),.Y(g3483),.A(g2716));
  NOT NOT1_1605(.VSS(VSS),.VDD(VDD),.Y(g3485),.A(g2986));
  NOT NOT1_1606(.VSS(VSS),.VDD(VDD),.Y(g3486),.A(g2869));
  NOT NOT1_1607(.VSS(VSS),.VDD(VDD),.Y(g3487),.A(g2622));
  NOT NOT1_1608(.VSS(VSS),.VDD(VDD),.Y(g3488),.A(g2728));
  NOT NOT1_1609(.VSS(VSS),.VDD(VDD),.Y(g3491),.A(g2608));
  NOT NOT1_1610(.VSS(VSS),.VDD(VDD),.Y(g3498),.A(g2634));
  NOT NOT1_1611(.VSS(VSS),.VDD(VDD),.Y(g3500),.A(g2647));
  NOT NOT1_1612(.VSS(VSS),.VDD(VDD),.Y(g3501),.A(g2650));
  NOT NOT1_1613(.VSS(VSS),.VDD(VDD),.Y(g3504),.A(g2675));
  NOT NOT1_1614(.VSS(VSS),.VDD(VDD),.Y(g3510),.A(g2709));
  NOT NOT1_1615(.VSS(VSS),.VDD(VDD),.Y(g3519),.A(g2740));
  NOT NOT1_1616(.VSS(VSS),.VDD(VDD),.Y(I4743),.A(g2594));
  NOT NOT1_1617(.VSS(VSS),.VDD(VDD),.Y(g3527),.A(I4743));
  NOT NOT1_1618(.VSS(VSS),.VDD(VDD),.Y(I4752),.A(g2859));
  NOT NOT1_1619(.VSS(VSS),.VDD(VDD),.Y(g3534),.A(I4752));
  NOT NOT1_1620(.VSS(VSS),.VDD(VDD),.Y(I4757),.A(g2861));
  NOT NOT1_1621(.VSS(VSS),.VDD(VDD),.Y(g3537),.A(I4757));
  NOT NOT1_1622(.VSS(VSS),.VDD(VDD),.Y(I4762),.A(g2862));
  NOT NOT1_1623(.VSS(VSS),.VDD(VDD),.Y(g3540),.A(I4762));
  NOT NOT1_1624(.VSS(VSS),.VDD(VDD),.Y(g3541),.A(g2643));
  NOT NOT1_1625(.VSS(VSS),.VDD(VDD),.Y(g3545),.A(g3085));
  NOT NOT1_1626(.VSS(VSS),.VDD(VDD),.Y(g3546),.A(g3095));
  NOT NOT1_1627(.VSS(VSS),.VDD(VDD),.Y(g3557),.A(g2598));
  NOT NOT1_1628(.VSS(VSS),.VDD(VDD),.Y(g3559),.A(g2603));
  NOT NOT1_1629(.VSS(VSS),.VDD(VDD),.Y(g3564),.A(g2618));
  NOT NOT1_1630(.VSS(VSS),.VDD(VDD),.Y(g3567),.A(g3074));
  NOT NOT1_1631(.VSS(VSS),.VDD(VDD),.Y(g3571),.A(g3084));
  NOT NOT1_1632(.VSS(VSS),.VDD(VDD),.Y(I4777),.A(g2962));
  NOT NOT1_1633(.VSS(VSS),.VDD(VDD),.Y(g3575),.A(I4777));
  NOT NOT1_1634(.VSS(VSS),.VDD(VDD),.Y(g3589),.A(g3094));
  NOT NOT1_1635(.VSS(VSS),.VDD(VDD),.Y(g3593),.A(g2997));
  NOT NOT1_1636(.VSS(VSS),.VDD(VDD),.Y(I4791),.A(g2814));
  NOT NOT1_1637(.VSS(VSS),.VDD(VDD),.Y(g3600),.A(I4791));
  NOT NOT1_1638(.VSS(VSS),.VDD(VDD),.Y(I4794),.A(g2814));
  NOT NOT1_1639(.VSS(VSS),.VDD(VDD),.Y(g3601),.A(I4794));
  NOT NOT1_1640(.VSS(VSS),.VDD(VDD),.Y(I4799),.A(g2967));
  NOT NOT1_1641(.VSS(VSS),.VDD(VDD),.Y(g3604),.A(I4799));
  NOT NOT1_1642(.VSS(VSS),.VDD(VDD),.Y(I4802),.A(g2877));
  NOT NOT1_1643(.VSS(VSS),.VDD(VDD),.Y(g3605),.A(I4802));
  NOT NOT1_1644(.VSS(VSS),.VDD(VDD),.Y(I4809),.A(g2974));
  NOT NOT1_1645(.VSS(VSS),.VDD(VDD),.Y(g3612),.A(I4809));
  NOT NOT1_1646(.VSS(VSS),.VDD(VDD),.Y(I4821),.A(g2877));
  NOT NOT1_1647(.VSS(VSS),.VDD(VDD),.Y(g3622),.A(I4821));
  NOT NOT1_1648(.VSS(VSS),.VDD(VDD),.Y(g3638),.A(g3108));
  NOT NOT1_1649(.VSS(VSS),.VDD(VDD),.Y(g3673),.A(g3075));
  NOT NOT1_1650(.VSS(VSS),.VDD(VDD),.Y(g3677),.A(g3140));
  NOT NOT1_1651(.VSS(VSS),.VDD(VDD),.Y(g3705),.A(g3014));
  NOT NOT1_1652(.VSS(VSS),.VDD(VDD),.Y(g3710),.A(g3029));
  NOT NOT1_1653(.VSS(VSS),.VDD(VDD),.Y(g3714),.A(g3041));
  NOT NOT1_1654(.VSS(VSS),.VDD(VDD),.Y(g3719),.A(g3053));
  NOT NOT1_1655(.VSS(VSS),.VDD(VDD),.Y(I4903),.A(g3223));
  NOT NOT1_1656(.VSS(VSS),.VDD(VDD),.Y(g3723),.A(I4903));
  NOT NOT1_1657(.VSS(VSS),.VDD(VDD),.Y(I4935),.A(g3369));
  NOT NOT1_1658(.VSS(VSS),.VDD(VDD),.Y(g3752),.A(I4935));
  NOT NOT1_1659(.VSS(VSS),.VDD(VDD),.Y(g3761),.A(g3605));
  NOT NOT1_1660(.VSS(VSS),.VDD(VDD),.Y(I4955),.A(g3673));
  NOT NOT1_1661(.VSS(VSS),.VDD(VDD),.Y(g3766),.A(I4955));
  NOT NOT1_1662(.VSS(VSS),.VDD(VDD),.Y(g3769),.A(g3622));
  NOT NOT1_1663(.VSS(VSS),.VDD(VDD),.Y(I4961),.A(g3597));
  NOT NOT1_1664(.VSS(VSS),.VDD(VDD),.Y(g3770),.A(I4961));
  NOT NOT1_1665(.VSS(VSS),.VDD(VDD),.Y(I4964),.A(g3673));
  NOT NOT1_1666(.VSS(VSS),.VDD(VDD),.Y(g3771),.A(I4964));
  NOT NOT1_1667(.VSS(VSS),.VDD(VDD),.Y(g3772),.A(g3466));
  NOT NOT1_1668(.VSS(VSS),.VDD(VDD),.Y(g3773),.A(g3466));
  NOT NOT1_1669(.VSS(VSS),.VDD(VDD),.Y(g3775),.A(g3388));
  NOT NOT1_1670(.VSS(VSS),.VDD(VDD),.Y(g3776),.A(g3466));
  NOT NOT1_1671(.VSS(VSS),.VDD(VDD),.Y(g3777),.A(g3388));
  NOT NOT1_1672(.VSS(VSS),.VDD(VDD),.Y(g3778),.A(g3388));
  NOT NOT1_1673(.VSS(VSS),.VDD(VDD),.Y(g3779),.A(g3466));
  NOT NOT1_1674(.VSS(VSS),.VDD(VDD),.Y(I4976),.A(g3575));
  NOT NOT1_1675(.VSS(VSS),.VDD(VDD),.Y(g3781),.A(I4976));
  NOT NOT1_1676(.VSS(VSS),.VDD(VDD),.Y(g3782),.A(g3388));
  NOT NOT1_1677(.VSS(VSS),.VDD(VDD),.Y(I4980),.A(g3546));
  NOT NOT1_1678(.VSS(VSS),.VDD(VDD),.Y(g3783),.A(I4980));
  NOT NOT1_1679(.VSS(VSS),.VDD(VDD),.Y(g3785),.A(g3466));
  NOT NOT1_1680(.VSS(VSS),.VDD(VDD),.Y(g3786),.A(g3388));
  NOT NOT1_1681(.VSS(VSS),.VDD(VDD),.Y(I4986),.A(g3638));
  NOT NOT1_1682(.VSS(VSS),.VDD(VDD),.Y(g3787),.A(I4986));
  NOT NOT1_1683(.VSS(VSS),.VDD(VDD),.Y(g3788),.A(g3466));
  NOT NOT1_1684(.VSS(VSS),.VDD(VDD),.Y(g3789),.A(g3388));
  NOT NOT1_1685(.VSS(VSS),.VDD(VDD),.Y(g3790),.A(g3388));
  NOT NOT1_1686(.VSS(VSS),.VDD(VDD),.Y(g3791),.A(g3388));
  NOT NOT1_1687(.VSS(VSS),.VDD(VDD),.Y(g3792),.A(g3388));
  NOT NOT1_1688(.VSS(VSS),.VDD(VDD),.Y(g3793),.A(g3491));
  NOT NOT1_1689(.VSS(VSS),.VDD(VDD),.Y(g3796),.A(g3388));
  NOT NOT1_1690(.VSS(VSS),.VDD(VDD),.Y(g3797),.A(g3388));
  NOT NOT1_1691(.VSS(VSS),.VDD(VDD),.Y(g3798),.A(g3388));
  NOT NOT1_1692(.VSS(VSS),.VDD(VDD),.Y(g3799),.A(g3388));
  NOT NOT1_1693(.VSS(VSS),.VDD(VDD),.Y(g3800),.A(g3388));
  NOT NOT1_1694(.VSS(VSS),.VDD(VDD),.Y(g3801),.A(g3388));
  NOT NOT1_1695(.VSS(VSS),.VDD(VDD),.Y(g3802),.A(g3388));
  NOT NOT1_1696(.VSS(VSS),.VDD(VDD),.Y(I5002),.A(g3612));
  NOT NOT1_1697(.VSS(VSS),.VDD(VDD),.Y(g3803),.A(I5002));
  NOT NOT1_1698(.VSS(VSS),.VDD(VDD),.Y(I5006),.A(g3604));
  NOT NOT1_1699(.VSS(VSS),.VDD(VDD),.Y(g3807),.A(I5006));
  NOT NOT1_1700(.VSS(VSS),.VDD(VDD),.Y(g3813),.A(g3258));
  NOT NOT1_1701(.VSS(VSS),.VDD(VDD),.Y(I5019),.A(g3318));
  NOT NOT1_1702(.VSS(VSS),.VDD(VDD),.Y(g3830),.A(I5019));
  NOT NOT1_1703(.VSS(VSS),.VDD(VDD),.Y(I5023),.A(g3263));
  NOT NOT1_1704(.VSS(VSS),.VDD(VDD),.Y(g3832),.A(I5023));
  NOT NOT1_1705(.VSS(VSS),.VDD(VDD),.Y(I5027),.A(g3267));
  NOT NOT1_1706(.VSS(VSS),.VDD(VDD),.Y(g3834),.A(I5027));
  NOT NOT1_1707(.VSS(VSS),.VDD(VDD),.Y(I5030),.A(g3242));
  NOT NOT1_1708(.VSS(VSS),.VDD(VDD),.Y(g3835),.A(I5030));
  NOT NOT1_1709(.VSS(VSS),.VDD(VDD),.Y(I5033),.A(g3527));
  NOT NOT1_1710(.VSS(VSS),.VDD(VDD),.Y(g3836),.A(I5033));
  NOT NOT1_1711(.VSS(VSS),.VDD(VDD),.Y(I5037),.A(g3705));
  NOT NOT1_1712(.VSS(VSS),.VDD(VDD),.Y(g3838),.A(I5037));
  NOT NOT1_1713(.VSS(VSS),.VDD(VDD),.Y(I5040),.A(g3271));
  NOT NOT1_1714(.VSS(VSS),.VDD(VDD),.Y(g3839),.A(I5040));
  NOT NOT1_1715(.VSS(VSS),.VDD(VDD),.Y(I5043),.A(g3247));
  NOT NOT1_1716(.VSS(VSS),.VDD(VDD),.Y(g3840),.A(I5043));
  NOT NOT1_1717(.VSS(VSS),.VDD(VDD),.Y(I5050),.A(g3246));
  NOT NOT1_1718(.VSS(VSS),.VDD(VDD),.Y(g3845),.A(I5050));
  NOT NOT1_1719(.VSS(VSS),.VDD(VDD),.Y(I5053),.A(g3710));
  NOT NOT1_1720(.VSS(VSS),.VDD(VDD),.Y(g3846),.A(I5053));
  NOT NOT1_1721(.VSS(VSS),.VDD(VDD),.Y(I5056),.A(g3567));
  NOT NOT1_1722(.VSS(VSS),.VDD(VDD),.Y(g3847),.A(I5056));
  NOT NOT1_1723(.VSS(VSS),.VDD(VDD),.Y(I5059),.A(g3259));
  NOT NOT1_1724(.VSS(VSS),.VDD(VDD),.Y(g3848),.A(I5059));
  NOT NOT1_1725(.VSS(VSS),.VDD(VDD),.Y(I5065),.A(g3714));
  NOT NOT1_1726(.VSS(VSS),.VDD(VDD),.Y(g3852),.A(I5065));
  NOT NOT1_1727(.VSS(VSS),.VDD(VDD),.Y(I5068),.A(g3571));
  NOT NOT1_1728(.VSS(VSS),.VDD(VDD),.Y(g3853),.A(I5068));
  NOT NOT1_1729(.VSS(VSS),.VDD(VDD),.Y(I5071),.A(g3263));
  NOT NOT1_1730(.VSS(VSS),.VDD(VDD),.Y(g3854),.A(I5071));
  NOT NOT1_1731(.VSS(VSS),.VDD(VDD),.Y(I5078),.A(g3719));
  NOT NOT1_1732(.VSS(VSS),.VDD(VDD),.Y(g3859),.A(I5078));
  NOT NOT1_1733(.VSS(VSS),.VDD(VDD),.Y(I5081),.A(g3589));
  NOT NOT1_1734(.VSS(VSS),.VDD(VDD),.Y(g3860),.A(I5081));
  NOT NOT1_1735(.VSS(VSS),.VDD(VDD),.Y(I5084),.A(g3593));
  NOT NOT1_1736(.VSS(VSS),.VDD(VDD),.Y(g3861),.A(I5084));
  NOT NOT1_1737(.VSS(VSS),.VDD(VDD),.Y(I5091),.A(g3242));
  NOT NOT1_1738(.VSS(VSS),.VDD(VDD),.Y(g3866),.A(I5091));
  NOT NOT1_1739(.VSS(VSS),.VDD(VDD),.Y(I5094),.A(g3705));
  NOT NOT1_1740(.VSS(VSS),.VDD(VDD),.Y(g3867),.A(I5094));
  NOT NOT1_1741(.VSS(VSS),.VDD(VDD),.Y(g3868),.A(g3491));
  NOT NOT1_1742(.VSS(VSS),.VDD(VDD),.Y(g3872),.A(g3312));
  NOT NOT1_1743(.VSS(VSS),.VDD(VDD),.Y(I5103),.A(g3440));
  NOT NOT1_1744(.VSS(VSS),.VDD(VDD),.Y(g3874),.A(I5103));
  NOT NOT1_1745(.VSS(VSS),.VDD(VDD),.Y(I5106),.A(g3247));
  NOT NOT1_1746(.VSS(VSS),.VDD(VDD),.Y(g3875),.A(I5106));
  NOT NOT1_1747(.VSS(VSS),.VDD(VDD),.Y(I5109),.A(g3710));
  NOT NOT1_1748(.VSS(VSS),.VDD(VDD),.Y(g3876),.A(I5109));
  NOT NOT1_1749(.VSS(VSS),.VDD(VDD),.Y(I5116),.A(g3259));
  NOT NOT1_1750(.VSS(VSS),.VDD(VDD),.Y(g3881),.A(I5116));
  NOT NOT1_1751(.VSS(VSS),.VDD(VDD),.Y(I5119),.A(g3714));
  NOT NOT1_1752(.VSS(VSS),.VDD(VDD),.Y(g3882),.A(I5119));
  NOT NOT1_1753(.VSS(VSS),.VDD(VDD),.Y(I5124),.A(g3719));
  NOT NOT1_1754(.VSS(VSS),.VDD(VDD),.Y(g3885),.A(I5124));
  NOT NOT1_1755(.VSS(VSS),.VDD(VDD),.Y(g3886),.A(g3346));
  NOT NOT1_1756(.VSS(VSS),.VDD(VDD),.Y(g3889),.A(g3575));
  NOT NOT1_1757(.VSS(VSS),.VDD(VDD),.Y(g3890),.A(g3575));
  NOT NOT1_1758(.VSS(VSS),.VDD(VDD),.Y(g3892),.A(g3575));
  NOT NOT1_1759(.VSS(VSS),.VDD(VDD),.Y(g3897),.A(g3251));
  NOT NOT1_1760(.VSS(VSS),.VDD(VDD),.Y(g3898),.A(g3575));
  NOT NOT1_1761(.VSS(VSS),.VDD(VDD),.Y(g3900),.A(g3575));
  NOT NOT1_1762(.VSS(VSS),.VDD(VDD),.Y(g3901),.A(g3575));
  NOT NOT1_1763(.VSS(VSS),.VDD(VDD),.Y(g3902),.A(g3575));
  NOT NOT1_1764(.VSS(VSS),.VDD(VDD),.Y(g3904),.A(g3575));
  NOT NOT1_1765(.VSS(VSS),.VDD(VDD),.Y(g3906),.A(g3575));
  NOT NOT1_1766(.VSS(VSS),.VDD(VDD),.Y(I5148),.A(g3450));
  NOT NOT1_1767(.VSS(VSS),.VDD(VDD),.Y(g3911),.A(I5148));
  NOT NOT1_1768(.VSS(VSS),.VDD(VDD),.Y(g3912),.A(g3505));
  NOT NOT1_1769(.VSS(VSS),.VDD(VDD),.Y(I5153),.A(g3330));
  NOT NOT1_1770(.VSS(VSS),.VDD(VDD),.Y(g3914),.A(I5153));
  NOT NOT1_1771(.VSS(VSS),.VDD(VDD),.Y(g3921),.A(g3512));
  NOT NOT1_1772(.VSS(VSS),.VDD(VDD),.Y(I5157),.A(g3454));
  NOT NOT1_1773(.VSS(VSS),.VDD(VDD),.Y(g3922),.A(I5157));
  NOT NOT1_1774(.VSS(VSS),.VDD(VDD),.Y(I5169),.A(g3593));
  NOT NOT1_1775(.VSS(VSS),.VDD(VDD),.Y(g3932),.A(I5169));
  NOT NOT1_1776(.VSS(VSS),.VDD(VDD),.Y(I5177),.A(g3267));
  NOT NOT1_1777(.VSS(VSS),.VDD(VDD),.Y(g3940),.A(I5177));
  NOT NOT1_1778(.VSS(VSS),.VDD(VDD),.Y(I5182),.A(g3271));
  NOT NOT1_1779(.VSS(VSS),.VDD(VDD),.Y(g3952),.A(I5182));
  NOT NOT1_1780(.VSS(VSS),.VDD(VDD),.Y(I5204),.A(g3534));
  NOT NOT1_1781(.VSS(VSS),.VDD(VDD),.Y(g3960),.A(I5204));
  NOT NOT1_1782(.VSS(VSS),.VDD(VDD),.Y(I5214),.A(g3567));
  NOT NOT1_1783(.VSS(VSS),.VDD(VDD),.Y(g3962),.A(I5214));
  NOT NOT1_1784(.VSS(VSS),.VDD(VDD),.Y(I5217),.A(g3673));
  NOT NOT1_1785(.VSS(VSS),.VDD(VDD),.Y(g3963),.A(I5217));
  NOT NOT1_1786(.VSS(VSS),.VDD(VDD),.Y(I5223),.A(g3537));
  NOT NOT1_1787(.VSS(VSS),.VDD(VDD),.Y(g3967),.A(I5223));
  NOT NOT1_1788(.VSS(VSS),.VDD(VDD),.Y(I5233),.A(g3571));
  NOT NOT1_1789(.VSS(VSS),.VDD(VDD),.Y(g3969),.A(I5233));
  NOT NOT1_1790(.VSS(VSS),.VDD(VDD),.Y(I5236),.A(g3545));
  NOT NOT1_1791(.VSS(VSS),.VDD(VDD),.Y(g3970),.A(I5236));
  NOT NOT1_1792(.VSS(VSS),.VDD(VDD),.Y(I5249),.A(g3589));
  NOT NOT1_1793(.VSS(VSS),.VDD(VDD),.Y(g3975),.A(I5249));
  NOT NOT1_1794(.VSS(VSS),.VDD(VDD),.Y(I5252),.A(g3546));
  NOT NOT1_1795(.VSS(VSS),.VDD(VDD),.Y(g3976),.A(I5252));
  NOT NOT1_1796(.VSS(VSS),.VDD(VDD),.Y(I5264),.A(g3638));
  NOT NOT1_1797(.VSS(VSS),.VDD(VDD),.Y(g3980),.A(I5264));
  NOT NOT1_1798(.VSS(VSS),.VDD(VDD),.Y(g3984),.A(g3564));
  NOT NOT1_1799(.VSS(VSS),.VDD(VDD),.Y(g4003),.A(g3441));
  NOT NOT1_1800(.VSS(VSS),.VDD(VDD),.Y(g4010),.A(g3601));
  NOT NOT1_1801(.VSS(VSS),.VDD(VDD),.Y(g4011),.A(g3486));
  NOT NOT1_1802(.VSS(VSS),.VDD(VDD),.Y(I5316),.A(g3557));
  NOT NOT1_1803(.VSS(VSS),.VDD(VDD),.Y(g4014),.A(I5316));
  NOT NOT1_1804(.VSS(VSS),.VDD(VDD),.Y(I5320),.A(g3559));
  NOT NOT1_1805(.VSS(VSS),.VDD(VDD),.Y(g4016),.A(I5320));
  NOT NOT1_1806(.VSS(VSS),.VDD(VDD),.Y(I5324),.A(g3466));
  NOT NOT1_1807(.VSS(VSS),.VDD(VDD),.Y(g4020),.A(I5324));
  NOT NOT1_1808(.VSS(VSS),.VDD(VDD),.Y(I5328),.A(g3502));
  NOT NOT1_1809(.VSS(VSS),.VDD(VDD),.Y(g4022),.A(I5328));
  NOT NOT1_1810(.VSS(VSS),.VDD(VDD),.Y(I5333),.A(g3491));
  NOT NOT1_1811(.VSS(VSS),.VDD(VDD),.Y(g4034),.A(I5333));
  NOT NOT1_1812(.VSS(VSS),.VDD(VDD),.Y(I5337),.A(g3564));
  NOT NOT1_1813(.VSS(VSS),.VDD(VDD),.Y(g4036),.A(I5337));
  NOT NOT1_1814(.VSS(VSS),.VDD(VDD),.Y(I5343),.A(g3599));
  NOT NOT1_1815(.VSS(VSS),.VDD(VDD),.Y(g4040),.A(I5343));
  NOT NOT1_1816(.VSS(VSS),.VDD(VDD),.Y(I5376),.A(g4014));
  NOT NOT1_1817(.VSS(VSS),.VDD(VDD),.Y(g4098),.A(I5376));
  NOT NOT1_1818(.VSS(VSS),.VDD(VDD),.Y(I5379),.A(g3940));
  NOT NOT1_1819(.VSS(VSS),.VDD(VDD),.Y(g4099),.A(I5379));
  NOT NOT1_1820(.VSS(VSS),.VDD(VDD),.Y(I5382),.A(g3952));
  NOT NOT1_1821(.VSS(VSS),.VDD(VDD),.Y(g4100),.A(I5382));
  NOT NOT1_1822(.VSS(VSS),.VDD(VDD),.Y(I5385),.A(g3962));
  NOT NOT1_1823(.VSS(VSS),.VDD(VDD),.Y(g4101),.A(I5385));
  NOT NOT1_1824(.VSS(VSS),.VDD(VDD),.Y(I5388),.A(g3969));
  NOT NOT1_1825(.VSS(VSS),.VDD(VDD),.Y(g4102),.A(I5388));
  NOT NOT1_1826(.VSS(VSS),.VDD(VDD),.Y(I5391),.A(g3975));
  NOT NOT1_1827(.VSS(VSS),.VDD(VDD),.Y(g4103),.A(I5391));
  NOT NOT1_1828(.VSS(VSS),.VDD(VDD),.Y(I5394),.A(g4016));
  NOT NOT1_1829(.VSS(VSS),.VDD(VDD),.Y(g4104),.A(I5394));
  NOT NOT1_1830(.VSS(VSS),.VDD(VDD),.Y(I5397),.A(g3932));
  NOT NOT1_1831(.VSS(VSS),.VDD(VDD),.Y(g4105),.A(I5397));
  NOT NOT1_1832(.VSS(VSS),.VDD(VDD),.Y(I5400),.A(g3963));
  NOT NOT1_1833(.VSS(VSS),.VDD(VDD),.Y(g4106),.A(I5400));
  NOT NOT1_1834(.VSS(VSS),.VDD(VDD),.Y(I5403),.A(g3970));
  NOT NOT1_1835(.VSS(VSS),.VDD(VDD),.Y(g4107),.A(I5403));
  NOT NOT1_1836(.VSS(VSS),.VDD(VDD),.Y(I5406),.A(g3976));
  NOT NOT1_1837(.VSS(VSS),.VDD(VDD),.Y(g4108),.A(I5406));
  NOT NOT1_1838(.VSS(VSS),.VDD(VDD),.Y(I5409),.A(g3980));
  NOT NOT1_1839(.VSS(VSS),.VDD(VDD),.Y(g4109),.A(I5409));
  NOT NOT1_1840(.VSS(VSS),.VDD(VDD),.Y(I5412),.A(g4034));
  NOT NOT1_1841(.VSS(VSS),.VDD(VDD),.Y(g4110),.A(I5412));
  NOT NOT1_1842(.VSS(VSS),.VDD(VDD),.Y(I5415),.A(g3723));
  NOT NOT1_1843(.VSS(VSS),.VDD(VDD),.Y(g4111),.A(I5415));
  NOT NOT1_1844(.VSS(VSS),.VDD(VDD),.Y(I5418),.A(g4036));
  NOT NOT1_1845(.VSS(VSS),.VDD(VDD),.Y(g4112),.A(I5418));
  NOT NOT1_1846(.VSS(VSS),.VDD(VDD),.Y(I5421),.A(g3724));
  NOT NOT1_1847(.VSS(VSS),.VDD(VDD),.Y(g4113),.A(I5421));
  NOT NOT1_1848(.VSS(VSS),.VDD(VDD),.Y(I5424),.A(g3725));
  NOT NOT1_1849(.VSS(VSS),.VDD(VDD),.Y(g4114),.A(I5424));
  NOT NOT1_1850(.VSS(VSS),.VDD(VDD),.Y(I5427),.A(g3726));
  NOT NOT1_1851(.VSS(VSS),.VDD(VDD),.Y(g4115),.A(I5427));
  NOT NOT1_1852(.VSS(VSS),.VDD(VDD),.Y(I5430),.A(g3727));
  NOT NOT1_1853(.VSS(VSS),.VDD(VDD),.Y(g4116),.A(I5430));
  NOT NOT1_1854(.VSS(VSS),.VDD(VDD),.Y(I5433),.A(g3728));
  NOT NOT1_1855(.VSS(VSS),.VDD(VDD),.Y(g4117),.A(I5433));
  NOT NOT1_1856(.VSS(VSS),.VDD(VDD),.Y(I5436),.A(g3729));
  NOT NOT1_1857(.VSS(VSS),.VDD(VDD),.Y(g4118),.A(I5436));
  NOT NOT1_1858(.VSS(VSS),.VDD(VDD),.Y(I5439),.A(g3730));
  NOT NOT1_1859(.VSS(VSS),.VDD(VDD),.Y(g4119),.A(I5439));
  NOT NOT1_1860(.VSS(VSS),.VDD(VDD),.Y(I5442),.A(g3731));
  NOT NOT1_1861(.VSS(VSS),.VDD(VDD),.Y(g4120),.A(I5442));
  NOT NOT1_1862(.VSS(VSS),.VDD(VDD),.Y(I5445),.A(g4040));
  NOT NOT1_1863(.VSS(VSS),.VDD(VDD),.Y(g4121),.A(I5445));
  NOT NOT1_1864(.VSS(VSS),.VDD(VDD),.Y(I5448),.A(g3960));
  NOT NOT1_1865(.VSS(VSS),.VDD(VDD),.Y(g4122),.A(I5448));
  NOT NOT1_1866(.VSS(VSS),.VDD(VDD),.Y(I5451),.A(g3967));
  NOT NOT1_1867(.VSS(VSS),.VDD(VDD),.Y(g4123),.A(I5451));
  NOT NOT1_1868(.VSS(VSS),.VDD(VDD),.Y(I5454),.A(g3874));
  NOT NOT1_1869(.VSS(VSS),.VDD(VDD),.Y(g4124),.A(I5454));
  NOT NOT1_1870(.VSS(VSS),.VDD(VDD),.Y(I5457),.A(g3766));
  NOT NOT1_1871(.VSS(VSS),.VDD(VDD),.Y(g4125),.A(I5457));
  NOT NOT1_1872(.VSS(VSS),.VDD(VDD),.Y(I5460),.A(g3771));
  NOT NOT1_1873(.VSS(VSS),.VDD(VDD),.Y(g4126),.A(I5460));
  NOT NOT1_1874(.VSS(VSS),.VDD(VDD),.Y(I5463),.A(g3783));
  NOT NOT1_1875(.VSS(VSS),.VDD(VDD),.Y(g4127),.A(I5463));
  NOT NOT1_1876(.VSS(VSS),.VDD(VDD),.Y(I5466),.A(g3787));
  NOT NOT1_1877(.VSS(VSS),.VDD(VDD),.Y(g4128),.A(I5466));
  NOT NOT1_1878(.VSS(VSS),.VDD(VDD),.Y(I5469),.A(g3838));
  NOT NOT1_1879(.VSS(VSS),.VDD(VDD),.Y(g4129),.A(I5469));
  NOT NOT1_1880(.VSS(VSS),.VDD(VDD),.Y(I5472),.A(g3846));
  NOT NOT1_1881(.VSS(VSS),.VDD(VDD),.Y(g4130),.A(I5472));
  NOT NOT1_1882(.VSS(VSS),.VDD(VDD),.Y(I5475),.A(g3852));
  NOT NOT1_1883(.VSS(VSS),.VDD(VDD),.Y(g4131),.A(I5475));
  NOT NOT1_1884(.VSS(VSS),.VDD(VDD),.Y(I5478),.A(g3859));
  NOT NOT1_1885(.VSS(VSS),.VDD(VDD),.Y(g4132),.A(I5478));
  NOT NOT1_1886(.VSS(VSS),.VDD(VDD),.Y(I5481),.A(g3866));
  NOT NOT1_1887(.VSS(VSS),.VDD(VDD),.Y(g4133),.A(I5481));
  NOT NOT1_1888(.VSS(VSS),.VDD(VDD),.Y(I5484),.A(g3875));
  NOT NOT1_1889(.VSS(VSS),.VDD(VDD),.Y(g4134),.A(I5484));
  NOT NOT1_1890(.VSS(VSS),.VDD(VDD),.Y(I5487),.A(g3881));
  NOT NOT1_1891(.VSS(VSS),.VDD(VDD),.Y(g4135),.A(I5487));
  NOT NOT1_1892(.VSS(VSS),.VDD(VDD),.Y(I5490),.A(g3832));
  NOT NOT1_1893(.VSS(VSS),.VDD(VDD),.Y(g4136),.A(I5490));
  NOT NOT1_1894(.VSS(VSS),.VDD(VDD),.Y(I5493),.A(g3834));
  NOT NOT1_1895(.VSS(VSS),.VDD(VDD),.Y(g4137),.A(I5493));
  NOT NOT1_1896(.VSS(VSS),.VDD(VDD),.Y(I5496),.A(g3839));
  NOT NOT1_1897(.VSS(VSS),.VDD(VDD),.Y(g4138),.A(I5496));
  NOT NOT1_1898(.VSS(VSS),.VDD(VDD),.Y(I5499),.A(g3847));
  NOT NOT1_1899(.VSS(VSS),.VDD(VDD),.Y(g4139),.A(I5499));
  NOT NOT1_1900(.VSS(VSS),.VDD(VDD),.Y(I5502),.A(g3853));
  NOT NOT1_1901(.VSS(VSS),.VDD(VDD),.Y(g4140),.A(I5502));
  NOT NOT1_1902(.VSS(VSS),.VDD(VDD),.Y(I5505),.A(g3860));
  NOT NOT1_1903(.VSS(VSS),.VDD(VDD),.Y(g4141),.A(I5505));
  NOT NOT1_1904(.VSS(VSS),.VDD(VDD),.Y(I5508),.A(g3867));
  NOT NOT1_1905(.VSS(VSS),.VDD(VDD),.Y(g4142),.A(I5508));
  NOT NOT1_1906(.VSS(VSS),.VDD(VDD),.Y(I5511),.A(g3876));
  NOT NOT1_1907(.VSS(VSS),.VDD(VDD),.Y(g4143),.A(I5511));
  NOT NOT1_1908(.VSS(VSS),.VDD(VDD),.Y(I5514),.A(g3882));
  NOT NOT1_1909(.VSS(VSS),.VDD(VDD),.Y(g4144),.A(I5514));
  NOT NOT1_1910(.VSS(VSS),.VDD(VDD),.Y(I5517),.A(g3885));
  NOT NOT1_1911(.VSS(VSS),.VDD(VDD),.Y(g4145),.A(I5517));
  NOT NOT1_1912(.VSS(VSS),.VDD(VDD),.Y(I5520),.A(g3835));
  NOT NOT1_1913(.VSS(VSS),.VDD(VDD),.Y(g4146),.A(I5520));
  NOT NOT1_1914(.VSS(VSS),.VDD(VDD),.Y(I5523),.A(g3840));
  NOT NOT1_1915(.VSS(VSS),.VDD(VDD),.Y(g4147),.A(I5523));
  NOT NOT1_1916(.VSS(VSS),.VDD(VDD),.Y(I5526),.A(g3848));
  NOT NOT1_1917(.VSS(VSS),.VDD(VDD),.Y(g4148),.A(I5526));
  NOT NOT1_1918(.VSS(VSS),.VDD(VDD),.Y(I5529),.A(g3854));
  NOT NOT1_1919(.VSS(VSS),.VDD(VDD),.Y(g4149),.A(I5529));
  NOT NOT1_1920(.VSS(VSS),.VDD(VDD),.Y(I5532),.A(g3861));
  NOT NOT1_1921(.VSS(VSS),.VDD(VDD),.Y(g4150),.A(I5532));
  NOT NOT1_1922(.VSS(VSS),.VDD(VDD),.Y(I5542),.A(g3984));
  NOT NOT1_1923(.VSS(VSS),.VDD(VDD),.Y(g4152),.A(I5542));
  NOT NOT1_1924(.VSS(VSS),.VDD(VDD),.Y(I5545),.A(g3814));
  NOT NOT1_1925(.VSS(VSS),.VDD(VDD),.Y(g4153),.A(I5545));
  NOT NOT1_1926(.VSS(VSS),.VDD(VDD),.Y(I5548),.A(g4059));
  NOT NOT1_1927(.VSS(VSS),.VDD(VDD),.Y(g4154),.A(I5548));
  NOT NOT1_1928(.VSS(VSS),.VDD(VDD),.Y(I5551),.A(g4059));
  NOT NOT1_1929(.VSS(VSS),.VDD(VDD),.Y(g4155),.A(I5551));
  NOT NOT1_1930(.VSS(VSS),.VDD(VDD),.Y(I5556),.A(g4059));
  NOT NOT1_1931(.VSS(VSS),.VDD(VDD),.Y(g4158),.A(I5556));
  NOT NOT1_1932(.VSS(VSS),.VDD(VDD),.Y(I5562),.A(g4002));
  NOT NOT1_1933(.VSS(VSS),.VDD(VDD),.Y(g4162),.A(I5562));
  NOT NOT1_1934(.VSS(VSS),.VDD(VDD),.Y(I5568),.A(g3897));
  NOT NOT1_1935(.VSS(VSS),.VDD(VDD),.Y(g4166),.A(I5568));
  NOT NOT1_1936(.VSS(VSS),.VDD(VDD),.Y(I5577),.A(g4022));
  NOT NOT1_1937(.VSS(VSS),.VDD(VDD),.Y(g4173),.A(I5577));
  NOT NOT1_1938(.VSS(VSS),.VDD(VDD),.Y(I5591),.A(g3821));
  NOT NOT1_1939(.VSS(VSS),.VDD(VDD),.Y(g4187),.A(I5591));
  NOT NOT1_1940(.VSS(VSS),.VDD(VDD),.Y(I5594),.A(g3821));
  NOT NOT1_1941(.VSS(VSS),.VDD(VDD),.Y(g4188),.A(I5594));
  NOT NOT1_1942(.VSS(VSS),.VDD(VDD),.Y(I5597),.A(g3821));
  NOT NOT1_1943(.VSS(VSS),.VDD(VDD),.Y(g4189),.A(I5597));
  NOT NOT1_1944(.VSS(VSS),.VDD(VDD),.Y(I5600),.A(g3821));
  NOT NOT1_1945(.VSS(VSS),.VDD(VDD),.Y(g4190),.A(I5600));
  NOT NOT1_1946(.VSS(VSS),.VDD(VDD),.Y(I5603),.A(g3893));
  NOT NOT1_1947(.VSS(VSS),.VDD(VDD),.Y(g4191),.A(I5603));
  NOT NOT1_1948(.VSS(VSS),.VDD(VDD),.Y(I5606),.A(g3821));
  NOT NOT1_1949(.VSS(VSS),.VDD(VDD),.Y(g4192),.A(I5606));
  NOT NOT1_1950(.VSS(VSS),.VDD(VDD),.Y(I5609),.A(g3893));
  NOT NOT1_1951(.VSS(VSS),.VDD(VDD),.Y(g4193),.A(I5609));
  NOT NOT1_1952(.VSS(VSS),.VDD(VDD),.Y(I5612),.A(g3910));
  NOT NOT1_1953(.VSS(VSS),.VDD(VDD),.Y(g4194),.A(I5612));
  NOT NOT1_1954(.VSS(VSS),.VDD(VDD),.Y(I5615),.A(g3914));
  NOT NOT1_1955(.VSS(VSS),.VDD(VDD),.Y(g4195),.A(I5615));
  NOT NOT1_1956(.VSS(VSS),.VDD(VDD),.Y(I5618),.A(g3821));
  NOT NOT1_1957(.VSS(VSS),.VDD(VDD),.Y(g4198),.A(I5618));
  NOT NOT1_1958(.VSS(VSS),.VDD(VDD),.Y(I5622),.A(g3914));
  NOT NOT1_1959(.VSS(VSS),.VDD(VDD),.Y(g4202),.A(I5622));
  NOT NOT1_1960(.VSS(VSS),.VDD(VDD),.Y(I5626),.A(g3914));
  NOT NOT1_1961(.VSS(VSS),.VDD(VDD),.Y(g4206),.A(I5626));
  NOT NOT1_1962(.VSS(VSS),.VDD(VDD),.Y(I5630),.A(g3914));
  NOT NOT1_1963(.VSS(VSS),.VDD(VDD),.Y(g4210),.A(I5630));
  NOT NOT1_1964(.VSS(VSS),.VDD(VDD),.Y(I5633),.A(g3768));
  NOT NOT1_1965(.VSS(VSS),.VDD(VDD),.Y(g4213),.A(I5633));
  NOT NOT1_1966(.VSS(VSS),.VDD(VDD),.Y(I5637),.A(g3914));
  NOT NOT1_1967(.VSS(VSS),.VDD(VDD),.Y(g4215),.A(I5637));
  NOT NOT1_1968(.VSS(VSS),.VDD(VDD),.Y(I5640),.A(g3770));
  NOT NOT1_1969(.VSS(VSS),.VDD(VDD),.Y(g4218),.A(I5640));
  NOT NOT1_1970(.VSS(VSS),.VDD(VDD),.Y(I5644),.A(g4059));
  NOT NOT1_1971(.VSS(VSS),.VDD(VDD),.Y(g4220),.A(I5644));
  NOT NOT1_1972(.VSS(VSS),.VDD(VDD),.Y(I5654),.A(g3742));
  NOT NOT1_1973(.VSS(VSS),.VDD(VDD),.Y(g4222),.A(I5654));
  NOT NOT1_1974(.VSS(VSS),.VDD(VDD),.Y(g4224),.A(g4046));
  NOT NOT1_1975(.VSS(VSS),.VDD(VDD),.Y(g4225),.A(g4059));
  NOT NOT1_1976(.VSS(VSS),.VDD(VDD),.Y(g4226),.A(g4050));
  NOT NOT1_1977(.VSS(VSS),.VDD(VDD),.Y(g4227),.A(g4059));
  NOT NOT1_1978(.VSS(VSS),.VDD(VDD),.Y(I5668),.A(g3828));
  NOT NOT1_1979(.VSS(VSS),.VDD(VDD),.Y(g4228),.A(I5668));
  NOT NOT1_1980(.VSS(VSS),.VDD(VDD),.Y(g4229),.A(g4059));
  NOT NOT1_1981(.VSS(VSS),.VDD(VDD),.Y(I5674),.A(g4003));
  NOT NOT1_1982(.VSS(VSS),.VDD(VDD),.Y(g4232),.A(I5674));
  NOT NOT1_1983(.VSS(VSS),.VDD(VDD),.Y(I5686),.A(g3942));
  NOT NOT1_1984(.VSS(VSS),.VDD(VDD),.Y(g4242),.A(I5686));
  NOT NOT1_1985(.VSS(VSS),.VDD(VDD),.Y(I5692),.A(g3942));
  NOT NOT1_1986(.VSS(VSS),.VDD(VDD),.Y(g4246),.A(I5692));
  NOT NOT1_1987(.VSS(VSS),.VDD(VDD),.Y(I5696),.A(g3942));
  NOT NOT1_1988(.VSS(VSS),.VDD(VDD),.Y(g4248),.A(I5696));
  NOT NOT1_1989(.VSS(VSS),.VDD(VDD),.Y(I5699),.A(g3844));
  NOT NOT1_1990(.VSS(VSS),.VDD(VDD),.Y(g4249),.A(I5699));
  NOT NOT1_1991(.VSS(VSS),.VDD(VDD),.Y(I5702),.A(g3845));
  NOT NOT1_1992(.VSS(VSS),.VDD(VDD),.Y(g4250),.A(I5702));
  NOT NOT1_1993(.VSS(VSS),.VDD(VDD),.Y(I5705),.A(g3942));
  NOT NOT1_1994(.VSS(VSS),.VDD(VDD),.Y(g4251),.A(I5705));
  NOT NOT1_1995(.VSS(VSS),.VDD(VDD),.Y(I5708),.A(g3942));
  NOT NOT1_1996(.VSS(VSS),.VDD(VDD),.Y(g4252),.A(I5708));
  NOT NOT1_1997(.VSS(VSS),.VDD(VDD),.Y(I5713),.A(g4022));
  NOT NOT1_1998(.VSS(VSS),.VDD(VDD),.Y(g4262),.A(I5713));
  NOT NOT1_1999(.VSS(VSS),.VDD(VDD),.Y(I5716),.A(g3942));
  NOT NOT1_2000(.VSS(VSS),.VDD(VDD),.Y(g4265),.A(I5716));
  NOT NOT1_2001(.VSS(VSS),.VDD(VDD),.Y(I5720),.A(g4022));
  NOT NOT1_2002(.VSS(VSS),.VDD(VDD),.Y(g4267),.A(I5720));
  NOT NOT1_2003(.VSS(VSS),.VDD(VDD),.Y(I5723),.A(g3942));
  NOT NOT1_2004(.VSS(VSS),.VDD(VDD),.Y(g4270),.A(I5723));
  NOT NOT1_2005(.VSS(VSS),.VDD(VDD),.Y(I5728),.A(g4022));
  NOT NOT1_2006(.VSS(VSS),.VDD(VDD),.Y(g4273),.A(I5728));
  NOT NOT1_2007(.VSS(VSS),.VDD(VDD),.Y(I5731),.A(g3942));
  NOT NOT1_2008(.VSS(VSS),.VDD(VDD),.Y(g4276),.A(I5731));
  NOT NOT1_2009(.VSS(VSS),.VDD(VDD),.Y(I5736),.A(g4022));
  NOT NOT1_2010(.VSS(VSS),.VDD(VDD),.Y(g4281),.A(I5736));
  NOT NOT1_2011(.VSS(VSS),.VDD(VDD),.Y(I5739),.A(g3942));
  NOT NOT1_2012(.VSS(VSS),.VDD(VDD),.Y(g4284),.A(I5739));
  NOT NOT1_2013(.VSS(VSS),.VDD(VDD),.Y(I5743),.A(g4022));
  NOT NOT1_2014(.VSS(VSS),.VDD(VDD),.Y(g4286),.A(I5743));
  NOT NOT1_2015(.VSS(VSS),.VDD(VDD),.Y(I5746),.A(g4022));
  NOT NOT1_2016(.VSS(VSS),.VDD(VDD),.Y(g4289),.A(I5746));
  NOT NOT1_2017(.VSS(VSS),.VDD(VDD),.Y(g4292),.A(g4059));
  NOT NOT1_2018(.VSS(VSS),.VDD(VDD),.Y(I5750),.A(g4022));
  NOT NOT1_2019(.VSS(VSS),.VDD(VDD),.Y(g4293),.A(I5750));
  NOT NOT1_2020(.VSS(VSS),.VDD(VDD),.Y(I5753),.A(g4022));
  NOT NOT1_2021(.VSS(VSS),.VDD(VDD),.Y(g4296),.A(I5753));
  NOT NOT1_2022(.VSS(VSS),.VDD(VDD),.Y(I5756),.A(g3922));
  NOT NOT1_2023(.VSS(VSS),.VDD(VDD),.Y(g4299),.A(I5756));
  NOT NOT1_2024(.VSS(VSS),.VDD(VDD),.Y(g4302),.A(g4068));
  NOT NOT1_2025(.VSS(VSS),.VDD(VDD),.Y(I5774),.A(g3807));
  NOT NOT1_2026(.VSS(VSS),.VDD(VDD),.Y(g4307),.A(I5774));
  NOT NOT1_2027(.VSS(VSS),.VDD(VDD),.Y(I5777),.A(g3807));
  NOT NOT1_2028(.VSS(VSS),.VDD(VDD),.Y(g4308),.A(I5777));
  NOT NOT1_2029(.VSS(VSS),.VDD(VDD),.Y(g4309),.A(g4074));
  NOT NOT1_2030(.VSS(VSS),.VDD(VDD),.Y(g4314),.A(g4080));
  NOT NOT1_2031(.VSS(VSS),.VDD(VDD),.Y(g4320),.A(g4011));
  NOT NOT1_2032(.VSS(VSS),.VDD(VDD),.Y(I5790),.A(g3803));
  NOT NOT1_2033(.VSS(VSS),.VDD(VDD),.Y(g4321),.A(I5790));
  NOT NOT1_2034(.VSS(VSS),.VDD(VDD),.Y(I5793),.A(g3803));
  NOT NOT1_2035(.VSS(VSS),.VDD(VDD),.Y(g4322),.A(I5793));
  NOT NOT1_2036(.VSS(VSS),.VDD(VDD),.Y(g4323),.A(g4086));
  NOT NOT1_2037(.VSS(VSS),.VDD(VDD),.Y(g4328),.A(g4092));
  NOT NOT1_2038(.VSS(VSS),.VDD(VDD),.Y(g4334),.A(g3733));
  NOT NOT1_2039(.VSS(VSS),.VDD(VDD),.Y(g4343),.A(g4011));
  NOT NOT1_2040(.VSS(VSS),.VDD(VDD),.Y(g4350),.A(g4010));
  NOT NOT1_2041(.VSS(VSS),.VDD(VDD),.Y(I5825),.A(g3914));
  NOT NOT1_2042(.VSS(VSS),.VDD(VDD),.Y(g4364),.A(I5825));
  NOT NOT1_2043(.VSS(VSS),.VDD(VDD),.Y(I5831),.A(g3842));
  NOT NOT1_2044(.VSS(VSS),.VDD(VDD),.Y(g4370),.A(I5831));
  NOT NOT1_2045(.VSS(VSS),.VDD(VDD),.Y(I5837),.A(g3850));
  NOT NOT1_2046(.VSS(VSS),.VDD(VDD),.Y(g4374),.A(I5837));
  NOT NOT1_2047(.VSS(VSS),.VDD(VDD),.Y(I5840),.A(g3732));
  NOT NOT1_2048(.VSS(VSS),.VDD(VDD),.Y(g4375),.A(I5840));
  NOT NOT1_2049(.VSS(VSS),.VDD(VDD),.Y(I5843),.A(g3851));
  NOT NOT1_2050(.VSS(VSS),.VDD(VDD),.Y(g4376),.A(I5843));
  NOT NOT1_2051(.VSS(VSS),.VDD(VDD),.Y(I5848),.A(g3856));
  NOT NOT1_2052(.VSS(VSS),.VDD(VDD),.Y(g4379),.A(I5848));
  NOT NOT1_2053(.VSS(VSS),.VDD(VDD),.Y(I5851),.A(g3739));
  NOT NOT1_2054(.VSS(VSS),.VDD(VDD),.Y(g4380),.A(I5851));
  NOT NOT1_2055(.VSS(VSS),.VDD(VDD),.Y(I5854),.A(g3857));
  NOT NOT1_2056(.VSS(VSS),.VDD(VDD),.Y(g4381),.A(I5854));
  NOT NOT1_2057(.VSS(VSS),.VDD(VDD),.Y(I5857),.A(g3740));
  NOT NOT1_2058(.VSS(VSS),.VDD(VDD),.Y(g4382),.A(I5857));
  NOT NOT1_2059(.VSS(VSS),.VDD(VDD),.Y(I5862),.A(g3863));
  NOT NOT1_2060(.VSS(VSS),.VDD(VDD),.Y(g4385),.A(I5862));
  NOT NOT1_2061(.VSS(VSS),.VDD(VDD),.Y(I5865),.A(g3743));
  NOT NOT1_2062(.VSS(VSS),.VDD(VDD),.Y(g4386),.A(I5865));
  NOT NOT1_2063(.VSS(VSS),.VDD(VDD),.Y(I5868),.A(g3864));
  NOT NOT1_2064(.VSS(VSS),.VDD(VDD),.Y(g4387),.A(I5868));
  NOT NOT1_2065(.VSS(VSS),.VDD(VDD),.Y(I5871),.A(g3744));
  NOT NOT1_2066(.VSS(VSS),.VDD(VDD),.Y(g4388),.A(I5871));
  NOT NOT1_2067(.VSS(VSS),.VDD(VDD),.Y(I5876),.A(g3870));
  NOT NOT1_2068(.VSS(VSS),.VDD(VDD),.Y(g4391),.A(I5876));
  NOT NOT1_2069(.VSS(VSS),.VDD(VDD),.Y(I5879),.A(g3745));
  NOT NOT1_2070(.VSS(VSS),.VDD(VDD),.Y(g4392),.A(I5879));
  NOT NOT1_2071(.VSS(VSS),.VDD(VDD),.Y(I5882),.A(g3871));
  NOT NOT1_2072(.VSS(VSS),.VDD(VDD),.Y(g4393),.A(I5882));
  NOT NOT1_2073(.VSS(VSS),.VDD(VDD),.Y(I5885),.A(g3746));
  NOT NOT1_2074(.VSS(VSS),.VDD(VDD),.Y(g4394),.A(I5885));
  NOT NOT1_2075(.VSS(VSS),.VDD(VDD),.Y(I5890),.A(g3878));
  NOT NOT1_2076(.VSS(VSS),.VDD(VDD),.Y(g4397),.A(I5890));
  NOT NOT1_2077(.VSS(VSS),.VDD(VDD),.Y(I5893),.A(g3747));
  NOT NOT1_2078(.VSS(VSS),.VDD(VDD),.Y(g4398),.A(I5893));
  NOT NOT1_2079(.VSS(VSS),.VDD(VDD),.Y(I5896),.A(g3879));
  NOT NOT1_2080(.VSS(VSS),.VDD(VDD),.Y(g4399),.A(I5896));
  NOT NOT1_2081(.VSS(VSS),.VDD(VDD),.Y(I5899),.A(g3748));
  NOT NOT1_2082(.VSS(VSS),.VDD(VDD),.Y(g4400),.A(I5899));
  NOT NOT1_2083(.VSS(VSS),.VDD(VDD),.Y(g4402),.A(g4017));
  NOT NOT1_2084(.VSS(VSS),.VDD(VDD),.Y(I5904),.A(g3749));
  NOT NOT1_2085(.VSS(VSS),.VDD(VDD),.Y(g4403),.A(I5904));
  NOT NOT1_2086(.VSS(VSS),.VDD(VDD),.Y(I5907),.A(g3883));
  NOT NOT1_2087(.VSS(VSS),.VDD(VDD),.Y(g4404),.A(I5907));
  NOT NOT1_2088(.VSS(VSS),.VDD(VDD),.Y(I5910),.A(g3750));
  NOT NOT1_2089(.VSS(VSS),.VDD(VDD),.Y(g4405),.A(I5910));
  NOT NOT1_2090(.VSS(VSS),.VDD(VDD),.Y(I5913),.A(g3751));
  NOT NOT1_2091(.VSS(VSS),.VDD(VDD),.Y(g4406),.A(I5913));
  NOT NOT1_2092(.VSS(VSS),.VDD(VDD),.Y(g4422),.A(g4111));
  NOT NOT1_2093(.VSS(VSS),.VDD(VDD),.Y(I5920),.A(g4228));
  NOT NOT1_2094(.VSS(VSS),.VDD(VDD),.Y(g4423),.A(I5920));
  NOT NOT1_2095(.VSS(VSS),.VDD(VDD),.Y(I5923),.A(g4299));
  NOT NOT1_2096(.VSS(VSS),.VDD(VDD),.Y(g4424),.A(I5923));
  NOT NOT1_2097(.VSS(VSS),.VDD(VDD),.Y(I5926),.A(g4153));
  NOT NOT1_2098(.VSS(VSS),.VDD(VDD),.Y(g4425),.A(I5926));
  NOT NOT1_2099(.VSS(VSS),.VDD(VDD),.Y(I5929),.A(g4152));
  NOT NOT1_2100(.VSS(VSS),.VDD(VDD),.Y(g4426),.A(I5929));
  NOT NOT1_2101(.VSS(VSS),.VDD(VDD),.Y(I5933),.A(g4346));
  NOT NOT1_2102(.VSS(VSS),.VDD(VDD),.Y(g4428),.A(I5933));
  NOT NOT1_2103(.VSS(VSS),.VDD(VDD),.Y(I5938),.A(g4351));
  NOT NOT1_2104(.VSS(VSS),.VDD(VDD),.Y(g4431),.A(I5938));
  NOT NOT1_2105(.VSS(VSS),.VDD(VDD),.Y(I5944),.A(g4356));
  NOT NOT1_2106(.VSS(VSS),.VDD(VDD),.Y(g4435),.A(I5944));
  NOT NOT1_2107(.VSS(VSS),.VDD(VDD),.Y(I5948),.A(g4360));
  NOT NOT1_2108(.VSS(VSS),.VDD(VDD),.Y(g4437),.A(I5948));
  NOT NOT1_2109(.VSS(VSS),.VDD(VDD),.Y(I5952),.A(g4367));
  NOT NOT1_2110(.VSS(VSS),.VDD(VDD),.Y(g4439),.A(I5952));
  NOT NOT1_2111(.VSS(VSS),.VDD(VDD),.Y(I5977),.A(g4319));
  NOT NOT1_2112(.VSS(VSS),.VDD(VDD),.Y(g4462),.A(I5977));
  NOT NOT1_2113(.VSS(VSS),.VDD(VDD),.Y(g4463),.A(g4364));
  NOT NOT1_2114(.VSS(VSS),.VDD(VDD),.Y(I5987),.A(g4224));
  NOT NOT1_2115(.VSS(VSS),.VDD(VDD),.Y(g4485),.A(I5987));
  NOT NOT1_2116(.VSS(VSS),.VDD(VDD),.Y(I5991),.A(g4226));
  NOT NOT1_2117(.VSS(VSS),.VDD(VDD),.Y(g4487),.A(I5991));
  NOT NOT1_2118(.VSS(VSS),.VDD(VDD),.Y(I5998),.A(g4157));
  NOT NOT1_2119(.VSS(VSS),.VDD(VDD),.Y(g4492),.A(I5998));
  NOT NOT1_2120(.VSS(VSS),.VDD(VDD),.Y(I6001),.A(g4162));
  NOT NOT1_2121(.VSS(VSS),.VDD(VDD),.Y(g4493),.A(I6001));
  NOT NOT1_2122(.VSS(VSS),.VDD(VDD),.Y(I6004),.A(g4159));
  NOT NOT1_2123(.VSS(VSS),.VDD(VDD),.Y(g4494),.A(I6004));
  NOT NOT1_2124(.VSS(VSS),.VDD(VDD),.Y(I6008),.A(g4163));
  NOT NOT1_2125(.VSS(VSS),.VDD(VDD),.Y(g4496),.A(I6008));
  NOT NOT1_2126(.VSS(VSS),.VDD(VDD),.Y(I6012),.A(g4167));
  NOT NOT1_2127(.VSS(VSS),.VDD(VDD),.Y(g4498),.A(I6012));
  NOT NOT1_2128(.VSS(VSS),.VDD(VDD),.Y(I6015),.A(g4170));
  NOT NOT1_2129(.VSS(VSS),.VDD(VDD),.Y(g4499),.A(I6015));
  NOT NOT1_2130(.VSS(VSS),.VDD(VDD),.Y(I6020),.A(g4176));
  NOT NOT1_2131(.VSS(VSS),.VDD(VDD),.Y(g4502),.A(I6020));
  NOT NOT1_2132(.VSS(VSS),.VDD(VDD),.Y(I6023),.A(g4151));
  NOT NOT1_2133(.VSS(VSS),.VDD(VDD),.Y(g4503),.A(I6023));
  NOT NOT1_2134(.VSS(VSS),.VDD(VDD),.Y(I6033),.A(g4179));
  NOT NOT1_2135(.VSS(VSS),.VDD(VDD),.Y(g4507),.A(I6033));
  NOT NOT1_2136(.VSS(VSS),.VDD(VDD),.Y(I6036),.A(g4370));
  NOT NOT1_2137(.VSS(VSS),.VDD(VDD),.Y(g4508),.A(I6036));
  NOT NOT1_2138(.VSS(VSS),.VDD(VDD),.Y(I6039),.A(g4182));
  NOT NOT1_2139(.VSS(VSS),.VDD(VDD),.Y(g4509),.A(I6039));
  NOT NOT1_2140(.VSS(VSS),.VDD(VDD),.Y(I6042),.A(g4374));
  NOT NOT1_2141(.VSS(VSS),.VDD(VDD),.Y(g4510),.A(I6042));
  NOT NOT1_2142(.VSS(VSS),.VDD(VDD),.Y(I6045),.A(g4375));
  NOT NOT1_2143(.VSS(VSS),.VDD(VDD),.Y(g4511),.A(I6045));
  NOT NOT1_2144(.VSS(VSS),.VDD(VDD),.Y(I6048),.A(g4376));
  NOT NOT1_2145(.VSS(VSS),.VDD(VDD),.Y(g4512),.A(I6048));
  NOT NOT1_2146(.VSS(VSS),.VDD(VDD),.Y(I6051),.A(g4185));
  NOT NOT1_2147(.VSS(VSS),.VDD(VDD),.Y(g4513),.A(I6051));
  NOT NOT1_2148(.VSS(VSS),.VDD(VDD),.Y(I6054),.A(g4194));
  NOT NOT1_2149(.VSS(VSS),.VDD(VDD),.Y(g4514),.A(I6054));
  NOT NOT1_2150(.VSS(VSS),.VDD(VDD),.Y(I6057),.A(g4379));
  NOT NOT1_2151(.VSS(VSS),.VDD(VDD),.Y(g4515),.A(I6057));
  NOT NOT1_2152(.VSS(VSS),.VDD(VDD),.Y(I6060),.A(g4380));
  NOT NOT1_2153(.VSS(VSS),.VDD(VDD),.Y(g4516),.A(I6060));
  NOT NOT1_2154(.VSS(VSS),.VDD(VDD),.Y(I6063),.A(g4381));
  NOT NOT1_2155(.VSS(VSS),.VDD(VDD),.Y(g4517),.A(I6063));
  NOT NOT1_2156(.VSS(VSS),.VDD(VDD),.Y(I6066),.A(g4382));
  NOT NOT1_2157(.VSS(VSS),.VDD(VDD),.Y(g4518),.A(I6066));
  NOT NOT1_2158(.VSS(VSS),.VDD(VDD),.Y(I6069),.A(g4213));
  NOT NOT1_2159(.VSS(VSS),.VDD(VDD),.Y(g4519),.A(I6069));
  NOT NOT1_2160(.VSS(VSS),.VDD(VDD),.Y(I6072),.A(g4385));
  NOT NOT1_2161(.VSS(VSS),.VDD(VDD),.Y(g4520),.A(I6072));
  NOT NOT1_2162(.VSS(VSS),.VDD(VDD),.Y(I6075),.A(g4386));
  NOT NOT1_2163(.VSS(VSS),.VDD(VDD),.Y(g4521),.A(I6075));
  NOT NOT1_2164(.VSS(VSS),.VDD(VDD),.Y(I6078),.A(g4387));
  NOT NOT1_2165(.VSS(VSS),.VDD(VDD),.Y(g4522),.A(I6078));
  NOT NOT1_2166(.VSS(VSS),.VDD(VDD),.Y(I6081),.A(g4388));
  NOT NOT1_2167(.VSS(VSS),.VDD(VDD),.Y(g4523),.A(I6081));
  NOT NOT1_2168(.VSS(VSS),.VDD(VDD),.Y(I6084),.A(g4391));
  NOT NOT1_2169(.VSS(VSS),.VDD(VDD),.Y(g4524),.A(I6084));
  NOT NOT1_2170(.VSS(VSS),.VDD(VDD),.Y(I6087),.A(g4392));
  NOT NOT1_2171(.VSS(VSS),.VDD(VDD),.Y(g4525),.A(I6087));
  NOT NOT1_2172(.VSS(VSS),.VDD(VDD),.Y(I6090),.A(g4393));
  NOT NOT1_2173(.VSS(VSS),.VDD(VDD),.Y(g4526),.A(I6090));
  NOT NOT1_2174(.VSS(VSS),.VDD(VDD),.Y(I6093),.A(g4394));
  NOT NOT1_2175(.VSS(VSS),.VDD(VDD),.Y(g4527),.A(I6093));
  NOT NOT1_2176(.VSS(VSS),.VDD(VDD),.Y(I6096),.A(g4397));
  NOT NOT1_2177(.VSS(VSS),.VDD(VDD),.Y(g4528),.A(I6096));
  NOT NOT1_2178(.VSS(VSS),.VDD(VDD),.Y(I6099),.A(g4398));
  NOT NOT1_2179(.VSS(VSS),.VDD(VDD),.Y(g4529),.A(I6099));
  NOT NOT1_2180(.VSS(VSS),.VDD(VDD),.Y(I6102),.A(g4399));
  NOT NOT1_2181(.VSS(VSS),.VDD(VDD),.Y(g4530),.A(I6102));
  NOT NOT1_2182(.VSS(VSS),.VDD(VDD),.Y(I6105),.A(g4400));
  NOT NOT1_2183(.VSS(VSS),.VDD(VDD),.Y(g4531),.A(I6105));
  NOT NOT1_2184(.VSS(VSS),.VDD(VDD),.Y(I6108),.A(g4403));
  NOT NOT1_2185(.VSS(VSS),.VDD(VDD),.Y(g4532),.A(I6108));
  NOT NOT1_2186(.VSS(VSS),.VDD(VDD),.Y(I6111),.A(g4404));
  NOT NOT1_2187(.VSS(VSS),.VDD(VDD),.Y(g4533),.A(I6111));
  NOT NOT1_2188(.VSS(VSS),.VDD(VDD),.Y(I6114),.A(g4405));
  NOT NOT1_2189(.VSS(VSS),.VDD(VDD),.Y(g4534),.A(I6114));
  NOT NOT1_2190(.VSS(VSS),.VDD(VDD),.Y(g4535),.A(g4173));
  NOT NOT1_2191(.VSS(VSS),.VDD(VDD),.Y(I6118),.A(g4406));
  NOT NOT1_2192(.VSS(VSS),.VDD(VDD),.Y(g4536),.A(I6118));
  NOT NOT1_2193(.VSS(VSS),.VDD(VDD),.Y(g4537),.A(g4410));
  NOT NOT1_2194(.VSS(VSS),.VDD(VDD),.Y(g4545),.A(g4416));
  NOT NOT1_2195(.VSS(VSS),.VDD(VDD),.Y(I6126),.A(g4240));
  NOT NOT1_2196(.VSS(VSS),.VDD(VDD),.Y(g4550),.A(I6126));
  NOT NOT1_2197(.VSS(VSS),.VDD(VDD),.Y(g4559),.A(g4187));
  NOT NOT1_2198(.VSS(VSS),.VDD(VDD),.Y(g4560),.A(g4188));
  NOT NOT1_2199(.VSS(VSS),.VDD(VDD),.Y(g4561),.A(g4189));
  NOT NOT1_2200(.VSS(VSS),.VDD(VDD),.Y(I6132),.A(g4219));
  NOT NOT1_2201(.VSS(VSS),.VDD(VDD),.Y(g4562),.A(I6132));
  NOT NOT1_2202(.VSS(VSS),.VDD(VDD),.Y(g4563),.A(g4190));
  NOT NOT1_2203(.VSS(VSS),.VDD(VDD),.Y(g4564),.A(g4192));
  NOT NOT1_2204(.VSS(VSS),.VDD(VDD),.Y(g4565),.A(g4195));
  NOT NOT1_2205(.VSS(VSS),.VDD(VDD),.Y(g4566),.A(g4198));
  NOT NOT1_2206(.VSS(VSS),.VDD(VDD),.Y(I6139),.A(g4222));
  NOT NOT1_2207(.VSS(VSS),.VDD(VDD),.Y(g4567),.A(I6139));
  NOT NOT1_2208(.VSS(VSS),.VDD(VDD),.Y(I6143),.A(g4237));
  NOT NOT1_2209(.VSS(VSS),.VDD(VDD),.Y(g4569),.A(I6143));
  NOT NOT1_2210(.VSS(VSS),.VDD(VDD),.Y(g4577),.A(g4202));
  NOT NOT1_2211(.VSS(VSS),.VDD(VDD),.Y(g4579),.A(g4206));
  NOT NOT1_2212(.VSS(VSS),.VDD(VDD),.Y(g4582),.A(g4210));
  NOT NOT1_2213(.VSS(VSS),.VDD(VDD),.Y(g4587),.A(g4215));
  NOT NOT1_2214(.VSS(VSS),.VDD(VDD),.Y(g4601),.A(g4191));
  NOT NOT1_2215(.VSS(VSS),.VDD(VDD),.Y(I6170),.A(g4343));
  NOT NOT1_2216(.VSS(VSS),.VDD(VDD),.Y(g4603),.A(I6170));
  NOT NOT1_2217(.VSS(VSS),.VDD(VDD),.Y(g4606),.A(g4193));
  NOT NOT1_2218(.VSS(VSS),.VDD(VDD),.Y(I6182),.A(g4249));
  NOT NOT1_2219(.VSS(VSS),.VDD(VDD),.Y(g4609),.A(I6182));
  NOT NOT1_2220(.VSS(VSS),.VDD(VDD),.Y(g4612),.A(g4320));
  NOT NOT1_2221(.VSS(VSS),.VDD(VDD),.Y(g4614),.A(g4308));
  NOT NOT1_2222(.VSS(VSS),.VDD(VDD),.Y(g4615),.A(g4322));
  NOT NOT1_2223(.VSS(VSS),.VDD(VDD),.Y(g4617),.A(g4242));
  NOT NOT1_2224(.VSS(VSS),.VDD(VDD),.Y(g4618),.A(g4246));
  NOT NOT1_2225(.VSS(VSS),.VDD(VDD),.Y(g4619),.A(g4248));
  NOT NOT1_2226(.VSS(VSS),.VDD(VDD),.Y(g4620),.A(g4251));
  NOT NOT1_2227(.VSS(VSS),.VDD(VDD),.Y(g4622),.A(g4252));
  NOT NOT1_2228(.VSS(VSS),.VDD(VDD),.Y(g4623),.A(g4262));
  NOT NOT1_2229(.VSS(VSS),.VDD(VDD),.Y(g4624),.A(g4265));
  NOT NOT1_2230(.VSS(VSS),.VDD(VDD),.Y(g4625),.A(g4267));
  NOT NOT1_2231(.VSS(VSS),.VDD(VDD),.Y(g4626),.A(g4270));
  NOT NOT1_2232(.VSS(VSS),.VDD(VDD),.Y(g4628),.A(g4273));
  NOT NOT1_2233(.VSS(VSS),.VDD(VDD),.Y(g4629),.A(g4276));
  NOT NOT1_2234(.VSS(VSS),.VDD(VDD),.Y(g4632),.A(g4281));
  NOT NOT1_2235(.VSS(VSS),.VDD(VDD),.Y(g4633),.A(g4284));
  NOT NOT1_2236(.VSS(VSS),.VDD(VDD),.Y(g4636),.A(g4286));
  NOT NOT1_2237(.VSS(VSS),.VDD(VDD),.Y(g4639),.A(g4289));
  NOT NOT1_2238(.VSS(VSS),.VDD(VDD),.Y(g4643),.A(g4293));
  NOT NOT1_2239(.VSS(VSS),.VDD(VDD),.Y(I6231),.A(g4350));
  NOT NOT1_2240(.VSS(VSS),.VDD(VDD),.Y(g4644),.A(I6231));
  NOT NOT1_2241(.VSS(VSS),.VDD(VDD),.Y(g4647),.A(g4296));
  NOT NOT1_2242(.VSS(VSS),.VDD(VDD),.Y(I6244),.A(g4519));
  NOT NOT1_2243(.VSS(VSS),.VDD(VDD),.Y(g4657),.A(I6244));
  NOT NOT1_2244(.VSS(VSS),.VDD(VDD),.Y(I6247),.A(g4609));
  NOT NOT1_2245(.VSS(VSS),.VDD(VDD),.Y(g4658),.A(I6247));
  NOT NOT1_2246(.VSS(VSS),.VDD(VDD),.Y(I6250),.A(g4514));
  NOT NOT1_2247(.VSS(VSS),.VDD(VDD),.Y(g4659),.A(I6250));
  NOT NOT1_2248(.VSS(VSS),.VDD(VDD),.Y(I6253),.A(g4608));
  NOT NOT1_2249(.VSS(VSS),.VDD(VDD),.Y(g4660),.A(I6253));
  NOT NOT1_2250(.VSS(VSS),.VDD(VDD),.Y(g4662),.A(g4640));
  NOT NOT1_2251(.VSS(VSS),.VDD(VDD),.Y(I6269),.A(g4655));
  NOT NOT1_2252(.VSS(VSS),.VDD(VDD),.Y(g4679),.A(I6269));
  NOT NOT1_2253(.VSS(VSS),.VDD(VDD),.Y(I6280),.A(g4430));
  NOT NOT1_2254(.VSS(VSS),.VDD(VDD),.Y(g4692),.A(I6280));
  NOT NOT1_2255(.VSS(VSS),.VDD(VDD),.Y(I6283),.A(g4613));
  NOT NOT1_2256(.VSS(VSS),.VDD(VDD),.Y(g4693),.A(I6283));
  NOT NOT1_2257(.VSS(VSS),.VDD(VDD),.Y(I6289),.A(g4433));
  NOT NOT1_2258(.VSS(VSS),.VDD(VDD),.Y(g4699),.A(I6289));
  NOT NOT1_2259(.VSS(VSS),.VDD(VDD),.Y(I6292),.A(g4434));
  NOT NOT1_2260(.VSS(VSS),.VDD(VDD),.Y(g4700),.A(I6292));
  NOT NOT1_2261(.VSS(VSS),.VDD(VDD),.Y(I6296),.A(g4436));
  NOT NOT1_2262(.VSS(VSS),.VDD(VDD),.Y(g4702),.A(I6296));
  NOT NOT1_2263(.VSS(VSS),.VDD(VDD),.Y(I6299),.A(g4438));
  NOT NOT1_2264(.VSS(VSS),.VDD(VDD),.Y(g4703),.A(I6299));
  NOT NOT1_2265(.VSS(VSS),.VDD(VDD),.Y(I6302),.A(g4440));
  NOT NOT1_2266(.VSS(VSS),.VDD(VDD),.Y(g4704),.A(I6302));
  NOT NOT1_2267(.VSS(VSS),.VDD(VDD),.Y(I6305),.A(g4441));
  NOT NOT1_2268(.VSS(VSS),.VDD(VDD),.Y(g4705),.A(I6305));
  NOT NOT1_2269(.VSS(VSS),.VDD(VDD),.Y(I6308),.A(g4443));
  NOT NOT1_2270(.VSS(VSS),.VDD(VDD),.Y(g4706),.A(I6308));
  NOT NOT1_2271(.VSS(VSS),.VDD(VDD),.Y(I6311),.A(g4444));
  NOT NOT1_2272(.VSS(VSS),.VDD(VDD),.Y(g4707),.A(I6311));
  NOT NOT1_2273(.VSS(VSS),.VDD(VDD),.Y(I6315),.A(g4446));
  NOT NOT1_2274(.VSS(VSS),.VDD(VDD),.Y(g4711),.A(I6315));
  NOT NOT1_2275(.VSS(VSS),.VDD(VDD),.Y(I6318),.A(g4447));
  NOT NOT1_2276(.VSS(VSS),.VDD(VDD),.Y(g4712),.A(I6318));
  NOT NOT1_2277(.VSS(VSS),.VDD(VDD),.Y(I6321),.A(g4559));
  NOT NOT1_2278(.VSS(VSS),.VDD(VDD),.Y(g4713),.A(I6321));
  NOT NOT1_2279(.VSS(VSS),.VDD(VDD),.Y(I6324),.A(g4450));
  NOT NOT1_2280(.VSS(VSS),.VDD(VDD),.Y(g4714),.A(I6324));
  NOT NOT1_2281(.VSS(VSS),.VDD(VDD),.Y(I6327),.A(g4451));
  NOT NOT1_2282(.VSS(VSS),.VDD(VDD),.Y(g4715),.A(I6327));
  NOT NOT1_2283(.VSS(VSS),.VDD(VDD),.Y(I6330),.A(g4560));
  NOT NOT1_2284(.VSS(VSS),.VDD(VDD),.Y(g4716),.A(I6330));
  NOT NOT1_2285(.VSS(VSS),.VDD(VDD),.Y(g4717),.A(g4465));
  NOT NOT1_2286(.VSS(VSS),.VDD(VDD),.Y(I6334),.A(g4454));
  NOT NOT1_2287(.VSS(VSS),.VDD(VDD),.Y(g4718),.A(I6334));
  NOT NOT1_2288(.VSS(VSS),.VDD(VDD),.Y(I6337),.A(g4455));
  NOT NOT1_2289(.VSS(VSS),.VDD(VDD),.Y(g4719),.A(I6337));
  NOT NOT1_2290(.VSS(VSS),.VDD(VDD),.Y(I6340),.A(g4561));
  NOT NOT1_2291(.VSS(VSS),.VDD(VDD),.Y(g4720),.A(I6340));
  NOT NOT1_2292(.VSS(VSS),.VDD(VDD),.Y(I6343),.A(g4458));
  NOT NOT1_2293(.VSS(VSS),.VDD(VDD),.Y(g4721),.A(I6343));
  NOT NOT1_2294(.VSS(VSS),.VDD(VDD),.Y(I6346),.A(g4563));
  NOT NOT1_2295(.VSS(VSS),.VDD(VDD),.Y(g4722),.A(I6346));
  NOT NOT1_2296(.VSS(VSS),.VDD(VDD),.Y(I6349),.A(g4569));
  NOT NOT1_2297(.VSS(VSS),.VDD(VDD),.Y(g4723),.A(I6349));
  NOT NOT1_2298(.VSS(VSS),.VDD(VDD),.Y(I6352),.A(g4564));
  NOT NOT1_2299(.VSS(VSS),.VDD(VDD),.Y(g4726),.A(I6352));
  NOT NOT1_2300(.VSS(VSS),.VDD(VDD),.Y(I6355),.A(g4569));
  NOT NOT1_2301(.VSS(VSS),.VDD(VDD),.Y(g4727),.A(I6355));
  NOT NOT1_2302(.VSS(VSS),.VDD(VDD),.Y(I6359),.A(g4566));
  NOT NOT1_2303(.VSS(VSS),.VDD(VDD),.Y(g4731),.A(I6359));
  NOT NOT1_2304(.VSS(VSS),.VDD(VDD),.Y(I6362),.A(g4569));
  NOT NOT1_2305(.VSS(VSS),.VDD(VDD),.Y(g4732),.A(I6362));
  NOT NOT1_2306(.VSS(VSS),.VDD(VDD),.Y(I6366),.A(g4569));
  NOT NOT1_2307(.VSS(VSS),.VDD(VDD),.Y(g4736),.A(I6366));
  NOT NOT1_2308(.VSS(VSS),.VDD(VDD),.Y(I6371),.A(g4569));
  NOT NOT1_2309(.VSS(VSS),.VDD(VDD),.Y(g4741),.A(I6371));
  NOT NOT1_2310(.VSS(VSS),.VDD(VDD),.Y(I6377),.A(g4569));
  NOT NOT1_2311(.VSS(VSS),.VDD(VDD),.Y(g4753),.A(I6377));
  NOT NOT1_2312(.VSS(VSS),.VDD(VDD),.Y(I6382),.A(g4460));
  NOT NOT1_2313(.VSS(VSS),.VDD(VDD),.Y(g4758),.A(I6382));
  NOT NOT1_2314(.VSS(VSS),.VDD(VDD),.Y(I6386),.A(g4462));
  NOT NOT1_2315(.VSS(VSS),.VDD(VDD),.Y(g4760),.A(I6386));
  NOT NOT1_2316(.VSS(VSS),.VDD(VDD),.Y(I6397),.A(g4473));
  NOT NOT1_2317(.VSS(VSS),.VDD(VDD),.Y(g4763),.A(I6397));
  NOT NOT1_2318(.VSS(VSS),.VDD(VDD),.Y(I6400),.A(g4473));
  NOT NOT1_2319(.VSS(VSS),.VDD(VDD),.Y(g4764),.A(I6400));
  NOT NOT1_2320(.VSS(VSS),.VDD(VDD),.Y(I6403),.A(g4492));
  NOT NOT1_2321(.VSS(VSS),.VDD(VDD),.Y(g4765),.A(I6403));
  NOT NOT1_2322(.VSS(VSS),.VDD(VDD),.Y(I6406),.A(g4473));
  NOT NOT1_2323(.VSS(VSS),.VDD(VDD),.Y(g4766),.A(I6406));
  NOT NOT1_2324(.VSS(VSS),.VDD(VDD),.Y(g4767),.A(g4601));
  NOT NOT1_2325(.VSS(VSS),.VDD(VDD),.Y(I6410),.A(g4473));
  NOT NOT1_2326(.VSS(VSS),.VDD(VDD),.Y(g4768),.A(I6410));
  NOT NOT1_2327(.VSS(VSS),.VDD(VDD),.Y(g4769),.A(g4606));
  NOT NOT1_2328(.VSS(VSS),.VDD(VDD),.Y(I6414),.A(g4497));
  NOT NOT1_2329(.VSS(VSS),.VDD(VDD),.Y(g4770),.A(I6414));
  NOT NOT1_2330(.VSS(VSS),.VDD(VDD),.Y(I6417),.A(g4617));
  NOT NOT1_2331(.VSS(VSS),.VDD(VDD),.Y(g4771),.A(I6417));
  NOT NOT1_2332(.VSS(VSS),.VDD(VDD),.Y(I6420),.A(g4618));
  NOT NOT1_2333(.VSS(VSS),.VDD(VDD),.Y(g4772),.A(I6420));
  NOT NOT1_2334(.VSS(VSS),.VDD(VDD),.Y(I6425),.A(g4619));
  NOT NOT1_2335(.VSS(VSS),.VDD(VDD),.Y(g4775),.A(I6425));
  NOT NOT1_2336(.VSS(VSS),.VDD(VDD),.Y(I6430),.A(g4620));
  NOT NOT1_2337(.VSS(VSS),.VDD(VDD),.Y(g4778),.A(I6430));
  NOT NOT1_2338(.VSS(VSS),.VDD(VDD),.Y(I6434),.A(g4622));
  NOT NOT1_2339(.VSS(VSS),.VDD(VDD),.Y(g4780),.A(I6434));
  NOT NOT1_2340(.VSS(VSS),.VDD(VDD),.Y(I6437),.A(g4501));
  NOT NOT1_2341(.VSS(VSS),.VDD(VDD),.Y(g4781),.A(I6437));
  NOT NOT1_2342(.VSS(VSS),.VDD(VDD),.Y(I6441),.A(g4624));
  NOT NOT1_2343(.VSS(VSS),.VDD(VDD),.Y(g4783),.A(I6441));
  NOT NOT1_2344(.VSS(VSS),.VDD(VDD),.Y(I6444),.A(g4503));
  NOT NOT1_2345(.VSS(VSS),.VDD(VDD),.Y(g4784),.A(I6444));
  NOT NOT1_2346(.VSS(VSS),.VDD(VDD),.Y(I6448),.A(g4626));
  NOT NOT1_2347(.VSS(VSS),.VDD(VDD),.Y(g4786),.A(I6448));
  NOT NOT1_2348(.VSS(VSS),.VDD(VDD),.Y(I6452),.A(g4629));
  NOT NOT1_2349(.VSS(VSS),.VDD(VDD),.Y(g4788),.A(I6452));
  NOT NOT1_2350(.VSS(VSS),.VDD(VDD),.Y(I6456),.A(g4633));
  NOT NOT1_2351(.VSS(VSS),.VDD(VDD),.Y(g4790),.A(I6456));
  NOT NOT1_2352(.VSS(VSS),.VDD(VDD),.Y(I6464),.A(g4562));
  NOT NOT1_2353(.VSS(VSS),.VDD(VDD),.Y(g4798),.A(I6464));
  NOT NOT1_2354(.VSS(VSS),.VDD(VDD),.Y(g4799),.A(g4485));
  NOT NOT1_2355(.VSS(VSS),.VDD(VDD),.Y(g4801),.A(g4487));
  NOT NOT1_2356(.VSS(VSS),.VDD(VDD),.Y(I6470),.A(g4473));
  NOT NOT1_2357(.VSS(VSS),.VDD(VDD),.Y(g4802),.A(I6470));
  NOT NOT1_2358(.VSS(VSS),.VDD(VDD),.Y(g4804),.A(g4473));
  NOT NOT1_2359(.VSS(VSS),.VDD(VDD),.Y(g4805),.A(g4473));
  NOT NOT1_2360(.VSS(VSS),.VDD(VDD),.Y(g4806),.A(g4473));
  NOT NOT1_2361(.VSS(VSS),.VDD(VDD),.Y(g4807),.A(g4473));
  NOT NOT1_2362(.VSS(VSS),.VDD(VDD),.Y(g4808),.A(g4473));
  NOT NOT1_2363(.VSS(VSS),.VDD(VDD),.Y(I6485),.A(g4603));
  NOT NOT1_2364(.VSS(VSS),.VDD(VDD),.Y(g4809),.A(I6485));
  NOT NOT1_2365(.VSS(VSS),.VDD(VDD),.Y(I6488),.A(g4603));
  NOT NOT1_2366(.VSS(VSS),.VDD(VDD),.Y(g4810),.A(I6488));
  NOT NOT1_2367(.VSS(VSS),.VDD(VDD),.Y(I6495),.A(g4607));
  NOT NOT1_2368(.VSS(VSS),.VDD(VDD),.Y(g4815),.A(I6495));
  NOT NOT1_2369(.VSS(VSS),.VDD(VDD),.Y(g4822),.A(g4614));
  NOT NOT1_2370(.VSS(VSS),.VDD(VDD),.Y(I6507),.A(g4644));
  NOT NOT1_2371(.VSS(VSS),.VDD(VDD),.Y(g4823),.A(I6507));
  NOT NOT1_2372(.VSS(VSS),.VDD(VDD),.Y(g4824),.A(g4615));
  NOT NOT1_2373(.VSS(VSS),.VDD(VDD),.Y(g4837),.A(g4473));
  NOT NOT1_2374(.VSS(VSS),.VDD(VDD),.Y(I6525),.A(g4770));
  NOT NOT1_2375(.VSS(VSS),.VDD(VDD),.Y(g4839),.A(I6525));
  NOT NOT1_2376(.VSS(VSS),.VDD(VDD),.Y(I6528),.A(g4815));
  NOT NOT1_2377(.VSS(VSS),.VDD(VDD),.Y(g4840),.A(I6528));
  NOT NOT1_2378(.VSS(VSS),.VDD(VDD),.Y(I6531),.A(g4704));
  NOT NOT1_2379(.VSS(VSS),.VDD(VDD),.Y(g4841),.A(I6531));
  NOT NOT1_2380(.VSS(VSS),.VDD(VDD),.Y(I6534),.A(g4706));
  NOT NOT1_2381(.VSS(VSS),.VDD(VDD),.Y(g4842),.A(I6534));
  NOT NOT1_2382(.VSS(VSS),.VDD(VDD),.Y(I6537),.A(g4711));
  NOT NOT1_2383(.VSS(VSS),.VDD(VDD),.Y(g4843),.A(I6537));
  NOT NOT1_2384(.VSS(VSS),.VDD(VDD),.Y(I6540),.A(g4714));
  NOT NOT1_2385(.VSS(VSS),.VDD(VDD),.Y(g4844),.A(I6540));
  NOT NOT1_2386(.VSS(VSS),.VDD(VDD),.Y(I6543),.A(g4718));
  NOT NOT1_2387(.VSS(VSS),.VDD(VDD),.Y(g4845),.A(I6543));
  NOT NOT1_2388(.VSS(VSS),.VDD(VDD),.Y(I6546),.A(g4692));
  NOT NOT1_2389(.VSS(VSS),.VDD(VDD),.Y(g4846),.A(I6546));
  NOT NOT1_2390(.VSS(VSS),.VDD(VDD),.Y(I6549),.A(g4699));
  NOT NOT1_2391(.VSS(VSS),.VDD(VDD),.Y(g4847),.A(I6549));
  NOT NOT1_2392(.VSS(VSS),.VDD(VDD),.Y(I6552),.A(g4702));
  NOT NOT1_2393(.VSS(VSS),.VDD(VDD),.Y(g4848),.A(I6552));
  NOT NOT1_2394(.VSS(VSS),.VDD(VDD),.Y(I6555),.A(g4703));
  NOT NOT1_2395(.VSS(VSS),.VDD(VDD),.Y(g4849),.A(I6555));
  NOT NOT1_2396(.VSS(VSS),.VDD(VDD),.Y(I6558),.A(g4705));
  NOT NOT1_2397(.VSS(VSS),.VDD(VDD),.Y(g4850),.A(I6558));
  NOT NOT1_2398(.VSS(VSS),.VDD(VDD),.Y(I6561),.A(g4707));
  NOT NOT1_2399(.VSS(VSS),.VDD(VDD),.Y(g4851),.A(I6561));
  NOT NOT1_2400(.VSS(VSS),.VDD(VDD),.Y(I6564),.A(g4712));
  NOT NOT1_2401(.VSS(VSS),.VDD(VDD),.Y(g4852),.A(I6564));
  NOT NOT1_2402(.VSS(VSS),.VDD(VDD),.Y(I6567),.A(g4715));
  NOT NOT1_2403(.VSS(VSS),.VDD(VDD),.Y(g4853),.A(I6567));
  NOT NOT1_2404(.VSS(VSS),.VDD(VDD),.Y(I6570),.A(g4719));
  NOT NOT1_2405(.VSS(VSS),.VDD(VDD),.Y(g4854),.A(I6570));
  NOT NOT1_2406(.VSS(VSS),.VDD(VDD),.Y(I6573),.A(g4721));
  NOT NOT1_2407(.VSS(VSS),.VDD(VDD),.Y(g4855),.A(I6573));
  NOT NOT1_2408(.VSS(VSS),.VDD(VDD),.Y(I6576),.A(g4700));
  NOT NOT1_2409(.VSS(VSS),.VDD(VDD),.Y(g4856),.A(I6576));
  NOT NOT1_2410(.VSS(VSS),.VDD(VDD),.Y(I6579),.A(g4798));
  NOT NOT1_2411(.VSS(VSS),.VDD(VDD),.Y(g4857),.A(I6579));
  NOT NOT1_2412(.VSS(VSS),.VDD(VDD),.Y(I6582),.A(g4765));
  NOT NOT1_2413(.VSS(VSS),.VDD(VDD),.Y(g4858),.A(I6582));
  NOT NOT1_2414(.VSS(VSS),.VDD(VDD),.Y(I6587),.A(g4803));
  NOT NOT1_2415(.VSS(VSS),.VDD(VDD),.Y(g4861),.A(I6587));
  NOT NOT1_2416(.VSS(VSS),.VDD(VDD),.Y(g4869),.A(g4662));
  NOT NOT1_2417(.VSS(VSS),.VDD(VDD),.Y(I6599),.A(g4823));
  NOT NOT1_2418(.VSS(VSS),.VDD(VDD),.Y(g4871),.A(I6599));
  NOT NOT1_2419(.VSS(VSS),.VDD(VDD),.Y(g4894),.A(g4813));
  NOT NOT1_2420(.VSS(VSS),.VDD(VDD),.Y(I6607),.A(g4745));
  NOT NOT1_2421(.VSS(VSS),.VDD(VDD),.Y(g4900),.A(I6607));
  NOT NOT1_2422(.VSS(VSS),.VDD(VDD),.Y(g4904),.A(g4812));
  NOT NOT1_2423(.VSS(VSS),.VDD(VDD),.Y(I6612),.A(g4660));
  NOT NOT1_2424(.VSS(VSS),.VDD(VDD),.Y(g4910),.A(I6612));
  NOT NOT1_2425(.VSS(VSS),.VDD(VDD),.Y(I6615),.A(g4745));
  NOT NOT1_2426(.VSS(VSS),.VDD(VDD),.Y(g4911),.A(I6615));
  NOT NOT1_2427(.VSS(VSS),.VDD(VDD),.Y(g4914),.A(g4816));
  NOT NOT1_2428(.VSS(VSS),.VDD(VDD),.Y(g4915),.A(g4669));
  NOT NOT1_2429(.VSS(VSS),.VDD(VDD),.Y(I6621),.A(g4745));
  NOT NOT1_2430(.VSS(VSS),.VDD(VDD),.Y(g4929),.A(I6621));
  NOT NOT1_2431(.VSS(VSS),.VDD(VDD),.Y(I6625),.A(g4745));
  NOT NOT1_2432(.VSS(VSS),.VDD(VDD),.Y(g4933),.A(I6625));
  NOT NOT1_2433(.VSS(VSS),.VDD(VDD),.Y(I6630),.A(g4745));
  NOT NOT1_2434(.VSS(VSS),.VDD(VDD),.Y(g4938),.A(I6630));
  NOT NOT1_2435(.VSS(VSS),.VDD(VDD),.Y(I6635),.A(g4745));
  NOT NOT1_2436(.VSS(VSS),.VDD(VDD),.Y(g4943),.A(I6635));
  NOT NOT1_2437(.VSS(VSS),.VDD(VDD),.Y(g4980),.A(g4678));
  NOT NOT1_2438(.VSS(VSS),.VDD(VDD),.Y(I6646),.A(g4687));
  NOT NOT1_2439(.VSS(VSS),.VDD(VDD),.Y(g5010),.A(I6646));
  NOT NOT1_2440(.VSS(VSS),.VDD(VDD),.Y(I6649),.A(g4693));
  NOT NOT1_2441(.VSS(VSS),.VDD(VDD),.Y(g5011),.A(I6649));
  NOT NOT1_2442(.VSS(VSS),.VDD(VDD),.Y(I6666),.A(g4740));
  NOT NOT1_2443(.VSS(VSS),.VDD(VDD),.Y(g5022),.A(I6666));
  NOT NOT1_2444(.VSS(VSS),.VDD(VDD),.Y(g5025),.A(g4814));
  NOT NOT1_2445(.VSS(VSS),.VDD(VDD),.Y(I6672),.A(g4752));
  NOT NOT1_2446(.VSS(VSS),.VDD(VDD),.Y(g5042),.A(I6672));
  NOT NOT1_2447(.VSS(VSS),.VDD(VDD),.Y(I6677),.A(g4757));
  NOT NOT1_2448(.VSS(VSS),.VDD(VDD),.Y(g5045),.A(I6677));
  NOT NOT1_2449(.VSS(VSS),.VDD(VDD),.Y(I6680),.A(g4713));
  NOT NOT1_2450(.VSS(VSS),.VDD(VDD),.Y(g5046),.A(I6680));
  NOT NOT1_2451(.VSS(VSS),.VDD(VDD),.Y(I6685),.A(g4716));
  NOT NOT1_2452(.VSS(VSS),.VDD(VDD),.Y(g5049),.A(I6685));
  NOT NOT1_2453(.VSS(VSS),.VDD(VDD),.Y(I6689),.A(g4758));
  NOT NOT1_2454(.VSS(VSS),.VDD(VDD),.Y(g5051),.A(I6689));
  NOT NOT1_2455(.VSS(VSS),.VDD(VDD),.Y(I6692),.A(g4720));
  NOT NOT1_2456(.VSS(VSS),.VDD(VDD),.Y(g5052),.A(I6692));
  NOT NOT1_2457(.VSS(VSS),.VDD(VDD),.Y(g5054),.A(g4816));
  NOT NOT1_2458(.VSS(VSS),.VDD(VDD),.Y(I6697),.A(g4722));
  NOT NOT1_2459(.VSS(VSS),.VDD(VDD),.Y(g5059),.A(I6697));
  NOT NOT1_2460(.VSS(VSS),.VDD(VDD),.Y(I6701),.A(g4726));
  NOT NOT1_2461(.VSS(VSS),.VDD(VDD),.Y(g5061),.A(I6701));
  NOT NOT1_2462(.VSS(VSS),.VDD(VDD),.Y(g5063),.A(g4799));
  NOT NOT1_2463(.VSS(VSS),.VDD(VDD),.Y(I6706),.A(g4731));
  NOT NOT1_2464(.VSS(VSS),.VDD(VDD),.Y(g5064),.A(I6706));
  NOT NOT1_2465(.VSS(VSS),.VDD(VDD),.Y(g5067),.A(g4801));
  NOT NOT1_2466(.VSS(VSS),.VDD(VDD),.Y(g5082),.A(g4723));
  NOT NOT1_2467(.VSS(VSS),.VDD(VDD),.Y(g5084),.A(g4727));
  NOT NOT1_2468(.VSS(VSS),.VDD(VDD),.Y(g5086),.A(g4732));
  NOT NOT1_2469(.VSS(VSS),.VDD(VDD),.Y(g5087),.A(g4736));
  NOT NOT1_2470(.VSS(VSS),.VDD(VDD),.Y(I6723),.A(g4761));
  NOT NOT1_2471(.VSS(VSS),.VDD(VDD),.Y(g5089),.A(I6723));
  NOT NOT1_2472(.VSS(VSS),.VDD(VDD),.Y(g5090),.A(g4741));
  NOT NOT1_2473(.VSS(VSS),.VDD(VDD),.Y(g5092),.A(g4753));
  NOT NOT1_2474(.VSS(VSS),.VDD(VDD),.Y(I6733),.A(g4773));
  NOT NOT1_2475(.VSS(VSS),.VDD(VDD),.Y(g5097),.A(I6733));
  NOT NOT1_2476(.VSS(VSS),.VDD(VDD),.Y(I6737),.A(g4662));
  NOT NOT1_2477(.VSS(VSS),.VDD(VDD),.Y(g5099),.A(I6737));
  NOT NOT1_2478(.VSS(VSS),.VDD(VDD),.Y(I6740),.A(g4781));
  NOT NOT1_2479(.VSS(VSS),.VDD(VDD),.Y(g5110),.A(I6740));
  NOT NOT1_2480(.VSS(VSS),.VDD(VDD),.Y(I6750),.A(g4771));
  NOT NOT1_2481(.VSS(VSS),.VDD(VDD),.Y(g5112),.A(I6750));
  NOT NOT1_2482(.VSS(VSS),.VDD(VDD),.Y(I6753),.A(g4772));
  NOT NOT1_2483(.VSS(VSS),.VDD(VDD),.Y(g5113),.A(I6753));
  NOT NOT1_2484(.VSS(VSS),.VDD(VDD),.Y(I6756),.A(g4775));
  NOT NOT1_2485(.VSS(VSS),.VDD(VDD),.Y(g5114),.A(I6756));
  NOT NOT1_2486(.VSS(VSS),.VDD(VDD),.Y(I6759),.A(g4778));
  NOT NOT1_2487(.VSS(VSS),.VDD(VDD),.Y(g5115),.A(I6759));
  NOT NOT1_2488(.VSS(VSS),.VDD(VDD),.Y(g5116),.A(g4810));
  NOT NOT1_2489(.VSS(VSS),.VDD(VDD),.Y(I6763),.A(g4780));
  NOT NOT1_2490(.VSS(VSS),.VDD(VDD),.Y(g5117),.A(I6763));
  NOT NOT1_2491(.VSS(VSS),.VDD(VDD),.Y(I6766),.A(g4783));
  NOT NOT1_2492(.VSS(VSS),.VDD(VDD),.Y(g5118),.A(I6766));
  NOT NOT1_2493(.VSS(VSS),.VDD(VDD),.Y(I6769),.A(g4786));
  NOT NOT1_2494(.VSS(VSS),.VDD(VDD),.Y(g5119),.A(I6769));
  NOT NOT1_2495(.VSS(VSS),.VDD(VDD),.Y(I6772),.A(g4788));
  NOT NOT1_2496(.VSS(VSS),.VDD(VDD),.Y(g5120),.A(I6772));
  NOT NOT1_2497(.VSS(VSS),.VDD(VDD),.Y(I6775),.A(g4790));
  NOT NOT1_2498(.VSS(VSS),.VDD(VDD),.Y(g5121),.A(I6775));
  NOT NOT1_2499(.VSS(VSS),.VDD(VDD),.Y(I6780),.A(g4825));
  NOT NOT1_2500(.VSS(VSS),.VDD(VDD),.Y(g5124),.A(I6780));
  NOT NOT1_2501(.VSS(VSS),.VDD(VDD),.Y(I6783),.A(g4822));
  NOT NOT1_2502(.VSS(VSS),.VDD(VDD),.Y(g5135),.A(I6783));
  NOT NOT1_2503(.VSS(VSS),.VDD(VDD),.Y(I6786),.A(g4824));
  NOT NOT1_2504(.VSS(VSS),.VDD(VDD),.Y(g5136),.A(I6786));
  NOT NOT1_2505(.VSS(VSS),.VDD(VDD),.Y(I6789),.A(g4871));
  NOT NOT1_2506(.VSS(VSS),.VDD(VDD),.Y(g5137),.A(I6789));
  NOT NOT1_2507(.VSS(VSS),.VDD(VDD),.Y(I6792),.A(g5097));
  NOT NOT1_2508(.VSS(VSS),.VDD(VDD),.Y(g5138),.A(I6792));
  NOT NOT1_2509(.VSS(VSS),.VDD(VDD),.Y(I6795),.A(g5022));
  NOT NOT1_2510(.VSS(VSS),.VDD(VDD),.Y(g5139),.A(I6795));
  NOT NOT1_2511(.VSS(VSS),.VDD(VDD),.Y(I6798),.A(g5042));
  NOT NOT1_2512(.VSS(VSS),.VDD(VDD),.Y(g5140),.A(I6798));
  NOT NOT1_2513(.VSS(VSS),.VDD(VDD),.Y(I6801),.A(g5045));
  NOT NOT1_2514(.VSS(VSS),.VDD(VDD),.Y(g5141),.A(I6801));
  NOT NOT1_2515(.VSS(VSS),.VDD(VDD),.Y(I6809),.A(g5051));
  NOT NOT1_2516(.VSS(VSS),.VDD(VDD),.Y(g5147),.A(I6809));
  NOT NOT1_2517(.VSS(VSS),.VDD(VDD),.Y(I6812),.A(g5110));
  NOT NOT1_2518(.VSS(VSS),.VDD(VDD),.Y(g5148),.A(I6812));
  NOT NOT1_2519(.VSS(VSS),.VDD(VDD),.Y(I6816),.A(g5111));
  NOT NOT1_2520(.VSS(VSS),.VDD(VDD),.Y(g5150),.A(I6816));
  NOT NOT1_2521(.VSS(VSS),.VDD(VDD),.Y(I6819),.A(g5019));
  NOT NOT1_2522(.VSS(VSS),.VDD(VDD),.Y(g5151),.A(I6819));
  NOT NOT1_2523(.VSS(VSS),.VDD(VDD),.Y(g5155),.A(g5099));
  NOT NOT1_2524(.VSS(VSS),.VDD(VDD),.Y(g5160),.A(g5099));
  NOT NOT1_2525(.VSS(VSS),.VDD(VDD),.Y(g5168),.A(g5099));
  NOT NOT1_2526(.VSS(VSS),.VDD(VDD),.Y(g5174),.A(g5099));
  NOT NOT1_2527(.VSS(VSS),.VDD(VDD),.Y(g5179),.A(g5099));
  NOT NOT1_2528(.VSS(VSS),.VDD(VDD),.Y(I6867),.A(g5082));
  NOT NOT1_2529(.VSS(VSS),.VDD(VDD),.Y(g5199),.A(I6867));
  NOT NOT1_2530(.VSS(VSS),.VDD(VDD),.Y(I6874),.A(g4861));
  NOT NOT1_2531(.VSS(VSS),.VDD(VDD),.Y(g5210),.A(I6874));
  NOT NOT1_2532(.VSS(VSS),.VDD(VDD),.Y(I6885),.A(g4872));
  NOT NOT1_2533(.VSS(VSS),.VDD(VDD),.Y(g5219),.A(I6885));
  NOT NOT1_2534(.VSS(VSS),.VDD(VDD),.Y(g5220),.A(g4903));
  NOT NOT1_2535(.VSS(VSS),.VDD(VDD),.Y(I6895),.A(g5010));
  NOT NOT1_2536(.VSS(VSS),.VDD(VDD),.Y(g5230),.A(I6895));
  NOT NOT1_2537(.VSS(VSS),.VDD(VDD),.Y(g5237),.A(g5083));
  NOT NOT1_2538(.VSS(VSS),.VDD(VDD),.Y(g5242),.A(g5085));
  NOT NOT1_2539(.VSS(VSS),.VDD(VDD),.Y(g5247),.A(g4900));
  NOT NOT1_2540(.VSS(VSS),.VDD(VDD),.Y(g5248),.A(g4911));
  NOT NOT1_2541(.VSS(VSS),.VDD(VDD),.Y(g5250),.A(g4929));
  NOT NOT1_2542(.VSS(VSS),.VDD(VDD),.Y(g5251),.A(g5069));
  NOT NOT1_2543(.VSS(VSS),.VDD(VDD),.Y(g5255),.A(g4933));
  NOT NOT1_2544(.VSS(VSS),.VDD(VDD),.Y(g5256),.A(g5077));
  NOT NOT1_2545(.VSS(VSS),.VDD(VDD),.Y(g5260),.A(g4938));
  NOT NOT1_2546(.VSS(VSS),.VDD(VDD),.Y(I6918),.A(g5124));
  NOT NOT1_2547(.VSS(VSS),.VDD(VDD),.Y(g5261),.A(I6918));
  NOT NOT1_2548(.VSS(VSS),.VDD(VDD),.Y(g5264),.A(g4943));
  NOT NOT1_2549(.VSS(VSS),.VDD(VDD),.Y(I6923),.A(g5124));
  NOT NOT1_2550(.VSS(VSS),.VDD(VDD),.Y(g5266),.A(I6923));
  NOT NOT1_2551(.VSS(VSS),.VDD(VDD),.Y(I6927),.A(g5124));
  NOT NOT1_2552(.VSS(VSS),.VDD(VDD),.Y(g5270),.A(I6927));
  NOT NOT1_2553(.VSS(VSS),.VDD(VDD),.Y(I6930),.A(g5017));
  NOT NOT1_2554(.VSS(VSS),.VDD(VDD),.Y(g5273),.A(I6930));
  NOT NOT1_2555(.VSS(VSS),.VDD(VDD),.Y(I6933),.A(g5124));
  NOT NOT1_2556(.VSS(VSS),.VDD(VDD),.Y(g5274),.A(I6933));
  NOT NOT1_2557(.VSS(VSS),.VDD(VDD),.Y(I6937),.A(g5124));
  NOT NOT1_2558(.VSS(VSS),.VDD(VDD),.Y(g5278),.A(I6937));
  NOT NOT1_2559(.VSS(VSS),.VDD(VDD),.Y(I6942),.A(g5124));
  NOT NOT1_2560(.VSS(VSS),.VDD(VDD),.Y(g5292),.A(I6942));
  NOT NOT1_2561(.VSS(VSS),.VDD(VDD),.Y(I6946),.A(g5124));
  NOT NOT1_2562(.VSS(VSS),.VDD(VDD),.Y(g5296),.A(I6946));
  NOT NOT1_2563(.VSS(VSS),.VDD(VDD),.Y(I6949),.A(g5050));
  NOT NOT1_2564(.VSS(VSS),.VDD(VDD),.Y(g5299),.A(I6949));
  NOT NOT1_2565(.VSS(VSS),.VDD(VDD),.Y(I6952),.A(g5124));
  NOT NOT1_2566(.VSS(VSS),.VDD(VDD),.Y(g5300),.A(I6952));
  NOT NOT1_2567(.VSS(VSS),.VDD(VDD),.Y(I6956),.A(g5124));
  NOT NOT1_2568(.VSS(VSS),.VDD(VDD),.Y(g5304),.A(I6956));
  NOT NOT1_2569(.VSS(VSS),.VDD(VDD),.Y(I6959),.A(g5089));
  NOT NOT1_2570(.VSS(VSS),.VDD(VDD),.Y(g5307),.A(I6959));
  NOT NOT1_2571(.VSS(VSS),.VDD(VDD),.Y(g5309),.A(g5063));
  NOT NOT1_2572(.VSS(VSS),.VDD(VDD),.Y(g5310),.A(g5067));
  NOT NOT1_2573(.VSS(VSS),.VDD(VDD),.Y(I6972),.A(g5135));
  NOT NOT1_2574(.VSS(VSS),.VDD(VDD),.Y(g5314),.A(I6972));
  NOT NOT1_2575(.VSS(VSS),.VDD(VDD),.Y(g5315),.A(g5116));
  NOT NOT1_2576(.VSS(VSS),.VDD(VDD),.Y(I6976),.A(g5136));
  NOT NOT1_2577(.VSS(VSS),.VDD(VDD),.Y(g5316),.A(I6976));
  NOT NOT1_2578(.VSS(VSS),.VDD(VDD),.Y(I6986),.A(g5230));
  NOT NOT1_2579(.VSS(VSS),.VDD(VDD),.Y(g5328),.A(I6986));
  NOT NOT1_2580(.VSS(VSS),.VDD(VDD),.Y(I6989),.A(g5307));
  NOT NOT1_2581(.VSS(VSS),.VDD(VDD),.Y(g5329),.A(I6989));
  NOT NOT1_2582(.VSS(VSS),.VDD(VDD),.Y(I6992),.A(g5151));
  NOT NOT1_2583(.VSS(VSS),.VDD(VDD),.Y(g5330),.A(I6992));
  NOT NOT1_2584(.VSS(VSS),.VDD(VDD),.Y(I6995),.A(g5220));
  NOT NOT1_2585(.VSS(VSS),.VDD(VDD),.Y(g5331),.A(I6995));
  NOT NOT1_2586(.VSS(VSS),.VDD(VDD),.Y(I7002),.A(g5308));
  NOT NOT1_2587(.VSS(VSS),.VDD(VDD),.Y(g5352),.A(I7002));
  NOT NOT1_2588(.VSS(VSS),.VDD(VDD),.Y(I7007),.A(g5314));
  NOT NOT1_2589(.VSS(VSS),.VDD(VDD),.Y(g5355),.A(I7007));
  NOT NOT1_2590(.VSS(VSS),.VDD(VDD),.Y(I7012),.A(g5316));
  NOT NOT1_2591(.VSS(VSS),.VDD(VDD),.Y(g5358),.A(I7012));
  NOT NOT1_2592(.VSS(VSS),.VDD(VDD),.Y(I7029),.A(g5149));
  NOT NOT1_2593(.VSS(VSS),.VDD(VDD),.Y(g5375),.A(I7029));
  NOT NOT1_2594(.VSS(VSS),.VDD(VDD),.Y(I7035),.A(g5150));
  NOT NOT1_2595(.VSS(VSS),.VDD(VDD),.Y(g5379),.A(I7035));
  NOT NOT1_2596(.VSS(VSS),.VDD(VDD),.Y(I7039),.A(g5309));
  NOT NOT1_2597(.VSS(VSS),.VDD(VDD),.Y(g5381),.A(I7039));
  NOT NOT1_2598(.VSS(VSS),.VDD(VDD),.Y(I7042),.A(g5310));
  NOT NOT1_2599(.VSS(VSS),.VDD(VDD),.Y(g5382),.A(I7042));
  NOT NOT1_2600(.VSS(VSS),.VDD(VDD),.Y(I7045),.A(g5167));
  NOT NOT1_2601(.VSS(VSS),.VDD(VDD),.Y(g5383),.A(I7045));
  NOT NOT1_2602(.VSS(VSS),.VDD(VDD),.Y(g5384),.A(g5220));
  NOT NOT1_2603(.VSS(VSS),.VDD(VDD),.Y(I7051),.A(g5219));
  NOT NOT1_2604(.VSS(VSS),.VDD(VDD),.Y(g5387),.A(I7051));
  NOT NOT1_2605(.VSS(VSS),.VDD(VDD),.Y(I7055),.A(g5318));
  NOT NOT1_2606(.VSS(VSS),.VDD(VDD),.Y(g5391),.A(I7055));
  NOT NOT1_2607(.VSS(VSS),.VDD(VDD),.Y(I7058),.A(g5281));
  NOT NOT1_2608(.VSS(VSS),.VDD(VDD),.Y(g5392),.A(I7058));
  NOT NOT1_2609(.VSS(VSS),.VDD(VDD),.Y(I7061),.A(g5281));
  NOT NOT1_2610(.VSS(VSS),.VDD(VDD),.Y(g5395),.A(I7061));
  NOT NOT1_2611(.VSS(VSS),.VDD(VDD),.Y(I7065),.A(g5281));
  NOT NOT1_2612(.VSS(VSS),.VDD(VDD),.Y(g5399),.A(I7065));
  NOT NOT1_2613(.VSS(VSS),.VDD(VDD),.Y(I7069),.A(g5281));
  NOT NOT1_2614(.VSS(VSS),.VDD(VDD),.Y(g5403),.A(I7069));
  NOT NOT1_2615(.VSS(VSS),.VDD(VDD),.Y(I7073),.A(g5281));
  NOT NOT1_2616(.VSS(VSS),.VDD(VDD),.Y(g5407),.A(I7073));
  NOT NOT1_2617(.VSS(VSS),.VDD(VDD),.Y(I7077),.A(g5281));
  NOT NOT1_2618(.VSS(VSS),.VDD(VDD),.Y(g5411),.A(I7077));
  NOT NOT1_2619(.VSS(VSS),.VDD(VDD),.Y(I7081),.A(g5281));
  NOT NOT1_2620(.VSS(VSS),.VDD(VDD),.Y(g5415),.A(I7081));
  NOT NOT1_2621(.VSS(VSS),.VDD(VDD),.Y(I7086),.A(g5281));
  NOT NOT1_2622(.VSS(VSS),.VDD(VDD),.Y(g5420),.A(I7086));
  NOT NOT1_2623(.VSS(VSS),.VDD(VDD),.Y(I7091),.A(g5281));
  NOT NOT1_2624(.VSS(VSS),.VDD(VDD),.Y(g5425),.A(I7091));
  NOT NOT1_2625(.VSS(VSS),.VDD(VDD),.Y(I7104),.A(g5273));
  NOT NOT1_2626(.VSS(VSS),.VDD(VDD),.Y(g5432),.A(I7104));
  NOT NOT1_2627(.VSS(VSS),.VDD(VDD),.Y(I7107),.A(g5277));
  NOT NOT1_2628(.VSS(VSS),.VDD(VDD),.Y(g5433),.A(I7107));
  NOT NOT1_2629(.VSS(VSS),.VDD(VDD),.Y(I7110),.A(g5291));
  NOT NOT1_2630(.VSS(VSS),.VDD(VDD),.Y(g5434),.A(I7110));
  NOT NOT1_2631(.VSS(VSS),.VDD(VDD),.Y(I7113),.A(g5295));
  NOT NOT1_2632(.VSS(VSS),.VDD(VDD),.Y(g5435),.A(I7113));
  NOT NOT1_2633(.VSS(VSS),.VDD(VDD),.Y(I7116),.A(g5299));
  NOT NOT1_2634(.VSS(VSS),.VDD(VDD),.Y(g5436),.A(I7116));
  NOT NOT1_2635(.VSS(VSS),.VDD(VDD),.Y(I7119),.A(g5303));
  NOT NOT1_2636(.VSS(VSS),.VDD(VDD),.Y(g5437),.A(I7119));
  NOT NOT1_2637(.VSS(VSS),.VDD(VDD),.Y(g5439),.A(g5261));
  NOT NOT1_2638(.VSS(VSS),.VDD(VDD),.Y(g5440),.A(g5266));
  NOT NOT1_2639(.VSS(VSS),.VDD(VDD),.Y(g5442),.A(g5270));
  NOT NOT1_2640(.VSS(VSS),.VDD(VDD),.Y(g5445),.A(g5274));
  NOT NOT1_2641(.VSS(VSS),.VDD(VDD),.Y(g5448),.A(g5278));
  NOT NOT1_2642(.VSS(VSS),.VDD(VDD),.Y(g5450),.A(g5292));
  NOT NOT1_2643(.VSS(VSS),.VDD(VDD),.Y(g5453),.A(g5296));
  NOT NOT1_2644(.VSS(VSS),.VDD(VDD),.Y(g5456),.A(g5300));
  NOT NOT1_2645(.VSS(VSS),.VDD(VDD),.Y(g5457),.A(g5304));
  NOT NOT1_2646(.VSS(VSS),.VDD(VDD),.Y(I7143),.A(g5323));
  NOT NOT1_2647(.VSS(VSS),.VDD(VDD),.Y(g5465),.A(I7143));
  NOT NOT1_2648(.VSS(VSS),.VDD(VDD),.Y(I7146),.A(g5231));
  NOT NOT1_2649(.VSS(VSS),.VDD(VDD),.Y(g5466),.A(I7146));
  NOT NOT1_2650(.VSS(VSS),.VDD(VDD),.Y(I7150),.A(g5355));
  NOT NOT1_2651(.VSS(VSS),.VDD(VDD),.Y(g5468),.A(I7150));
  NOT NOT1_2652(.VSS(VSS),.VDD(VDD),.Y(I7153),.A(g5358));
  NOT NOT1_2653(.VSS(VSS),.VDD(VDD),.Y(g5469),.A(I7153));
  NOT NOT1_2654(.VSS(VSS),.VDD(VDD),.Y(I7161),.A(g5465));
  NOT NOT1_2655(.VSS(VSS),.VDD(VDD),.Y(g5475),.A(I7161));
  NOT NOT1_2656(.VSS(VSS),.VDD(VDD),.Y(I7164),.A(g5433));
  NOT NOT1_2657(.VSS(VSS),.VDD(VDD),.Y(g5476),.A(I7164));
  NOT NOT1_2658(.VSS(VSS),.VDD(VDD),.Y(I7167),.A(g5434));
  NOT NOT1_2659(.VSS(VSS),.VDD(VDD),.Y(g5477),.A(I7167));
  NOT NOT1_2660(.VSS(VSS),.VDD(VDD),.Y(I7170),.A(g5435));
  NOT NOT1_2661(.VSS(VSS),.VDD(VDD),.Y(g5478),.A(I7170));
  NOT NOT1_2662(.VSS(VSS),.VDD(VDD),.Y(I7173),.A(g5436));
  NOT NOT1_2663(.VSS(VSS),.VDD(VDD),.Y(g5479),.A(I7173));
  NOT NOT1_2664(.VSS(VSS),.VDD(VDD),.Y(I7176),.A(g5437));
  NOT NOT1_2665(.VSS(VSS),.VDD(VDD),.Y(g5480),.A(I7176));
  NOT NOT1_2666(.VSS(VSS),.VDD(VDD),.Y(I7187),.A(g5387));
  NOT NOT1_2667(.VSS(VSS),.VDD(VDD),.Y(g5489),.A(I7187));
  NOT NOT1_2668(.VSS(VSS),.VDD(VDD),.Y(I7190),.A(g5432));
  NOT NOT1_2669(.VSS(VSS),.VDD(VDD),.Y(g5490),.A(I7190));
  NOT NOT1_2670(.VSS(VSS),.VDD(VDD),.Y(I7193),.A(g5466));
  NOT NOT1_2671(.VSS(VSS),.VDD(VDD),.Y(g5491),.A(I7193));
  NOT NOT1_2672(.VSS(VSS),.VDD(VDD),.Y(I7197),.A(g5431));
  NOT NOT1_2673(.VSS(VSS),.VDD(VDD),.Y(g5493),.A(I7197));
  NOT NOT1_2674(.VSS(VSS),.VDD(VDD),.Y(I7251),.A(g5458));
  NOT NOT1_2675(.VSS(VSS),.VDD(VDD),.Y(g5509),.A(I7251));
  NOT NOT1_2676(.VSS(VSS),.VDD(VDD),.Y(I7254),.A(g5458));
  NOT NOT1_2677(.VSS(VSS),.VDD(VDD),.Y(g5512),.A(I7254));
  NOT NOT1_2678(.VSS(VSS),.VDD(VDD),.Y(I7258),.A(g5458));
  NOT NOT1_2679(.VSS(VSS),.VDD(VDD),.Y(g5518),.A(I7258));
  NOT NOT1_2680(.VSS(VSS),.VDD(VDD),.Y(I7261),.A(g5458));
  NOT NOT1_2681(.VSS(VSS),.VDD(VDD),.Y(g5521),.A(I7261));
  NOT NOT1_2682(.VSS(VSS),.VDD(VDD),.Y(I7264),.A(g5458));
  NOT NOT1_2683(.VSS(VSS),.VDD(VDD),.Y(g5524),.A(I7264));
  NOT NOT1_2684(.VSS(VSS),.VDD(VDD),.Y(I7267),.A(g5458));
  NOT NOT1_2685(.VSS(VSS),.VDD(VDD),.Y(g5527),.A(I7267));
  NOT NOT1_2686(.VSS(VSS),.VDD(VDD),.Y(I7270),.A(g5352));
  NOT NOT1_2687(.VSS(VSS),.VDD(VDD),.Y(g5530),.A(I7270));
  NOT NOT1_2688(.VSS(VSS),.VDD(VDD),.Y(I7276),.A(g5375));
  NOT NOT1_2689(.VSS(VSS),.VDD(VDD),.Y(g5534),.A(I7276));
  NOT NOT1_2690(.VSS(VSS),.VDD(VDD),.Y(g5536),.A(g5467));
  NOT NOT1_2691(.VSS(VSS),.VDD(VDD),.Y(g5537),.A(g5385));
  NOT NOT1_2692(.VSS(VSS),.VDD(VDD),.Y(g5538),.A(g5331));
  NOT NOT1_2693(.VSS(VSS),.VDD(VDD),.Y(g5539),.A(g5331));
  NOT NOT1_2694(.VSS(VSS),.VDD(VDD),.Y(I7284),.A(g5383));
  NOT NOT1_2695(.VSS(VSS),.VDD(VDD),.Y(g5540),.A(I7284));
  NOT NOT1_2696(.VSS(VSS),.VDD(VDD),.Y(g5542),.A(g5331));
  NOT NOT1_2697(.VSS(VSS),.VDD(VDD),.Y(g5543),.A(g5331));
  NOT NOT1_2698(.VSS(VSS),.VDD(VDD),.Y(g5544),.A(g5331));
  NOT NOT1_2699(.VSS(VSS),.VDD(VDD),.Y(g5545),.A(g5331));
  NOT NOT1_2700(.VSS(VSS),.VDD(VDD),.Y(g5546),.A(g5388));
  NOT NOT1_2701(.VSS(VSS),.VDD(VDD),.Y(g5549),.A(g5331));
  NOT NOT1_2702(.VSS(VSS),.VDD(VDD),.Y(g5550),.A(g5331));
  NOT NOT1_2703(.VSS(VSS),.VDD(VDD),.Y(I7295),.A(g5439));
  NOT NOT1_2704(.VSS(VSS),.VDD(VDD),.Y(g5551),.A(I7295));
  NOT NOT1_2705(.VSS(VSS),.VDD(VDD),.Y(g5554),.A(g5455));
  NOT NOT1_2706(.VSS(VSS),.VDD(VDD),.Y(g5563),.A(g5381));
  NOT NOT1_2707(.VSS(VSS),.VDD(VDD),.Y(g5564),.A(g5382));
  NOT NOT1_2708(.VSS(VSS),.VDD(VDD),.Y(I7318),.A(g5452));
  NOT NOT1_2709(.VSS(VSS),.VDD(VDD),.Y(g5566),.A(I7318));
  NOT NOT1_2710(.VSS(VSS),.VDD(VDD),.Y(g5567),.A(g5418));
  NOT NOT1_2711(.VSS(VSS),.VDD(VDD),.Y(g5568),.A(g5423));
  NOT NOT1_2712(.VSS(VSS),.VDD(VDD),.Y(g5570),.A(g5392));
  NOT NOT1_2713(.VSS(VSS),.VDD(VDD),.Y(g5571),.A(g5395));
  NOT NOT1_2714(.VSS(VSS),.VDD(VDD),.Y(g5572),.A(g5399));
  NOT NOT1_2715(.VSS(VSS),.VDD(VDD),.Y(g5573),.A(g5403));
  NOT NOT1_2716(.VSS(VSS),.VDD(VDD),.Y(g5574),.A(g5407));
  NOT NOT1_2717(.VSS(VSS),.VDD(VDD),.Y(g5575),.A(g5411));
  NOT NOT1_2718(.VSS(VSS),.VDD(VDD),.Y(g5576),.A(g5415));
  NOT NOT1_2719(.VSS(VSS),.VDD(VDD),.Y(g5577),.A(g5420));
  NOT NOT1_2720(.VSS(VSS),.VDD(VDD),.Y(g5578),.A(g5425));
  NOT NOT1_2721(.VSS(VSS),.VDD(VDD),.Y(I7333),.A(g5386));
  NOT NOT1_2722(.VSS(VSS),.VDD(VDD),.Y(g5579),.A(I7333));
  NOT NOT1_2723(.VSS(VSS),.VDD(VDD),.Y(I7336),.A(g5534));
  NOT NOT1_2724(.VSS(VSS),.VDD(VDD),.Y(g5580),.A(I7336));
  NOT NOT1_2725(.VSS(VSS),.VDD(VDD),.Y(I7339),.A(g5540));
  NOT NOT1_2726(.VSS(VSS),.VDD(VDD),.Y(g5581),.A(I7339));
  NOT NOT1_2727(.VSS(VSS),.VDD(VDD),.Y(I7342),.A(g5579));
  NOT NOT1_2728(.VSS(VSS),.VDD(VDD),.Y(g5582),.A(I7342));
  NOT NOT1_2729(.VSS(VSS),.VDD(VDD),.Y(I7346),.A(g5531));
  NOT NOT1_2730(.VSS(VSS),.VDD(VDD),.Y(g5584),.A(I7346));
  NOT NOT1_2731(.VSS(VSS),.VDD(VDD),.Y(I7349),.A(g5532));
  NOT NOT1_2732(.VSS(VSS),.VDD(VDD),.Y(g5587),.A(I7349));
  NOT NOT1_2733(.VSS(VSS),.VDD(VDD),.Y(I7352),.A(g5533));
  NOT NOT1_2734(.VSS(VSS),.VDD(VDD),.Y(g5590),.A(I7352));
  NOT NOT1_2735(.VSS(VSS),.VDD(VDD),.Y(I7355),.A(g5535));
  NOT NOT1_2736(.VSS(VSS),.VDD(VDD),.Y(g5593),.A(I7355));
  NOT NOT1_2737(.VSS(VSS),.VDD(VDD),.Y(I7358),.A(g5565));
  NOT NOT1_2738(.VSS(VSS),.VDD(VDD),.Y(g5596),.A(I7358));
  NOT NOT1_2739(.VSS(VSS),.VDD(VDD),.Y(I7361),.A(g5566));
  NOT NOT1_2740(.VSS(VSS),.VDD(VDD),.Y(g5597),.A(I7361));
  NOT NOT1_2741(.VSS(VSS),.VDD(VDD),.Y(I7372),.A(g5493));
  NOT NOT1_2742(.VSS(VSS),.VDD(VDD),.Y(g5615),.A(I7372));
  NOT NOT1_2743(.VSS(VSS),.VDD(VDD),.Y(g5631),.A(g5536));
  NOT NOT1_2744(.VSS(VSS),.VDD(VDD),.Y(I7397),.A(g5561));
  NOT NOT1_2745(.VSS(VSS),.VDD(VDD),.Y(g5638),.A(I7397));
  NOT NOT1_2746(.VSS(VSS),.VDD(VDD),.Y(g5645),.A(g5537));
  NOT NOT1_2747(.VSS(VSS),.VDD(VDD),.Y(g5647),.A(g5509));
  NOT NOT1_2748(.VSS(VSS),.VDD(VDD),.Y(I7404),.A(g5541));
  NOT NOT1_2749(.VSS(VSS),.VDD(VDD),.Y(g5649),.A(I7404));
  NOT NOT1_2750(.VSS(VSS),.VDD(VDD),.Y(g5658),.A(g5512));
  NOT NOT1_2751(.VSS(VSS),.VDD(VDD),.Y(g5661),.A(g5518));
  NOT NOT1_2752(.VSS(VSS),.VDD(VDD),.Y(g5664),.A(g5521));
  NOT NOT1_2753(.VSS(VSS),.VDD(VDD),.Y(g5667),.A(g5524));
  NOT NOT1_2754(.VSS(VSS),.VDD(VDD),.Y(g5670),.A(g5527));
  NOT NOT1_2755(.VSS(VSS),.VDD(VDD),.Y(g5685),.A(g5552));
  NOT NOT1_2756(.VSS(VSS),.VDD(VDD),.Y(g5687),.A(g5567));
  NOT NOT1_2757(.VSS(VSS),.VDD(VDD),.Y(g5691),.A(g5568));
  NOT NOT1_2758(.VSS(VSS),.VDD(VDD),.Y(I7451),.A(g5597));
  NOT NOT1_2759(.VSS(VSS),.VDD(VDD),.Y(g5692),.A(I7451));
  NOT NOT1_2760(.VSS(VSS),.VDD(VDD),.Y(I7463),.A(g5622));
  NOT NOT1_2761(.VSS(VSS),.VDD(VDD),.Y(g5702),.A(I7463));
  NOT NOT1_2762(.VSS(VSS),.VDD(VDD),.Y(I7466),.A(g5624));
  NOT NOT1_2763(.VSS(VSS),.VDD(VDD),.Y(g5705),.A(I7466));
  NOT NOT1_2764(.VSS(VSS),.VDD(VDD),.Y(I7469),.A(g5625));
  NOT NOT1_2765(.VSS(VSS),.VDD(VDD),.Y(g5708),.A(I7469));
  NOT NOT1_2766(.VSS(VSS),.VDD(VDD),.Y(I7472),.A(g5626));
  NOT NOT1_2767(.VSS(VSS),.VDD(VDD),.Y(g5711),.A(I7472));
  NOT NOT1_2768(.VSS(VSS),.VDD(VDD),.Y(I7475),.A(g5627));
  NOT NOT1_2769(.VSS(VSS),.VDD(VDD),.Y(g5714),.A(I7475));
  NOT NOT1_2770(.VSS(VSS),.VDD(VDD),.Y(I7478),.A(g5628));
  NOT NOT1_2771(.VSS(VSS),.VDD(VDD),.Y(g5717),.A(I7478));
  NOT NOT1_2772(.VSS(VSS),.VDD(VDD),.Y(I7481),.A(g5629));
  NOT NOT1_2773(.VSS(VSS),.VDD(VDD),.Y(g5720),.A(I7481));
  NOT NOT1_2774(.VSS(VSS),.VDD(VDD),.Y(I7484),.A(g5630));
  NOT NOT1_2775(.VSS(VSS),.VDD(VDD),.Y(g5723),.A(I7484));
  NOT NOT1_2776(.VSS(VSS),.VDD(VDD),.Y(I7487),.A(g5684));
  NOT NOT1_2777(.VSS(VSS),.VDD(VDD),.Y(g5726),.A(I7487));
  NOT NOT1_2778(.VSS(VSS),.VDD(VDD),.Y(I7490),.A(g5583));
  NOT NOT1_2779(.VSS(VSS),.VDD(VDD),.Y(g5727),.A(I7490));
  NOT NOT1_2780(.VSS(VSS),.VDD(VDD),.Y(I7494),.A(g5691));
  NOT NOT1_2781(.VSS(VSS),.VDD(VDD),.Y(g5729),.A(I7494));
  NOT NOT1_2782(.VSS(VSS),.VDD(VDD),.Y(I7497),.A(g5687));
  NOT NOT1_2783(.VSS(VSS),.VDD(VDD),.Y(g5730),.A(I7497));
  NOT NOT1_2784(.VSS(VSS),.VDD(VDD),.Y(I7501),.A(g5596));
  NOT NOT1_2785(.VSS(VSS),.VDD(VDD),.Y(g5740),.A(I7501));
  NOT NOT1_2786(.VSS(VSS),.VDD(VDD),.Y(g5741),.A(g5602));
  NOT NOT1_2787(.VSS(VSS),.VDD(VDD),.Y(g5742),.A(g5686));
  NOT NOT1_2788(.VSS(VSS),.VDD(VDD),.Y(I7506),.A(g5584));
  NOT NOT1_2789(.VSS(VSS),.VDD(VDD),.Y(g5751),.A(I7506));
  NOT NOT1_2790(.VSS(VSS),.VDD(VDD),.Y(I7509),.A(g5587));
  NOT NOT1_2791(.VSS(VSS),.VDD(VDD),.Y(g5752),.A(I7509));
  NOT NOT1_2792(.VSS(VSS),.VDD(VDD),.Y(g5770),.A(g5645));
  NOT NOT1_2793(.VSS(VSS),.VDD(VDD),.Y(I7514),.A(g5590));
  NOT NOT1_2794(.VSS(VSS),.VDD(VDD),.Y(g5773),.A(I7514));
  NOT NOT1_2795(.VSS(VSS),.VDD(VDD),.Y(I7517),.A(g5593));
  NOT NOT1_2796(.VSS(VSS),.VDD(VDD),.Y(g5774),.A(I7517));
  NOT NOT1_2797(.VSS(VSS),.VDD(VDD),.Y(I7583),.A(g5605));
  NOT NOT1_2798(.VSS(VSS),.VDD(VDD),.Y(g5784),.A(I7583));
  NOT NOT1_2799(.VSS(VSS),.VDD(VDD),.Y(g5787),.A(g5685));
  NOT NOT1_2800(.VSS(VSS),.VDD(VDD),.Y(I7587),.A(g5605));
  NOT NOT1_2801(.VSS(VSS),.VDD(VDD),.Y(g5788),.A(I7587));
  NOT NOT1_2802(.VSS(VSS),.VDD(VDD),.Y(I7590),.A(g5605));
  NOT NOT1_2803(.VSS(VSS),.VDD(VDD),.Y(g5791),.A(I7590));
  NOT NOT1_2804(.VSS(VSS),.VDD(VDD),.Y(I7593),.A(g5605));
  NOT NOT1_2805(.VSS(VSS),.VDD(VDD),.Y(g5794),.A(I7593));
  NOT NOT1_2806(.VSS(VSS),.VDD(VDD),.Y(I7596),.A(g5605));
  NOT NOT1_2807(.VSS(VSS),.VDD(VDD),.Y(g5797),.A(I7596));
  NOT NOT1_2808(.VSS(VSS),.VDD(VDD),.Y(I7600),.A(g5605));
  NOT NOT1_2809(.VSS(VSS),.VDD(VDD),.Y(g5801),.A(I7600));
  NOT NOT1_2810(.VSS(VSS),.VDD(VDD),.Y(I7604),.A(g5605));
  NOT NOT1_2811(.VSS(VSS),.VDD(VDD),.Y(g5805),.A(I7604));
  NOT NOT1_2812(.VSS(VSS),.VDD(VDD),.Y(I7608),.A(g5605));
  NOT NOT1_2813(.VSS(VSS),.VDD(VDD),.Y(g5809),.A(I7608));
  NOT NOT1_2814(.VSS(VSS),.VDD(VDD),.Y(I7612),.A(g5605));
  NOT NOT1_2815(.VSS(VSS),.VDD(VDD),.Y(g5813),.A(I7612));
  NOT NOT1_2816(.VSS(VSS),.VDD(VDD),.Y(g5824),.A(g5631));
  NOT NOT1_2817(.VSS(VSS),.VDD(VDD),.Y(g5860),.A(g5634));
  NOT NOT1_2818(.VSS(VSS),.VDD(VDD),.Y(g5861),.A(g5636));
  NOT NOT1_2819(.VSS(VSS),.VDD(VDD),.Y(I7634),.A(g5727));
  NOT NOT1_2820(.VSS(VSS),.VDD(VDD),.Y(g5874),.A(I7634));
  NOT NOT1_2821(.VSS(VSS),.VDD(VDD),.Y(I7637),.A(g5751));
  NOT NOT1_2822(.VSS(VSS),.VDD(VDD),.Y(g5875),.A(I7637));
  NOT NOT1_2823(.VSS(VSS),.VDD(VDD),.Y(I7640),.A(g5773));
  NOT NOT1_2824(.VSS(VSS),.VDD(VDD),.Y(g5876),.A(I7640));
  NOT NOT1_2825(.VSS(VSS),.VDD(VDD),.Y(I7643),.A(g5752));
  NOT NOT1_2826(.VSS(VSS),.VDD(VDD),.Y(g5877),.A(I7643));
  NOT NOT1_2827(.VSS(VSS),.VDD(VDD),.Y(I7646),.A(g5774));
  NOT NOT1_2828(.VSS(VSS),.VDD(VDD),.Y(g5878),.A(I7646));
  NOT NOT1_2829(.VSS(VSS),.VDD(VDD),.Y(g5879),.A(g5770));
  NOT NOT1_2830(.VSS(VSS),.VDD(VDD),.Y(g5880),.A(g5824));
  NOT NOT1_2831(.VSS(VSS),.VDD(VDD),.Y(g5884),.A(g5864));
  NOT NOT1_2832(.VSS(VSS),.VDD(VDD),.Y(g5885),.A(g5865));
  NOT NOT1_2833(.VSS(VSS),.VDD(VDD),.Y(g5886),.A(g5753));
  NOT NOT1_2834(.VSS(VSS),.VDD(VDD),.Y(g5887),.A(g5742));
  NOT NOT1_2835(.VSS(VSS),.VDD(VDD),.Y(g5888),.A(g5731));
  NOT NOT1_2836(.VSS(VSS),.VDD(VDD),.Y(g5889),.A(g5742));
  NOT NOT1_2837(.VSS(VSS),.VDD(VDD),.Y(g5890),.A(g5753));
  NOT NOT1_2838(.VSS(VSS),.VDD(VDD),.Y(g5891),.A(g5731));
  NOT NOT1_2839(.VSS(VSS),.VDD(VDD),.Y(g5892),.A(g5742));
  NOT NOT1_2840(.VSS(VSS),.VDD(VDD),.Y(g5893),.A(g5753));
  NOT NOT1_2841(.VSS(VSS),.VDD(VDD),.Y(g5894),.A(g5731));
  NOT NOT1_2842(.VSS(VSS),.VDD(VDD),.Y(g5895),.A(g5742));
  NOT NOT1_2843(.VSS(VSS),.VDD(VDD),.Y(g5896),.A(g5753));
  NOT NOT1_2844(.VSS(VSS),.VDD(VDD),.Y(g5897),.A(g5731));
  NOT NOT1_2845(.VSS(VSS),.VDD(VDD),.Y(g5899),.A(g5753));
  NOT NOT1_2846(.VSS(VSS),.VDD(VDD),.Y(g5901),.A(g5753));
  NOT NOT1_2847(.VSS(VSS),.VDD(VDD),.Y(g5903),.A(g5753));
  NOT NOT1_2848(.VSS(VSS),.VDD(VDD),.Y(g5905),.A(g5852));
  NOT NOT1_2849(.VSS(VSS),.VDD(VDD),.Y(g5908),.A(g5753));
  NOT NOT1_2850(.VSS(VSS),.VDD(VDD),.Y(g5912),.A(g5853));
  NOT NOT1_2851(.VSS(VSS),.VDD(VDD),.Y(I7679),.A(g5726));
  NOT NOT1_2852(.VSS(VSS),.VDD(VDD),.Y(g5915),.A(I7679));
  NOT NOT1_2853(.VSS(VSS),.VDD(VDD),.Y(I7683),.A(g5702));
  NOT NOT1_2854(.VSS(VSS),.VDD(VDD),.Y(g5917),.A(I7683));
  NOT NOT1_2855(.VSS(VSS),.VDD(VDD),.Y(I7686),.A(g5705));
  NOT NOT1_2856(.VSS(VSS),.VDD(VDD),.Y(g5918),.A(I7686));
  NOT NOT1_2857(.VSS(VSS),.VDD(VDD),.Y(I7689),.A(g5708));
  NOT NOT1_2858(.VSS(VSS),.VDD(VDD),.Y(g5919),.A(I7689));
  NOT NOT1_2859(.VSS(VSS),.VDD(VDD),.Y(I7692),.A(g5711));
  NOT NOT1_2860(.VSS(VSS),.VDD(VDD),.Y(g5920),.A(I7692));
  NOT NOT1_2861(.VSS(VSS),.VDD(VDD),.Y(I7695),.A(g5714));
  NOT NOT1_2862(.VSS(VSS),.VDD(VDD),.Y(g5921),.A(I7695));
  NOT NOT1_2863(.VSS(VSS),.VDD(VDD),.Y(I7698),.A(g5717));
  NOT NOT1_2864(.VSS(VSS),.VDD(VDD),.Y(g5922),.A(I7698));
  NOT NOT1_2865(.VSS(VSS),.VDD(VDD),.Y(I7701),.A(g5720));
  NOT NOT1_2866(.VSS(VSS),.VDD(VDD),.Y(g5923),.A(I7701));
  NOT NOT1_2867(.VSS(VSS),.VDD(VDD),.Y(I7704),.A(g5723));
  NOT NOT1_2868(.VSS(VSS),.VDD(VDD),.Y(g5924),.A(I7704));
  NOT NOT1_2869(.VSS(VSS),.VDD(VDD),.Y(I7707),.A(g5701));
  NOT NOT1_2870(.VSS(VSS),.VDD(VDD),.Y(g5925),.A(I7707));
  NOT NOT1_2871(.VSS(VSS),.VDD(VDD),.Y(g5946),.A(g5729));
  NOT NOT1_2872(.VSS(VSS),.VDD(VDD),.Y(g5950),.A(g5730));
  NOT NOT1_2873(.VSS(VSS),.VDD(VDD),.Y(g5957),.A(g5866));
  NOT NOT1_2874(.VSS(VSS),.VDD(VDD),.Y(g5958),.A(g5818));
  NOT NOT1_2875(.VSS(VSS),.VDD(VDD),.Y(g5975),.A(g5821));
  NOT NOT1_2876(.VSS(VSS),.VDD(VDD),.Y(g5992),.A(g5869));
  NOT NOT1_2877(.VSS(VSS),.VDD(VDD),.Y(g5993),.A(g5872));
  NOT NOT1_2878(.VSS(VSS),.VDD(VDD),.Y(g5994),.A(g5873));
  NOT NOT1_2879(.VSS(VSS),.VDD(VDD),.Y(g5995),.A(g5824));
  NOT NOT1_2880(.VSS(VSS),.VDD(VDD),.Y(g5996),.A(g5824));
  NOT NOT1_2881(.VSS(VSS),.VDD(VDD),.Y(g5997),.A(g5854));
  NOT NOT1_2882(.VSS(VSS),.VDD(VDD),.Y(g6014),.A(g5824));
  NOT NOT1_2883(.VSS(VSS),.VDD(VDD),.Y(g6015),.A(g5857));
  NOT NOT1_2884(.VSS(VSS),.VDD(VDD),.Y(g6032),.A(g5770));
  NOT NOT1_2885(.VSS(VSS),.VDD(VDD),.Y(g6033),.A(g5824));
  NOT NOT1_2886(.VSS(VSS),.VDD(VDD),.Y(g6034),.A(g5824));
  NOT NOT1_2887(.VSS(VSS),.VDD(VDD),.Y(g6035),.A(g5824));
  NOT NOT1_2888(.VSS(VSS),.VDD(VDD),.Y(g6036),.A(g5824));
  NOT NOT1_2889(.VSS(VSS),.VDD(VDD),.Y(g6039),.A(g5824));
  NOT NOT1_2890(.VSS(VSS),.VDD(VDD),.Y(g6040),.A(g5824));
  NOT NOT1_2891(.VSS(VSS),.VDD(VDD),.Y(g6043),.A(g5824));
  NOT NOT1_2892(.VSS(VSS),.VDD(VDD),.Y(g6044),.A(g5824));
  NOT NOT1_2893(.VSS(VSS),.VDD(VDD),.Y(g6048),.A(g5824));
  NOT NOT1_2894(.VSS(VSS),.VDD(VDD),.Y(g6051),.A(g5824));
  NOT NOT1_2895(.VSS(VSS),.VDD(VDD),.Y(g6052),.A(g5824));
  NOT NOT1_2896(.VSS(VSS),.VDD(VDD),.Y(g6057),.A(g5824));
  NOT NOT1_2897(.VSS(VSS),.VDD(VDD),.Y(g6062),.A(g5824));
  NOT NOT1_2898(.VSS(VSS),.VDD(VDD),.Y(g6065),.A(g5784));
  NOT NOT1_2899(.VSS(VSS),.VDD(VDD),.Y(g6067),.A(g5788));
  NOT NOT1_2900(.VSS(VSS),.VDD(VDD),.Y(g6069),.A(g5791));
  NOT NOT1_2901(.VSS(VSS),.VDD(VDD),.Y(g6070),.A(g5824));
  NOT NOT1_2902(.VSS(VSS),.VDD(VDD),.Y(g6074),.A(g5794));
  NOT NOT1_2903(.VSS(VSS),.VDD(VDD),.Y(g6076),.A(g5797));
  NOT NOT1_2904(.VSS(VSS),.VDD(VDD),.Y(g6078),.A(g5801));
  NOT NOT1_2905(.VSS(VSS),.VDD(VDD),.Y(g6080),.A(g5805));
  NOT NOT1_2906(.VSS(VSS),.VDD(VDD),.Y(g6083),.A(g5809));
  NOT NOT1_2907(.VSS(VSS),.VDD(VDD),.Y(g6087),.A(g5813));
  NOT NOT1_2908(.VSS(VSS),.VDD(VDD),.Y(I7796),.A(g5917));
  NOT NOT1_2909(.VSS(VSS),.VDD(VDD),.Y(g6100),.A(I7796));
  NOT NOT1_2910(.VSS(VSS),.VDD(VDD),.Y(I7799),.A(g5918));
  NOT NOT1_2911(.VSS(VSS),.VDD(VDD),.Y(g6101),.A(I7799));
  NOT NOT1_2912(.VSS(VSS),.VDD(VDD),.Y(I7802),.A(g5920));
  NOT NOT1_2913(.VSS(VSS),.VDD(VDD),.Y(g6102),.A(I7802));
  NOT NOT1_2914(.VSS(VSS),.VDD(VDD),.Y(I7805),.A(g5923));
  NOT NOT1_2915(.VSS(VSS),.VDD(VDD),.Y(g6103),.A(I7805));
  NOT NOT1_2916(.VSS(VSS),.VDD(VDD),.Y(I7808),.A(g5919));
  NOT NOT1_2917(.VSS(VSS),.VDD(VDD),.Y(g6104),.A(I7808));
  NOT NOT1_2918(.VSS(VSS),.VDD(VDD),.Y(I7811),.A(g5921));
  NOT NOT1_2919(.VSS(VSS),.VDD(VDD),.Y(g6105),.A(I7811));
  NOT NOT1_2920(.VSS(VSS),.VDD(VDD),.Y(I7814),.A(g5922));
  NOT NOT1_2921(.VSS(VSS),.VDD(VDD),.Y(g6106),.A(I7814));
  NOT NOT1_2922(.VSS(VSS),.VDD(VDD),.Y(I7817),.A(g5924));
  NOT NOT1_2923(.VSS(VSS),.VDD(VDD),.Y(g6107),.A(I7817));
  NOT NOT1_2924(.VSS(VSS),.VDD(VDD),.Y(g6115),.A(g5879));
  NOT NOT1_2925(.VSS(VSS),.VDD(VDD),.Y(g6117),.A(g5880));
  NOT NOT1_2926(.VSS(VSS),.VDD(VDD),.Y(I7829),.A(g5926));
  NOT NOT1_2927(.VSS(VSS),.VDD(VDD),.Y(g6119),.A(I7829));
  NOT NOT1_2928(.VSS(VSS),.VDD(VDD),.Y(I7832),.A(g5943));
  NOT NOT1_2929(.VSS(VSS),.VDD(VDD),.Y(g6120),.A(I7832));
  NOT NOT1_2930(.VSS(VSS),.VDD(VDD),.Y(I7835),.A(g5926));
  NOT NOT1_2931(.VSS(VSS),.VDD(VDD),.Y(g6121),.A(I7835));
  NOT NOT1_2932(.VSS(VSS),.VDD(VDD),.Y(I7838),.A(g5947));
  NOT NOT1_2933(.VSS(VSS),.VDD(VDD),.Y(g6122),.A(I7838));
  NOT NOT1_2934(.VSS(VSS),.VDD(VDD),.Y(I7852),.A(g5993));
  NOT NOT1_2935(.VSS(VSS),.VDD(VDD),.Y(g6134),.A(I7852));
  NOT NOT1_2936(.VSS(VSS),.VDD(VDD),.Y(I7856),.A(g5994));
  NOT NOT1_2937(.VSS(VSS),.VDD(VDD),.Y(g6136),.A(I7856));
  NOT NOT1_2938(.VSS(VSS),.VDD(VDD),.Y(I7859),.A(g6032));
  NOT NOT1_2939(.VSS(VSS),.VDD(VDD),.Y(g6137),.A(I7859));
  NOT NOT1_2940(.VSS(VSS),.VDD(VDD),.Y(I7865),.A(g6095));
  NOT NOT1_2941(.VSS(VSS),.VDD(VDD),.Y(g6143),.A(I7865));
  NOT NOT1_2942(.VSS(VSS),.VDD(VDD),.Y(I7871),.A(g6097));
  NOT NOT1_2943(.VSS(VSS),.VDD(VDD),.Y(g6147),.A(I7871));
  NOT NOT1_2944(.VSS(VSS),.VDD(VDD),.Y(g6160),.A(g5926));
  NOT NOT1_2945(.VSS(VSS),.VDD(VDD),.Y(g6161),.A(g5926));
  NOT NOT1_2946(.VSS(VSS),.VDD(VDD),.Y(g6162),.A(g5926));
  NOT NOT1_2947(.VSS(VSS),.VDD(VDD),.Y(g6163),.A(g5926));
  NOT NOT1_2948(.VSS(VSS),.VDD(VDD),.Y(g6164),.A(g5926));
  NOT NOT1_2949(.VSS(VSS),.VDD(VDD),.Y(g6165),.A(g5926));
  NOT NOT1_2950(.VSS(VSS),.VDD(VDD),.Y(I7892),.A(g5916));
  NOT NOT1_2951(.VSS(VSS),.VDD(VDD),.Y(g6166),.A(I7892));
  NOT NOT1_2952(.VSS(VSS),.VDD(VDD),.Y(g6188),.A(g5950));
  NOT NOT1_2953(.VSS(VSS),.VDD(VDD),.Y(g6192),.A(g5946));
  NOT NOT1_2954(.VSS(VSS),.VDD(VDD),.Y(g6193),.A(g5957));
  NOT NOT1_2955(.VSS(VSS),.VDD(VDD),.Y(I7906),.A(g5912));
  NOT NOT1_2956(.VSS(VSS),.VDD(VDD),.Y(g6194),.A(I7906));
  NOT NOT1_2957(.VSS(VSS),.VDD(VDD),.Y(g6211),.A(g5992));
  NOT NOT1_2958(.VSS(VSS),.VDD(VDD),.Y(I7910),.A(g5905));
  NOT NOT1_2959(.VSS(VSS),.VDD(VDD),.Y(g6212),.A(I7910));
  NOT NOT1_2960(.VSS(VSS),.VDD(VDD),.Y(g6229),.A(g6036));
  NOT NOT1_2961(.VSS(VSS),.VDD(VDD),.Y(g6230),.A(g6040));
  NOT NOT1_2962(.VSS(VSS),.VDD(VDD),.Y(g6231),.A(g6044));
  NOT NOT1_2963(.VSS(VSS),.VDD(VDD),.Y(g6232),.A(g6048));
  NOT NOT1_2964(.VSS(VSS),.VDD(VDD),.Y(g6233),.A(g6052));
  NOT NOT1_2965(.VSS(VSS),.VDD(VDD),.Y(g6234),.A(g6057));
  NOT NOT1_2966(.VSS(VSS),.VDD(VDD),.Y(g6235),.A(g6062));
  NOT NOT1_2967(.VSS(VSS),.VDD(VDD),.Y(g6236),.A(g6070));
  NOT NOT1_2968(.VSS(VSS),.VDD(VDD),.Y(I7960),.A(g5925));
  NOT NOT1_2969(.VSS(VSS),.VDD(VDD),.Y(g6276),.A(I7960));
  NOT NOT1_2970(.VSS(VSS),.VDD(VDD),.Y(I7963),.A(g6276));
  NOT NOT1_2971(.VSS(VSS),.VDD(VDD),.Y(g6277),.A(I7963));
  NOT NOT1_2972(.VSS(VSS),.VDD(VDD),.Y(I7966),.A(g6166));
  NOT NOT1_2973(.VSS(VSS),.VDD(VDD),.Y(g6278),.A(I7966));
  NOT NOT1_2974(.VSS(VSS),.VDD(VDD),.Y(I7996),.A(g6137));
  NOT NOT1_2975(.VSS(VSS),.VDD(VDD),.Y(g6282),.A(I7996));
  NOT NOT1_2976(.VSS(VSS),.VDD(VDD),.Y(I7999),.A(g6137));
  NOT NOT1_2977(.VSS(VSS),.VDD(VDD),.Y(g6283),.A(I7999));
  NOT NOT1_2978(.VSS(VSS),.VDD(VDD),.Y(I8002),.A(g6110));
  NOT NOT1_2979(.VSS(VSS),.VDD(VDD),.Y(g6284),.A(I8002));
  NOT NOT1_2980(.VSS(VSS),.VDD(VDD),.Y(I8005),.A(g6110));
  NOT NOT1_2981(.VSS(VSS),.VDD(VDD),.Y(g6285),.A(I8005));
  NOT NOT1_2982(.VSS(VSS),.VDD(VDD),.Y(I8027),.A(g6237));
  NOT NOT1_2983(.VSS(VSS),.VDD(VDD),.Y(g6305),.A(I8027));
  NOT NOT1_2984(.VSS(VSS),.VDD(VDD),.Y(I8030),.A(g6239));
  NOT NOT1_2985(.VSS(VSS),.VDD(VDD),.Y(g6306),.A(I8030));
  NOT NOT1_2986(.VSS(VSS),.VDD(VDD),.Y(I8034),.A(g6242));
  NOT NOT1_2987(.VSS(VSS),.VDD(VDD),.Y(g6308),.A(I8034));
  NOT NOT1_2988(.VSS(VSS),.VDD(VDD),.Y(I8040),.A(g6142));
  NOT NOT1_2989(.VSS(VSS),.VDD(VDD),.Y(g6312),.A(I8040));
  NOT NOT1_2990(.VSS(VSS),.VDD(VDD),.Y(I8044),.A(g6252));
  NOT NOT1_2991(.VSS(VSS),.VDD(VDD),.Y(g6314),.A(I8044));
  NOT NOT1_2992(.VSS(VSS),.VDD(VDD),.Y(I8051),.A(g6108));
  NOT NOT1_2993(.VSS(VSS),.VDD(VDD),.Y(g6319),.A(I8051));
  NOT NOT1_2994(.VSS(VSS),.VDD(VDD),.Y(I8056),.A(g6109));
  NOT NOT1_2995(.VSS(VSS),.VDD(VDD),.Y(g6322),.A(I8056));
  NOT NOT1_2996(.VSS(VSS),.VDD(VDD),.Y(I8061),.A(g6113));
  NOT NOT1_2997(.VSS(VSS),.VDD(VDD),.Y(g6325),.A(I8061));
  NOT NOT1_2998(.VSS(VSS),.VDD(VDD),.Y(I8066),.A(g6114));
  NOT NOT1_2999(.VSS(VSS),.VDD(VDD),.Y(g6328),.A(I8066));
  NOT NOT1_3000(.VSS(VSS),.VDD(VDD),.Y(I8070),.A(g6116));
  NOT NOT1_3001(.VSS(VSS),.VDD(VDD),.Y(g6330),.A(I8070));
  NOT NOT1_3002(.VSS(VSS),.VDD(VDD),.Y(I8074),.A(g6118));
  NOT NOT1_3003(.VSS(VSS),.VDD(VDD),.Y(g6332),.A(I8074));
  NOT NOT1_3004(.VSS(VSS),.VDD(VDD),.Y(I8089),.A(g6120));
  NOT NOT1_3005(.VSS(VSS),.VDD(VDD),.Y(g6337),.A(I8089));
  NOT NOT1_3006(.VSS(VSS),.VDD(VDD),.Y(I8093),.A(g6122));
  NOT NOT1_3007(.VSS(VSS),.VDD(VDD),.Y(g6339),.A(I8093));
  NOT NOT1_3008(.VSS(VSS),.VDD(VDD),.Y(I8103),.A(g6134));
  NOT NOT1_3009(.VSS(VSS),.VDD(VDD),.Y(g6347),.A(I8103));
  NOT NOT1_3010(.VSS(VSS),.VDD(VDD),.Y(I8107),.A(g6136));
  NOT NOT1_3011(.VSS(VSS),.VDD(VDD),.Y(g6351),.A(I8107));
  NOT NOT1_3012(.VSS(VSS),.VDD(VDD),.Y(I8110),.A(g6143));
  NOT NOT1_3013(.VSS(VSS),.VDD(VDD),.Y(g6352),.A(I8110));
  NOT NOT1_3014(.VSS(VSS),.VDD(VDD),.Y(I8113),.A(g6147));
  NOT NOT1_3015(.VSS(VSS),.VDD(VDD),.Y(g6353),.A(I8113));
  NOT NOT1_3016(.VSS(VSS),.VDD(VDD),.Y(I8144),.A(g6182));
  NOT NOT1_3017(.VSS(VSS),.VDD(VDD),.Y(g6360),.A(I8144));
  NOT NOT1_3018(.VSS(VSS),.VDD(VDD),.Y(I8147),.A(g6182));
  NOT NOT1_3019(.VSS(VSS),.VDD(VDD),.Y(g6361),.A(I8147));
  NOT NOT1_3020(.VSS(VSS),.VDD(VDD),.Y(I8150),.A(g6185));
  NOT NOT1_3021(.VSS(VSS),.VDD(VDD),.Y(g6362),.A(I8150));
  NOT NOT1_3022(.VSS(VSS),.VDD(VDD),.Y(I8153),.A(g6185));
  NOT NOT1_3023(.VSS(VSS),.VDD(VDD),.Y(g6363),.A(I8153));
  NOT NOT1_3024(.VSS(VSS),.VDD(VDD),.Y(I8156),.A(g6167));
  NOT NOT1_3025(.VSS(VSS),.VDD(VDD),.Y(g6364),.A(I8156));
  NOT NOT1_3026(.VSS(VSS),.VDD(VDD),.Y(I8159),.A(g6167));
  NOT NOT1_3027(.VSS(VSS),.VDD(VDD),.Y(g6365),.A(I8159));
  NOT NOT1_3028(.VSS(VSS),.VDD(VDD),.Y(I8162),.A(g6189));
  NOT NOT1_3029(.VSS(VSS),.VDD(VDD),.Y(g6366),.A(I8162));
  NOT NOT1_3030(.VSS(VSS),.VDD(VDD),.Y(I8165),.A(g6189));
  NOT NOT1_3031(.VSS(VSS),.VDD(VDD),.Y(g6367),.A(I8165));
  NOT NOT1_3032(.VSS(VSS),.VDD(VDD),.Y(I8168),.A(g6170));
  NOT NOT1_3033(.VSS(VSS),.VDD(VDD),.Y(g6368),.A(I8168));
  NOT NOT1_3034(.VSS(VSS),.VDD(VDD),.Y(I8171),.A(g6170));
  NOT NOT1_3035(.VSS(VSS),.VDD(VDD),.Y(g6369),.A(I8171));
  NOT NOT1_3036(.VSS(VSS),.VDD(VDD),.Y(I8174),.A(g6173));
  NOT NOT1_3037(.VSS(VSS),.VDD(VDD),.Y(g6370),.A(I8174));
  NOT NOT1_3038(.VSS(VSS),.VDD(VDD),.Y(I8177),.A(g6173));
  NOT NOT1_3039(.VSS(VSS),.VDD(VDD),.Y(g6371),.A(I8177));
  NOT NOT1_3040(.VSS(VSS),.VDD(VDD),.Y(I8180),.A(g6176));
  NOT NOT1_3041(.VSS(VSS),.VDD(VDD),.Y(g6372),.A(I8180));
  NOT NOT1_3042(.VSS(VSS),.VDD(VDD),.Y(I8183),.A(g6176));
  NOT NOT1_3043(.VSS(VSS),.VDD(VDD),.Y(g6373),.A(I8183));
  NOT NOT1_3044(.VSS(VSS),.VDD(VDD),.Y(I8186),.A(g6179));
  NOT NOT1_3045(.VSS(VSS),.VDD(VDD),.Y(g6374),.A(I8186));
  NOT NOT1_3046(.VSS(VSS),.VDD(VDD),.Y(I8189),.A(g6179));
  NOT NOT1_3047(.VSS(VSS),.VDD(VDD),.Y(g6375),.A(I8189));
  NOT NOT1_3048(.VSS(VSS),.VDD(VDD),.Y(g6376),.A(g6267));
  NOT NOT1_3049(.VSS(VSS),.VDD(VDD),.Y(g6385),.A(g6271));
  NOT NOT1_3050(.VSS(VSS),.VDD(VDD),.Y(I8217),.A(g6319));
  NOT NOT1_3051(.VSS(VSS),.VDD(VDD),.Y(g6401),.A(I8217));
  NOT NOT1_3052(.VSS(VSS),.VDD(VDD),.Y(I8220),.A(g6322));
  NOT NOT1_3053(.VSS(VSS),.VDD(VDD),.Y(g6402),.A(I8220));
  NOT NOT1_3054(.VSS(VSS),.VDD(VDD),.Y(I8223),.A(g6325));
  NOT NOT1_3055(.VSS(VSS),.VDD(VDD),.Y(g6403),.A(I8223));
  NOT NOT1_3056(.VSS(VSS),.VDD(VDD),.Y(I8226),.A(g6328));
  NOT NOT1_3057(.VSS(VSS),.VDD(VDD),.Y(g6404),.A(I8226));
  NOT NOT1_3058(.VSS(VSS),.VDD(VDD),.Y(I8229),.A(g6330));
  NOT NOT1_3059(.VSS(VSS),.VDD(VDD),.Y(g6405),.A(I8229));
  NOT NOT1_3060(.VSS(VSS),.VDD(VDD),.Y(I8232),.A(g6332));
  NOT NOT1_3061(.VSS(VSS),.VDD(VDD),.Y(g6406),.A(I8232));
  NOT NOT1_3062(.VSS(VSS),.VDD(VDD),.Y(I8235),.A(g6312));
  NOT NOT1_3063(.VSS(VSS),.VDD(VDD),.Y(g6407),.A(I8235));
  NOT NOT1_3064(.VSS(VSS),.VDD(VDD),.Y(g6408),.A(g6283));
  NOT NOT1_3065(.VSS(VSS),.VDD(VDD),.Y(g6409),.A(g6285));
  NOT NOT1_3066(.VSS(VSS),.VDD(VDD),.Y(I8240),.A(g6287));
  NOT NOT1_3067(.VSS(VSS),.VDD(VDD),.Y(g6410),.A(I8240));
  NOT NOT1_3068(.VSS(VSS),.VDD(VDD),.Y(I8243),.A(g6286));
  NOT NOT1_3069(.VSS(VSS),.VDD(VDD),.Y(g6411),.A(I8243));
  NOT NOT1_3070(.VSS(VSS),.VDD(VDD),.Y(I8246),.A(g6290));
  NOT NOT1_3071(.VSS(VSS),.VDD(VDD),.Y(g6412),.A(I8246));
  NOT NOT1_3072(.VSS(VSS),.VDD(VDD),.Y(I8249),.A(g6289));
  NOT NOT1_3073(.VSS(VSS),.VDD(VDD),.Y(g6413),.A(I8249));
  NOT NOT1_3074(.VSS(VSS),.VDD(VDD),.Y(I8252),.A(g6294));
  NOT NOT1_3075(.VSS(VSS),.VDD(VDD),.Y(g6414),.A(I8252));
  NOT NOT1_3076(.VSS(VSS),.VDD(VDD),.Y(I8255),.A(g6292));
  NOT NOT1_3077(.VSS(VSS),.VDD(VDD),.Y(g6415),.A(I8255));
  NOT NOT1_3078(.VSS(VSS),.VDD(VDD),.Y(I8258),.A(g6293));
  NOT NOT1_3079(.VSS(VSS),.VDD(VDD),.Y(g6416),.A(I8258));
  NOT NOT1_3080(.VSS(VSS),.VDD(VDD),.Y(I8261),.A(g6298));
  NOT NOT1_3081(.VSS(VSS),.VDD(VDD),.Y(g6417),.A(I8261));
  NOT NOT1_3082(.VSS(VSS),.VDD(VDD),.Y(I8264),.A(g6296));
  NOT NOT1_3083(.VSS(VSS),.VDD(VDD),.Y(g6418),.A(I8264));
  NOT NOT1_3084(.VSS(VSS),.VDD(VDD),.Y(I8267),.A(g6297));
  NOT NOT1_3085(.VSS(VSS),.VDD(VDD),.Y(g6419),.A(I8267));
  NOT NOT1_3086(.VSS(VSS),.VDD(VDD),.Y(I8270),.A(g6300));
  NOT NOT1_3087(.VSS(VSS),.VDD(VDD),.Y(g6420),.A(I8270));
  NOT NOT1_3088(.VSS(VSS),.VDD(VDD),.Y(I8273),.A(g6301));
  NOT NOT1_3089(.VSS(VSS),.VDD(VDD),.Y(g6421),.A(I8273));
  NOT NOT1_3090(.VSS(VSS),.VDD(VDD),.Y(I8276),.A(g6303));
  NOT NOT1_3091(.VSS(VSS),.VDD(VDD),.Y(g6422),.A(I8276));
  NOT NOT1_3092(.VSS(VSS),.VDD(VDD),.Y(I8279),.A(g6307));
  NOT NOT1_3093(.VSS(VSS),.VDD(VDD),.Y(g6423),.A(I8279));
  NOT NOT1_3094(.VSS(VSS),.VDD(VDD),.Y(I8282),.A(g6309));
  NOT NOT1_3095(.VSS(VSS),.VDD(VDD),.Y(g6424),.A(I8282));
  NOT NOT1_3096(.VSS(VSS),.VDD(VDD),.Y(I8285),.A(g6310));
  NOT NOT1_3097(.VSS(VSS),.VDD(VDD),.Y(g6425),.A(I8285));
  NOT NOT1_3098(.VSS(VSS),.VDD(VDD),.Y(I8290),.A(g6291));
  NOT NOT1_3099(.VSS(VSS),.VDD(VDD),.Y(g6428),.A(I8290));
  NOT NOT1_3100(.VSS(VSS),.VDD(VDD),.Y(I8295),.A(g6295));
  NOT NOT1_3101(.VSS(VSS),.VDD(VDD),.Y(g6431),.A(I8295));
  NOT NOT1_3102(.VSS(VSS),.VDD(VDD),.Y(I8300),.A(g6299));
  NOT NOT1_3103(.VSS(VSS),.VDD(VDD),.Y(g6434),.A(I8300));
  NOT NOT1_3104(.VSS(VSS),.VDD(VDD),.Y(I8309),.A(g6304));
  NOT NOT1_3105(.VSS(VSS),.VDD(VDD),.Y(g6441),.A(I8309));
  NOT NOT1_3106(.VSS(VSS),.VDD(VDD),.Y(I8329),.A(g6305));
  NOT NOT1_3107(.VSS(VSS),.VDD(VDD),.Y(g6465),.A(I8329));
  NOT NOT1_3108(.VSS(VSS),.VDD(VDD),.Y(I8332),.A(g6306));
  NOT NOT1_3109(.VSS(VSS),.VDD(VDD),.Y(g6466),.A(I8332));
  NOT NOT1_3110(.VSS(VSS),.VDD(VDD),.Y(I8335),.A(g6308));
  NOT NOT1_3111(.VSS(VSS),.VDD(VDD),.Y(g6467),.A(I8335));
  NOT NOT1_3112(.VSS(VSS),.VDD(VDD),.Y(I8342),.A(g6314));
  NOT NOT1_3113(.VSS(VSS),.VDD(VDD),.Y(g6478),.A(I8342));
  NOT NOT1_3114(.VSS(VSS),.VDD(VDD),.Y(g6484),.A(g6361));
  NOT NOT1_3115(.VSS(VSS),.VDD(VDD),.Y(g6486),.A(g6363));
  NOT NOT1_3116(.VSS(VSS),.VDD(VDD),.Y(g6487),.A(g6365));
  NOT NOT1_3117(.VSS(VSS),.VDD(VDD),.Y(g6488),.A(g6367));
  NOT NOT1_3118(.VSS(VSS),.VDD(VDD),.Y(g6489),.A(g6369));
  NOT NOT1_3119(.VSS(VSS),.VDD(VDD),.Y(g6490),.A(g6371));
  NOT NOT1_3120(.VSS(VSS),.VDD(VDD),.Y(g6491),.A(g6373));
  NOT NOT1_3121(.VSS(VSS),.VDD(VDD),.Y(g6493),.A(g6375));
  NOT NOT1_3122(.VSS(VSS),.VDD(VDD),.Y(I8411),.A(g6415));
  NOT NOT1_3123(.VSS(VSS),.VDD(VDD),.Y(g6497),.A(I8411));
  NOT NOT1_3124(.VSS(VSS),.VDD(VDD),.Y(I8414),.A(g6418));
  NOT NOT1_3125(.VSS(VSS),.VDD(VDD),.Y(g6498),.A(I8414));
  NOT NOT1_3126(.VSS(VSS),.VDD(VDD),.Y(I8417),.A(g6420));
  NOT NOT1_3127(.VSS(VSS),.VDD(VDD),.Y(g6499),.A(I8417));
  NOT NOT1_3128(.VSS(VSS),.VDD(VDD),.Y(I8420),.A(g6422));
  NOT NOT1_3129(.VSS(VSS),.VDD(VDD),.Y(g6500),.A(I8420));
  NOT NOT1_3130(.VSS(VSS),.VDD(VDD),.Y(I8423),.A(g6423));
  NOT NOT1_3131(.VSS(VSS),.VDD(VDD),.Y(g6501),.A(I8423));
  NOT NOT1_3132(.VSS(VSS),.VDD(VDD),.Y(I8426),.A(g6424));
  NOT NOT1_3133(.VSS(VSS),.VDD(VDD),.Y(g6502),.A(I8426));
  NOT NOT1_3134(.VSS(VSS),.VDD(VDD),.Y(I8429),.A(g6425));
  NOT NOT1_3135(.VSS(VSS),.VDD(VDD),.Y(g6503),.A(I8429));
  NOT NOT1_3136(.VSS(VSS),.VDD(VDD),.Y(I8432),.A(g6411));
  NOT NOT1_3137(.VSS(VSS),.VDD(VDD),.Y(g6504),.A(I8432));
  NOT NOT1_3138(.VSS(VSS),.VDD(VDD),.Y(I8435),.A(g6413));
  NOT NOT1_3139(.VSS(VSS),.VDD(VDD),.Y(g6505),.A(I8435));
  NOT NOT1_3140(.VSS(VSS),.VDD(VDD),.Y(I8438),.A(g6416));
  NOT NOT1_3141(.VSS(VSS),.VDD(VDD),.Y(g6506),.A(I8438));
  NOT NOT1_3142(.VSS(VSS),.VDD(VDD),.Y(I8441),.A(g6419));
  NOT NOT1_3143(.VSS(VSS),.VDD(VDD),.Y(g6507),.A(I8441));
  NOT NOT1_3144(.VSS(VSS),.VDD(VDD),.Y(I8444),.A(g6421));
  NOT NOT1_3145(.VSS(VSS),.VDD(VDD),.Y(g6508),.A(I8444));
  NOT NOT1_3146(.VSS(VSS),.VDD(VDD),.Y(I8447),.A(g6410));
  NOT NOT1_3147(.VSS(VSS),.VDD(VDD),.Y(g6509),.A(I8447));
  NOT NOT1_3148(.VSS(VSS),.VDD(VDD),.Y(I8450),.A(g6412));
  NOT NOT1_3149(.VSS(VSS),.VDD(VDD),.Y(g6510),.A(I8450));
  NOT NOT1_3150(.VSS(VSS),.VDD(VDD),.Y(I8453),.A(g6414));
  NOT NOT1_3151(.VSS(VSS),.VDD(VDD),.Y(g6511),.A(I8453));
  NOT NOT1_3152(.VSS(VSS),.VDD(VDD),.Y(I8456),.A(g6417));
  NOT NOT1_3153(.VSS(VSS),.VDD(VDD),.Y(g6512),.A(I8456));
  NOT NOT1_3154(.VSS(VSS),.VDD(VDD),.Y(I8459),.A(g6427));
  NOT NOT1_3155(.VSS(VSS),.VDD(VDD),.Y(g6513),.A(I8459));
  NOT NOT1_3156(.VSS(VSS),.VDD(VDD),.Y(I8462),.A(g6430));
  NOT NOT1_3157(.VSS(VSS),.VDD(VDD),.Y(g6514),.A(I8462));
  NOT NOT1_3158(.VSS(VSS),.VDD(VDD),.Y(g6515),.A(g6408));
  NOT NOT1_3159(.VSS(VSS),.VDD(VDD),.Y(g6516),.A(g6409));
  NOT NOT1_3160(.VSS(VSS),.VDD(VDD),.Y(I8467),.A(g6457));
  NOT NOT1_3161(.VSS(VSS),.VDD(VDD),.Y(g6517),.A(I8467));
  NOT NOT1_3162(.VSS(VSS),.VDD(VDD),.Y(I8470),.A(g6461));
  NOT NOT1_3163(.VSS(VSS),.VDD(VDD),.Y(g6518),.A(I8470));
  NOT NOT1_3164(.VSS(VSS),.VDD(VDD),.Y(I8473),.A(g6485));
  NOT NOT1_3165(.VSS(VSS),.VDD(VDD),.Y(g6519),.A(I8473));
  NOT NOT1_3166(.VSS(VSS),.VDD(VDD),.Y(I8476),.A(g6457));
  NOT NOT1_3167(.VSS(VSS),.VDD(VDD),.Y(g6520),.A(I8476));
  NOT NOT1_3168(.VSS(VSS),.VDD(VDD),.Y(I8479),.A(g6482));
  NOT NOT1_3169(.VSS(VSS),.VDD(VDD),.Y(g6521),.A(I8479));
  NOT NOT1_3170(.VSS(VSS),.VDD(VDD),.Y(I8482),.A(g6461));
  NOT NOT1_3171(.VSS(VSS),.VDD(VDD),.Y(g6522),.A(I8482));
  NOT NOT1_3172(.VSS(VSS),.VDD(VDD),.Y(I8485),.A(g6479));
  NOT NOT1_3173(.VSS(VSS),.VDD(VDD),.Y(g6523),.A(I8485));
  NOT NOT1_3174(.VSS(VSS),.VDD(VDD),.Y(I8488),.A(g6426));
  NOT NOT1_3175(.VSS(VSS),.VDD(VDD),.Y(g6524),.A(I8488));
  NOT NOT1_3176(.VSS(VSS),.VDD(VDD),.Y(I8491),.A(g6480));
  NOT NOT1_3177(.VSS(VSS),.VDD(VDD),.Y(g6525),.A(I8491));
  NOT NOT1_3178(.VSS(VSS),.VDD(VDD),.Y(I8494),.A(g6428));
  NOT NOT1_3179(.VSS(VSS),.VDD(VDD),.Y(g6526),.A(I8494));
  NOT NOT1_3180(.VSS(VSS),.VDD(VDD),.Y(I8497),.A(g6481));
  NOT NOT1_3181(.VSS(VSS),.VDD(VDD),.Y(g6527),.A(I8497));
  NOT NOT1_3182(.VSS(VSS),.VDD(VDD),.Y(I8500),.A(g6431));
  NOT NOT1_3183(.VSS(VSS),.VDD(VDD),.Y(g6528),.A(I8500));
  NOT NOT1_3184(.VSS(VSS),.VDD(VDD),.Y(I8503),.A(g6434));
  NOT NOT1_3185(.VSS(VSS),.VDD(VDD),.Y(g6529),.A(I8503));
  NOT NOT1_3186(.VSS(VSS),.VDD(VDD),.Y(I8506),.A(g6483));
  NOT NOT1_3187(.VSS(VSS),.VDD(VDD),.Y(g6530),.A(I8506));
  NOT NOT1_3188(.VSS(VSS),.VDD(VDD),.Y(I8509),.A(g6437));
  NOT NOT1_3189(.VSS(VSS),.VDD(VDD),.Y(g6531),.A(I8509));
  NOT NOT1_3190(.VSS(VSS),.VDD(VDD),.Y(I8512),.A(g6441));
  NOT NOT1_3191(.VSS(VSS),.VDD(VDD),.Y(g6532),.A(I8512));
  NOT NOT1_3192(.VSS(VSS),.VDD(VDD),.Y(I8515),.A(g6492));
  NOT NOT1_3193(.VSS(VSS),.VDD(VDD),.Y(g6533),.A(I8515));
  NOT NOT1_3194(.VSS(VSS),.VDD(VDD),.Y(I8518),.A(g6494));
  NOT NOT1_3195(.VSS(VSS),.VDD(VDD),.Y(g6534),.A(I8518));
  NOT NOT1_3196(.VSS(VSS),.VDD(VDD),.Y(I8521),.A(g6495));
  NOT NOT1_3197(.VSS(VSS),.VDD(VDD),.Y(g6535),.A(I8521));
  NOT NOT1_3198(.VSS(VSS),.VDD(VDD),.Y(I8524),.A(g6496));
  NOT NOT1_3199(.VSS(VSS),.VDD(VDD),.Y(g6536),.A(I8524));
  NOT NOT1_3200(.VSS(VSS),.VDD(VDD),.Y(I8527),.A(g6440));
  NOT NOT1_3201(.VSS(VSS),.VDD(VDD),.Y(g6537),.A(I8527));
  NOT NOT1_3202(.VSS(VSS),.VDD(VDD),.Y(g6538),.A(g6469));
  NOT NOT1_3203(.VSS(VSS),.VDD(VDD),.Y(I8531),.A(g6444));
  NOT NOT1_3204(.VSS(VSS),.VDD(VDD),.Y(g6539),.A(I8531));
  NOT NOT1_3205(.VSS(VSS),.VDD(VDD),.Y(g6540),.A(g6474));
  NOT NOT1_3206(.VSS(VSS),.VDD(VDD),.Y(I8535),.A(g6447));
  NOT NOT1_3207(.VSS(VSS),.VDD(VDD),.Y(g6541),.A(I8535));
  NOT NOT1_3208(.VSS(VSS),.VDD(VDD),.Y(I8538),.A(g6450));
  NOT NOT1_3209(.VSS(VSS),.VDD(VDD),.Y(g6542),.A(I8538));
  NOT NOT1_3210(.VSS(VSS),.VDD(VDD),.Y(I8541),.A(g6452));
  NOT NOT1_3211(.VSS(VSS),.VDD(VDD),.Y(g6543),.A(I8541));
  NOT NOT1_3212(.VSS(VSS),.VDD(VDD),.Y(I8544),.A(g6453));
  NOT NOT1_3213(.VSS(VSS),.VDD(VDD),.Y(g6544),.A(I8544));
  NOT NOT1_3214(.VSS(VSS),.VDD(VDD),.Y(I8548),.A(g6454));
  NOT NOT1_3215(.VSS(VSS),.VDD(VDD),.Y(g6548),.A(I8548));
  NOT NOT1_3216(.VSS(VSS),.VDD(VDD),.Y(I8552),.A(g6455));
  NOT NOT1_3217(.VSS(VSS),.VDD(VDD),.Y(g6552),.A(I8552));
  NOT NOT1_3218(.VSS(VSS),.VDD(VDD),.Y(I8555),.A(g6456));
  NOT NOT1_3219(.VSS(VSS),.VDD(VDD),.Y(g6553),.A(I8555));
  NOT NOT1_3220(.VSS(VSS),.VDD(VDD),.Y(I8564),.A(g6429));
  NOT NOT1_3221(.VSS(VSS),.VDD(VDD),.Y(g6560),.A(I8564));
  NOT NOT1_3222(.VSS(VSS),.VDD(VDD),.Y(I8567),.A(g6432));
  NOT NOT1_3223(.VSS(VSS),.VDD(VDD),.Y(g6561),.A(I8567));
  NOT NOT1_3224(.VSS(VSS),.VDD(VDD),.Y(I8570),.A(g6433));
  NOT NOT1_3225(.VSS(VSS),.VDD(VDD),.Y(g6562),.A(I8570));
  NOT NOT1_3226(.VSS(VSS),.VDD(VDD),.Y(I8573),.A(g6435));
  NOT NOT1_3227(.VSS(VSS),.VDD(VDD),.Y(g6563),.A(I8573));
  NOT NOT1_3228(.VSS(VSS),.VDD(VDD),.Y(I8576),.A(g6436));
  NOT NOT1_3229(.VSS(VSS),.VDD(VDD),.Y(g6564),.A(I8576));
  NOT NOT1_3230(.VSS(VSS),.VDD(VDD),.Y(I8579),.A(g6438));
  NOT NOT1_3231(.VSS(VSS),.VDD(VDD),.Y(g6565),.A(I8579));
  NOT NOT1_3232(.VSS(VSS),.VDD(VDD),.Y(I8582),.A(g6439));
  NOT NOT1_3233(.VSS(VSS),.VDD(VDD),.Y(g6566),.A(I8582));
  NOT NOT1_3234(.VSS(VSS),.VDD(VDD),.Y(I8585),.A(g6442));
  NOT NOT1_3235(.VSS(VSS),.VDD(VDD),.Y(g6567),.A(I8585));
  NOT NOT1_3236(.VSS(VSS),.VDD(VDD),.Y(I8588),.A(g6443));
  NOT NOT1_3237(.VSS(VSS),.VDD(VDD),.Y(g6568),.A(I8588));
  NOT NOT1_3238(.VSS(VSS),.VDD(VDD),.Y(I8591),.A(g6448));
  NOT NOT1_3239(.VSS(VSS),.VDD(VDD),.Y(g6569),.A(I8591));
  NOT NOT1_3240(.VSS(VSS),.VDD(VDD),.Y(I8594),.A(g6446));
  NOT NOT1_3241(.VSS(VSS),.VDD(VDD),.Y(g6570),.A(I8594));
  NOT NOT1_3242(.VSS(VSS),.VDD(VDD),.Y(I8597),.A(g6445));
  NOT NOT1_3243(.VSS(VSS),.VDD(VDD),.Y(g6571),.A(I8597));
  NOT NOT1_3244(.VSS(VSS),.VDD(VDD),.Y(I8600),.A(g6451));
  NOT NOT1_3245(.VSS(VSS),.VDD(VDD),.Y(g6572),.A(I8600));
  NOT NOT1_3246(.VSS(VSS),.VDD(VDD),.Y(I8603),.A(g6449));
  NOT NOT1_3247(.VSS(VSS),.VDD(VDD),.Y(g6573),.A(I8603));
  NOT NOT1_3248(.VSS(VSS),.VDD(VDD),.Y(g6574),.A(g6484));
  NOT NOT1_3249(.VSS(VSS),.VDD(VDD),.Y(g6575),.A(g6486));
  NOT NOT1_3250(.VSS(VSS),.VDD(VDD),.Y(g6576),.A(g6487));
  NOT NOT1_3251(.VSS(VSS),.VDD(VDD),.Y(g6577),.A(g6488));
  NOT NOT1_3252(.VSS(VSS),.VDD(VDD),.Y(g6578),.A(g6489));
  NOT NOT1_3253(.VSS(VSS),.VDD(VDD),.Y(g6579),.A(g6490));
  NOT NOT1_3254(.VSS(VSS),.VDD(VDD),.Y(g6580),.A(g6491));
  NOT NOT1_3255(.VSS(VSS),.VDD(VDD),.Y(g6581),.A(g6493));
  NOT NOT1_3256(.VSS(VSS),.VDD(VDD),.Y(I8614),.A(g6537));
  NOT NOT1_3257(.VSS(VSS),.VDD(VDD),.Y(g6582),.A(I8614));
  NOT NOT1_3258(.VSS(VSS),.VDD(VDD),.Y(I8617),.A(g6539));
  NOT NOT1_3259(.VSS(VSS),.VDD(VDD),.Y(g6583),.A(I8617));
  NOT NOT1_3260(.VSS(VSS),.VDD(VDD),.Y(I8620),.A(g6541));
  NOT NOT1_3261(.VSS(VSS),.VDD(VDD),.Y(g6584),.A(I8620));
  NOT NOT1_3262(.VSS(VSS),.VDD(VDD),.Y(I8623),.A(g6542));
  NOT NOT1_3263(.VSS(VSS),.VDD(VDD),.Y(g6585),.A(I8623));
  NOT NOT1_3264(.VSS(VSS),.VDD(VDD),.Y(I8626),.A(g6543));
  NOT NOT1_3265(.VSS(VSS),.VDD(VDD),.Y(g6586),.A(I8626));
  NOT NOT1_3266(.VSS(VSS),.VDD(VDD),.Y(I8629),.A(g6544));
  NOT NOT1_3267(.VSS(VSS),.VDD(VDD),.Y(g6587),.A(I8629));
  NOT NOT1_3268(.VSS(VSS),.VDD(VDD),.Y(I8632),.A(g6548));
  NOT NOT1_3269(.VSS(VSS),.VDD(VDD),.Y(g6588),.A(I8632));
  NOT NOT1_3270(.VSS(VSS),.VDD(VDD),.Y(I8635),.A(g6552));
  NOT NOT1_3271(.VSS(VSS),.VDD(VDD),.Y(g6589),.A(I8635));
  NOT NOT1_3272(.VSS(VSS),.VDD(VDD),.Y(I8638),.A(g6553));
  NOT NOT1_3273(.VSS(VSS),.VDD(VDD),.Y(g6590),.A(I8638));
  NOT NOT1_3274(.VSS(VSS),.VDD(VDD),.Y(I8641),.A(g6524));
  NOT NOT1_3275(.VSS(VSS),.VDD(VDD),.Y(g6591),.A(I8641));
  NOT NOT1_3276(.VSS(VSS),.VDD(VDD),.Y(I8644),.A(g6526));
  NOT NOT1_3277(.VSS(VSS),.VDD(VDD),.Y(g6592),.A(I8644));
  NOT NOT1_3278(.VSS(VSS),.VDD(VDD),.Y(I8647),.A(g6528));
  NOT NOT1_3279(.VSS(VSS),.VDD(VDD),.Y(g6593),.A(I8647));
  NOT NOT1_3280(.VSS(VSS),.VDD(VDD),.Y(I8650),.A(g6529));
  NOT NOT1_3281(.VSS(VSS),.VDD(VDD),.Y(g6594),.A(I8650));
  NOT NOT1_3282(.VSS(VSS),.VDD(VDD),.Y(I8653),.A(g6531));
  NOT NOT1_3283(.VSS(VSS),.VDD(VDD),.Y(g6595),.A(I8653));
  NOT NOT1_3284(.VSS(VSS),.VDD(VDD),.Y(I8656),.A(g6532));
  NOT NOT1_3285(.VSS(VSS),.VDD(VDD),.Y(g6596),.A(I8656));
  NOT NOT1_3286(.VSS(VSS),.VDD(VDD),.Y(I8659),.A(g6523));
  NOT NOT1_3287(.VSS(VSS),.VDD(VDD),.Y(g6597),.A(I8659));
  NOT NOT1_3288(.VSS(VSS),.VDD(VDD),.Y(I8662),.A(g6525));
  NOT NOT1_3289(.VSS(VSS),.VDD(VDD),.Y(g6598),.A(I8662));
  NOT NOT1_3290(.VSS(VSS),.VDD(VDD),.Y(I8665),.A(g6527));
  NOT NOT1_3291(.VSS(VSS),.VDD(VDD),.Y(g6599),.A(I8665));
  NOT NOT1_3292(.VSS(VSS),.VDD(VDD),.Y(I8668),.A(g6530));
  NOT NOT1_3293(.VSS(VSS),.VDD(VDD),.Y(g6600),.A(I8668));
  NOT NOT1_3294(.VSS(VSS),.VDD(VDD),.Y(I8671),.A(g6519));
  NOT NOT1_3295(.VSS(VSS),.VDD(VDD),.Y(g6601),.A(I8671));
  NOT NOT1_3296(.VSS(VSS),.VDD(VDD),.Y(I8674),.A(g6521));
  NOT NOT1_3297(.VSS(VSS),.VDD(VDD),.Y(g6602),.A(I8674));
  NOT NOT1_3298(.VSS(VSS),.VDD(VDD),.Y(I8678),.A(g6565));
  NOT NOT1_3299(.VSS(VSS),.VDD(VDD),.Y(g6604),.A(I8678));
  NOT NOT1_3300(.VSS(VSS),.VDD(VDD),.Y(I8681),.A(g6566));
  NOT NOT1_3301(.VSS(VSS),.VDD(VDD),.Y(g6605),.A(I8681));
  NOT NOT1_3302(.VSS(VSS),.VDD(VDD),.Y(I8684),.A(g6567));
  NOT NOT1_3303(.VSS(VSS),.VDD(VDD),.Y(g6606),.A(I8684));
  NOT NOT1_3304(.VSS(VSS),.VDD(VDD),.Y(I8687),.A(g6568));
  NOT NOT1_3305(.VSS(VSS),.VDD(VDD),.Y(g6607),.A(I8687));
  NOT NOT1_3306(.VSS(VSS),.VDD(VDD),.Y(I8690),.A(g6571));
  NOT NOT1_3307(.VSS(VSS),.VDD(VDD),.Y(g6608),.A(I8690));
  NOT NOT1_3308(.VSS(VSS),.VDD(VDD),.Y(I8693),.A(g6570));
  NOT NOT1_3309(.VSS(VSS),.VDD(VDD),.Y(g6609),.A(I8693));
  NOT NOT1_3310(.VSS(VSS),.VDD(VDD),.Y(I8696),.A(g6569));
  NOT NOT1_3311(.VSS(VSS),.VDD(VDD),.Y(g6610),.A(I8696));
  NOT NOT1_3312(.VSS(VSS),.VDD(VDD),.Y(I8699),.A(g6573));
  NOT NOT1_3313(.VSS(VSS),.VDD(VDD),.Y(g6611),.A(I8699));
  NOT NOT1_3314(.VSS(VSS),.VDD(VDD),.Y(I8702),.A(g6572));
  NOT NOT1_3315(.VSS(VSS),.VDD(VDD),.Y(g6612),.A(I8702));
  NOT NOT1_3316(.VSS(VSS),.VDD(VDD),.Y(I8707),.A(g6520));
  NOT NOT1_3317(.VSS(VSS),.VDD(VDD),.Y(g6615),.A(I8707));
  NOT NOT1_3318(.VSS(VSS),.VDD(VDD),.Y(I8710),.A(g6517));
  NOT NOT1_3319(.VSS(VSS),.VDD(VDD),.Y(g6616),.A(I8710));
  NOT NOT1_3320(.VSS(VSS),.VDD(VDD),.Y(I8713),.A(g6522));
  NOT NOT1_3321(.VSS(VSS),.VDD(VDD),.Y(g6617),.A(I8713));
  NOT NOT1_3322(.VSS(VSS),.VDD(VDD),.Y(I8716),.A(g6518));
  NOT NOT1_3323(.VSS(VSS),.VDD(VDD),.Y(g6618),.A(I8716));
  NOT NOT1_3324(.VSS(VSS),.VDD(VDD),.Y(I8721),.A(g6534));
  NOT NOT1_3325(.VSS(VSS),.VDD(VDD),.Y(g6621),.A(I8721));
  NOT NOT1_3326(.VSS(VSS),.VDD(VDD),.Y(I8724),.A(g6533));
  NOT NOT1_3327(.VSS(VSS),.VDD(VDD),.Y(g6622),.A(I8724));
  NOT NOT1_3328(.VSS(VSS),.VDD(VDD),.Y(I8727),.A(g6536));
  NOT NOT1_3329(.VSS(VSS),.VDD(VDD),.Y(g6623),.A(I8727));
  NOT NOT1_3330(.VSS(VSS),.VDD(VDD),.Y(I8730),.A(g6535));
  NOT NOT1_3331(.VSS(VSS),.VDD(VDD),.Y(g6624),.A(I8730));
  NOT NOT1_3332(.VSS(VSS),.VDD(VDD),.Y(I8745),.A(g6513));
  NOT NOT1_3333(.VSS(VSS),.VDD(VDD),.Y(g6649),.A(I8745));
  NOT NOT1_3334(.VSS(VSS),.VDD(VDD),.Y(I8749),.A(g6560));
  NOT NOT1_3335(.VSS(VSS),.VDD(VDD),.Y(g6651),.A(I8749));
  NOT NOT1_3336(.VSS(VSS),.VDD(VDD),.Y(I8752),.A(g6514));
  NOT NOT1_3337(.VSS(VSS),.VDD(VDD),.Y(g6652),.A(I8752));
  NOT NOT1_3338(.VSS(VSS),.VDD(VDD),.Y(I8755),.A(g6561));
  NOT NOT1_3339(.VSS(VSS),.VDD(VDD),.Y(g6653),.A(I8755));
  NOT NOT1_3340(.VSS(VSS),.VDD(VDD),.Y(I8758),.A(g6562));
  NOT NOT1_3341(.VSS(VSS),.VDD(VDD),.Y(g6654),.A(I8758));
  NOT NOT1_3342(.VSS(VSS),.VDD(VDD),.Y(I8761),.A(g6563));
  NOT NOT1_3343(.VSS(VSS),.VDD(VDD),.Y(g6655),.A(I8761));
  NOT NOT1_3344(.VSS(VSS),.VDD(VDD),.Y(I8764),.A(g6564));
  NOT NOT1_3345(.VSS(VSS),.VDD(VDD),.Y(g6656),.A(I8764));
  NOT NOT1_3346(.VSS(VSS),.VDD(VDD),.Y(I8767),.A(g6619));
  NOT NOT1_3347(.VSS(VSS),.VDD(VDD),.Y(g6657),.A(I8767));
  NOT NOT1_3348(.VSS(VSS),.VDD(VDD),.Y(I8800),.A(g6684));
  NOT NOT1_3349(.VSS(VSS),.VDD(VDD),.Y(g6694),.A(I8800));
  NOT NOT1_3350(.VSS(VSS),.VDD(VDD),.Y(I8803),.A(g6685));
  NOT NOT1_3351(.VSS(VSS),.VDD(VDD),.Y(g6695),.A(I8803));
  NOT NOT1_3352(.VSS(VSS),.VDD(VDD),.Y(I8806),.A(g6686));
  NOT NOT1_3353(.VSS(VSS),.VDD(VDD),.Y(g6696),.A(I8806));
  NOT NOT1_3354(.VSS(VSS),.VDD(VDD),.Y(I8809),.A(g6687));
  NOT NOT1_3355(.VSS(VSS),.VDD(VDD),.Y(g6697),.A(I8809));
  NOT NOT1_3356(.VSS(VSS),.VDD(VDD),.Y(I8812),.A(g6688));
  NOT NOT1_3357(.VSS(VSS),.VDD(VDD),.Y(g6698),.A(I8812));
  NOT NOT1_3358(.VSS(VSS),.VDD(VDD),.Y(I8815),.A(g6689));
  NOT NOT1_3359(.VSS(VSS),.VDD(VDD),.Y(g6699),.A(I8815));
  NOT NOT1_3360(.VSS(VSS),.VDD(VDD),.Y(I8818),.A(g6690));
  NOT NOT1_3361(.VSS(VSS),.VDD(VDD),.Y(g6700),.A(I8818));
  NOT NOT1_3362(.VSS(VSS),.VDD(VDD),.Y(I8821),.A(g6691));
  NOT NOT1_3363(.VSS(VSS),.VDD(VDD),.Y(g6701),.A(I8821));
  NOT NOT1_3364(.VSS(VSS),.VDD(VDD),.Y(I8828),.A(g6661));
  NOT NOT1_3365(.VSS(VSS),.VDD(VDD),.Y(g6706),.A(I8828));
  NOT NOT1_3366(.VSS(VSS),.VDD(VDD),.Y(I8831),.A(g6665));
  NOT NOT1_3367(.VSS(VSS),.VDD(VDD),.Y(g6707),.A(I8831));
  NOT NOT1_3368(.VSS(VSS),.VDD(VDD),.Y(I8834),.A(g6661));
  NOT NOT1_3369(.VSS(VSS),.VDD(VDD),.Y(g6708),.A(I8834));
  NOT NOT1_3370(.VSS(VSS),.VDD(VDD),.Y(I8837),.A(g6665));
  NOT NOT1_3371(.VSS(VSS),.VDD(VDD),.Y(g6709),.A(I8837));
  NOT NOT1_3372(.VSS(VSS),.VDD(VDD),.Y(I8840),.A(g6657));
  NOT NOT1_3373(.VSS(VSS),.VDD(VDD),.Y(g6710),.A(I8840));
  NOT NOT1_3374(.VSS(VSS),.VDD(VDD),.Y(I8843),.A(g6658));
  NOT NOT1_3375(.VSS(VSS),.VDD(VDD),.Y(g6711),.A(I8843));
  NOT NOT1_3376(.VSS(VSS),.VDD(VDD),.Y(g6712),.A(g6676));
  NOT NOT1_3377(.VSS(VSS),.VDD(VDD),.Y(g6713),.A(g6679));
  NOT NOT1_3378(.VSS(VSS),.VDD(VDD),.Y(g6714),.A(g6670));
  NOT NOT1_3379(.VSS(VSS),.VDD(VDD),.Y(g6715),.A(g6673));
  NOT NOT1_3380(.VSS(VSS),.VDD(VDD),.Y(I8854),.A(g6696));
  NOT NOT1_3381(.VSS(VSS),.VDD(VDD),.Y(g6720),.A(I8854));
  NOT NOT1_3382(.VSS(VSS),.VDD(VDD),.Y(I8857),.A(g6698));
  NOT NOT1_3383(.VSS(VSS),.VDD(VDD),.Y(g6721),.A(I8857));
  NOT NOT1_3384(.VSS(VSS),.VDD(VDD),.Y(I8860),.A(g6699));
  NOT NOT1_3385(.VSS(VSS),.VDD(VDD),.Y(g6722),.A(I8860));
  NOT NOT1_3386(.VSS(VSS),.VDD(VDD),.Y(I8863),.A(g6700));
  NOT NOT1_3387(.VSS(VSS),.VDD(VDD),.Y(g6723),.A(I8863));
  NOT NOT1_3388(.VSS(VSS),.VDD(VDD),.Y(I8866),.A(g6701));
  NOT NOT1_3389(.VSS(VSS),.VDD(VDD),.Y(g6724),.A(I8866));
  NOT NOT1_3390(.VSS(VSS),.VDD(VDD),.Y(I8869),.A(g6694));
  NOT NOT1_3391(.VSS(VSS),.VDD(VDD),.Y(g6725),.A(I8869));
  NOT NOT1_3392(.VSS(VSS),.VDD(VDD),.Y(I8872),.A(g6695));
  NOT NOT1_3393(.VSS(VSS),.VDD(VDD),.Y(g6726),.A(I8872));
  NOT NOT1_3394(.VSS(VSS),.VDD(VDD),.Y(I8875),.A(g6697));
  NOT NOT1_3395(.VSS(VSS),.VDD(VDD),.Y(g6727),.A(I8875));
  NOT NOT1_3396(.VSS(VSS),.VDD(VDD),.Y(I8878),.A(g6710));
  NOT NOT1_3397(.VSS(VSS),.VDD(VDD),.Y(g6728),.A(I8878));
  NOT NOT1_3398(.VSS(VSS),.VDD(VDD),.Y(I8881),.A(g6711));
  NOT NOT1_3399(.VSS(VSS),.VDD(VDD),.Y(g6729),.A(I8881));
  NOT NOT1_3400(.VSS(VSS),.VDD(VDD),.Y(I8884),.A(g6704));
  NOT NOT1_3401(.VSS(VSS),.VDD(VDD),.Y(g6730),.A(I8884));
  NOT NOT1_3402(.VSS(VSS),.VDD(VDD),.Y(I8888),.A(g6708));
  NOT NOT1_3403(.VSS(VSS),.VDD(VDD),.Y(g6732),.A(I8888));
  NOT NOT1_3404(.VSS(VSS),.VDD(VDD),.Y(I8891),.A(g6706));
  NOT NOT1_3405(.VSS(VSS),.VDD(VDD),.Y(g6733),.A(I8891));
  NOT NOT1_3406(.VSS(VSS),.VDD(VDD),.Y(I8894),.A(g6709));
  NOT NOT1_3407(.VSS(VSS),.VDD(VDD),.Y(g6734),.A(I8894));
  NOT NOT1_3408(.VSS(VSS),.VDD(VDD),.Y(I8897),.A(g6707));
  NOT NOT1_3409(.VSS(VSS),.VDD(VDD),.Y(g6735),.A(I8897));
  NOT NOT1_3410(.VSS(VSS),.VDD(VDD),.Y(I8907),.A(g6702));
  NOT NOT1_3411(.VSS(VSS),.VDD(VDD),.Y(g6743),.A(I8907));
  NOT NOT1_3412(.VSS(VSS),.VDD(VDD),.Y(I8910),.A(g6730));
  NOT NOT1_3413(.VSS(VSS),.VDD(VDD),.Y(g6744),.A(I8910));
  NOT NOT1_3414(.VSS(VSS),.VDD(VDD),.Y(I8913),.A(g6743));
  NOT NOT1_3415(.VSS(VSS),.VDD(VDD),.Y(g6745),.A(I8913));
  NOT NOT1_3416(.VSS(VSS),.VDD(VDD),.Y(I8916),.A(g6742));
  NOT NOT1_3417(.VSS(VSS),.VDD(VDD),.Y(g6746),.A(I8916));
  NOT NOT1_3418(.VSS(VSS),.VDD(VDD),.Y(I8940),.A(g6783));
  NOT NOT1_3419(.VSS(VSS),.VDD(VDD),.Y(g6784),.A(I8940));
  NOT NOT1_3420(.VSS(VSS),.VDD(VDD),.Y(I8943),.A(g6774));
  NOT NOT1_3421(.VSS(VSS),.VDD(VDD),.Y(g6785),.A(I8943));
  NOT NOT1_3422(.VSS(VSS),.VDD(VDD),.Y(I8946),.A(g6778));
  NOT NOT1_3423(.VSS(VSS),.VDD(VDD),.Y(g6786),.A(I8946));
  NOT NOT1_3424(.VSS(VSS),.VDD(VDD),.Y(I8958),.A(g6774));
  NOT NOT1_3425(.VSS(VSS),.VDD(VDD),.Y(g6796),.A(I8958));
  NOT NOT1_3426(.VSS(VSS),.VDD(VDD),.Y(I8961),.A(g6778));
  NOT NOT1_3427(.VSS(VSS),.VDD(VDD),.Y(g6797),.A(I8961));
  NOT NOT1_3428(.VSS(VSS),.VDD(VDD),.Y(I8966),.A(g6796));
  NOT NOT1_3429(.VSS(VSS),.VDD(VDD),.Y(g6800),.A(I8966));
  NOT NOT1_3430(.VSS(VSS),.VDD(VDD),.Y(I8969),.A(g6797));
  NOT NOT1_3431(.VSS(VSS),.VDD(VDD),.Y(g6801),.A(I8969));
  NOT NOT1_3432(.VSS(VSS),.VDD(VDD),.Y(I8972),.A(g6795));
  NOT NOT1_3433(.VSS(VSS),.VDD(VDD),.Y(g6802),.A(I8972));
  NOT NOT1_3434(.VSS(VSS),.VDD(VDD),.Y(I8975),.A(g6791));
  NOT NOT1_3435(.VSS(VSS),.VDD(VDD),.Y(g6803),.A(I8975));
  NOT NOT1_3436(.VSS(VSS),.VDD(VDD),.Y(I8978),.A(g6792));
  NOT NOT1_3437(.VSS(VSS),.VDD(VDD),.Y(g6806),.A(I8978));
  NOT NOT1_3438(.VSS(VSS),.VDD(VDD),.Y(I8981),.A(g6793));
  NOT NOT1_3439(.VSS(VSS),.VDD(VDD),.Y(g6809),.A(I8981));
  NOT NOT1_3440(.VSS(VSS),.VDD(VDD),.Y(I8984),.A(g6794));
  NOT NOT1_3441(.VSS(VSS),.VDD(VDD),.Y(g6812),.A(I8984));
  NOT NOT1_3442(.VSS(VSS),.VDD(VDD),.Y(I8988),.A(g6787));
  NOT NOT1_3443(.VSS(VSS),.VDD(VDD),.Y(g6817),.A(I8988));
  NOT NOT1_3444(.VSS(VSS),.VDD(VDD),.Y(I8991),.A(g6788));
  NOT NOT1_3445(.VSS(VSS),.VDD(VDD),.Y(g6818),.A(I8991));
  NOT NOT1_3446(.VSS(VSS),.VDD(VDD),.Y(I8994),.A(g6789));
  NOT NOT1_3447(.VSS(VSS),.VDD(VDD),.Y(g6819),.A(I8994));
  NOT NOT1_3448(.VSS(VSS),.VDD(VDD),.Y(I8997),.A(g6790));
  NOT NOT1_3449(.VSS(VSS),.VDD(VDD),.Y(g6820),.A(I8997));
  NOT NOT1_3450(.VSS(VSS),.VDD(VDD),.Y(g6821),.A(g6785));
  NOT NOT1_3451(.VSS(VSS),.VDD(VDD),.Y(g6822),.A(g6786));
  NOT NOT1_3452(.VSS(VSS),.VDD(VDD),.Y(I9002),.A(g6802));
  NOT NOT1_3453(.VSS(VSS),.VDD(VDD),.Y(g6823),.A(I9002));
  NOT NOT1_3454(.VSS(VSS),.VDD(VDD),.Y(I9005),.A(g6817));
  NOT NOT1_3455(.VSS(VSS),.VDD(VDD),.Y(g6824),.A(I9005));
  NOT NOT1_3456(.VSS(VSS),.VDD(VDD),.Y(I9008),.A(g6818));
  NOT NOT1_3457(.VSS(VSS),.VDD(VDD),.Y(g6825),.A(I9008));
  NOT NOT1_3458(.VSS(VSS),.VDD(VDD),.Y(I9011),.A(g6819));
  NOT NOT1_3459(.VSS(VSS),.VDD(VDD),.Y(g6826),.A(I9011));
  NOT NOT1_3460(.VSS(VSS),.VDD(VDD),.Y(I9014),.A(g6820));
  NOT NOT1_3461(.VSS(VSS),.VDD(VDD),.Y(g6827),.A(I9014));
  NOT NOT1_3462(.VSS(VSS),.VDD(VDD),.Y(I9021),.A(g6812));
  NOT NOT1_3463(.VSS(VSS),.VDD(VDD),.Y(g6832),.A(I9021));
  NOT NOT1_3464(.VSS(VSS),.VDD(VDD),.Y(I9024),.A(g6803));
  NOT NOT1_3465(.VSS(VSS),.VDD(VDD),.Y(g6833),.A(I9024));
  NOT NOT1_3466(.VSS(VSS),.VDD(VDD),.Y(g6834),.A(g6821));
  NOT NOT1_3467(.VSS(VSS),.VDD(VDD),.Y(I9028),.A(g6806));
  NOT NOT1_3468(.VSS(VSS),.VDD(VDD),.Y(g6835),.A(I9028));
  NOT NOT1_3469(.VSS(VSS),.VDD(VDD),.Y(I9031),.A(g6809));
  NOT NOT1_3470(.VSS(VSS),.VDD(VDD),.Y(g6836),.A(I9031));
  NOT NOT1_3471(.VSS(VSS),.VDD(VDD),.Y(g6837),.A(g6822));
  NOT NOT1_3472(.VSS(VSS),.VDD(VDD),.Y(I9035),.A(g6812));
  NOT NOT1_3473(.VSS(VSS),.VDD(VDD),.Y(g6838),.A(I9035));
  NOT NOT1_3474(.VSS(VSS),.VDD(VDD),.Y(I9038),.A(g6833));
  NOT NOT1_3475(.VSS(VSS),.VDD(VDD),.Y(g6839),.A(I9038));
  NOT NOT1_3476(.VSS(VSS),.VDD(VDD),.Y(I9041),.A(g6835));
  NOT NOT1_3477(.VSS(VSS),.VDD(VDD),.Y(g6840),.A(I9041));
  NOT NOT1_3478(.VSS(VSS),.VDD(VDD),.Y(I9044),.A(g6836));
  NOT NOT1_3479(.VSS(VSS),.VDD(VDD),.Y(g6841),.A(I9044));
  NOT NOT1_3480(.VSS(VSS),.VDD(VDD),.Y(I9047),.A(g6838));
  NOT NOT1_3481(.VSS(VSS),.VDD(VDD),.Y(g6842),.A(I9047));
  NOT NOT1_3482(.VSS(VSS),.VDD(VDD),.Y(I9074),.A(g6844));
  NOT NOT1_3483(.VSS(VSS),.VDD(VDD),.Y(g6849),.A(I9074));
  NOT NOT1_3484(.VSS(VSS),.VDD(VDD),.Y(I9077),.A(g6845));
  NOT NOT1_3485(.VSS(VSS),.VDD(VDD),.Y(g6850),.A(I9077));
  NOT NOT1_3486(.VSS(VSS),.VDD(VDD),.Y(I9082),.A(g6849));
  NOT NOT1_3487(.VSS(VSS),.VDD(VDD),.Y(g6853),.A(I9082));
  NOT NOT1_3488(.VSS(VSS),.VDD(VDD),.Y(I9085),.A(g6850));
  NOT NOT1_3489(.VSS(VSS),.VDD(VDD),.Y(g6854),.A(I9085));
  NOT NOT1_3490(.VSS(VSS),.VDD(VDD),.Y(I9092),.A(g6855));
  NOT NOT1_3491(.VSS(VSS),.VDD(VDD),.Y(g6875),.A(I9092));
  NOT NOT1_3492(.VSS(VSS),.VDD(VDD),.Y(I9095),.A(g6855));
  NOT NOT1_3493(.VSS(VSS),.VDD(VDD),.Y(g6876),.A(I9095));
  NOT NOT1_3494(.VSS(VSS),.VDD(VDD),.Y(I9098),.A(g6864));
  NOT NOT1_3495(.VSS(VSS),.VDD(VDD),.Y(g6877),.A(I9098));
  NOT NOT1_3496(.VSS(VSS),.VDD(VDD),.Y(I9101),.A(g6855));
  NOT NOT1_3497(.VSS(VSS),.VDD(VDD),.Y(g6878),.A(I9101));
  NOT NOT1_3498(.VSS(VSS),.VDD(VDD),.Y(I9104),.A(g6864));
  NOT NOT1_3499(.VSS(VSS),.VDD(VDD),.Y(g6879),.A(I9104));
  NOT NOT1_3500(.VSS(VSS),.VDD(VDD),.Y(I9107),.A(g6855));
  NOT NOT1_3501(.VSS(VSS),.VDD(VDD),.Y(g6880),.A(I9107));
  NOT NOT1_3502(.VSS(VSS),.VDD(VDD),.Y(I9110),.A(g6864));
  NOT NOT1_3503(.VSS(VSS),.VDD(VDD),.Y(g6881),.A(I9110));
  NOT NOT1_3504(.VSS(VSS),.VDD(VDD),.Y(I9113),.A(g6855));
  NOT NOT1_3505(.VSS(VSS),.VDD(VDD),.Y(g6882),.A(I9113));
  NOT NOT1_3506(.VSS(VSS),.VDD(VDD),.Y(I9116),.A(g6864));
  NOT NOT1_3507(.VSS(VSS),.VDD(VDD),.Y(g6883),.A(I9116));
  NOT NOT1_3508(.VSS(VSS),.VDD(VDD),.Y(I9119),.A(g6855));
  NOT NOT1_3509(.VSS(VSS),.VDD(VDD),.Y(g6884),.A(I9119));
  NOT NOT1_3510(.VSS(VSS),.VDD(VDD),.Y(I9122),.A(g6864));
  NOT NOT1_3511(.VSS(VSS),.VDD(VDD),.Y(g6885),.A(I9122));
  NOT NOT1_3512(.VSS(VSS),.VDD(VDD),.Y(I9125),.A(g6855));
  NOT NOT1_3513(.VSS(VSS),.VDD(VDD),.Y(g6886),.A(I9125));
  NOT NOT1_3514(.VSS(VSS),.VDD(VDD),.Y(I9128),.A(g6864));
  NOT NOT1_3515(.VSS(VSS),.VDD(VDD),.Y(g6887),.A(I9128));
  NOT NOT1_3516(.VSS(VSS),.VDD(VDD),.Y(I9131),.A(g6855));
  NOT NOT1_3517(.VSS(VSS),.VDD(VDD),.Y(g6888),.A(I9131));
  NOT NOT1_3518(.VSS(VSS),.VDD(VDD),.Y(I9134),.A(g6864));
  NOT NOT1_3519(.VSS(VSS),.VDD(VDD),.Y(g6889),.A(I9134));
  NOT NOT1_3520(.VSS(VSS),.VDD(VDD),.Y(I9137),.A(g6864));
  NOT NOT1_3521(.VSS(VSS),.VDD(VDD),.Y(g6890),.A(I9137));
  NOT NOT1_3522(.VSS(VSS),.VDD(VDD),.Y(I9140),.A(g6888));
  NOT NOT1_3523(.VSS(VSS),.VDD(VDD),.Y(g6891),.A(I9140));
  NOT NOT1_3524(.VSS(VSS),.VDD(VDD),.Y(I9143),.A(g6886));
  NOT NOT1_3525(.VSS(VSS),.VDD(VDD),.Y(g6892),.A(I9143));
  NOT NOT1_3526(.VSS(VSS),.VDD(VDD),.Y(I9146),.A(g6890));
  NOT NOT1_3527(.VSS(VSS),.VDD(VDD),.Y(g6893),.A(I9146));
  NOT NOT1_3528(.VSS(VSS),.VDD(VDD),.Y(I9149),.A(g6884));
  NOT NOT1_3529(.VSS(VSS),.VDD(VDD),.Y(g6894),.A(I9149));
  NOT NOT1_3530(.VSS(VSS),.VDD(VDD),.Y(I9152),.A(g6889));
  NOT NOT1_3531(.VSS(VSS),.VDD(VDD),.Y(g6895),.A(I9152));
  NOT NOT1_3532(.VSS(VSS),.VDD(VDD),.Y(I9155),.A(g6882));
  NOT NOT1_3533(.VSS(VSS),.VDD(VDD),.Y(g6896),.A(I9155));
  NOT NOT1_3534(.VSS(VSS),.VDD(VDD),.Y(I9158),.A(g6887));
  NOT NOT1_3535(.VSS(VSS),.VDD(VDD),.Y(g6897),.A(I9158));
  NOT NOT1_3536(.VSS(VSS),.VDD(VDD),.Y(I9161),.A(g6880));
  NOT NOT1_3537(.VSS(VSS),.VDD(VDD),.Y(g6898),.A(I9161));
  NOT NOT1_3538(.VSS(VSS),.VDD(VDD),.Y(I9164),.A(g6885));
  NOT NOT1_3539(.VSS(VSS),.VDD(VDD),.Y(g6899),.A(I9164));
  NOT NOT1_3540(.VSS(VSS),.VDD(VDD),.Y(I9167),.A(g6878));
  NOT NOT1_3541(.VSS(VSS),.VDD(VDD),.Y(g6900),.A(I9167));
  NOT NOT1_3542(.VSS(VSS),.VDD(VDD),.Y(I9170),.A(g6883));
  NOT NOT1_3543(.VSS(VSS),.VDD(VDD),.Y(g6901),.A(I9170));
  NOT NOT1_3544(.VSS(VSS),.VDD(VDD),.Y(I9173),.A(g6876));
  NOT NOT1_3545(.VSS(VSS),.VDD(VDD),.Y(g6902),.A(I9173));
  NOT NOT1_3546(.VSS(VSS),.VDD(VDD),.Y(I9176),.A(g6881));
  NOT NOT1_3547(.VSS(VSS),.VDD(VDD),.Y(g6903),.A(I9176));
  NOT NOT1_3548(.VSS(VSS),.VDD(VDD),.Y(I9179),.A(g6875));
  NOT NOT1_3549(.VSS(VSS),.VDD(VDD),.Y(g6904),.A(I9179));
  NOT NOT1_3550(.VSS(VSS),.VDD(VDD),.Y(I9182),.A(g6879));
  NOT NOT1_3551(.VSS(VSS),.VDD(VDD),.Y(g6905),.A(I9182));
  NOT NOT1_3552(.VSS(VSS),.VDD(VDD),.Y(I9185),.A(g6877));
  NOT NOT1_3553(.VSS(VSS),.VDD(VDD),.Y(g6906),.A(I9185));
  NOT NOT1_3554(.VSS(VSS),.VDD(VDD),.Y(I9203),.A(g6921));
  NOT NOT1_3555(.VSS(VSS),.VDD(VDD),.Y(g6922),.A(I9203));
  NOT NOT1_3556(.VSS(VSS),.VDD(VDD),.Y(I9208),.A(g6922));
  NOT NOT1_3557(.VSS(VSS),.VDD(VDD),.Y(g6925),.A(I9208));
  NOT NOT1_3558(.VSS(VSS),.VDD(VDD),.Y(I9217),.A(g6931));
  NOT NOT1_3559(.VSS(VSS),.VDD(VDD),.Y(g6932),.A(I9217));
  NOT NOT1_3560(.VSS(VSS),.VDD(VDD),.Y(I9220),.A(g6930));
  NOT NOT1_3561(.VSS(VSS),.VDD(VDD),.Y(g6933),.A(I9220));
  NOT NOT1_3562(.VSS(VSS),.VDD(VDD),.Y(I9227),.A(g6937));
  NOT NOT1_3563(.VSS(VSS),.VDD(VDD),.Y(g6938),.A(I9227));
  NOT NOT1_3564(.VSS(VSS),.VDD(VDD),.Y(I9230),.A(g6936));
  NOT NOT1_3565(.VSS(VSS),.VDD(VDD),.Y(g6939),.A(I9230));
  NOT NOT1_3566(.VSS(VSS),.VDD(VDD),.Y(I9233),.A(g6938));
  NOT NOT1_3567(.VSS(VSS),.VDD(VDD),.Y(g6940),.A(I9233));
  NOT NOT1_3568(.VSS(VSS),.VDD(VDD),.Y(I9236),.A(g6939));
  NOT NOT1_3569(.VSS(VSS),.VDD(VDD),.Y(g6941),.A(I9236));
//
  AND2 AND2_0(.VSS(VSS),.VDD(VDD),.Y(g918),.A(g610),.B(g602));
  AND2 AND2_1(.VSS(VSS),.VDD(VDD),.Y(g1027),.A(g598),.B(g567));
  AND2 AND2_2(.VSS(VSS),.VDD(VDD),.Y(g1407),.A(g301),.B(g866));
  AND2 AND2_3(.VSS(VSS),.VDD(VDD),.Y(g1416),.A(g913),.B(g266));
  AND2 AND2_4(.VSS(VSS),.VDD(VDD),.Y(g1419),.A(g613),.B(g918));
  AND2 AND2_5(.VSS(VSS),.VDD(VDD),.Y(g1436),.A(g834),.B(g830));
  AND2 AND2_6(.VSS(VSS),.VDD(VDD),.Y(g1499),.A(g1101),.B(g1094));
  AND2 AND2_7(.VSS(VSS),.VDD(VDD),.Y(g1514),.A(g1017),.B(g1011));
  AND2 AND2_8(.VSS(VSS),.VDD(VDD),.Y(g1570),.A(g634),.B(g1027));
  AND2 AND2_9(.VSS(VSS),.VDD(VDD),.Y(g1575),.A(g980),.B(g965));
  AND2 AND2_10(.VSS(VSS),.VDD(VDD),.Y(g1576),.A(g1101),.B(g1094));
  AND2 AND2_11(.VSS(VSS),.VDD(VDD),.Y(g1585),.A(g1017),.B(g1011));
  AND3 AND3_0(.VSS(VSS),.VDD(VDD),.Y(I2566),.A(g749),.B(g743),.C(g736));
  AND4 AND4_0(.VSS(VSS),.VDD(VDD),.Y(g1595),.A(g729),.B(g719),.C(g766),.D(I2566));
  AND2 AND2_12(.VSS(VSS),.VDD(VDD),.Y(g1609),.A(g760),.B(g754));
  AND3 AND3_1(.VSS(VSS),.VDD(VDD),.Y(I2574),.A(g804),.B(g798),.C(g791));
  AND4 AND4_1(.VSS(VSS),.VDD(VDD),.Y(g1612),.A(g784),.B(g774),.C(g821),.D(I2574));
  AND2 AND2_13(.VSS(VSS),.VDD(VDD),.Y(g1620),.A(g1056),.B(g1084));
  AND2 AND2_14(.VSS(VSS),.VDD(VDD),.Y(g1628),.A(g815),.B(g809));
  AND2 AND2_15(.VSS(VSS),.VDD(VDD),.Y(g1633),.A(g716),.B(g152));
  AND2 AND2_16(.VSS(VSS),.VDD(VDD),.Y(g1689),.A(g766),.B(g719));
  AND2 AND2_17(.VSS(VSS),.VDD(VDD),.Y(g1691),.A(g821),.B(g774));
  AND3 AND3_2(.VSS(VSS),.VDD(VDD),.Y(g1706),.A(g766),.B(g719),.C(g729));
  AND3 AND3_3(.VSS(VSS),.VDD(VDD),.Y(g1716),.A(g821),.B(g774),.C(g784));
  AND2 AND2_18(.VSS(VSS),.VDD(VDD),.Y(g1763),.A(g478),.B(g1119));
  AND2 AND2_19(.VSS(VSS),.VDD(VDD),.Y(g1784),.A(g858),.B(g889));
  AND2 AND2_20(.VSS(VSS),.VDD(VDD),.Y(g1802),.A(g89),.B(g1064));
  AND2 AND2_21(.VSS(VSS),.VDD(VDD),.Y(g1808),.A(g706),.B(g49));
  AND2 AND2_22(.VSS(VSS),.VDD(VDD),.Y(g1826),.A(g714),.B(g710));
  AND2 AND2_23(.VSS(VSS),.VDD(VDD),.Y(g2015),.A(g616),.B(g1419));
  AND2 AND2_24(.VSS(VSS),.VDD(VDD),.Y(g2018),.A(g1423),.B(g1254));
  AND2 AND2_25(.VSS(VSS),.VDD(VDD),.Y(g2021),.A(g835),.B(g1436));
  AND4 AND4_2(.VSS(VSS),.VDD(VDD),.Y(g2026),.A(g1359),.B(g1402),.C(g1398),.D(g901));
  AND2 AND2_26(.VSS(VSS),.VDD(VDD),.Y(g2053),.A(g1094),.B(g1675));
  AND2 AND2_27(.VSS(VSS),.VDD(VDD),.Y(g2056),.A(g1672),.B(g1675));
  AND2 AND2_28(.VSS(VSS),.VDD(VDD),.Y(g2062),.A(g1499),.B(g1666));
  AND2 AND2_29(.VSS(VSS),.VDD(VDD),.Y(g2068),.A(g1541),.B(g1546));
  AND2 AND2_30(.VSS(VSS),.VDD(VDD),.Y(g2073),.A(g1088),.B(g1499));
  AND2 AND2_31(.VSS(VSS),.VDD(VDD),.Y(g2081),.A(g1094),.B(g1546));
  AND2 AND2_32(.VSS(VSS),.VDD(VDD),.Y(g2084),.A(g1577),.B(g1563));
  AND2 AND2_33(.VSS(VSS),.VDD(VDD),.Y(g2085),.A(g1123),.B(g1567));
  AND2 AND2_34(.VSS(VSS),.VDD(VDD),.Y(g2089),.A(g1123),.B(g1578));
  AND2 AND2_35(.VSS(VSS),.VDD(VDD),.Y(g2092),.A(g642),.B(g1570));
  AND2 AND2_36(.VSS(VSS),.VDD(VDD),.Y(g2101),.A(g1001),.B(g1543));
  AND2 AND2_37(.VSS(VSS),.VDD(VDD),.Y(g2107),.A(g1583),.B(g1543));
  AND2 AND2_38(.VSS(VSS),.VDD(VDD),.Y(g2113),.A(g1576),.B(g1535));
  AND2 AND2_39(.VSS(VSS),.VDD(VDD),.Y(g2121),.A(g1632),.B(g754));
  AND2 AND2_40(.VSS(VSS),.VDD(VDD),.Y(g2137),.A(g760),.B(g1638));
  AND2 AND2_41(.VSS(VSS),.VDD(VDD),.Y(g2138),.A(g1639),.B(g809));
  AND2 AND2_42(.VSS(VSS),.VDD(VDD),.Y(g2142),.A(g1793),.B(g1777));
  AND2 AND2_43(.VSS(VSS),.VDD(VDD),.Y(g2156),.A(g815),.B(g1642));
  AND2 AND2_44(.VSS(VSS),.VDD(VDD),.Y(g2160),.A(g1624),.B(g929));
  AND2 AND2_45(.VSS(VSS),.VDD(VDD),.Y(g2166),.A(g1633),.B(g161));
  AND2 AND2_46(.VSS(VSS),.VDD(VDD),.Y(g2255),.A(g1706),.B(g736));
  AND2 AND2_47(.VSS(VSS),.VDD(VDD),.Y(g2267),.A(g1716),.B(g791));
  AND3 AND3_4(.VSS(VSS),.VDD(VDD),.Y(g2292),.A(g1706),.B(g736),.C(g743));
  AND3 AND3_5(.VSS(VSS),.VDD(VDD),.Y(g2294),.A(g1716),.B(g791),.C(g798));
  AND2 AND2_48(.VSS(VSS),.VDD(VDD),.Y(g2323),.A(g471),.B(g1358));
  AND2 AND2_49(.VSS(VSS),.VDD(VDD),.Y(g2339),.A(g1603),.B(g197));
  AND2 AND2_50(.VSS(VSS),.VDD(VDD),.Y(g2340),.A(g1398),.B(g1387));
  AND2 AND2_51(.VSS(VSS),.VDD(VDD),.Y(g2356),.A(g1603),.B(g269));
  AND2 AND2_52(.VSS(VSS),.VDD(VDD),.Y(g2419),.A(g1808),.B(g54));
  AND2 AND2_53(.VSS(VSS),.VDD(VDD),.Y(g2551),.A(g715),.B(g1826));
  AND4 AND4_3(.VSS(VSS),.VDD(VDD),.Y(g2577),.A(g1743),.B(g1797),.C(g1793),.D(g1138));
  AND2 AND2_54(.VSS(VSS),.VDD(VDD),.Y(g2659),.A(g1686),.B(g2296));
  AND2 AND2_55(.VSS(VSS),.VDD(VDD),.Y(g2670),.A(g2029),.B(g1503));
  AND2 AND2_56(.VSS(VSS),.VDD(VDD),.Y(g2671),.A(g2263),.B(g2296));
  AND2 AND2_57(.VSS(VSS),.VDD(VDD),.Y(g2685),.A(g2370),.B(g1887));
  AND2 AND2_58(.VSS(VSS),.VDD(VDD),.Y(g2699),.A(g2397),.B(g1905));
  AND2 AND2_59(.VSS(VSS),.VDD(VDD),.Y(g2700),.A(g2370),.B(g1908));
  AND2 AND2_60(.VSS(VSS),.VDD(VDD),.Y(g2720),.A(g2422),.B(g1919));
  AND2 AND2_61(.VSS(VSS),.VDD(VDD),.Y(g2721),.A(g2397),.B(g1922));
  AND2 AND2_62(.VSS(VSS),.VDD(VDD),.Y(g2732),.A(g2449),.B(g1940));
  AND2 AND2_63(.VSS(VSS),.VDD(VDD),.Y(g2733),.A(g2422),.B(g1943));
  AND2 AND2_64(.VSS(VSS),.VDD(VDD),.Y(g2746),.A(g2473),.B(g1954));
  AND2 AND2_65(.VSS(VSS),.VDD(VDD),.Y(g2747),.A(g2449),.B(g1957));
  AND2 AND2_66(.VSS(VSS),.VDD(VDD),.Y(g2758),.A(g2497),.B(g1963));
  AND2 AND2_67(.VSS(VSS),.VDD(VDD),.Y(g2759),.A(g2473),.B(g1966));
  AND2 AND2_68(.VSS(VSS),.VDD(VDD),.Y(g2770),.A(g2518),.B(g1972));
  AND2 AND2_69(.VSS(VSS),.VDD(VDD),.Y(g2771),.A(g2497),.B(g1975));
  AND2 AND2_70(.VSS(VSS),.VDD(VDD),.Y(g2781),.A(g2544),.B(g1982));
  AND2 AND2_71(.VSS(VSS),.VDD(VDD),.Y(g2782),.A(g2518),.B(g1985));
  AND2 AND2_72(.VSS(VSS),.VDD(VDD),.Y(g2793),.A(g2568),.B(g1991));
  AND2 AND2_73(.VSS(VSS),.VDD(VDD),.Y(g2794),.A(g2544),.B(g1994));
  AND2 AND2_74(.VSS(VSS),.VDD(VDD),.Y(g2807),.A(g2568),.B(g2001));
  AND2 AND2_75(.VSS(VSS),.VDD(VDD),.Y(g2808),.A(g2009),.B(g1581));
  AND2 AND2_76(.VSS(VSS),.VDD(VDD),.Y(g2821),.A(g1890),.B(g910));
  AND3 AND3_6(.VSS(VSS),.VDD(VDD),.Y(I4040),.A(g1279),.B(g2025),.C(g1267));
  AND4 AND4_4(.VSS(VSS),.VDD(VDD),.Y(g2834),.A(g1263),.B(g1257),.C(g1270),.D(I4040));
  AND2 AND2_77(.VSS(VSS),.VDD(VDD),.Y(g2846),.A(g619),.B(g2015));
  AND2 AND2_78(.VSS(VSS),.VDD(VDD),.Y(g2850),.A(g2018),.B(g1255));
  AND2 AND2_79(.VSS(VSS),.VDD(VDD),.Y(g2853),.A(g836),.B(g2021));
  AND2 AND2_80(.VSS(VSS),.VDD(VDD),.Y(g2859),.A(g2112),.B(g1649));
  AND2 AND2_81(.VSS(VSS),.VDD(VDD),.Y(g2860),.A(g710),.B(g2296));
  AND2 AND2_82(.VSS(VSS),.VDD(VDD),.Y(g2861),.A(g2120),.B(g1654));
  AND2 AND2_83(.VSS(VSS),.VDD(VDD),.Y(g2868),.A(g1316),.B(g1861));
  AND2 AND2_84(.VSS(VSS),.VDD(VDD),.Y(g2873),.A(g1845),.B(g1861));
  AND2 AND2_85(.VSS(VSS),.VDD(VDD),.Y(g2897),.A(g1030),.B(g2062));
  AND2 AND2_86(.VSS(VSS),.VDD(VDD),.Y(g2909),.A(g606),.B(g2092));
  AND2 AND2_87(.VSS(VSS),.VDD(VDD),.Y(g2916),.A(g1030),.B(g2113));
  AND2 AND2_88(.VSS(VSS),.VDD(VDD),.Y(g2935),.A(g2291),.B(g1788));
  AND2 AND2_89(.VSS(VSS),.VDD(VDD),.Y(g2937),.A(g2160),.B(g931));
  AND2 AND2_90(.VSS(VSS),.VDD(VDD),.Y(g2941),.A(g2166),.B(g170));
  AND2 AND2_91(.VSS(VSS),.VDD(VDD),.Y(g2948),.A(g2137),.B(g1595));
  AND2 AND2_92(.VSS(VSS),.VDD(VDD),.Y(g2949),.A(g830),.B(g1861));
  AND2 AND2_93(.VSS(VSS),.VDD(VDD),.Y(g2950),.A(g2156),.B(g1612));
  AND2 AND2_94(.VSS(VSS),.VDD(VDD),.Y(g2953),.A(g2381),.B(g293));
  AND2 AND2_95(.VSS(VSS),.VDD(VDD),.Y(g2955),.A(g2381),.B(g297));
  AND2 AND2_96(.VSS(VSS),.VDD(VDD),.Y(g3089),.A(g212),.B(g2336));
  AND2 AND2_97(.VSS(VSS),.VDD(VDD),.Y(g3099),.A(g218),.B(g2350));
  AND2 AND2_98(.VSS(VSS),.VDD(VDD),.Y(g3103),.A(g212),.B(g2353));
  AND2 AND2_99(.VSS(VSS),.VDD(VDD),.Y(g3113),.A(g224),.B(g2364));
  AND2 AND2_100(.VSS(VSS),.VDD(VDD),.Y(g3117),.A(g218),.B(g2367));
  AND2 AND2_101(.VSS(VSS),.VDD(VDD),.Y(g3122),.A(g2435),.B(g1394));
  AND2 AND2_102(.VSS(VSS),.VDD(VDD),.Y(g3123),.A(g230),.B(g2391));
  AND2 AND2_103(.VSS(VSS),.VDD(VDD),.Y(g3127),.A(g224),.B(g2394));
  AND2 AND2_104(.VSS(VSS),.VDD(VDD),.Y(g3132),.A(g2306),.B(g1206));
  AND2 AND2_105(.VSS(VSS),.VDD(VDD),.Y(g3133),.A(g236),.B(g2410));
  AND2 AND2_106(.VSS(VSS),.VDD(VDD),.Y(g3134),.A(g230),.B(g2413));
  AND2 AND2_107(.VSS(VSS),.VDD(VDD),.Y(g3135),.A(g2370),.B(g2416));
  AND2 AND2_108(.VSS(VSS),.VDD(VDD),.Y(g3143),.A(g242),.B(g2437));
  AND2 AND2_109(.VSS(VSS),.VDD(VDD),.Y(g3144),.A(g236),.B(g2440));
  AND2 AND2_110(.VSS(VSS),.VDD(VDD),.Y(g3145),.A(g2397),.B(g2443));
  AND2 AND2_111(.VSS(VSS),.VDD(VDD),.Y(g3146),.A(g2370),.B(g2446));
  AND2 AND2_112(.VSS(VSS),.VDD(VDD),.Y(g3147),.A(g2419),.B(g59));
  AND2 AND2_113(.VSS(VSS),.VDD(VDD),.Y(g3154),.A(g2039),.B(g1410));
  AND2 AND2_114(.VSS(VSS),.VDD(VDD),.Y(g3155),.A(g248),.B(g2461));
  AND2 AND2_115(.VSS(VSS),.VDD(VDD),.Y(g3156),.A(g242),.B(g2464));
  AND2 AND2_116(.VSS(VSS),.VDD(VDD),.Y(g3157),.A(g2422),.B(g2467));
  AND2 AND2_117(.VSS(VSS),.VDD(VDD),.Y(g3161),.A(g2397),.B(g2470));
  AND2 AND2_118(.VSS(VSS),.VDD(VDD),.Y(g3166),.A(g2042),.B(g1233));
  AND2 AND2_119(.VSS(VSS),.VDD(VDD),.Y(g3167),.A(g1883),.B(g921));
  AND2 AND2_120(.VSS(VSS),.VDD(VDD),.Y(g3170),.A(g254),.B(g2485));
  AND2 AND2_121(.VSS(VSS),.VDD(VDD),.Y(g3171),.A(g248),.B(g2488));
  AND2 AND2_122(.VSS(VSS),.VDD(VDD),.Y(g3172),.A(g2449),.B(g2491));
  AND2 AND2_123(.VSS(VSS),.VDD(VDD),.Y(g3176),.A(g2422),.B(g2494));
  AND2 AND2_124(.VSS(VSS),.VDD(VDD),.Y(g3180),.A(g260),.B(g2506));
  AND2 AND2_125(.VSS(VSS),.VDD(VDD),.Y(g3181),.A(g254),.B(g2509));
  AND2 AND2_126(.VSS(VSS),.VDD(VDD),.Y(g3182),.A(g2473),.B(g2512));
  AND2 AND2_127(.VSS(VSS),.VDD(VDD),.Y(g3186),.A(g2449),.B(g2515));
  AND2 AND2_128(.VSS(VSS),.VDD(VDD),.Y(g3190),.A(g260),.B(g2535));
  AND2 AND2_129(.VSS(VSS),.VDD(VDD),.Y(g3191),.A(g2497),.B(g2538));
  AND2 AND2_130(.VSS(VSS),.VDD(VDD),.Y(g3195),.A(g2473),.B(g2541));
  AND2 AND2_131(.VSS(VSS),.VDD(VDD),.Y(g3203),.A(g2497),.B(g2565));
  AND2 AND2_132(.VSS(VSS),.VDD(VDD),.Y(g3208),.A(g895),.B(g2551));
  AND2 AND2_133(.VSS(VSS),.VDD(VDD),.Y(g3275),.A(g2172),.B(g2615));
  AND2 AND2_134(.VSS(VSS),.VDD(VDD),.Y(g3277),.A(g2174),.B(g2625));
  AND2 AND2_135(.VSS(VSS),.VDD(VDD),.Y(g3278),.A(g2175),.B(g2628));
  AND2 AND2_136(.VSS(VSS),.VDD(VDD),.Y(g3279),.A(g2599),.B(g2612));
  AND2 AND2_137(.VSS(VSS),.VDD(VDD),.Y(g3280),.A(g2177),.B(g2637));
  AND2 AND2_138(.VSS(VSS),.VDD(VDD),.Y(g3281),.A(g2178),.B(g2640));
  AND2 AND2_139(.VSS(VSS),.VDD(VDD),.Y(g3282),.A(g131),.B(g2863));
  AND2 AND2_140(.VSS(VSS),.VDD(VDD),.Y(g3283),.A(g2609),.B(g2622));
  AND2 AND2_141(.VSS(VSS),.VDD(VDD),.Y(g3285),.A(g2195),.B(g2653));
  AND2 AND2_142(.VSS(VSS),.VDD(VDD),.Y(g3286),.A(g2196),.B(g2656));
  AND2 AND2_143(.VSS(VSS),.VDD(VDD),.Y(g3287),.A(g135),.B(g2865));
  AND2 AND2_144(.VSS(VSS),.VDD(VDD),.Y(g3288),.A(g2631),.B(g2634));
  AND2 AND2_145(.VSS(VSS),.VDD(VDD),.Y(g3290),.A(g2213),.B(g2664));
  AND2 AND2_146(.VSS(VSS),.VDD(VDD),.Y(g3292),.A(g2214),.B(g2667));
  AND2 AND2_147(.VSS(VSS),.VDD(VDD),.Y(g3293),.A(g212),.B(g2864));
  AND2 AND2_148(.VSS(VSS),.VDD(VDD),.Y(g3294),.A(g139),.B(g2870));
  AND2 AND2_149(.VSS(VSS),.VDD(VDD),.Y(g3295),.A(g2660),.B(g2647));
  AND2 AND2_150(.VSS(VSS),.VDD(VDD),.Y(g3296),.A(g3054),.B(g2650));
  AND2 AND2_151(.VSS(VSS),.VDD(VDD),.Y(g3298),.A(g2231),.B(g2679));
  AND2 AND2_152(.VSS(VSS),.VDD(VDD),.Y(g3300),.A(g2232),.B(g2682));
  AND2 AND2_153(.VSS(VSS),.VDD(VDD),.Y(g3301),.A(g218),.B(g2866));
  AND2 AND2_154(.VSS(VSS),.VDD(VDD),.Y(g3302),.A(g212),.B(g2867));
  AND2 AND2_155(.VSS(VSS),.VDD(VDD),.Y(g3303),.A(g2722),.B(g2890));
  AND2 AND2_156(.VSS(VSS),.VDD(VDD),.Y(g3304),.A(g2857),.B(g1513));
  AND2 AND2_157(.VSS(VSS),.VDD(VDD),.Y(g3305),.A(g2960),.B(g2296));
  AND2 AND2_158(.VSS(VSS),.VDD(VDD),.Y(g3307),.A(g2242),.B(g2692));
  AND2 AND2_159(.VSS(VSS),.VDD(VDD),.Y(g3309),.A(g2243),.B(g2695));
  AND2 AND2_160(.VSS(VSS),.VDD(VDD),.Y(g3310),.A(g224),.B(g2871));
  AND2 AND2_161(.VSS(VSS),.VDD(VDD),.Y(g3311),.A(g218),.B(g2872));
  AND2 AND2_162(.VSS(VSS),.VDD(VDD),.Y(g3315),.A(g2701),.B(g1875));
  AND2 AND2_163(.VSS(VSS),.VDD(VDD),.Y(g3316),.A(g2748),.B(g2894));
  AND2 AND2_164(.VSS(VSS),.VDD(VDD),.Y(g3317),.A(g2722),.B(g2895));
  AND2 AND2_165(.VSS(VSS),.VDD(VDD),.Y(g3319),.A(g2688),.B(g2675));
  AND2 AND2_166(.VSS(VSS),.VDD(VDD),.Y(g3321),.A(g2252),.B(g2713));
  AND2 AND2_167(.VSS(VSS),.VDD(VDD),.Y(g3323),.A(g2253),.B(g2716));
  AND2 AND2_168(.VSS(VSS),.VDD(VDD),.Y(g3324),.A(g230),.B(g2875));
  AND2 AND2_169(.VSS(VSS),.VDD(VDD),.Y(g3325),.A(g224),.B(g2876));
  AND2 AND2_170(.VSS(VSS),.VDD(VDD),.Y(g3326),.A(g2734),.B(g1891));
  AND2 AND2_171(.VSS(VSS),.VDD(VDD),.Y(g3327),.A(g2772),.B(g2906));
  AND2 AND2_172(.VSS(VSS),.VDD(VDD),.Y(g3328),.A(g2701),.B(g1894));
  AND2 AND2_173(.VSS(VSS),.VDD(VDD),.Y(g3329),.A(g2748),.B(g2907));
  AND2 AND2_174(.VSS(VSS),.VDD(VDD),.Y(g3333),.A(g2264),.B(g2728));
  AND2 AND2_175(.VSS(VSS),.VDD(VDD),.Y(g3334),.A(g236),.B(g2883));
  AND2 AND2_176(.VSS(VSS),.VDD(VDD),.Y(g3335),.A(g230),.B(g2884));
  AND2 AND2_177(.VSS(VSS),.VDD(VDD),.Y(g3336),.A(g2760),.B(g1911));
  AND2 AND2_178(.VSS(VSS),.VDD(VDD),.Y(g3337),.A(g2796),.B(g2913));
  AND2 AND2_179(.VSS(VSS),.VDD(VDD),.Y(g3338),.A(g3162),.B(g2914));
  AND2 AND2_180(.VSS(VSS),.VDD(VDD),.Y(g3339),.A(g2734),.B(g1914));
  AND2 AND2_181(.VSS(VSS),.VDD(VDD),.Y(g3340),.A(g2772),.B(g2915));
  AND2 AND2_182(.VSS(VSS),.VDD(VDD),.Y(g3341),.A(g2998),.B(g2709));
  AND2 AND2_183(.VSS(VSS),.VDD(VDD),.Y(g3344),.A(g242),.B(g2885));
  AND2 AND2_184(.VSS(VSS),.VDD(VDD),.Y(g3345),.A(g236),.B(g2886));
  AND2 AND2_185(.VSS(VSS),.VDD(VDD),.Y(g3349),.A(g2783),.B(g1925));
  AND2 AND2_186(.VSS(VSS),.VDD(VDD),.Y(g3350),.A(g3150),.B(g1928));
  AND2 AND2_187(.VSS(VSS),.VDD(VDD),.Y(g3351),.A(g2760),.B(g1931));
  AND2 AND2_188(.VSS(VSS),.VDD(VDD),.Y(g3352),.A(g2796),.B(g2920));
  AND2 AND2_189(.VSS(VSS),.VDD(VDD),.Y(g3353),.A(g3162),.B(g2921));
  AND2 AND2_190(.VSS(VSS),.VDD(VDD),.Y(g3356),.A(g248),.B(g2888));
  AND2 AND2_191(.VSS(VSS),.VDD(VDD),.Y(g3357),.A(g242),.B(g2889));
  AND2 AND2_192(.VSS(VSS),.VDD(VDD),.Y(g3358),.A(g2842),.B(g1369));
  AND2 AND2_193(.VSS(VSS),.VDD(VDD),.Y(g3359),.A(g2822),.B(g2922));
  AND2 AND2_194(.VSS(VSS),.VDD(VDD),.Y(g3360),.A(g2783),.B(g1947));
  AND2 AND2_195(.VSS(VSS),.VDD(VDD),.Y(g3361),.A(g3150),.B(g1950));
  AND2 AND2_196(.VSS(VSS),.VDD(VDD),.Y(g3362),.A(g3031),.B(g2740));
  AND2 AND2_197(.VSS(VSS),.VDD(VDD),.Y(g3365),.A(g254),.B(g2892));
  AND2 AND2_198(.VSS(VSS),.VDD(VDD),.Y(g3366),.A(g248),.B(g2893));
  AND2 AND2_199(.VSS(VSS),.VDD(VDD),.Y(g3367),.A(g2809),.B(g1960));
  AND2 AND2_200(.VSS(VSS),.VDD(VDD),.Y(g3368),.A(g2822),.B(g2923));
  AND2 AND2_201(.VSS(VSS),.VDD(VDD),.Y(g3371),.A(g260),.B(g2904));
  AND2 AND2_202(.VSS(VSS),.VDD(VDD),.Y(g3372),.A(g254),.B(g2905));
  AND2 AND2_203(.VSS(VSS),.VDD(VDD),.Y(g3373),.A(g3118),.B(g2927));
  AND2 AND2_204(.VSS(VSS),.VDD(VDD),.Y(g3374),.A(g2809),.B(g1969));
  AND2 AND2_205(.VSS(VSS),.VDD(VDD),.Y(g3375),.A(g260),.B(g2912));
  AND2 AND2_206(.VSS(VSS),.VDD(VDD),.Y(g3376),.A(g3104),.B(g1979));
  AND2 AND2_207(.VSS(VSS),.VDD(VDD),.Y(g3377),.A(g3118),.B(g2931));
  AND2 AND2_208(.VSS(VSS),.VDD(VDD),.Y(g3378),.A(g3136),.B(g2932));
  AND2 AND2_209(.VSS(VSS),.VDD(VDD),.Y(g3379),.A(g3104),.B(g1988));
  AND2 AND2_210(.VSS(VSS),.VDD(VDD),.Y(g3381),.A(g3128),.B(g1998));
  AND2 AND2_211(.VSS(VSS),.VDD(VDD),.Y(g3382),.A(g3136),.B(g2934));
  AND2 AND2_212(.VSS(VSS),.VDD(VDD),.Y(g3383),.A(g3128),.B(g2004));
  AND2 AND2_213(.VSS(VSS),.VDD(VDD),.Y(g3421),.A(g622),.B(g2846));
  AND2 AND2_214(.VSS(VSS),.VDD(VDD),.Y(g3425),.A(g2296),.B(g3208));
  AND3 AND3_7(.VSS(VSS),.VDD(VDD),.Y(g3433),.A(g1359),.B(g2831),.C(g905));
  AND2 AND2_215(.VSS(VSS),.VDD(VDD),.Y(g3434),.A(g2850),.B(g857));
  AND2 AND2_216(.VSS(VSS),.VDD(VDD),.Y(g3437),.A(g837),.B(g2853));
  AND2 AND2_217(.VSS(VSS),.VDD(VDD),.Y(g3449),.A(g128),.B(g2946));
  AND2 AND2_218(.VSS(VSS),.VDD(VDD),.Y(g3454),.A(g2933),.B(g1660));
  AND2 AND2_219(.VSS(VSS),.VDD(VDD),.Y(g3464),.A(g341),.B(g2956));
  AND2 AND2_220(.VSS(VSS),.VDD(VDD),.Y(g3479),.A(g345),.B(g2957));
  AND2 AND2_221(.VSS(VSS),.VDD(VDD),.Y(g3484),.A(g349),.B(g2958));
  AND2 AND2_222(.VSS(VSS),.VDD(VDD),.Y(g3489),.A(g2607),.B(g1861));
  AND2 AND2_223(.VSS(VSS),.VDD(VDD),.Y(g3490),.A(g353),.B(g2959));
  AND2 AND2_224(.VSS(VSS),.VDD(VDD),.Y(g3499),.A(g357),.B(g2961));
  AND2 AND2_225(.VSS(VSS),.VDD(VDD),.Y(g3505),.A(g2924),.B(g1749));
  AND2 AND2_226(.VSS(VSS),.VDD(VDD),.Y(g3512),.A(g2928),.B(g1764));
  AND2 AND2_227(.VSS(VSS),.VDD(VDD),.Y(g3522),.A(g646),.B(g2909));
  AND2 AND2_228(.VSS(VSS),.VDD(VDD),.Y(g3551),.A(g2937),.B(g938));
  AND2 AND2_229(.VSS(VSS),.VDD(VDD),.Y(g3554),.A(g2941),.B(g179));
  AND2 AND2_230(.VSS(VSS),.VDD(VDD),.Y(g3558),.A(g338),.B(g3199));
  AND2 AND2_231(.VSS(VSS),.VDD(VDD),.Y(g3602),.A(g2688),.B(g2663));
  AND2 AND2_232(.VSS(VSS),.VDD(VDD),.Y(g3603),.A(g2370),.B(g3019));
  AND2 AND2_233(.VSS(VSS),.VDD(VDD),.Y(g3608),.A(g2599),.B(g2308));
  AND2 AND2_234(.VSS(VSS),.VDD(VDD),.Y(g3609),.A(g2706),.B(g2678));
  AND2 AND2_235(.VSS(VSS),.VDD(VDD),.Y(g3610),.A(g2397),.B(g3034));
  AND2 AND2_236(.VSS(VSS),.VDD(VDD),.Y(g3611),.A(g2370),.B(g3037));
  AND2 AND2_237(.VSS(VSS),.VDD(VDD),.Y(g3613),.A(g2604),.B(g2312));
  AND2 AND2_238(.VSS(VSS),.VDD(VDD),.Y(g3614),.A(g2998),.B(g2691));
  AND2 AND2_239(.VSS(VSS),.VDD(VDD),.Y(g3615),.A(g2422),.B(g3046));
  AND2 AND2_240(.VSS(VSS),.VDD(VDD),.Y(g3616),.A(g2397),.B(g3049));
  AND2 AND2_241(.VSS(VSS),.VDD(VDD),.Y(g3617),.A(g2609),.B(g2317));
  AND2 AND2_242(.VSS(VSS),.VDD(VDD),.Y(g3618),.A(g3016),.B(g2712));
  AND2 AND2_243(.VSS(VSS),.VDD(VDD),.Y(g3619),.A(g2449),.B(g3057));
  AND2 AND2_244(.VSS(VSS),.VDD(VDD),.Y(g3620),.A(g2422),.B(g3060));
  AND2 AND2_245(.VSS(VSS),.VDD(VDD),.Y(g3625),.A(g2619),.B(g2320));
  AND2 AND2_246(.VSS(VSS),.VDD(VDD),.Y(g3626),.A(g3031),.B(g2727));
  AND2 AND2_247(.VSS(VSS),.VDD(VDD),.Y(g3627),.A(g2473),.B(g3067));
  AND2 AND2_248(.VSS(VSS),.VDD(VDD),.Y(g3628),.A(g2449),.B(g3070));
  AND2 AND2_249(.VSS(VSS),.VDD(VDD),.Y(g3629),.A(g2809),.B(g2738));
  AND2 AND2_250(.VSS(VSS),.VDD(VDD),.Y(g3630),.A(g3167),.B(g1756));
  AND2 AND2_251(.VSS(VSS),.VDD(VDD),.Y(g3631),.A(g2631),.B(g2324));
  AND2 AND2_252(.VSS(VSS),.VDD(VDD),.Y(g3632),.A(g3043),.B(g2743));
  AND2 AND2_253(.VSS(VSS),.VDD(VDD),.Y(g3633),.A(g2497),.B(g3076));
  AND2 AND2_254(.VSS(VSS),.VDD(VDD),.Y(g3634),.A(g2179),.B(g2744));
  AND2 AND2_255(.VSS(VSS),.VDD(VDD),.Y(g3635),.A(g2473),.B(g3079));
  AND2 AND2_256(.VSS(VSS),.VDD(VDD),.Y(g3636),.A(g2701),.B(g2327));
  AND2 AND2_257(.VSS(VSS),.VDD(VDD),.Y(g3637),.A(g2822),.B(g2752));
  AND2 AND2_258(.VSS(VSS),.VDD(VDD),.Y(g3641),.A(g2644),.B(g2333));
  AND2 AND2_259(.VSS(VSS),.VDD(VDD),.Y(g3642),.A(g3054),.B(g2754));
  AND2 AND2_260(.VSS(VSS),.VDD(VDD),.Y(g3643),.A(g2518),.B(g3086));
  AND2 AND2_261(.VSS(VSS),.VDD(VDD),.Y(g3644),.A(g2197),.B(g2755));
  AND2 AND2_262(.VSS(VSS),.VDD(VDD),.Y(g3645),.A(g2497),.B(g3090));
  AND2 AND2_263(.VSS(VSS),.VDD(VDD),.Y(g3646),.A(g2179),.B(g2756));
  AND2 AND2_264(.VSS(VSS),.VDD(VDD),.Y(g3648),.A(g2722),.B(g2343));
  AND2 AND2_265(.VSS(VSS),.VDD(VDD),.Y(g3649),.A(g3104),.B(g2764));
  AND2 AND2_266(.VSS(VSS),.VDD(VDD),.Y(g3650),.A(g2660),.B(g2347));
  AND2 AND2_267(.VSS(VSS),.VDD(VDD),.Y(g3651),.A(g3064),.B(g2766));
  AND2 AND2_268(.VSS(VSS),.VDD(VDD),.Y(g3652),.A(g2544),.B(g3096));
  AND2 AND2_269(.VSS(VSS),.VDD(VDD),.Y(g3653),.A(g2215),.B(g2767));
  AND2 AND2_270(.VSS(VSS),.VDD(VDD),.Y(g3654),.A(g2518),.B(g3100));
  AND2 AND2_271(.VSS(VSS),.VDD(VDD),.Y(g3655),.A(g2197),.B(g2768));
  AND2 AND2_272(.VSS(VSS),.VDD(VDD),.Y(g3657),.A(g2734),.B(g2357));
  AND2 AND2_273(.VSS(VSS),.VDD(VDD),.Y(g3658),.A(g3118),.B(g2776));
  AND2 AND2_274(.VSS(VSS),.VDD(VDD),.Y(g3659),.A(g2672),.B(g2361));
  AND2 AND2_275(.VSS(VSS),.VDD(VDD),.Y(g3660),.A(g2568),.B(g3110));
  AND2 AND2_276(.VSS(VSS),.VDD(VDD),.Y(g3661),.A(g2234),.B(g2778));
  AND2 AND2_277(.VSS(VSS),.VDD(VDD),.Y(g3662),.A(g2544),.B(g3114));
  AND2 AND2_278(.VSS(VSS),.VDD(VDD),.Y(g3663),.A(g2215),.B(g2779));
  AND2 AND2_279(.VSS(VSS),.VDD(VDD),.Y(g3665),.A(g2748),.B(g2378));
  AND2 AND2_280(.VSS(VSS),.VDD(VDD),.Y(g3666),.A(g3128),.B(g2787));
  AND2 AND2_281(.VSS(VSS),.VDD(VDD),.Y(g3667),.A(g2245),.B(g2789));
  AND2 AND2_282(.VSS(VSS),.VDD(VDD),.Y(g3668),.A(g2568),.B(g3124));
  AND2 AND2_283(.VSS(VSS),.VDD(VDD),.Y(g3669),.A(g2234),.B(g2790));
  AND2 AND2_284(.VSS(VSS),.VDD(VDD),.Y(g3670),.A(g2234),.B(g2792));
  AND2 AND2_285(.VSS(VSS),.VDD(VDD),.Y(g3671),.A(g2760),.B(g2405));
  AND2 AND2_286(.VSS(VSS),.VDD(VDD),.Y(g3672),.A(g3136),.B(g2800));
  AND2 AND2_287(.VSS(VSS),.VDD(VDD),.Y(g3678),.A(g2256),.B(g2802));
  AND2 AND2_288(.VSS(VSS),.VDD(VDD),.Y(g3679),.A(g2245),.B(g2803));
  AND2 AND2_289(.VSS(VSS),.VDD(VDD),.Y(g3680),.A(g2245),.B(g2805));
  AND2 AND2_290(.VSS(VSS),.VDD(VDD),.Y(g3681),.A(g2234),.B(g2806));
  AND2 AND2_291(.VSS(VSS),.VDD(VDD),.Y(g3682),.A(g2772),.B(g2430));
  AND2 AND2_292(.VSS(VSS),.VDD(VDD),.Y(g3683),.A(g3150),.B(g2813));
  AND2 AND2_293(.VSS(VSS),.VDD(VDD),.Y(g3684),.A(g2268),.B(g2817));
  AND2 AND2_294(.VSS(VSS),.VDD(VDD),.Y(g3685),.A(g2256),.B(g2818));
  AND2 AND2_295(.VSS(VSS),.VDD(VDD),.Y(g3686),.A(g2256),.B(g2819));
  AND2 AND2_296(.VSS(VSS),.VDD(VDD),.Y(g3687),.A(g2245),.B(g2820));
  AND2 AND2_297(.VSS(VSS),.VDD(VDD),.Y(g3688),.A(g2783),.B(g2457));
  AND2 AND2_298(.VSS(VSS),.VDD(VDD),.Y(g3689),.A(g3162),.B(g2826));
  AND2 AND2_299(.VSS(VSS),.VDD(VDD),.Y(g3690),.A(g2276),.B(g2827));
  AND2 AND2_300(.VSS(VSS),.VDD(VDD),.Y(g3691),.A(g2268),.B(g2828));
  AND2 AND2_301(.VSS(VSS),.VDD(VDD),.Y(g3692),.A(g2268),.B(g2829));
  AND2 AND2_302(.VSS(VSS),.VDD(VDD),.Y(g3693),.A(g2256),.B(g2830));
  AND2 AND2_303(.VSS(VSS),.VDD(VDD),.Y(g3694),.A(g3147),.B(g64));
  AND2 AND2_304(.VSS(VSS),.VDD(VDD),.Y(g3697),.A(g2796),.B(g2481));
  AND2 AND2_305(.VSS(VSS),.VDD(VDD),.Y(g3698),.A(g2284),.B(g2835));
  AND2 AND2_306(.VSS(VSS),.VDD(VDD),.Y(g3699),.A(g2276),.B(g2836));
  AND2 AND2_307(.VSS(VSS),.VDD(VDD),.Y(g3700),.A(g2276),.B(g2837));
  AND2 AND2_308(.VSS(VSS),.VDD(VDD),.Y(g3701),.A(g2268),.B(g2838));
  AND2 AND2_309(.VSS(VSS),.VDD(VDD),.Y(g3702),.A(g2284),.B(g2839));
  AND2 AND2_310(.VSS(VSS),.VDD(VDD),.Y(g3703),.A(g2284),.B(g2840));
  AND2 AND2_311(.VSS(VSS),.VDD(VDD),.Y(g3704),.A(g2276),.B(g2841));
  AND2 AND2_312(.VSS(VSS),.VDD(VDD),.Y(g3709),.A(g2284),.B(g2845));
  AND3 AND3_8(.VSS(VSS),.VDD(VDD),.Y(g3718),.A(g1743),.B(g3140),.C(g1157));
  AND2 AND2_313(.VSS(VSS),.VDD(VDD),.Y(g3724),.A(g117),.B(g3251));
  AND2 AND2_314(.VSS(VSS),.VDD(VDD),.Y(g3725),.A(g118),.B(g3251));
  AND2 AND2_315(.VSS(VSS),.VDD(VDD),.Y(g3726),.A(g119),.B(g3251));
  AND2 AND2_316(.VSS(VSS),.VDD(VDD),.Y(g3727),.A(g122),.B(g3251));
  AND2 AND2_317(.VSS(VSS),.VDD(VDD),.Y(g3728),.A(g326),.B(g3441));
  AND2 AND2_318(.VSS(VSS),.VDD(VDD),.Y(g3729),.A(g327),.B(g3441));
  AND2 AND2_319(.VSS(VSS),.VDD(VDD),.Y(g3730),.A(g328),.B(g3441));
  AND2 AND2_320(.VSS(VSS),.VDD(VDD),.Y(g3731),.A(g331),.B(g3441));
  AND2 AND2_321(.VSS(VSS),.VDD(VDD),.Y(g3755),.A(g2604),.B(g3481));
  AND2 AND2_322(.VSS(VSS),.VDD(VDD),.Y(g3757),.A(g2619),.B(g3487));
  AND2 AND2_323(.VSS(VSS),.VDD(VDD),.Y(g3758),.A(g545),.B(g3461));
  AND2 AND2_324(.VSS(VSS),.VDD(VDD),.Y(g3759),.A(g2644),.B(g3498));
  AND2 AND2_325(.VSS(VSS),.VDD(VDD),.Y(g3760),.A(g548),.B(g3465));
  AND2 AND2_326(.VSS(VSS),.VDD(VDD),.Y(g3762),.A(g2672),.B(g3500));
  AND2 AND2_327(.VSS(VSS),.VDD(VDD),.Y(g3763),.A(g3064),.B(g3501));
  AND2 AND2_328(.VSS(VSS),.VDD(VDD),.Y(g3764),.A(g551),.B(g3480));
  AND2 AND2_329(.VSS(VSS),.VDD(VDD),.Y(g3765),.A(g554),.B(g3485));
  AND2 AND2_330(.VSS(VSS),.VDD(VDD),.Y(g3767),.A(g2706),.B(g3504));
  AND2 AND2_331(.VSS(VSS),.VDD(VDD),.Y(g3768),.A(g3448),.B(g1528));
  AND2 AND2_332(.VSS(VSS),.VDD(VDD),.Y(g3774),.A(g3016),.B(g3510));
  AND2 AND2_333(.VSS(VSS),.VDD(VDD),.Y(g3780),.A(g3043),.B(g3519));
  AND2 AND2_334(.VSS(VSS),.VDD(VDD),.Y(g3784),.A(g114),.B(g3251));
  AND2 AND2_335(.VSS(VSS),.VDD(VDD),.Y(g3806),.A(g3384),.B(g2024));
  AND2 AND2_336(.VSS(VSS),.VDD(VDD),.Y(g3810),.A(g625),.B(g3421));
  AND2 AND2_337(.VSS(VSS),.VDD(VDD),.Y(g3814),.A(g913),.B(g3546));
  AND2 AND2_338(.VSS(VSS),.VDD(VDD),.Y(g3816),.A(g3434),.B(g861));
  AND2 AND2_339(.VSS(VSS),.VDD(VDD),.Y(g3819),.A(g964),.B(g3437));
  AND2 AND2_340(.VSS(VSS),.VDD(VDD),.Y(g3831),.A(g2330),.B(g3425));
  AND3 AND3_9(.VSS(VSS),.VDD(VDD),.Y(g3843),.A(g2856),.B(g945),.C(g3533));
  AND2 AND2_341(.VSS(VSS),.VDD(VDD),.Y(g3844),.A(g3540),.B(g1665));
  AND2 AND2_342(.VSS(VSS),.VDD(VDD),.Y(g3887),.A(g3276),.B(g1861));
  AND2 AND2_343(.VSS(VSS),.VDD(VDD),.Y(g3899),.A(g323),.B(g3441));
  AND2 AND2_344(.VSS(VSS),.VDD(VDD),.Y(g3907),.A(g650),.B(g3522));
  AND2 AND2_345(.VSS(VSS),.VDD(VDD),.Y(g3910),.A(g3546),.B(g1049));
  AND2 AND2_346(.VSS(VSS),.VDD(VDD),.Y(g3924),.A(g3505),.B(g471));
  AND2 AND2_347(.VSS(VSS),.VDD(VDD),.Y(g3928),.A(g3512),.B(g478));
  AND2 AND2_348(.VSS(VSS),.VDD(VDD),.Y(g3936),.A(g3551),.B(g940));
  AND2 AND2_349(.VSS(VSS),.VDD(VDD),.Y(g3953),.A(g3554),.B(g188));
  AND3 AND3_10(.VSS(VSS),.VDD(VDD),.Y(g3997),.A(g1250),.B(g3425),.C(g2849));
  AND2 AND2_350(.VSS(VSS),.VDD(VDD),.Y(g4015),.A(g445),.B(g3388));
  AND2 AND2_351(.VSS(VSS),.VDD(VDD),.Y(g4032),.A(g441),.B(g3388));
  AND2 AND2_352(.VSS(VSS),.VDD(VDD),.Y(g4033),.A(g426),.B(g3388));
  AND2 AND2_353(.VSS(VSS),.VDD(VDD),.Y(g4035),.A(g437),.B(g3388));
  AND2 AND2_354(.VSS(VSS),.VDD(VDD),.Y(g4037),.A(g2896),.B(g3388));
  AND2 AND2_355(.VSS(VSS),.VDD(VDD),.Y(g4038),.A(g430),.B(g3388));
  AND2 AND2_356(.VSS(VSS),.VDD(VDD),.Y(g4039),.A(g402),.B(g3388));
  AND2 AND2_357(.VSS(VSS),.VDD(VDD),.Y(g4041),.A(g461),.B(g3388));
  AND2 AND2_358(.VSS(VSS),.VDD(VDD),.Y(g4042),.A(g406),.B(g3388));
  AND2 AND2_359(.VSS(VSS),.VDD(VDD),.Y(g4043),.A(g457),.B(g3388));
  AND2 AND2_360(.VSS(VSS),.VDD(VDD),.Y(g4044),.A(g410),.B(g3388));
  AND2 AND2_361(.VSS(VSS),.VDD(VDD),.Y(g4045),.A(g3425),.B(g123));
  AND4 AND4_5(.VSS(VSS),.VDD(VDD),.Y(I5351),.A(g3511),.B(g3517),.C(g3520),.D(g3525));
  AND4 AND4_6(.VSS(VSS),.VDD(VDD),.Y(I5352),.A(g3529),.B(g3531),.C(g3535),.D(g3538));
  AND2 AND2_362(.VSS(VSS),.VDD(VDD),.Y(g4046),.A(I5351),.B(I5352));
  AND2 AND2_363(.VSS(VSS),.VDD(VDD),.Y(g4047),.A(g453),.B(g3388));
  AND2 AND2_364(.VSS(VSS),.VDD(VDD),.Y(g4048),.A(g414),.B(g3388));
  AND4 AND4_7(.VSS(VSS),.VDD(VDD),.Y(I5359),.A(g3518),.B(g3521),.C(g3526),.D(g3530));
  AND4 AND4_8(.VSS(VSS),.VDD(VDD),.Y(I5360),.A(g3532),.B(g3536),.C(g3539),.D(g3544));
  AND2 AND2_365(.VSS(VSS),.VDD(VDD),.Y(g4050),.A(I5359),.B(I5360));
  AND2 AND2_366(.VSS(VSS),.VDD(VDD),.Y(g4051),.A(g449),.B(g3388));
  AND2 AND2_367(.VSS(VSS),.VDD(VDD),.Y(g4052),.A(g418),.B(g3388));
  AND2 AND2_368(.VSS(VSS),.VDD(VDD),.Y(g4053),.A(g3387),.B(g1415));
  AND2 AND2_369(.VSS(VSS),.VDD(VDD),.Y(g4054),.A(g3694),.B(g69));
  AND2 AND2_370(.VSS(VSS),.VDD(VDD),.Y(g4057),.A(g422),.B(g3388));
  AND2 AND2_371(.VSS(VSS),.VDD(VDD),.Y(g4058),.A(g3424),.B(g1246));
  AND2 AND2_372(.VSS(VSS),.VDD(VDD),.Y(g4156),.A(g3926),.B(g2078));
  AND2 AND2_373(.VSS(VSS),.VDD(VDD),.Y(g4157),.A(g3830),.B(g1533));
  AND2 AND2_374(.VSS(VSS),.VDD(VDD),.Y(g4159),.A(g370),.B(g3890));
  AND2 AND2_375(.VSS(VSS),.VDD(VDD),.Y(g4160),.A(g3923),.B(g1345));
  AND2 AND2_376(.VSS(VSS),.VDD(VDD),.Y(g4161),.A(g3931),.B(g2087));
  AND2 AND2_377(.VSS(VSS),.VDD(VDD),.Y(g4163),.A(g374),.B(g3892));
  AND2 AND2_378(.VSS(VSS),.VDD(VDD),.Y(g4164),.A(g3958),.B(g2091));
  AND2 AND2_379(.VSS(VSS),.VDD(VDD),.Y(g4165),.A(g3927),.B(g1352));
  AND2 AND2_380(.VSS(VSS),.VDD(VDD),.Y(g4167),.A(g378),.B(g3898));
  AND2 AND2_381(.VSS(VSS),.VDD(VDD),.Y(g4168),.A(g3925),.B(g1355));
  AND2 AND2_382(.VSS(VSS),.VDD(VDD),.Y(g4169),.A(g3966),.B(g2099));
  AND2 AND2_383(.VSS(VSS),.VDD(VDD),.Y(g4170),.A(g382),.B(g3900));
  AND2 AND2_384(.VSS(VSS),.VDD(VDD),.Y(g4171),.A(g3956),.B(g2104));
  AND2 AND2_385(.VSS(VSS),.VDD(VDD),.Y(g4172),.A(g3930),.B(g1366));
  AND2 AND2_386(.VSS(VSS),.VDD(VDD),.Y(g4176),.A(g386),.B(g3901));
  AND2 AND2_387(.VSS(VSS),.VDD(VDD),.Y(g4177),.A(g3933),.B(g1372));
  AND2 AND2_388(.VSS(VSS),.VDD(VDD),.Y(g4178),.A(g3959),.B(g2110));
  AND2 AND2_389(.VSS(VSS),.VDD(VDD),.Y(g4179),.A(g390),.B(g3902));
  AND2 AND2_390(.VSS(VSS),.VDD(VDD),.Y(g4180),.A(g3929),.B(g2119));
  AND2 AND2_391(.VSS(VSS),.VDD(VDD),.Y(g4181),.A(g3939),.B(g1381));
  AND2 AND2_392(.VSS(VSS),.VDD(VDD),.Y(g4182),.A(g394),.B(g3904));
  AND2 AND2_393(.VSS(VSS),.VDD(VDD),.Y(g4183),.A(g3965),.B(g1391));
  AND2 AND2_394(.VSS(VSS),.VDD(VDD),.Y(g4184),.A(g3934),.B(g2136));
  AND2 AND2_395(.VSS(VSS),.VDD(VDD),.Y(g4185),.A(g398),.B(g3906));
  AND2 AND2_396(.VSS(VSS),.VDD(VDD),.Y(g4186),.A(g3973),.B(g1395));
  AND2 AND2_397(.VSS(VSS),.VDD(VDD),.Y(g4199),.A(g628),.B(g3810));
  AND2 AND2_398(.VSS(VSS),.VDD(VDD),.Y(g4209),.A(g3816),.B(g865));
  AND2 AND2_399(.VSS(VSS),.VDD(VDD),.Y(g4214),.A(g1822),.B(g4045));
  AND2 AND2_400(.VSS(VSS),.VDD(VDD),.Y(g4219),.A(g3911),.B(g1655));
  AND2 AND2_401(.VSS(VSS),.VDD(VDD),.Y(g4230),.A(g3756),.B(g1861));
  AND2 AND2_402(.VSS(VSS),.VDD(VDD),.Y(g4236),.A(g654),.B(g3907));
  AND3 AND3_11(.VSS(VSS),.VDD(VDD),.Y(g4244),.A(g1749),.B(g4004),.C(g1609));
  AND3 AND3_12(.VSS(VSS),.VDD(VDD),.Y(g4247),.A(g1764),.B(g4007),.C(g1628));
  AND2 AND2_403(.VSS(VSS),.VDD(VDD),.Y(g4253),.A(g1861),.B(g3819));
  AND3 AND3_13(.VSS(VSS),.VDD(VDD),.Y(g4271),.A(g2121),.B(g1749),.C(g4004));
  AND2 AND2_404(.VSS(VSS),.VDD(VDD),.Y(g4277),.A(g3936),.B(g942));
  AND3 AND3_14(.VSS(VSS),.VDD(VDD),.Y(g4280),.A(g2138),.B(g1764),.C(g4007));
  AND2 AND2_405(.VSS(VSS),.VDD(VDD),.Y(g4333),.A(g3964),.B(g3284));
  AND2 AND2_406(.VSS(VSS),.VDD(VDD),.Y(g4339),.A(g3971),.B(g3289));
  AND2 AND2_407(.VSS(VSS),.VDD(VDD),.Y(g4340),.A(g3972),.B(g3291));
  AND2 AND2_408(.VSS(VSS),.VDD(VDD),.Y(g4341),.A(g3977),.B(g3297));
  AND2 AND2_409(.VSS(VSS),.VDD(VDD),.Y(g4342),.A(g3978),.B(g3299));
  AND2 AND2_410(.VSS(VSS),.VDD(VDD),.Y(g4344),.A(g3981),.B(g3306));
  AND2 AND2_411(.VSS(VSS),.VDD(VDD),.Y(g4345),.A(g3982),.B(g3308));
  AND2 AND2_412(.VSS(VSS),.VDD(VDD),.Y(g4346),.A(g157),.B(g3773));
  AND2 AND2_413(.VSS(VSS),.VDD(VDD),.Y(g4347),.A(g3986),.B(g3320));
  AND2 AND2_414(.VSS(VSS),.VDD(VDD),.Y(g4348),.A(g3987),.B(g3322));
  AND2 AND2_415(.VSS(VSS),.VDD(VDD),.Y(g4349),.A(g441),.B(g3775));
  AND2 AND2_416(.VSS(VSS),.VDD(VDD),.Y(g4351),.A(g166),.B(g3776));
  AND2 AND2_417(.VSS(VSS),.VDD(VDD),.Y(g4352),.A(g3988),.B(g3331));
  AND2 AND2_418(.VSS(VSS),.VDD(VDD),.Y(g4353),.A(g3989),.B(g3332));
  AND2 AND2_419(.VSS(VSS),.VDD(VDD),.Y(g4354),.A(g437),.B(g3777));
  AND2 AND2_420(.VSS(VSS),.VDD(VDD),.Y(g4355),.A(g430),.B(g3778));
  AND2 AND2_421(.VSS(VSS),.VDD(VDD),.Y(g4356),.A(g175),.B(g3779));
  AND2 AND2_422(.VSS(VSS),.VDD(VDD),.Y(g4357),.A(g3990),.B(g3342));
  AND2 AND2_423(.VSS(VSS),.VDD(VDD),.Y(g4358),.A(g3991),.B(g3343));
  AND2 AND2_424(.VSS(VSS),.VDD(VDD),.Y(g4359),.A(g434),.B(g3782));
  AND2 AND2_425(.VSS(VSS),.VDD(VDD),.Y(g4360),.A(g184),.B(g3785));
  AND2 AND2_426(.VSS(VSS),.VDD(VDD),.Y(g4361),.A(g3995),.B(g3354));
  AND2 AND2_427(.VSS(VSS),.VDD(VDD),.Y(g4362),.A(g3996),.B(g3355));
  AND2 AND2_428(.VSS(VSS),.VDD(VDD),.Y(g4363),.A(g402),.B(g3786));
  AND2 AND2_429(.VSS(VSS),.VDD(VDD),.Y(g4367),.A(g193),.B(g3788));
  AND2 AND2_430(.VSS(VSS),.VDD(VDD),.Y(g4368),.A(g3998),.B(g3363));
  AND2 AND2_431(.VSS(VSS),.VDD(VDD),.Y(g4369),.A(g3999),.B(g3364));
  AND2 AND2_432(.VSS(VSS),.VDD(VDD),.Y(g4371),.A(g461),.B(g3789));
  AND2 AND2_433(.VSS(VSS),.VDD(VDD),.Y(g4372),.A(g406),.B(g3790));
  AND2 AND2_434(.VSS(VSS),.VDD(VDD),.Y(g4373),.A(g4001),.B(g3370));
  AND2 AND2_435(.VSS(VSS),.VDD(VDD),.Y(g4377),.A(g457),.B(g3791));
  AND2 AND2_436(.VSS(VSS),.VDD(VDD),.Y(g4378),.A(g410),.B(g3792));
  AND2 AND2_437(.VSS(VSS),.VDD(VDD),.Y(g4383),.A(g453),.B(g3796));
  AND2 AND2_438(.VSS(VSS),.VDD(VDD),.Y(g4384),.A(g414),.B(g3797));
  AND2 AND2_439(.VSS(VSS),.VDD(VDD),.Y(g4389),.A(g449),.B(g3798));
  AND2 AND2_440(.VSS(VSS),.VDD(VDD),.Y(g4390),.A(g418),.B(g3799));
  AND2 AND2_441(.VSS(VSS),.VDD(VDD),.Y(g4395),.A(g445),.B(g3800));
  AND2 AND2_442(.VSS(VSS),.VDD(VDD),.Y(g4396),.A(g422),.B(g3801));
  AND2 AND2_443(.VSS(VSS),.VDD(VDD),.Y(g4401),.A(g426),.B(g3802));
  AND2 AND2_444(.VSS(VSS),.VDD(VDD),.Y(g4407),.A(g4054),.B(g74));
  AND2 AND2_445(.VSS(VSS),.VDD(VDD),.Y(g4410),.A(g3903),.B(g1474));
  AND2 AND2_446(.VSS(VSS),.VDD(VDD),.Y(g4416),.A(g3905),.B(g1481));
  AND3 AND3_15(.VSS(VSS),.VDD(VDD),.Y(g4429),.A(g923),.B(g4253),.C(g2936));
  AND2 AND2_447(.VSS(VSS),.VDD(VDD),.Y(g4442),.A(g4239),.B(g2882));
  AND2 AND2_448(.VSS(VSS),.VDD(VDD),.Y(g4445),.A(g4235),.B(g1854));
  AND2 AND2_449(.VSS(VSS),.VDD(VDD),.Y(g4448),.A(g3815),.B(g4225));
  AND2 AND2_450(.VSS(VSS),.VDD(VDD),.Y(g4449),.A(g4266),.B(g2887));
  AND2 AND2_451(.VSS(VSS),.VDD(VDD),.Y(g4452),.A(g3820),.B(g4227));
  AND2 AND2_452(.VSS(VSS),.VDD(VDD),.Y(g4453),.A(g4238),.B(g1858));
  AND2 AND2_453(.VSS(VSS),.VDD(VDD),.Y(g4456),.A(g3829),.B(g4229));
  AND2 AND2_454(.VSS(VSS),.VDD(VDD),.Y(g4457),.A(g4261),.B(g2902));
  AND2 AND2_455(.VSS(VSS),.VDD(VDD),.Y(g4459),.A(g4245),.B(g1899));
  AND2 AND2_456(.VSS(VSS),.VDD(VDD),.Y(g4460),.A(g4218),.B(g1539));
  AND2 AND2_457(.VSS(VSS),.VDD(VDD),.Y(g4461),.A(g4241),.B(g2919));
  AND2 AND2_458(.VSS(VSS),.VDD(VDD),.Y(g4464),.A(g4272),.B(g1937));
  AND2 AND2_459(.VSS(VSS),.VDD(VDD),.Y(g4471),.A(g4253),.B(g332));
  AND2 AND2_460(.VSS(VSS),.VDD(VDD),.Y(g4486),.A(g716),.B(g4195));
  AND2 AND2_461(.VSS(VSS),.VDD(VDD),.Y(g4488),.A(g1633),.B(g4202));
  AND2 AND2_462(.VSS(VSS),.VDD(VDD),.Y(g4489),.A(g2166),.B(g4206));
  AND2 AND2_463(.VSS(VSS),.VDD(VDD),.Y(g4490),.A(g2941),.B(g4210));
  AND2 AND2_464(.VSS(VSS),.VDD(VDD),.Y(g4491),.A(g3554),.B(g4215));
  AND2 AND2_465(.VSS(VSS),.VDD(VDD),.Y(g4495),.A(g3913),.B(g4292));
  AND2 AND2_466(.VSS(VSS),.VDD(VDD),.Y(g4501),.A(g4250),.B(g1671));
  AND2 AND2_467(.VSS(VSS),.VDD(VDD),.Y(g4541),.A(g631),.B(g4199));
  AND2 AND2_468(.VSS(VSS),.VDD(VDD),.Y(g4580),.A(g706),.B(g4262));
  AND2 AND2_469(.VSS(VSS),.VDD(VDD),.Y(g4583),.A(g1808),.B(g4267));
  AND2 AND2_470(.VSS(VSS),.VDD(VDD),.Y(g4588),.A(g2419),.B(g4273));
  AND2 AND2_471(.VSS(VSS),.VDD(VDD),.Y(g4592),.A(g3147),.B(g4281));
  AND2 AND2_472(.VSS(VSS),.VDD(VDD),.Y(g4593),.A(g4277),.B(g947));
  AND2 AND2_473(.VSS(VSS),.VDD(VDD),.Y(g4597),.A(g3694),.B(g4286));
  AND2 AND2_474(.VSS(VSS),.VDD(VDD),.Y(g4598),.A(g1978),.B(g4253));
  AND2 AND2_475(.VSS(VSS),.VDD(VDD),.Y(g4600),.A(g4054),.B(g4289));
  AND2 AND2_476(.VSS(VSS),.VDD(VDD),.Y(g4602),.A(g4407),.B(g4293));
  AND3 AND3_16(.VSS(VSS),.VDD(VDD),.Y(g4611),.A(g3985),.B(g119),.C(g4300));
  AND2 AND2_477(.VSS(VSS),.VDD(VDD),.Y(g4616),.A(g4231),.B(g3761));
  AND2 AND2_478(.VSS(VSS),.VDD(VDD),.Y(g4621),.A(g3953),.B(g4364));
  AND2 AND2_479(.VSS(VSS),.VDD(VDD),.Y(g4648),.A(g4407),.B(g79));
  AND2 AND2_480(.VSS(VSS),.VDD(VDD),.Y(g4661),.A(g4637),.B(g4634));
  AND2 AND2_481(.VSS(VSS),.VDD(VDD),.Y(g4666),.A(g4630),.B(g4627));
  AND2 AND2_482(.VSS(VSS),.VDD(VDD),.Y(g4667),.A(g4653),.B(g4651));
  AND2 AND2_483(.VSS(VSS),.VDD(VDD),.Y(g4668),.A(g4642),.B(g4638));
  AND2 AND2_484(.VSS(VSS),.VDD(VDD),.Y(g4671),.A(g4645),.B(g4641));
  AND2 AND2_485(.VSS(VSS),.VDD(VDD),.Y(g4672),.A(g4635),.B(g4631));
  AND2 AND2_486(.VSS(VSS),.VDD(VDD),.Y(g4673),.A(g4656),.B(g4654));
  AND2 AND2_487(.VSS(VSS),.VDD(VDD),.Y(g4677),.A(g4652),.B(g4646));
  AND2 AND2_488(.VSS(VSS),.VDD(VDD),.Y(g4683),.A(g4585),.B(g2066));
  AND2 AND2_489(.VSS(VSS),.VDD(VDD),.Y(g4684),.A(g4584),.B(g1341));
  AND2 AND2_490(.VSS(VSS),.VDD(VDD),.Y(g4685),.A(g4591),.B(g2079));
  AND2 AND2_491(.VSS(VSS),.VDD(VDD),.Y(g4686),.A(g4590),.B(g1348));
  AND2 AND2_492(.VSS(VSS),.VDD(VDD),.Y(g4687),.A(g4493),.B(g1542));
  AND2 AND2_493(.VSS(VSS),.VDD(VDD),.Y(g4688),.A(g1474),.B(g4568));
  AND2 AND2_494(.VSS(VSS),.VDD(VDD),.Y(g4691),.A(g4581),.B(g2098));
  AND2 AND2_495(.VSS(VSS),.VDD(VDD),.Y(g4694),.A(g1481),.B(g4578));
  AND2 AND2_496(.VSS(VSS),.VDD(VDD),.Y(g4697),.A(g4589),.B(g1363));
  AND2 AND2_497(.VSS(VSS),.VDD(VDD),.Y(g4698),.A(g4586),.B(g2106));
  AND2 AND2_498(.VSS(VSS),.VDD(VDD),.Y(g4701),.A(g4596),.B(g1378));
  AND2 AND2_499(.VSS(VSS),.VDD(VDD),.Y(g4708),.A(g578),.B(g4541));
  AND2 AND2_500(.VSS(VSS),.VDD(VDD),.Y(g4730),.A(g1423),.B(g4565));
  AND2 AND2_501(.VSS(VSS),.VDD(VDD),.Y(g4735),.A(g2018),.B(g4577));
  AND2 AND2_502(.VSS(VSS),.VDD(VDD),.Y(g4739),.A(g2850),.B(g4579));
  AND2 AND2_503(.VSS(VSS),.VDD(VDD),.Y(g4744),.A(g3434),.B(g4582));
  AND2 AND2_504(.VSS(VSS),.VDD(VDD),.Y(g4756),.A(g3816),.B(g4587));
  AND2 AND2_505(.VSS(VSS),.VDD(VDD),.Y(g4759),.A(g536),.B(g4500));
  AND2 AND2_506(.VSS(VSS),.VDD(VDD),.Y(g4761),.A(g4567),.B(g1674));
  AND2 AND2_507(.VSS(VSS),.VDD(VDD),.Y(g4782),.A(g1624),.B(g4623));
  AND2 AND2_508(.VSS(VSS),.VDD(VDD),.Y(g4785),.A(g2160),.B(g4625));
  AND2 AND2_509(.VSS(VSS),.VDD(VDD),.Y(g4787),.A(g2937),.B(g4628));
  AND2 AND2_510(.VSS(VSS),.VDD(VDD),.Y(g4789),.A(g3551),.B(g4632));
  AND2 AND2_511(.VSS(VSS),.VDD(VDD),.Y(g4791),.A(g3936),.B(g4636));
  AND2 AND2_512(.VSS(VSS),.VDD(VDD),.Y(g4792),.A(g1417),.B(g4471));
  AND2 AND2_513(.VSS(VSS),.VDD(VDD),.Y(g4793),.A(g4277),.B(g4639));
  AND2 AND2_514(.VSS(VSS),.VDD(VDD),.Y(g4794),.A(g4593),.B(g949));
  AND2 AND2_515(.VSS(VSS),.VDD(VDD),.Y(g4797),.A(g4593),.B(g4643));
  AND2 AND2_516(.VSS(VSS),.VDD(VDD),.Y(g4800),.A(g4648),.B(g4296));
  AND2 AND2_517(.VSS(VSS),.VDD(VDD),.Y(g4826),.A(g4209),.B(g4463));
  AND2 AND2_518(.VSS(VSS),.VDD(VDD),.Y(g4827),.A(g4520),.B(g4515));
  AND2 AND2_519(.VSS(VSS),.VDD(VDD),.Y(g4828),.A(g4510),.B(g4508));
  AND2 AND2_520(.VSS(VSS),.VDD(VDD),.Y(g4829),.A(g4526),.B(g4522));
  AND2 AND2_521(.VSS(VSS),.VDD(VDD),.Y(g4830),.A(g4529),.B(g4525));
  AND2 AND2_522(.VSS(VSS),.VDD(VDD),.Y(g4831),.A(g4528),.B(g4524));
  AND2 AND2_523(.VSS(VSS),.VDD(VDD),.Y(g4832),.A(g4517),.B(g4512));
  AND2 AND2_524(.VSS(VSS),.VDD(VDD),.Y(g4833),.A(g4521),.B(g4516));
  AND2 AND2_525(.VSS(VSS),.VDD(VDD),.Y(g4834),.A(g4534),.B(g4531));
  AND2 AND2_526(.VSS(VSS),.VDD(VDD),.Y(g4835),.A(g4533),.B(g4530));
  AND2 AND2_527(.VSS(VSS),.VDD(VDD),.Y(g4836),.A(g4527),.B(g4523));
  AND2 AND2_528(.VSS(VSS),.VDD(VDD),.Y(g4838),.A(g4648),.B(g84));
  AND2 AND2_529(.VSS(VSS),.VDD(VDD),.Y(g4863),.A(g4777),.B(g2874));
  AND2 AND2_530(.VSS(VSS),.VDD(VDD),.Y(g4865),.A(g4776),.B(g1849));
  AND2 AND2_531(.VSS(VSS),.VDD(VDD),.Y(g4867),.A(g4811),.B(g3872));
  AND2 AND2_532(.VSS(VSS),.VDD(VDD),.Y(g4868),.A(g4774),.B(g2891));
  AND2 AND2_533(.VSS(VSS),.VDD(VDD),.Y(g4870),.A(g4779),.B(g1884));
  AND2 AND2_534(.VSS(VSS),.VDD(VDD),.Y(g4872),.A(g4760),.B(g1549));
  AND2 AND2_535(.VSS(VSS),.VDD(VDD),.Y(g4873),.A(g4838),.B(g4173));
  AND2 AND2_536(.VSS(VSS),.VDD(VDD),.Y(g4874),.A(g582),.B(g4708));
  AND2 AND2_537(.VSS(VSS),.VDD(VDD),.Y(g4928),.A(g148),.B(g4723));
  AND2 AND2_538(.VSS(VSS),.VDD(VDD),.Y(g4932),.A(g157),.B(g4727));
  AND2 AND2_539(.VSS(VSS),.VDD(VDD),.Y(g4937),.A(g166),.B(g4732));
  AND2 AND2_540(.VSS(VSS),.VDD(VDD),.Y(g4942),.A(g175),.B(g4736));
  AND2 AND2_541(.VSS(VSS),.VDD(VDD),.Y(g4947),.A(g184),.B(g4741));
  AND2 AND2_542(.VSS(VSS),.VDD(VDD),.Y(g4949),.A(g193),.B(g4753));
  AND2 AND2_543(.VSS(VSS),.VDD(VDD),.Y(g5017),.A(g4784),.B(g1679));
  AND2 AND2_544(.VSS(VSS),.VDD(VDD),.Y(g5023),.A(g3935),.B(g4804));
  AND2 AND2_545(.VSS(VSS),.VDD(VDD),.Y(g5043),.A(g3941),.B(g4805));
  AND2 AND2_546(.VSS(VSS),.VDD(VDD),.Y(g5047),.A(g3954),.B(g4806));
  AND2 AND2_547(.VSS(VSS),.VDD(VDD),.Y(g5050),.A(g4285),.B(g4807));
  AND2 AND2_548(.VSS(VSS),.VDD(VDD),.Y(g5053),.A(g4599),.B(g4808));
  AND2 AND2_549(.VSS(VSS),.VDD(VDD),.Y(g5095),.A(g4794),.B(g951));
  AND2 AND2_550(.VSS(VSS),.VDD(VDD),.Y(g5096),.A(g4794),.B(g4647));
  AND2 AND2_551(.VSS(VSS),.VDD(VDD),.Y(g5098),.A(g4021),.B(g4837));
  AND2 AND2_552(.VSS(VSS),.VDD(VDD),.Y(g5122),.A(g193),.B(g4662));
  AND2 AND2_553(.VSS(VSS),.VDD(VDD),.Y(g5123),.A(g4670),.B(g1936));
  AND2 AND2_554(.VSS(VSS),.VDD(VDD),.Y(g5142),.A(g148),.B(g5099));
  AND2 AND2_555(.VSS(VSS),.VDD(VDD),.Y(g5143),.A(g157),.B(g5099));
  AND2 AND2_556(.VSS(VSS),.VDD(VDD),.Y(g5144),.A(g166),.B(g5099));
  AND2 AND2_557(.VSS(VSS),.VDD(VDD),.Y(g5145),.A(g175),.B(g5099));
  AND2 AND2_558(.VSS(VSS),.VDD(VDD),.Y(g5146),.A(g184),.B(g5099));
  AND2 AND2_559(.VSS(VSS),.VDD(VDD),.Y(g5149),.A(g4910),.B(g1480));
  AND2 AND2_560(.VSS(VSS),.VDD(VDD),.Y(g5152),.A(g430),.B(g4950));
  AND2 AND2_561(.VSS(VSS),.VDD(VDD),.Y(g5153),.A(g492),.B(g4904));
  AND2 AND2_562(.VSS(VSS),.VDD(VDD),.Y(g5154),.A(g500),.B(g4993));
  AND2 AND2_563(.VSS(VSS),.VDD(VDD),.Y(g5156),.A(g434),.B(g4877));
  AND2 AND2_564(.VSS(VSS),.VDD(VDD),.Y(g5157),.A(g496),.B(g4904));
  AND2 AND2_565(.VSS(VSS),.VDD(VDD),.Y(g5158),.A(g504),.B(g4993));
  AND2 AND2_566(.VSS(VSS),.VDD(VDD),.Y(g5159),.A(g536),.B(g4967));
  AND2 AND2_567(.VSS(VSS),.VDD(VDD),.Y(g5161),.A(g5095),.B(g4535));
  AND2 AND2_568(.VSS(VSS),.VDD(VDD),.Y(g5162),.A(g5088),.B(g2105));
  AND2 AND2_569(.VSS(VSS),.VDD(VDD),.Y(g5163),.A(g402),.B(g4950));
  AND2 AND2_570(.VSS(VSS),.VDD(VDD),.Y(g5164),.A(g437),.B(g4877));
  AND2 AND2_571(.VSS(VSS),.VDD(VDD),.Y(g5165),.A(g508),.B(g4993));
  AND2 AND2_572(.VSS(VSS),.VDD(VDD),.Y(g5166),.A(g541),.B(g4967));
  AND2 AND2_573(.VSS(VSS),.VDD(VDD),.Y(g5167),.A(g5011),.B(g1556));
  AND2 AND2_574(.VSS(VSS),.VDD(VDD),.Y(g5169),.A(g5093),.B(g1375));
  AND2 AND2_575(.VSS(VSS),.VDD(VDD),.Y(g5170),.A(g5091),.B(g2111));
  AND2 AND2_576(.VSS(VSS),.VDD(VDD),.Y(g5171),.A(g406),.B(g4950));
  AND2 AND2_577(.VSS(VSS),.VDD(VDD),.Y(g5172),.A(g441),.B(g4877));
  AND2 AND2_578(.VSS(VSS),.VDD(VDD),.Y(g5173),.A(g512),.B(g4993));
  AND2 AND2_579(.VSS(VSS),.VDD(VDD),.Y(g5175),.A(g5094),.B(g1384));
  AND2 AND2_580(.VSS(VSS),.VDD(VDD),.Y(g5176),.A(g410),.B(g4950));
  AND2 AND2_581(.VSS(VSS),.VDD(VDD),.Y(g5177),.A(g445),.B(g4877));
  AND2 AND2_582(.VSS(VSS),.VDD(VDD),.Y(g5178),.A(g516),.B(g4993));
  AND2 AND2_583(.VSS(VSS),.VDD(VDD),.Y(g5180),.A(g414),.B(g4950));
  AND2 AND2_584(.VSS(VSS),.VDD(VDD),.Y(g5181),.A(g449),.B(g4877));
  AND2 AND2_585(.VSS(VSS),.VDD(VDD),.Y(g5182),.A(g520),.B(g4993));
  AND2 AND2_586(.VSS(VSS),.VDD(VDD),.Y(g5183),.A(g418),.B(g4950));
  AND2 AND2_587(.VSS(VSS),.VDD(VDD),.Y(g5184),.A(g453),.B(g4877));
  AND2 AND2_588(.VSS(VSS),.VDD(VDD),.Y(g5185),.A(g524),.B(g4993));
  AND2 AND2_589(.VSS(VSS),.VDD(VDD),.Y(g5186),.A(g422),.B(g4950));
  AND2 AND2_590(.VSS(VSS),.VDD(VDD),.Y(g5187),.A(g457),.B(g4877));
  AND2 AND2_591(.VSS(VSS),.VDD(VDD),.Y(g5188),.A(g1043),.B(g4894));
  AND2 AND2_592(.VSS(VSS),.VDD(VDD),.Y(g5189),.A(g528),.B(g4993));
  AND2 AND2_593(.VSS(VSS),.VDD(VDD),.Y(g5190),.A(g426),.B(g4950));
  AND2 AND2_594(.VSS(VSS),.VDD(VDD),.Y(g5191),.A(g461),.B(g4877));
  AND2 AND2_595(.VSS(VSS),.VDD(VDD),.Y(g5192),.A(g1046),.B(g4894));
  AND2 AND2_596(.VSS(VSS),.VDD(VDD),.Y(g5193),.A(g532),.B(g4967));
  AND2 AND2_597(.VSS(VSS),.VDD(VDD),.Y(g5194),.A(g586),.B(g4874));
  AND2 AND2_598(.VSS(VSS),.VDD(VDD),.Y(g5197),.A(g465),.B(g4967));
  AND2 AND2_599(.VSS(VSS),.VDD(VDD),.Y(g5198),.A(g558),.B(g5025));
  AND2 AND2_600(.VSS(VSS),.VDD(VDD),.Y(g5200),.A(g559),.B(g5025));
  AND2 AND2_601(.VSS(VSS),.VDD(VDD),.Y(g5201),.A(g4859),.B(g5084));
  AND2 AND2_602(.VSS(VSS),.VDD(VDD),.Y(g5209),.A(g560),.B(g5025));
  AND2 AND2_603(.VSS(VSS),.VDD(VDD),.Y(g5211),.A(g4860),.B(g5086));
  AND2 AND2_604(.VSS(VSS),.VDD(VDD),.Y(g5212),.A(g561),.B(g5025));
  AND2 AND2_605(.VSS(VSS),.VDD(VDD),.Y(g5213),.A(g4862),.B(g5087));
  AND2 AND2_606(.VSS(VSS),.VDD(VDD),.Y(g5214),.A(g562),.B(g5025));
  AND2 AND2_607(.VSS(VSS),.VDD(VDD),.Y(g5215),.A(g4864),.B(g5090));
  AND2 AND2_608(.VSS(VSS),.VDD(VDD),.Y(g5216),.A(g563),.B(g5025));
  AND2 AND2_609(.VSS(VSS),.VDD(VDD),.Y(g5217),.A(g4866),.B(g5092));
  AND2 AND2_610(.VSS(VSS),.VDD(VDD),.Y(g5218),.A(g564),.B(g5025));
  AND2 AND2_611(.VSS(VSS),.VDD(VDD),.Y(g5225),.A(g669),.B(g5054));
  AND2 AND2_612(.VSS(VSS),.VDD(VDD),.Y(g5226),.A(g672),.B(g5054));
  AND2 AND2_613(.VSS(VSS),.VDD(VDD),.Y(g5229),.A(g545),.B(g4980));
  AND2 AND2_614(.VSS(VSS),.VDD(VDD),.Y(g5232),.A(g548),.B(g4980));
  AND2 AND2_615(.VSS(VSS),.VDD(VDD),.Y(g5233),.A(g551),.B(g4980));
  AND2 AND2_616(.VSS(VSS),.VDD(VDD),.Y(g5234),.A(g197),.B(g4915));
  AND2 AND2_617(.VSS(VSS),.VDD(VDD),.Y(g5235),.A(g554),.B(g4980));
  AND2 AND2_618(.VSS(VSS),.VDD(VDD),.Y(g5236),.A(g269),.B(g4915));
  AND2 AND2_619(.VSS(VSS),.VDD(VDD),.Y(g5240),.A(g293),.B(g4915));
  AND2 AND2_620(.VSS(VSS),.VDD(VDD),.Y(g5245),.A(g297),.B(g4915));
  AND2 AND2_621(.VSS(VSS),.VDD(VDD),.Y(g5269),.A(g557),.B(g5025));
  AND2 AND2_622(.VSS(VSS),.VDD(VDD),.Y(g5311),.A(g5013),.B(g4468));
  AND2 AND2_623(.VSS(VSS),.VDD(VDD),.Y(g5317),.A(g148),.B(g4869));
  AND2 AND2_624(.VSS(VSS),.VDD(VDD),.Y(g5349),.A(g5324),.B(g3451));
  AND2 AND2_625(.VSS(VSS),.VDD(VDD),.Y(g5350),.A(g5325),.B(g3453));
  AND2 AND2_626(.VSS(VSS),.VDD(VDD),.Y(g5351),.A(g5326),.B(g3459));
  AND2 AND2_627(.VSS(VSS),.VDD(VDD),.Y(g5353),.A(g5327),.B(g3463));
  AND2 AND2_628(.VSS(VSS),.VDD(VDD),.Y(g5354),.A(g5249),.B(g2903));
  AND2 AND2_629(.VSS(VSS),.VDD(VDD),.Y(g5356),.A(g5265),.B(g1902));
  AND2 AND2_630(.VSS(VSS),.VDD(VDD),.Y(g5357),.A(g398),.B(g5220));
  AND2 AND2_631(.VSS(VSS),.VDD(VDD),.Y(g5359),.A(g4428),.B(g5155));
  AND2 AND2_632(.VSS(VSS),.VDD(VDD),.Y(g5360),.A(g4431),.B(g5160));
  AND2 AND2_633(.VSS(VSS),.VDD(VDD),.Y(g5361),.A(g4435),.B(g5168));
  AND2 AND2_634(.VSS(VSS),.VDD(VDD),.Y(g5362),.A(g4437),.B(g5174));
  AND2 AND2_635(.VSS(VSS),.VDD(VDD),.Y(g5363),.A(g4439),.B(g5179));
  AND2 AND2_636(.VSS(VSS),.VDD(VDD),.Y(g5364),.A(g574),.B(g5194));
  AND2 AND2_637(.VSS(VSS),.VDD(VDD),.Y(g5369),.A(g143),.B(g5247));
  AND2 AND2_638(.VSS(VSS),.VDD(VDD),.Y(g5371),.A(g152),.B(g5248));
  AND2 AND2_639(.VSS(VSS),.VDD(VDD),.Y(g5373),.A(g161),.B(g5250));
  AND2 AND2_640(.VSS(VSS),.VDD(VDD),.Y(g5376),.A(g170),.B(g5255));
  AND2 AND2_641(.VSS(VSS),.VDD(VDD),.Y(g5378),.A(g179),.B(g5260));
  AND2 AND2_642(.VSS(VSS),.VDD(VDD),.Y(g5380),.A(g188),.B(g5264));
  AND2 AND2_643(.VSS(VSS),.VDD(VDD),.Y(g5398),.A(g366),.B(g5261));
  AND2 AND2_644(.VSS(VSS),.VDD(VDD),.Y(g5402),.A(g370),.B(g5266));
  AND2 AND2_645(.VSS(VSS),.VDD(VDD),.Y(g5406),.A(g374),.B(g5270));
  AND2 AND2_646(.VSS(VSS),.VDD(VDD),.Y(g5410),.A(g378),.B(g5274));
  AND2 AND2_647(.VSS(VSS),.VDD(VDD),.Y(g5414),.A(g382),.B(g5278));
  AND2 AND2_648(.VSS(VSS),.VDD(VDD),.Y(g5419),.A(g386),.B(g5292));
  AND2 AND2_649(.VSS(VSS),.VDD(VDD),.Y(g5424),.A(g390),.B(g5296));
  AND2 AND2_650(.VSS(VSS),.VDD(VDD),.Y(g5428),.A(g394),.B(g5300));
  AND2 AND2_651(.VSS(VSS),.VDD(VDD),.Y(g5429),.A(g398),.B(g5304));
  AND2 AND2_652(.VSS(VSS),.VDD(VDD),.Y(g5438),.A(g5224),.B(g3769));
  AND3 AND3_17(.VSS(VSS),.VDD(VDD),.Y(g5441),.A(g4537),.B(g5251),.C(g1558));
  AND3 AND3_18(.VSS(VSS),.VDD(VDD),.Y(g5443),.A(g4537),.B(g5251),.C(g2307));
  AND3 AND3_19(.VSS(VSS),.VDD(VDD),.Y(g5444),.A(g4545),.B(g5256),.C(g1574));
  AND2 AND2_653(.VSS(VSS),.VDD(VDD),.Y(g5446),.A(g4537),.B(g5241));
  AND3 AND3_20(.VSS(VSS),.VDD(VDD),.Y(g5447),.A(g4545),.B(g5256),.C(g2311));
  AND2 AND2_654(.VSS(VSS),.VDD(VDD),.Y(g5449),.A(g4545),.B(g5246));
  AND2 AND2_655(.VSS(VSS),.VDD(VDD),.Y(g5451),.A(g5251),.B(g4544));
  AND2 AND2_656(.VSS(VSS),.VDD(VDD),.Y(g5452),.A(g5315),.B(g4612));
  AND2 AND2_657(.VSS(VSS),.VDD(VDD),.Y(g5454),.A(g5256),.B(g4549));
  AND2 AND2_658(.VSS(VSS),.VDD(VDD),.Y(g5481),.A(g366),.B(g5331));
  AND2 AND2_659(.VSS(VSS),.VDD(VDD),.Y(g5482),.A(g370),.B(g5331));
  AND2 AND2_660(.VSS(VSS),.VDD(VDD),.Y(g5483),.A(g374),.B(g5331));
  AND2 AND2_661(.VSS(VSS),.VDD(VDD),.Y(g5484),.A(g378),.B(g5331));
  AND2 AND2_662(.VSS(VSS),.VDD(VDD),.Y(g5485),.A(g382),.B(g5331));
  AND2 AND2_663(.VSS(VSS),.VDD(VDD),.Y(g5486),.A(g386),.B(g5331));
  AND2 AND2_664(.VSS(VSS),.VDD(VDD),.Y(g5487),.A(g390),.B(g5331));
  AND2 AND2_665(.VSS(VSS),.VDD(VDD),.Y(g5488),.A(g394),.B(g5331));
  AND2 AND2_666(.VSS(VSS),.VDD(VDD),.Y(g5492),.A(g5441),.B(g3452));
  AND2 AND2_667(.VSS(VSS),.VDD(VDD),.Y(g5494),.A(g5443),.B(g3455));
  AND2 AND2_668(.VSS(VSS),.VDD(VDD),.Y(g5495),.A(g5444),.B(g3456));
  AND2 AND2_669(.VSS(VSS),.VDD(VDD),.Y(g5496),.A(g5446),.B(g3457));
  AND2 AND2_670(.VSS(VSS),.VDD(VDD),.Y(g5497),.A(g5447),.B(g3458));
  AND2 AND2_671(.VSS(VSS),.VDD(VDD),.Y(g5498),.A(g5449),.B(g3460));
  AND2 AND2_672(.VSS(VSS),.VDD(VDD),.Y(g5499),.A(g5451),.B(g3462));
  AND2 AND2_673(.VSS(VSS),.VDD(VDD),.Y(g5500),.A(g5430),.B(g5074));
  AND2 AND2_674(.VSS(VSS),.VDD(VDD),.Y(g5501),.A(g5454),.B(g3478));
  AND2 AND2_675(.VSS(VSS),.VDD(VDD),.Y(g5503),.A(g366),.B(g5384));
  AND2 AND2_676(.VSS(VSS),.VDD(VDD),.Y(g5515),.A(g590),.B(g5364));
  AND2 AND2_677(.VSS(VSS),.VDD(VDD),.Y(g5553),.A(g5012),.B(g5440));
  AND2 AND2_678(.VSS(VSS),.VDD(VDD),.Y(g5555),.A(g5014),.B(g5442));
  AND2 AND2_679(.VSS(VSS),.VDD(VDD),.Y(g5556),.A(g5015),.B(g5445));
  AND2 AND2_680(.VSS(VSS),.VDD(VDD),.Y(g5557),.A(g5016),.B(g5448));
  AND2 AND2_681(.VSS(VSS),.VDD(VDD),.Y(g5558),.A(g5018),.B(g5450));
  AND2 AND2_682(.VSS(VSS),.VDD(VDD),.Y(g5559),.A(g5024),.B(g5453));
  AND2 AND2_683(.VSS(VSS),.VDD(VDD),.Y(g5560),.A(g5044),.B(g5456));
  AND2 AND2_684(.VSS(VSS),.VDD(VDD),.Y(g5562),.A(g5228),.B(g5457));
  AND2 AND2_685(.VSS(VSS),.VDD(VDD),.Y(g5569),.A(g5348),.B(g3772));
  AND2 AND2_686(.VSS(VSS),.VDD(VDD),.Y(g5598),.A(g5046),.B(g5509));
  AND2 AND2_687(.VSS(VSS),.VDD(VDD),.Y(g5599),.A(g5049),.B(g5512));
  AND2 AND2_688(.VSS(VSS),.VDD(VDD),.Y(g5600),.A(g5502),.B(g4900));
  AND2 AND2_689(.VSS(VSS),.VDD(VDD),.Y(g5601),.A(g5052),.B(g5518));
  AND2 AND2_690(.VSS(VSS),.VDD(VDD),.Y(g5602),.A(g594),.B(g5515));
  AND2 AND2_691(.VSS(VSS),.VDD(VDD),.Y(g5603),.A(g5504),.B(g4911));
  AND2 AND2_692(.VSS(VSS),.VDD(VDD),.Y(g5604),.A(g5059),.B(g5521));
  AND2 AND2_693(.VSS(VSS),.VDD(VDD),.Y(g5616),.A(g5505),.B(g4929));
  AND2 AND2_694(.VSS(VSS),.VDD(VDD),.Y(g5617),.A(g5061),.B(g5524));
  AND2 AND2_695(.VSS(VSS),.VDD(VDD),.Y(g5618),.A(g5506),.B(g4933));
  AND2 AND2_696(.VSS(VSS),.VDD(VDD),.Y(g5619),.A(g5064),.B(g5527));
  AND2 AND2_697(.VSS(VSS),.VDD(VDD),.Y(g5620),.A(g5507),.B(g4938));
  AND2 AND2_698(.VSS(VSS),.VDD(VDD),.Y(g5621),.A(g5508),.B(g4943));
  AND2 AND2_699(.VSS(VSS),.VDD(VDD),.Y(g5632),.A(g4494),.B(g5538));
  AND2 AND2_700(.VSS(VSS),.VDD(VDD),.Y(g5633),.A(g4496),.B(g5539));
  AND2 AND2_701(.VSS(VSS),.VDD(VDD),.Y(g5635),.A(g4498),.B(g5542));
  AND2 AND2_702(.VSS(VSS),.VDD(VDD),.Y(g5637),.A(g4499),.B(g5543));
  AND2 AND2_703(.VSS(VSS),.VDD(VDD),.Y(g5646),.A(g4502),.B(g5544));
  AND2 AND2_704(.VSS(VSS),.VDD(VDD),.Y(g5648),.A(g4507),.B(g5545));
  AND2 AND2_705(.VSS(VSS),.VDD(VDD),.Y(g5660),.A(g4509),.B(g5549));
  AND2 AND2_706(.VSS(VSS),.VDD(VDD),.Y(g5663),.A(g4513),.B(g5550));
  AND2 AND2_707(.VSS(VSS),.VDD(VDD),.Y(g5665),.A(g361),.B(g5570));
  AND2 AND2_708(.VSS(VSS),.VDD(VDD),.Y(g5668),.A(g49),.B(g5571));
  AND2 AND2_709(.VSS(VSS),.VDD(VDD),.Y(g5671),.A(g54),.B(g5572));
  AND2 AND2_710(.VSS(VSS),.VDD(VDD),.Y(g5673),.A(g59),.B(g5573));
  AND2 AND2_711(.VSS(VSS),.VDD(VDD),.Y(g5675),.A(g64),.B(g5574));
  AND2 AND2_712(.VSS(VSS),.VDD(VDD),.Y(g5677),.A(g69),.B(g5575));
  AND2 AND2_713(.VSS(VSS),.VDD(VDD),.Y(g5679),.A(g74),.B(g5576));
  AND2 AND2_714(.VSS(VSS),.VDD(VDD),.Y(g5681),.A(g79),.B(g5577));
  AND2 AND2_715(.VSS(VSS),.VDD(VDD),.Y(g5682),.A(g84),.B(g5578));
  AND2 AND2_716(.VSS(VSS),.VDD(VDD),.Y(g5701),.A(g5683),.B(g3813));
  AND2 AND2_717(.VSS(VSS),.VDD(VDD),.Y(g5728),.A(g5623),.B(g3889));
  AND2 AND2_718(.VSS(VSS),.VDD(VDD),.Y(g5883),.A(g5824),.B(g3752));
  AND2 AND2_719(.VSS(VSS),.VDD(VDD),.Y(g5898),.A(g5800),.B(g5647));
  AND2 AND2_720(.VSS(VSS),.VDD(VDD),.Y(g5900),.A(g5804),.B(g5658));
  AND2 AND2_721(.VSS(VSS),.VDD(VDD),.Y(g5902),.A(g5808),.B(g5661));
  AND2 AND2_722(.VSS(VSS),.VDD(VDD),.Y(g5904),.A(g5812),.B(g5664));
  AND2 AND2_723(.VSS(VSS),.VDD(VDD),.Y(g5909),.A(g5787),.B(g3384));
  AND2 AND2_724(.VSS(VSS),.VDD(VDD),.Y(g5910),.A(g5816),.B(g5667));
  AND2 AND2_725(.VSS(VSS),.VDD(VDD),.Y(g5911),.A(g5817),.B(g5670));
  AND2 AND2_726(.VSS(VSS),.VDD(VDD),.Y(g5935),.A(g5112),.B(g5784));
  AND2 AND2_727(.VSS(VSS),.VDD(VDD),.Y(g5936),.A(g5113),.B(g5788));
  AND2 AND2_728(.VSS(VSS),.VDD(VDD),.Y(g5937),.A(g5775),.B(g5392));
  AND2 AND2_729(.VSS(VSS),.VDD(VDD),.Y(g5938),.A(g5114),.B(g5791));
  AND2 AND2_730(.VSS(VSS),.VDD(VDD),.Y(g5939),.A(g5776),.B(g5395));
  AND2 AND2_731(.VSS(VSS),.VDD(VDD),.Y(g5940),.A(g5115),.B(g5794));
  AND2 AND2_732(.VSS(VSS),.VDD(VDD),.Y(g5941),.A(g5777),.B(g5399));
  AND2 AND2_733(.VSS(VSS),.VDD(VDD),.Y(g5942),.A(g5117),.B(g5797));
  AND2 AND2_734(.VSS(VSS),.VDD(VDD),.Y(g5944),.A(g5778),.B(g5403));
  AND2 AND2_735(.VSS(VSS),.VDD(VDD),.Y(g5945),.A(g5118),.B(g5801));
  AND2 AND2_736(.VSS(VSS),.VDD(VDD),.Y(g5948),.A(g5779),.B(g5407));
  AND2 AND2_737(.VSS(VSS),.VDD(VDD),.Y(g5949),.A(g5119),.B(g5805));
  AND2 AND2_738(.VSS(VSS),.VDD(VDD),.Y(g5951),.A(g5780),.B(g5411));
  AND2 AND2_739(.VSS(VSS),.VDD(VDD),.Y(g5952),.A(g5120),.B(g5809));
  AND2 AND2_740(.VSS(VSS),.VDD(VDD),.Y(g5953),.A(g5781),.B(g5415));
  AND2 AND2_741(.VSS(VSS),.VDD(VDD),.Y(g5954),.A(g5121),.B(g5813));
  AND2 AND2_742(.VSS(VSS),.VDD(VDD),.Y(g5955),.A(g5782),.B(g5420));
  AND2 AND2_743(.VSS(VSS),.VDD(VDD),.Y(g5956),.A(g5783),.B(g5425));
  AND2 AND2_744(.VSS(VSS),.VDD(VDD),.Y(g6047),.A(g5824),.B(g1692));
  AND2 AND2_745(.VSS(VSS),.VDD(VDD),.Y(g6055),.A(g5824),.B(g1696));
  AND2 AND2_746(.VSS(VSS),.VDD(VDD),.Y(g6056),.A(g5824),.B(g1699));
  AND2 AND2_747(.VSS(VSS),.VDD(VDD),.Y(g6060),.A(g5824),.B(g1703));
  AND2 AND2_748(.VSS(VSS),.VDD(VDD),.Y(g6061),.A(g5824),.B(g1711));
  AND2 AND2_749(.VSS(VSS),.VDD(VDD),.Y(g6066),.A(g5824),.B(g1721));
  AND2 AND2_750(.VSS(VSS),.VDD(VDD),.Y(g6068),.A(g5824),.B(g1726));
  AND2 AND2_751(.VSS(VSS),.VDD(VDD),.Y(g6077),.A(g5824),.B(g1735));
  AND2 AND2_752(.VSS(VSS),.VDD(VDD),.Y(g6079),.A(g1236),.B(g5753));
  AND2 AND2_753(.VSS(VSS),.VDD(VDD),.Y(g6081),.A(g1177),.B(g5731));
  AND2 AND2_754(.VSS(VSS),.VDD(VDD),.Y(g6082),.A(g1123),.B(g5742));
  AND2 AND2_755(.VSS(VSS),.VDD(VDD),.Y(g6084),.A(g1123),.B(g5753));
  AND2 AND2_756(.VSS(VSS),.VDD(VDD),.Y(g6085),.A(g1161),.B(g5731));
  AND2 AND2_757(.VSS(VSS),.VDD(VDD),.Y(g6086),.A(g1143),.B(g5742));
  AND2 AND2_758(.VSS(VSS),.VDD(VDD),.Y(g6088),.A(g1143),.B(g5753));
  AND2 AND2_759(.VSS(VSS),.VDD(VDD),.Y(g6089),.A(g1143),.B(g5731));
  AND2 AND2_760(.VSS(VSS),.VDD(VDD),.Y(g6090),.A(g1161),.B(g5742));
  AND2 AND2_761(.VSS(VSS),.VDD(VDD),.Y(g6091),.A(g1161),.B(g5753));
  AND2 AND2_762(.VSS(VSS),.VDD(VDD),.Y(g6092),.A(g1123),.B(g5731));
  AND2 AND2_763(.VSS(VSS),.VDD(VDD),.Y(g6093),.A(g1177),.B(g5742));
  AND2 AND2_764(.VSS(VSS),.VDD(VDD),.Y(g6094),.A(g1177),.B(g5753));
  AND2 AND2_765(.VSS(VSS),.VDD(VDD),.Y(g6096),.A(g1193),.B(g5753));
  AND2 AND2_766(.VSS(VSS),.VDD(VDD),.Y(g6098),.A(g1209),.B(g5753));
  AND2 AND2_767(.VSS(VSS),.VDD(VDD),.Y(g6099),.A(g1222),.B(g5753));
  AND2 AND2_768(.VSS(VSS),.VDD(VDD),.Y(g6123),.A(g5702),.B(g5958));
  AND2 AND2_769(.VSS(VSS),.VDD(VDD),.Y(g6124),.A(g5705),.B(g5958));
  AND2 AND2_770(.VSS(VSS),.VDD(VDD),.Y(g6125),.A(g5708),.B(g5975));
  AND2 AND2_771(.VSS(VSS),.VDD(VDD),.Y(g6126),.A(g5711),.B(g5958));
  AND2 AND2_772(.VSS(VSS),.VDD(VDD),.Y(g6127),.A(g5714),.B(g5975));
  AND2 AND2_773(.VSS(VSS),.VDD(VDD),.Y(g6128),.A(g5590),.B(g5958));
  AND2 AND2_774(.VSS(VSS),.VDD(VDD),.Y(g6129),.A(g5717),.B(g5975));
  AND2 AND2_775(.VSS(VSS),.VDD(VDD),.Y(g6130),.A(g5720),.B(g5958));
  AND2 AND2_776(.VSS(VSS),.VDD(VDD),.Y(g6131),.A(g5593),.B(g5975));
  AND2 AND2_777(.VSS(VSS),.VDD(VDD),.Y(g6132),.A(g3752),.B(g5880));
  AND2 AND2_778(.VSS(VSS),.VDD(VDD),.Y(g6133),.A(g5723),.B(g5975));
  AND2 AND2_779(.VSS(VSS),.VDD(VDD),.Y(g6135),.A(g5584),.B(g5958));
  AND2 AND2_780(.VSS(VSS),.VDD(VDD),.Y(g6140),.A(g5587),.B(g5975));
  AND2 AND2_781(.VSS(VSS),.VDD(VDD),.Y(g6141),.A(g3173),.B(g5997));
  AND2 AND2_782(.VSS(VSS),.VDD(VDD),.Y(g6144),.A(g3183),.B(g5997));
  AND2 AND2_783(.VSS(VSS),.VDD(VDD),.Y(g6145),.A(g3187),.B(g6015));
  AND2 AND2_784(.VSS(VSS),.VDD(VDD),.Y(g6146),.A(g3192),.B(g5997));
  AND2 AND2_785(.VSS(VSS),.VDD(VDD),.Y(g6148),.A(g3196),.B(g6015));
  AND2 AND2_786(.VSS(VSS),.VDD(VDD),.Y(g6149),.A(g3200),.B(g5997));
  AND2 AND2_787(.VSS(VSS),.VDD(VDD),.Y(g6150),.A(g3204),.B(g6015));
  AND2 AND2_788(.VSS(VSS),.VDD(VDD),.Y(g6151),.A(g3209),.B(g5997));
  AND2 AND2_789(.VSS(VSS),.VDD(VDD),.Y(g6152),.A(g3212),.B(g6015));
  AND2 AND2_790(.VSS(VSS),.VDD(VDD),.Y(g6153),.A(g3216),.B(g5997));
  AND2 AND2_791(.VSS(VSS),.VDD(VDD),.Y(g6154),.A(g3219),.B(g6015));
  AND2 AND2_792(.VSS(VSS),.VDD(VDD),.Y(g6155),.A(g2588),.B(g5997));
  AND2 AND2_793(.VSS(VSS),.VDD(VDD),.Y(g6156),.A(g2591),.B(g6015));
  AND2 AND2_794(.VSS(VSS),.VDD(VDD),.Y(g6157),.A(g3158),.B(g5997));
  AND2 AND2_795(.VSS(VSS),.VDD(VDD),.Y(g6158),.A(g2594),.B(g6015));
  AND2 AND2_796(.VSS(VSS),.VDD(VDD),.Y(g6159),.A(g3177),.B(g6015));
  AND2 AND2_797(.VSS(VSS),.VDD(VDD),.Y(g6238),.A(g528),.B(g5886));
  AND2 AND2_798(.VSS(VSS),.VDD(VDD),.Y(g6240),.A(g4205),.B(g5888));
  AND2 AND2_799(.VSS(VSS),.VDD(VDD),.Y(g6241),.A(g1325),.B(g5887));
  AND2 AND2_800(.VSS(VSS),.VDD(VDD),.Y(g6243),.A(g500),.B(g5890));
  AND2 AND2_801(.VSS(VSS),.VDD(VDD),.Y(g6244),.A(g4759),.B(g5891));
  AND2 AND2_802(.VSS(VSS),.VDD(VDD),.Y(g6245),.A(g1329),.B(g5889));
  AND2 AND2_803(.VSS(VSS),.VDD(VDD),.Y(g6247),.A(g504),.B(g5893));
  AND2 AND2_804(.VSS(VSS),.VDD(VDD),.Y(g6248),.A(g465),.B(g5894));
  AND2 AND2_805(.VSS(VSS),.VDD(VDD),.Y(g6249),.A(g1332),.B(g5892));
  AND2 AND2_806(.VSS(VSS),.VDD(VDD),.Y(g6250),.A(g1692),.B(g6036));
  AND2 AND2_807(.VSS(VSS),.VDD(VDD),.Y(g6253),.A(g508),.B(g5896));
  AND2 AND2_808(.VSS(VSS),.VDD(VDD),.Y(g6254),.A(g532),.B(g5897));
  AND2 AND2_809(.VSS(VSS),.VDD(VDD),.Y(g6255),.A(g1335),.B(g5895));
  AND2 AND2_810(.VSS(VSS),.VDD(VDD),.Y(g6256),.A(g1696),.B(g6040));
  AND2 AND2_811(.VSS(VSS),.VDD(VDD),.Y(g6258),.A(g512),.B(g5899));
  AND2 AND2_812(.VSS(VSS),.VDD(VDD),.Y(g6259),.A(g1699),.B(g6044));
  AND2 AND2_813(.VSS(VSS),.VDD(VDD),.Y(g6260),.A(g1703),.B(g6048));
  AND2 AND2_814(.VSS(VSS),.VDD(VDD),.Y(g6262),.A(g516),.B(g5901));
  AND2 AND2_815(.VSS(VSS),.VDD(VDD),.Y(g6263),.A(g1711),.B(g6052));
  AND2 AND2_816(.VSS(VSS),.VDD(VDD),.Y(g6265),.A(g520),.B(g5903));
  AND2 AND2_817(.VSS(VSS),.VDD(VDD),.Y(g6266),.A(g1721),.B(g6057));
  AND2 AND2_818(.VSS(VSS),.VDD(VDD),.Y(g6269),.A(g524),.B(g5908));
  AND2 AND2_819(.VSS(VSS),.VDD(VDD),.Y(g6270),.A(g1726),.B(g6062));
  AND2 AND2_820(.VSS(VSS),.VDD(VDD),.Y(g6275),.A(g1735),.B(g6070));
  AND2 AND2_821(.VSS(VSS),.VDD(VDD),.Y(g6288),.A(g5615),.B(g6160));
  AND2 AND2_822(.VSS(VSS),.VDD(VDD),.Y(g6291),.A(g5210),.B(g6161));
  AND2 AND2_823(.VSS(VSS),.VDD(VDD),.Y(g6295),.A(g5379),.B(g6162));
  AND2 AND2_824(.VSS(VSS),.VDD(VDD),.Y(g6299),.A(g5530),.B(g6163));
  AND2 AND2_825(.VSS(VSS),.VDD(VDD),.Y(g6302),.A(g5740),.B(g6164));
  AND2 AND2_826(.VSS(VSS),.VDD(VDD),.Y(g6304),.A(g5915),.B(g6165));
  AND2 AND2_827(.VSS(VSS),.VDD(VDD),.Y(g6311),.A(g3837),.B(g6194));
  AND2 AND2_828(.VSS(VSS),.VDD(VDD),.Y(g6313),.A(g3841),.B(g6194));
  AND2 AND2_829(.VSS(VSS),.VDD(VDD),.Y(g6315),.A(g3849),.B(g6194));
  AND2 AND2_830(.VSS(VSS),.VDD(VDD),.Y(g6316),.A(g3855),.B(g6194));
  AND2 AND2_831(.VSS(VSS),.VDD(VDD),.Y(g6317),.A(g3862),.B(g6194));
  AND2 AND2_832(.VSS(VSS),.VDD(VDD),.Y(g6318),.A(g3865),.B(g6212));
  AND2 AND2_833(.VSS(VSS),.VDD(VDD),.Y(g6320),.A(g3869),.B(g6194));
  AND2 AND2_834(.VSS(VSS),.VDD(VDD),.Y(g6321),.A(g3873),.B(g6212));
  AND2 AND2_835(.VSS(VSS),.VDD(VDD),.Y(g6323),.A(g3877),.B(g6194));
  AND2 AND2_836(.VSS(VSS),.VDD(VDD),.Y(g6324),.A(g3880),.B(g6212));
  AND2 AND2_837(.VSS(VSS),.VDD(VDD),.Y(g6326),.A(g3833),.B(g6194));
  AND2 AND2_838(.VSS(VSS),.VDD(VDD),.Y(g6327),.A(g3884),.B(g6212));
  AND2 AND2_839(.VSS(VSS),.VDD(VDD),.Y(g6329),.A(g3888),.B(g6212));
  AND2 AND2_840(.VSS(VSS),.VDD(VDD),.Y(g6331),.A(g3891),.B(g6212));
  AND2 AND2_841(.VSS(VSS),.VDD(VDD),.Y(g6333),.A(g3896),.B(g6212));
  AND2 AND2_842(.VSS(VSS),.VDD(VDD),.Y(g6334),.A(g3858),.B(g6212));
  AND2 AND2_843(.VSS(VSS),.VDD(VDD),.Y(g6336),.A(g6246),.B(g6065));
  AND2 AND2_844(.VSS(VSS),.VDD(VDD),.Y(g6338),.A(g6251),.B(g6067));
  AND2 AND2_845(.VSS(VSS),.VDD(VDD),.Y(g6340),.A(g6257),.B(g6069));
  AND2 AND2_846(.VSS(VSS),.VDD(VDD),.Y(g6341),.A(g6261),.B(g6074));
  AND2 AND2_847(.VSS(VSS),.VDD(VDD),.Y(g6342),.A(g6264),.B(g6076));
  AND2 AND2_848(.VSS(VSS),.VDD(VDD),.Y(g6343),.A(g6268),.B(g6078));
  AND2 AND2_849(.VSS(VSS),.VDD(VDD),.Y(g6344),.A(g6272),.B(g6080));
  AND2 AND2_850(.VSS(VSS),.VDD(VDD),.Y(g6345),.A(g6273),.B(g6083));
  AND2 AND2_851(.VSS(VSS),.VDD(VDD),.Y(g6346),.A(g6274),.B(g6087));
  AND2 AND2_852(.VSS(VSS),.VDD(VDD),.Y(g6348),.A(g5869),.B(g6211));
  AND2 AND2_853(.VSS(VSS),.VDD(VDD),.Y(g6354),.A(g5866),.B(g6193));
  AND3 AND3_21(.VSS(VSS),.VDD(VDD),.Y(g6468),.A(g2032),.B(g6394),.C(g1609));
  AND3 AND3_22(.VSS(VSS),.VDD(VDD),.Y(g6469),.A(g2121),.B(g2032),.C(g6394));
  AND3 AND3_23(.VSS(VSS),.VDD(VDD),.Y(g6473),.A(g2036),.B(g6397),.C(g1628));
  AND3 AND3_24(.VSS(VSS),.VDD(VDD),.Y(g6474),.A(g2138),.B(g2036),.C(g6397));
  AND2 AND2_854(.VSS(VSS),.VDD(VDD),.Y(g6555),.A(g1838),.B(g6469));
  AND2 AND2_855(.VSS(VSS),.VDD(VDD),.Y(g6557),.A(g1595),.B(g6469));
  AND2 AND2_856(.VSS(VSS),.VDD(VDD),.Y(g6558),.A(g1842),.B(g6474));
  AND2 AND2_857(.VSS(VSS),.VDD(VDD),.Y(g6559),.A(g1612),.B(g6474));
  AND2 AND2_858(.VSS(VSS),.VDD(VDD),.Y(g6603),.A(g6581),.B(g6236));
  AND2 AND2_859(.VSS(VSS),.VDD(VDD),.Y(g6613),.A(g932),.B(g6554));
  AND2 AND2_860(.VSS(VSS),.VDD(VDD),.Y(g6614),.A(g932),.B(g6556));
  AND2 AND2_861(.VSS(VSS),.VDD(VDD),.Y(g6619),.A(g6515),.B(g6115));
  AND2 AND2_862(.VSS(VSS),.VDD(VDD),.Y(g6620),.A(g6516),.B(g6117));
  AND3 AND3_25(.VSS(VSS),.VDD(VDD),.Y(g6625),.A(g2121),.B(g1595),.C(g6538));
  AND3 AND3_26(.VSS(VSS),.VDD(VDD),.Y(g6628),.A(g2138),.B(g1612),.C(g6540));
  AND2 AND2_863(.VSS(VSS),.VDD(VDD),.Y(g6631),.A(g1838),.B(g6545));
  AND2 AND2_864(.VSS(VSS),.VDD(VDD),.Y(g6634),.A(g1595),.B(g6545));
  AND2 AND2_865(.VSS(VSS),.VDD(VDD),.Y(g6637),.A(g1842),.B(g6549));
  AND2 AND2_866(.VSS(VSS),.VDD(VDD),.Y(g6640),.A(g1612),.B(g6549));
  AND2 AND2_867(.VSS(VSS),.VDD(VDD),.Y(g6643),.A(g6574),.B(g6229));
  AND2 AND2_868(.VSS(VSS),.VDD(VDD),.Y(g6644),.A(g6575),.B(g6230));
  AND2 AND2_869(.VSS(VSS),.VDD(VDD),.Y(g6645),.A(g6576),.B(g6231));
  AND2 AND2_870(.VSS(VSS),.VDD(VDD),.Y(g6646),.A(g6577),.B(g6232));
  AND2 AND2_871(.VSS(VSS),.VDD(VDD),.Y(g6647),.A(g6578),.B(g6233));
  AND2 AND2_872(.VSS(VSS),.VDD(VDD),.Y(g6648),.A(g6579),.B(g6234));
  AND2 AND2_873(.VSS(VSS),.VDD(VDD),.Y(g6650),.A(g6580),.B(g6235));
  AND2 AND2_874(.VSS(VSS),.VDD(VDD),.Y(g6692),.A(g6616),.B(g6615));
  AND2 AND2_875(.VSS(VSS),.VDD(VDD),.Y(g6693),.A(g6618),.B(g6617));
  AND2 AND2_876(.VSS(VSS),.VDD(VDD),.Y(g6716),.A(g6682),.B(g932));
  AND2 AND2_877(.VSS(VSS),.VDD(VDD),.Y(g6718),.A(g4511),.B(g6661));
  AND2 AND2_878(.VSS(VSS),.VDD(VDD),.Y(g6719),.A(g4518),.B(g6665));
  AND2 AND2_879(.VSS(VSS),.VDD(VDD),.Y(g6731),.A(g6717),.B(g4427));
  AND3 AND3_27(.VSS(VSS),.VDD(VDD),.Y(g6736),.A(g6712),.B(g754),.C(g5237));
  AND3 AND3_28(.VSS(VSS),.VDD(VDD),.Y(g6737),.A(g6714),.B(g760),.C(g5237));
  AND3 AND3_29(.VSS(VSS),.VDD(VDD),.Y(g6738),.A(g6713),.B(g809),.C(g5242));
  AND3 AND3_30(.VSS(VSS),.VDD(VDD),.Y(g6739),.A(g6715),.B(g815),.C(g5242));
  AND2 AND2_880(.VSS(VSS),.VDD(VDD),.Y(g6748),.A(g6733),.B(g6732));
  AND2 AND2_881(.VSS(VSS),.VDD(VDD),.Y(g6749),.A(g6735),.B(g6734));
  AND2 AND2_882(.VSS(VSS),.VDD(VDD),.Y(g6766),.A(g6750),.B(g2986));
  AND2 AND2_883(.VSS(VSS),.VDD(VDD),.Y(g6767),.A(g6754),.B(g2986));
  AND2 AND2_884(.VSS(VSS),.VDD(VDD),.Y(g6768),.A(g6750),.B(g3477));
  AND2 AND2_885(.VSS(VSS),.VDD(VDD),.Y(g6769),.A(g6758),.B(g2986));
  AND2 AND2_886(.VSS(VSS),.VDD(VDD),.Y(g6770),.A(g6754),.B(g3482));
  AND2 AND2_887(.VSS(VSS),.VDD(VDD),.Y(g6771),.A(g6758),.B(g3483));
  AND2 AND2_888(.VSS(VSS),.VDD(VDD),.Y(g6772),.A(g6746),.B(g3312));
  AND2 AND2_889(.VSS(VSS),.VDD(VDD),.Y(g6773),.A(g6762),.B(g2986));
  AND2 AND2_890(.VSS(VSS),.VDD(VDD),.Y(g6777),.A(g6762),.B(g3488));
  AND2 AND2_891(.VSS(VSS),.VDD(VDD),.Y(g6798),.A(g4946),.B(g6781));
  AND2 AND2_892(.VSS(VSS),.VDD(VDD),.Y(g6799),.A(g4948),.B(g6782));
  AND2 AND2_893(.VSS(VSS),.VDD(VDD),.Y(g6816),.A(g6784),.B(g3346));
  AND2 AND2_894(.VSS(VSS),.VDD(VDD),.Y(g6828),.A(g6803),.B(g5958));
  AND2 AND2_895(.VSS(VSS),.VDD(VDD),.Y(g6829),.A(g6806),.B(g5958));
  AND2 AND2_896(.VSS(VSS),.VDD(VDD),.Y(g6830),.A(g6809),.B(g5975));
  AND2 AND2_897(.VSS(VSS),.VDD(VDD),.Y(g6831),.A(g6812),.B(g5975));
  AND3 AND3_31(.VSS(VSS),.VDD(VDD),.Y(g6848),.A(g3741),.B(g328),.C(g6843));
  AND2 AND2_898(.VSS(VSS),.VDD(VDD),.Y(g6851),.A(g6846),.B(g2293));
  AND2 AND2_899(.VSS(VSS),.VDD(VDD),.Y(g6852),.A(g6847),.B(g2295));
  AND2 AND2_900(.VSS(VSS),.VDD(VDD),.Y(g6874),.A(g6873),.B(g2060));
  AND2 AND2_901(.VSS(VSS),.VDD(VDD),.Y(g6908),.A(g6907),.B(g3886));
  AND2 AND2_902(.VSS(VSS),.VDD(VDD),.Y(g6909),.A(g6896),.B(g6894));
  AND2 AND2_903(.VSS(VSS),.VDD(VDD),.Y(g6910),.A(g6892),.B(g6891));
  AND2 AND2_904(.VSS(VSS),.VDD(VDD),.Y(g6911),.A(g6904),.B(g6902));
  AND2 AND2_905(.VSS(VSS),.VDD(VDD),.Y(g6912),.A(g6899),.B(g6897));
  AND2 AND2_906(.VSS(VSS),.VDD(VDD),.Y(g6913),.A(g6900),.B(g6898));
  AND2 AND2_907(.VSS(VSS),.VDD(VDD),.Y(g6914),.A(g6895),.B(g6893));
  AND2 AND2_908(.VSS(VSS),.VDD(VDD),.Y(g6915),.A(g6906),.B(g6905));
  AND2 AND2_909(.VSS(VSS),.VDD(VDD),.Y(g6916),.A(g6903),.B(g6901));
  AND2 AND2_910(.VSS(VSS),.VDD(VDD),.Y(g6923),.A(g6918),.B(g6917));
  AND2 AND2_911(.VSS(VSS),.VDD(VDD),.Y(g6924),.A(g6920),.B(g6919));
  AND2 AND2_912(.VSS(VSS),.VDD(VDD),.Y(g6934),.A(g6932),.B(g3605));
  AND2 AND2_913(.VSS(VSS),.VDD(VDD),.Y(g6935),.A(g6933),.B(g3622));
//
  OR2 OR2_0(.VSS(VSS),.VDD(VDD),.Y(g1589),.A(g1059),.B(g1045));
  OR2 OR2_1(.VSS(VSS),.VDD(VDD),.Y(g2896),.A(g2323),.B(g1763));
  OR2 OR2_2(.VSS(VSS),.VDD(VDD),.Y(g2924),.A(g2095),.B(g1573));
  OR2 OR2_3(.VSS(VSS),.VDD(VDD),.Y(g2928),.A(g2100),.B(g1582));
  OR2 OR2_4(.VSS(VSS),.VDD(VDD),.Y(g3503),.A(g3122),.B(g3132));
  OR2 OR2_5(.VSS(VSS),.VDD(VDD),.Y(g3533),.A(g3154),.B(g3166));
  OR2 OR2_6(.VSS(VSS),.VDD(VDD),.Y(g3598),.A(g2808),.B(g2821));
  OR2 OR2_7(.VSS(VSS),.VDD(VDD),.Y(g3599),.A(g2935),.B(g1637));
  OR2 OR2_8(.VSS(VSS),.VDD(VDD),.Y(g3732),.A(g3324),.B(g2732));
  OR2 OR2_9(.VSS(VSS),.VDD(VDD),.Y(g3733),.A(g3325),.B(g2733));
  OR2 OR2_10(.VSS(VSS),.VDD(VDD),.Y(g3739),.A(g3334),.B(g2746));
  OR2 OR2_11(.VSS(VSS),.VDD(VDD),.Y(g3740),.A(g3335),.B(g2747));
  OR2 OR2_12(.VSS(VSS),.VDD(VDD),.Y(g3743),.A(g3344),.B(g2758));
  OR2 OR2_13(.VSS(VSS),.VDD(VDD),.Y(g3744),.A(g3345),.B(g2759));
  OR2 OR2_14(.VSS(VSS),.VDD(VDD),.Y(g3745),.A(g3356),.B(g2770));
  OR2 OR2_15(.VSS(VSS),.VDD(VDD),.Y(g3746),.A(g3357),.B(g2771));
  OR2 OR2_16(.VSS(VSS),.VDD(VDD),.Y(g3747),.A(g3365),.B(g2781));
  OR2 OR2_17(.VSS(VSS),.VDD(VDD),.Y(g3748),.A(g3366),.B(g2782));
  OR2 OR2_18(.VSS(VSS),.VDD(VDD),.Y(g3749),.A(g3371),.B(g2793));
  OR2 OR2_19(.VSS(VSS),.VDD(VDD),.Y(g3750),.A(g3372),.B(g2794));
  OR2 OR2_20(.VSS(VSS),.VDD(VDD),.Y(g3751),.A(g3375),.B(g2807));
  OR2 OR2_21(.VSS(VSS),.VDD(VDD),.Y(g3815),.A(g3282),.B(g2659));
  OR2 OR2_22(.VSS(VSS),.VDD(VDD),.Y(g3820),.A(g3287),.B(g2671));
  OR2 OR2_23(.VSS(VSS),.VDD(VDD),.Y(g3821),.A(g2951),.B(g3466));
  OR2 OR2_24(.VSS(VSS),.VDD(VDD),.Y(g3828),.A(g3304),.B(g1351));
  OR2 OR2_25(.VSS(VSS),.VDD(VDD),.Y(g3829),.A(g3294),.B(g3305));
  OR2 OR2_26(.VSS(VSS),.VDD(VDD),.Y(g3833),.A(g3602),.B(g3608));
  OR2 OR2_27(.VSS(VSS),.VDD(VDD),.Y(g3837),.A(g3609),.B(g3613));
  OR2 OR2_28(.VSS(VSS),.VDD(VDD),.Y(g3841),.A(g3614),.B(g3617));
  OR2 OR2_29(.VSS(VSS),.VDD(VDD),.Y(g3842),.A(g3670),.B(g3135));
  OR2 OR2_30(.VSS(VSS),.VDD(VDD),.Y(g3849),.A(g3618),.B(g3625));
  OR2 OR2_31(.VSS(VSS),.VDD(VDD),.Y(g3850),.A(g3680),.B(g3145));
  OR2 OR2_32(.VSS(VSS),.VDD(VDD),.Y(g3851),.A(g3681),.B(g3146));
  OR2 OR2_33(.VSS(VSS),.VDD(VDD),.Y(g3855),.A(g3626),.B(g3631));
  OR2 OR2_34(.VSS(VSS),.VDD(VDD),.Y(g3856),.A(g3686),.B(g3157));
  OR2 OR2_35(.VSS(VSS),.VDD(VDD),.Y(g3857),.A(g3687),.B(g3161));
  OR2 OR2_36(.VSS(VSS),.VDD(VDD),.Y(g3858),.A(g3629),.B(g3636));
  OR2 OR2_37(.VSS(VSS),.VDD(VDD),.Y(g3862),.A(g3632),.B(g3641));
  OR2 OR2_38(.VSS(VSS),.VDD(VDD),.Y(g3863),.A(g3692),.B(g3172));
  OR2 OR2_39(.VSS(VSS),.VDD(VDD),.Y(g3864),.A(g3693),.B(g3176));
  OR2 OR2_40(.VSS(VSS),.VDD(VDD),.Y(g3865),.A(g3637),.B(g3648));
  OR2 OR2_41(.VSS(VSS),.VDD(VDD),.Y(g3869),.A(g3642),.B(g3650));
  OR2 OR2_42(.VSS(VSS),.VDD(VDD),.Y(g3870),.A(g3700),.B(g3182));
  OR2 OR2_43(.VSS(VSS),.VDD(VDD),.Y(g3871),.A(g3701),.B(g3186));
  OR2 OR2_44(.VSS(VSS),.VDD(VDD),.Y(g3873),.A(g3649),.B(g3657));
  OR2 OR2_45(.VSS(VSS),.VDD(VDD),.Y(g3877),.A(g3651),.B(g3659));
  OR2 OR2_46(.VSS(VSS),.VDD(VDD),.Y(g3878),.A(g3703),.B(g3191));
  OR2 OR2_47(.VSS(VSS),.VDD(VDD),.Y(g3879),.A(g3704),.B(g3195));
  OR2 OR2_48(.VSS(VSS),.VDD(VDD),.Y(g3880),.A(g3658),.B(g3665));
  OR2 OR2_49(.VSS(VSS),.VDD(VDD),.Y(g3883),.A(g3709),.B(g3203));
  OR2 OR2_50(.VSS(VSS),.VDD(VDD),.Y(g3884),.A(g3666),.B(g3671));
  OR2 OR2_51(.VSS(VSS),.VDD(VDD),.Y(g3888),.A(g3672),.B(g3682));
  OR2 OR2_52(.VSS(VSS),.VDD(VDD),.Y(g3891),.A(g3683),.B(g3688));
  OR2 OR2_53(.VSS(VSS),.VDD(VDD),.Y(g3896),.A(g3689),.B(g3697));
  OR2 OR2_54(.VSS(VSS),.VDD(VDD),.Y(g3913),.A(g3449),.B(g2860));
  OR2 OR2_55(.VSS(VSS),.VDD(VDD),.Y(g3935),.A(g3464),.B(g2868));
  OR2 OR2_56(.VSS(VSS),.VDD(VDD),.Y(g3941),.A(g3479),.B(g2873));
  OR2 OR2_57(.VSS(VSS),.VDD(VDD),.Y(g3942),.A(g3215),.B(g3575));
  OR2 OR2_58(.VSS(VSS),.VDD(VDD),.Y(g3954),.A(g3484),.B(g3489));
  OR2 OR2_59(.VSS(VSS),.VDD(VDD),.Y(g3964),.A(g3634),.B(g3089));
  OR2 OR2_60(.VSS(VSS),.VDD(VDD),.Y(g3971),.A(g3644),.B(g3099));
  OR2 OR2_61(.VSS(VSS),.VDD(VDD),.Y(g3972),.A(g3646),.B(g3103));
  OR2 OR2_62(.VSS(VSS),.VDD(VDD),.Y(g3977),.A(g3653),.B(g3113));
  OR2 OR2_63(.VSS(VSS),.VDD(VDD),.Y(g3978),.A(g3655),.B(g3117));
  OR2 OR2_64(.VSS(VSS),.VDD(VDD),.Y(g3981),.A(g3661),.B(g3123));
  OR2 OR2_65(.VSS(VSS),.VDD(VDD),.Y(g3982),.A(g3663),.B(g3127));
  OR2 OR2_66(.VSS(VSS),.VDD(VDD),.Y(g3986),.A(g3667),.B(g3133));
  OR2 OR2_67(.VSS(VSS),.VDD(VDD),.Y(g3987),.A(g3669),.B(g3134));
  OR2 OR2_68(.VSS(VSS),.VDD(VDD),.Y(g3988),.A(g3678),.B(g3143));
  OR2 OR2_69(.VSS(VSS),.VDD(VDD),.Y(g3989),.A(g3679),.B(g3144));
  OR2 OR2_70(.VSS(VSS),.VDD(VDD),.Y(g3990),.A(g3684),.B(g3155));
  OR2 OR2_71(.VSS(VSS),.VDD(VDD),.Y(g3991),.A(g3685),.B(g3156));
  OR2 OR2_72(.VSS(VSS),.VDD(VDD),.Y(g3992),.A(g1555),.B(g3559));
  OR2 OR2_73(.VSS(VSS),.VDD(VDD),.Y(g3995),.A(g3690),.B(g3170));
  OR2 OR2_74(.VSS(VSS),.VDD(VDD),.Y(g3996),.A(g3691),.B(g3171));
  OR2 OR2_75(.VSS(VSS),.VDD(VDD),.Y(g3998),.A(g3698),.B(g3180));
  OR2 OR2_76(.VSS(VSS),.VDD(VDD),.Y(g3999),.A(g3699),.B(g3181));
  OR2 OR2_77(.VSS(VSS),.VDD(VDD),.Y(g4001),.A(g3702),.B(g3190));
  OR2 OR2_78(.VSS(VSS),.VDD(VDD),.Y(g4021),.A(g3558),.B(g2949));
  OR2 OR2_79(.VSS(VSS),.VDD(VDD),.Y(g4059),.A(g3466),.B(g3425));
  OR2 OR2_80(.VSS(VSS),.VDD(VDD),.Y(g4068),.A(g3293),.B(g2685));
  OR2 OR2_81(.VSS(VSS),.VDD(VDD),.Y(g4074),.A(g3301),.B(g2699));
  OR2 OR2_82(.VSS(VSS),.VDD(VDD),.Y(g4080),.A(g3302),.B(g2700));
  OR2 OR2_83(.VSS(VSS),.VDD(VDD),.Y(g4086),.A(g3310),.B(g2720));
  OR2 OR2_84(.VSS(VSS),.VDD(VDD),.Y(g4092),.A(g3311),.B(g2721));
  OR2 OR2_85(.VSS(VSS),.VDD(VDD),.Y(g4205),.A(g3843),.B(g541));
  OR2 OR2_86(.VSS(VSS),.VDD(VDD),.Y(g4231),.A(g3997),.B(g4000));
  OR2 OR2_87(.VSS(VSS),.VDD(VDD),.Y(g4233),.A(g3912),.B(g471));
  OR2 OR2_88(.VSS(VSS),.VDD(VDD),.Y(g4234),.A(g3921),.B(g478));
  OR2 OR2_89(.VSS(VSS),.VDD(VDD),.Y(g4243),.A(g4053),.B(g4058));
  OR2 OR2_90(.VSS(VSS),.VDD(VDD),.Y(g4285),.A(g3490),.B(g3887));
  OR2 OR2_91(.VSS(VSS),.VDD(VDD),.Y(g4427),.A(g4373),.B(g3668));
  OR2 OR2_92(.VSS(VSS),.VDD(VDD),.Y(g4430),.A(g4349),.B(g4015));
  OR2 OR2_93(.VSS(VSS),.VDD(VDD),.Y(g4433),.A(g4354),.B(g4032));
  OR2 OR2_94(.VSS(VSS),.VDD(VDD),.Y(g4434),.A(g4355),.B(g4033));
  OR2 OR2_95(.VSS(VSS),.VDD(VDD),.Y(g4436),.A(g4359),.B(g4035));
  OR2 OR2_96(.VSS(VSS),.VDD(VDD),.Y(g4438),.A(g4363),.B(g4037));
  OR2 OR2_97(.VSS(VSS),.VDD(VDD),.Y(g4440),.A(g4371),.B(g4038));
  OR2 OR2_98(.VSS(VSS),.VDD(VDD),.Y(g4441),.A(g4372),.B(g4039));
  OR2 OR2_99(.VSS(VSS),.VDD(VDD),.Y(g4443),.A(g4377),.B(g4041));
  OR2 OR2_100(.VSS(VSS),.VDD(VDD),.Y(g4444),.A(g4378),.B(g4042));
  OR2 OR2_101(.VSS(VSS),.VDD(VDD),.Y(g4446),.A(g4383),.B(g4043));
  OR2 OR2_102(.VSS(VSS),.VDD(VDD),.Y(g4447),.A(g4384),.B(g4044));
  OR2 OR2_103(.VSS(VSS),.VDD(VDD),.Y(g4450),.A(g4389),.B(g4047));
  OR2 OR2_104(.VSS(VSS),.VDD(VDD),.Y(g4451),.A(g4390),.B(g4048));
  OR2 OR2_105(.VSS(VSS),.VDD(VDD),.Y(g4454),.A(g4395),.B(g4051));
  OR2 OR2_106(.VSS(VSS),.VDD(VDD),.Y(g4455),.A(g4396),.B(g4052));
  OR2 OR2_107(.VSS(VSS),.VDD(VDD),.Y(g4458),.A(g4401),.B(g4057));
  OR2 OR2_108(.VSS(VSS),.VDD(VDD),.Y(g4468),.A(g4214),.B(g3831));
  OR2 OR2_109(.VSS(VSS),.VDD(VDD),.Y(g4473),.A(g3575),.B(g4253));
  OR2 OR2_110(.VSS(VSS),.VDD(VDD),.Y(g4497),.A(g4166),.B(g3784));
  OR2 OR2_111(.VSS(VSS),.VDD(VDD),.Y(g4500),.A(g4243),.B(g2010));
  OR2 OR2_112(.VSS(VSS),.VDD(VDD),.Y(g4544),.A(g4410),.B(g2995));
  OR2 OR2_113(.VSS(VSS),.VDD(VDD),.Y(g4549),.A(g4416),.B(g3013));
  OR2 OR2_114(.VSS(VSS),.VDD(VDD),.Y(g4599),.A(g3499),.B(g4230));
  OR2 OR2_115(.VSS(VSS),.VDD(VDD),.Y(g4607),.A(g4232),.B(g3899));
  OR2 OR2_116(.VSS(VSS),.VDD(VDD),.Y(g4627),.A(g4333),.B(g3603));
  OR2 OR2_117(.VSS(VSS),.VDD(VDD),.Y(g4630),.A(g4339),.B(g3610));
  OR2 OR2_118(.VSS(VSS),.VDD(VDD),.Y(g4631),.A(g4340),.B(g3611));
  OR2 OR2_119(.VSS(VSS),.VDD(VDD),.Y(g4634),.A(g4341),.B(g3615));
  OR2 OR2_120(.VSS(VSS),.VDD(VDD),.Y(g4635),.A(g4342),.B(g3616));
  OR2 OR2_121(.VSS(VSS),.VDD(VDD),.Y(g4637),.A(g4344),.B(g3619));
  OR2 OR2_122(.VSS(VSS),.VDD(VDD),.Y(g4638),.A(g4345),.B(g3620));
  OR2 OR2_123(.VSS(VSS),.VDD(VDD),.Y(g4641),.A(g4347),.B(g3627));
  OR2 OR2_124(.VSS(VSS),.VDD(VDD),.Y(g4642),.A(g4348),.B(g3628));
  OR2 OR2_125(.VSS(VSS),.VDD(VDD),.Y(g4645),.A(g4352),.B(g3633));
  OR2 OR2_126(.VSS(VSS),.VDD(VDD),.Y(g4646),.A(g4353),.B(g3635));
  OR2 OR2_127(.VSS(VSS),.VDD(VDD),.Y(g4651),.A(g4357),.B(g3643));
  OR2 OR2_128(.VSS(VSS),.VDD(VDD),.Y(g4652),.A(g4358),.B(g3645));
  OR2 OR2_129(.VSS(VSS),.VDD(VDD),.Y(g4653),.A(g4361),.B(g3652));
  OR2 OR2_130(.VSS(VSS),.VDD(VDD),.Y(g4654),.A(g4362),.B(g3654));
  OR2 OR2_131(.VSS(VSS),.VDD(VDD),.Y(g4655),.A(g4368),.B(g3660));
  OR2 OR2_132(.VSS(VSS),.VDD(VDD),.Y(g4656),.A(g4369),.B(g3662));
  OR2 OR2_133(.VSS(VSS),.VDD(VDD),.Y(g4740),.A(g4448),.B(g4154));
  OR2 OR2_134(.VSS(VSS),.VDD(VDD),.Y(g4745),.A(g4468),.B(g4569));
  OR2 OR2_135(.VSS(VSS),.VDD(VDD),.Y(g4752),.A(g4452),.B(g4155));
  OR2 OR2_136(.VSS(VSS),.VDD(VDD),.Y(g4757),.A(g4456),.B(g4158));
  OR2 OR2_137(.VSS(VSS),.VDD(VDD),.Y(g4773),.A(g4495),.B(g4220));
  OR2 OR2_138(.VSS(VSS),.VDD(VDD),.Y(g4811),.A(g4429),.B(g4432));
  OR2 OR2_139(.VSS(VSS),.VDD(VDD),.Y(g4859),.A(g4730),.B(g4486));
  OR2 OR2_140(.VSS(VSS),.VDD(VDD),.Y(g4860),.A(g4735),.B(g4488));
  OR2 OR2_141(.VSS(VSS),.VDD(VDD),.Y(g4862),.A(g4739),.B(g4489));
  OR2 OR2_142(.VSS(VSS),.VDD(VDD),.Y(g4864),.A(g4744),.B(g4490));
  OR2 OR2_143(.VSS(VSS),.VDD(VDD),.Y(g4866),.A(g4756),.B(g4491));
  OR2 OR2_144(.VSS(VSS),.VDD(VDD),.Y(g4936),.A(g4827),.B(g4828));
  OR2 OR2_145(.VSS(VSS),.VDD(VDD),.Y(g4941),.A(g4829),.B(g4832));
  OR2 OR2_146(.VSS(VSS),.VDD(VDD),.Y(g4946),.A(g4830),.B(g4833));
  OR2 OR2_147(.VSS(VSS),.VDD(VDD),.Y(g4948),.A(g4834),.B(g4836));
  OR2 OR2_148(.VSS(VSS),.VDD(VDD),.Y(g5012),.A(g4782),.B(g4580));
  OR2 OR2_149(.VSS(VSS),.VDD(VDD),.Y(g5013),.A(g4826),.B(g4621));
  OR2 OR2_150(.VSS(VSS),.VDD(VDD),.Y(g5014),.A(g4785),.B(g4583));
  OR2 OR2_151(.VSS(VSS),.VDD(VDD),.Y(g5015),.A(g4787),.B(g4588));
  OR2 OR2_152(.VSS(VSS),.VDD(VDD),.Y(g5016),.A(g4789),.B(g4592));
  OR2 OR2_153(.VSS(VSS),.VDD(VDD),.Y(g5018),.A(g4791),.B(g4597));
  OR2 OR2_154(.VSS(VSS),.VDD(VDD),.Y(g5024),.A(g4793),.B(g4600));
  OR2 OR2_155(.VSS(VSS),.VDD(VDD),.Y(g5044),.A(g4797),.B(g4602));
  OR2 OR2_156(.VSS(VSS),.VDD(VDD),.Y(g5060),.A(g3491),.B(g4819));
  OR2 OR2_157(.VSS(VSS),.VDD(VDD),.Y(g5062),.A(g4661),.B(g4666));
  OR2 OR2_158(.VSS(VSS),.VDD(VDD),.Y(g5065),.A(g4667),.B(g4671));
  OR2 OR2_159(.VSS(VSS),.VDD(VDD),.Y(g5066),.A(g4668),.B(g4672));
  OR2 OR2_160(.VSS(VSS),.VDD(VDD),.Y(g5068),.A(g4673),.B(g4677));
  OR2 OR2_161(.VSS(VSS),.VDD(VDD),.Y(g5069),.A(g1595),.B(g4688));
  OR2 OR2_162(.VSS(VSS),.VDD(VDD),.Y(g5074),.A(g4792),.B(g4598));
  OR2 OR2_163(.VSS(VSS),.VDD(VDD),.Y(g5077),.A(g1612),.B(g4694));
  OR2 OR2_164(.VSS(VSS),.VDD(VDD),.Y(g5083),.A(g4688),.B(g4271));
  OR2 OR2_165(.VSS(VSS),.VDD(VDD),.Y(g5085),.A(g4694),.B(g4280));
  OR3 OR3_0(.VSS(VSS),.VDD(VDD),.Y(g5202),.A(g4904),.B(g4914),.C(g4894));
  OR2 OR2_166(.VSS(VSS),.VDD(VDD),.Y(g5224),.A(g5123),.B(g3630));
  OR2 OR2_167(.VSS(VSS),.VDD(VDD),.Y(g5228),.A(g5096),.B(g4800));
  OR2 OR2_168(.VSS(VSS),.VDD(VDD),.Y(g5231),.A(g5048),.B(g672));
  OR2 OR2_169(.VSS(VSS),.VDD(VDD),.Y(g5241),.A(g5069),.B(g2067));
  OR2 OR2_170(.VSS(VSS),.VDD(VDD),.Y(g5246),.A(g5077),.B(g2080));
  OR2 OR2_171(.VSS(VSS),.VDD(VDD),.Y(g5277),.A(g5023),.B(g4763));
  OR2 OR2_172(.VSS(VSS),.VDD(VDD),.Y(g5281),.A(g5074),.B(g5124));
  OR2 OR2_173(.VSS(VSS),.VDD(VDD),.Y(g5291),.A(g5043),.B(g4764));
  OR2 OR2_174(.VSS(VSS),.VDD(VDD),.Y(g5295),.A(g5047),.B(g4766));
  OR2 OR2_175(.VSS(VSS),.VDD(VDD),.Y(g5303),.A(g5053),.B(g4768));
  OR2 OR2_176(.VSS(VSS),.VDD(VDD),.Y(g5323),.A(g5098),.B(g4802));
  OR3 OR3_1(.VSS(VSS),.VDD(VDD),.Y(g5326),.A(g5069),.B(g4410),.C(g3012));
  OR3 OR3_2(.VSS(VSS),.VDD(VDD),.Y(g5327),.A(g5077),.B(g4416),.C(g3028));
  OR2 OR2_177(.VSS(VSS),.VDD(VDD),.Y(g5348),.A(g5317),.B(g5122));
  OR2 OR2_178(.VSS(VSS),.VDD(VDD),.Y(g5367),.A(g5199),.B(g4928));
  OR2 OR2_179(.VSS(VSS),.VDD(VDD),.Y(g5368),.A(g5201),.B(g4932));
  OR2 OR2_180(.VSS(VSS),.VDD(VDD),.Y(g5370),.A(g5211),.B(g4937));
  OR2 OR2_181(.VSS(VSS),.VDD(VDD),.Y(g5372),.A(g5213),.B(g4942));
  OR2 OR2_182(.VSS(VSS),.VDD(VDD),.Y(g5374),.A(g5215),.B(g4947));
  OR2 OR2_183(.VSS(VSS),.VDD(VDD),.Y(g5377),.A(g5217),.B(g4949));
  OR2 OR2_184(.VSS(VSS),.VDD(VDD),.Y(g5385),.A(g3992),.B(g5318));
  OR2 OR2_185(.VSS(VSS),.VDD(VDD),.Y(g5386),.A(g5227),.B(g669));
  OR3 OR3_3(.VSS(VSS),.VDD(VDD),.Y(g5388),.A(g5318),.B(g1589),.C(g3491));
  OR2 OR2_186(.VSS(VSS),.VDD(VDD),.Y(g5430),.A(g5161),.B(g4873));
  OR2 OR2_187(.VSS(VSS),.VDD(VDD),.Y(g5458),.A(g3466),.B(g5311));
  OR3 OR3_4(.VSS(VSS),.VDD(VDD),.Y(g5467),.A(g3868),.B(g5318),.C(g3992));
  OR2 OR2_188(.VSS(VSS),.VDD(VDD),.Y(g5470),.A(g5359),.B(g5142));
  OR2 OR2_189(.VSS(VSS),.VDD(VDD),.Y(g5471),.A(g5360),.B(g5143));
  OR2 OR2_190(.VSS(VSS),.VDD(VDD),.Y(g5472),.A(g5361),.B(g5144));
  OR2 OR2_191(.VSS(VSS),.VDD(VDD),.Y(g5473),.A(g5362),.B(g5145));
  OR2 OR2_192(.VSS(VSS),.VDD(VDD),.Y(g5474),.A(g5363),.B(g5146));
  OR2 OR2_193(.VSS(VSS),.VDD(VDD),.Y(g5531),.A(g5349),.B(g3275));
  OR2 OR2_194(.VSS(VSS),.VDD(VDD),.Y(g5532),.A(g5350),.B(g3278));
  OR2 OR2_195(.VSS(VSS),.VDD(VDD),.Y(g5533),.A(g5351),.B(g3290));
  OR2 OR2_196(.VSS(VSS),.VDD(VDD),.Y(g5535),.A(g5353),.B(g3300));
  OR2 OR2_197(.VSS(VSS),.VDD(VDD),.Y(g5583),.A(g5569),.B(g4020));
  OR2 OR2_198(.VSS(VSS),.VDD(VDD),.Y(g5605),.A(g3575),.B(g5500));
  OR2 OR2_199(.VSS(VSS),.VDD(VDD),.Y(g5622),.A(g5492),.B(g3277));
  OR2 OR2_200(.VSS(VSS),.VDD(VDD),.Y(g5623),.A(g5503),.B(g5357));
  OR2 OR2_201(.VSS(VSS),.VDD(VDD),.Y(g5624),.A(g5494),.B(g3280));
  OR2 OR2_202(.VSS(VSS),.VDD(VDD),.Y(g5625),.A(g5495),.B(g3281));
  OR2 OR2_203(.VSS(VSS),.VDD(VDD),.Y(g5626),.A(g5496),.B(g3285));
  OR2 OR2_204(.VSS(VSS),.VDD(VDD),.Y(g5627),.A(g5497),.B(g3286));
  OR2 OR2_205(.VSS(VSS),.VDD(VDD),.Y(g5628),.A(g5498),.B(g3292));
  OR2 OR2_206(.VSS(VSS),.VDD(VDD),.Y(g5629),.A(g5499),.B(g3298));
  OR2 OR2_207(.VSS(VSS),.VDD(VDD),.Y(g5630),.A(g5501),.B(g3309));
  OR2 OR2_208(.VSS(VSS),.VDD(VDD),.Y(g5659),.A(g5551),.B(g5398));
  OR2 OR2_209(.VSS(VSS),.VDD(VDD),.Y(g5662),.A(g5553),.B(g5402));
  OR2 OR2_210(.VSS(VSS),.VDD(VDD),.Y(g5666),.A(g5555),.B(g5406));
  OR2 OR2_211(.VSS(VSS),.VDD(VDD),.Y(g5669),.A(g5556),.B(g5410));
  OR2 OR2_212(.VSS(VSS),.VDD(VDD),.Y(g5672),.A(g5557),.B(g5414));
  OR2 OR2_213(.VSS(VSS),.VDD(VDD),.Y(g5674),.A(g5558),.B(g5419));
  OR2 OR2_214(.VSS(VSS),.VDD(VDD),.Y(g5676),.A(g5559),.B(g5424));
  OR2 OR2_215(.VSS(VSS),.VDD(VDD),.Y(g5678),.A(g5560),.B(g5428));
  OR2 OR2_216(.VSS(VSS),.VDD(VDD),.Y(g5680),.A(g5562),.B(g5429));
  OR2 OR2_217(.VSS(VSS),.VDD(VDD),.Y(g5693),.A(g5632),.B(g5481));
  OR2 OR2_218(.VSS(VSS),.VDD(VDD),.Y(g5694),.A(g5633),.B(g5482));
  OR2 OR2_219(.VSS(VSS),.VDD(VDD),.Y(g5695),.A(g5635),.B(g5483));
  OR2 OR2_220(.VSS(VSS),.VDD(VDD),.Y(g5696),.A(g5637),.B(g5484));
  OR2 OR2_221(.VSS(VSS),.VDD(VDD),.Y(g5697),.A(g5646),.B(g5485));
  OR2 OR2_222(.VSS(VSS),.VDD(VDD),.Y(g5698),.A(g5648),.B(g5486));
  OR2 OR2_223(.VSS(VSS),.VDD(VDD),.Y(g5699),.A(g5660),.B(g5487));
  OR2 OR2_224(.VSS(VSS),.VDD(VDD),.Y(g5700),.A(g5663),.B(g5488));
  OR2 OR2_225(.VSS(VSS),.VDD(VDD),.Y(g5800),.A(g5369),.B(g5600));
  OR2 OR2_226(.VSS(VSS),.VDD(VDD),.Y(g5804),.A(g5371),.B(g5603));
  OR2 OR2_227(.VSS(VSS),.VDD(VDD),.Y(g5808),.A(g5373),.B(g5616));
  OR2 OR2_228(.VSS(VSS),.VDD(VDD),.Y(g5812),.A(g5376),.B(g5618));
  OR2 OR2_229(.VSS(VSS),.VDD(VDD),.Y(g5816),.A(g5378),.B(g5620));
  OR2 OR2_230(.VSS(VSS),.VDD(VDD),.Y(g5817),.A(g5380),.B(g5621));
  OR2 OR2_231(.VSS(VSS),.VDD(VDD),.Y(g5916),.A(g5728),.B(g3781));
  OR2 OR2_232(.VSS(VSS),.VDD(VDD),.Y(g6108),.A(g5898),.B(g5598));
  OR2 OR2_233(.VSS(VSS),.VDD(VDD),.Y(g6109),.A(g5900),.B(g5599));
  OR2 OR2_234(.VSS(VSS),.VDD(VDD),.Y(g6110),.A(g5883),.B(g5996));
  OR2 OR2_235(.VSS(VSS),.VDD(VDD),.Y(g6113),.A(g5902),.B(g5601));
  OR2 OR2_236(.VSS(VSS),.VDD(VDD),.Y(g6114),.A(g5904),.B(g5604));
  OR2 OR2_237(.VSS(VSS),.VDD(VDD),.Y(g6116),.A(g5910),.B(g5617));
  OR2 OR2_238(.VSS(VSS),.VDD(VDD),.Y(g6118),.A(g5911),.B(g5619));
  OR2 OR2_239(.VSS(VSS),.VDD(VDD),.Y(g6142),.A(g5909),.B(g3806));
  OR2 OR2_240(.VSS(VSS),.VDD(VDD),.Y(g6167),.A(g6056),.B(g6039));
  OR2 OR2_241(.VSS(VSS),.VDD(VDD),.Y(g6170),.A(g6061),.B(g6014));
  OR2 OR2_242(.VSS(VSS),.VDD(VDD),.Y(g6173),.A(g6066),.B(g6043));
  OR2 OR2_243(.VSS(VSS),.VDD(VDD),.Y(g6176),.A(g6068),.B(g6033));
  OR2 OR2_244(.VSS(VSS),.VDD(VDD),.Y(g6179),.A(g6077),.B(g6051));
  OR2 OR2_245(.VSS(VSS),.VDD(VDD),.Y(g6182),.A(g6047),.B(g6034));
  OR2 OR2_246(.VSS(VSS),.VDD(VDD),.Y(g6185),.A(g6055),.B(g5995));
  OR2 OR2_247(.VSS(VSS),.VDD(VDD),.Y(g6189),.A(g6060),.B(g6035));
  OR2 OR2_248(.VSS(VSS),.VDD(VDD),.Y(g6237),.A(g5912),.B(g2381));
  OR2 OR2_249(.VSS(VSS),.VDD(VDD),.Y(g6239),.A(g2339),.B(g6073));
  OR2 OR2_250(.VSS(VSS),.VDD(VDD),.Y(g6242),.A(g2356),.B(g6075));
  OR2 OR2_251(.VSS(VSS),.VDD(VDD),.Y(g6246),.A(g5665),.B(g5937));
  OR2 OR2_252(.VSS(VSS),.VDD(VDD),.Y(g6251),.A(g5668),.B(g5939));
  OR2 OR2_253(.VSS(VSS),.VDD(VDD),.Y(g6252),.A(g5905),.B(g2381));
  OR2 OR2_254(.VSS(VSS),.VDD(VDD),.Y(g6257),.A(g5671),.B(g5941));
  OR2 OR2_255(.VSS(VSS),.VDD(VDD),.Y(g6261),.A(g5673),.B(g5944));
  OR2 OR2_256(.VSS(VSS),.VDD(VDD),.Y(g6264),.A(g5675),.B(g5948));
  OR2 OR2_257(.VSS(VSS),.VDD(VDD),.Y(g6267),.A(g2953),.B(g5884));
  OR2 OR2_258(.VSS(VSS),.VDD(VDD),.Y(g6268),.A(g5677),.B(g5951));
  OR2 OR2_259(.VSS(VSS),.VDD(VDD),.Y(g6271),.A(g2955),.B(g5885));
  OR2 OR2_260(.VSS(VSS),.VDD(VDD),.Y(g6272),.A(g5679),.B(g5953));
  OR2 OR2_261(.VSS(VSS),.VDD(VDD),.Y(g6273),.A(g5681),.B(g5955));
  OR2 OR2_262(.VSS(VSS),.VDD(VDD),.Y(g6274),.A(g5682),.B(g5956));
  OR4 OR4_0(.VSS(VSS),.VDD(VDD),.Y(I7969),.A(g6194),.B(g5958),.C(g5975),.D(g5997));
  OR4 OR4_1(.VSS(VSS),.VDD(VDD),.Y(I7970),.A(g6015),.B(g6212),.C(g4950),.D(g4877));
  OR4 OR4_2(.VSS(VSS),.VDD(VDD),.Y(I7971),.A(g5202),.B(g4993),.C(g4967),.D(g4980));
  OR2 OR2_263(.VSS(VSS),.VDD(VDD),.Y(I7972),.A(g4915),.B(g5025));
  OR4 OR4_3(.VSS(VSS),.VDD(VDD),.Y(I7978),.A(g6194),.B(g5958),.C(g5975),.D(g5997));
  OR4 OR4_4(.VSS(VSS),.VDD(VDD),.Y(I7979),.A(g6015),.B(g6212),.C(g4950),.D(g4877));
  OR4 OR4_5(.VSS(VSS),.VDD(VDD),.Y(I7980),.A(g5202),.B(g4993),.C(g4967),.D(g4980));
  OR2 OR2_264(.VSS(VSS),.VDD(VDD),.Y(I7981),.A(g4915),.B(g5025));
  OR4 OR4_6(.VSS(VSS),.VDD(VDD),.Y(I7987),.A(g6194),.B(g5958),.C(g5975),.D(g5997));
  OR4 OR4_7(.VSS(VSS),.VDD(VDD),.Y(I7988),.A(g6015),.B(g6212),.C(g4950),.D(g4877));
  OR4 OR4_8(.VSS(VSS),.VDD(VDD),.Y(I7989),.A(g5202),.B(g4993),.C(g4967),.D(g4980));
  OR2 OR2_265(.VSS(VSS),.VDD(VDD),.Y(I7990),.A(g4915),.B(g5025));
  OR2 OR2_266(.VSS(VSS),.VDD(VDD),.Y(g6286),.A(g6238),.B(g6079));
  OR2 OR2_267(.VSS(VSS),.VDD(VDD),.Y(g6287),.A(g6241),.B(g6082));
  OR2 OR2_268(.VSS(VSS),.VDD(VDD),.Y(g6289),.A(g6240),.B(g6081));
  OR2 OR2_269(.VSS(VSS),.VDD(VDD),.Y(g6290),.A(g6245),.B(g6086));
  OR2 OR2_270(.VSS(VSS),.VDD(VDD),.Y(g6292),.A(g6243),.B(g6084));
  OR2 OR2_271(.VSS(VSS),.VDD(VDD),.Y(g6293),.A(g6244),.B(g6085));
  OR2 OR2_272(.VSS(VSS),.VDD(VDD),.Y(g6294),.A(g6249),.B(g6090));
  OR2 OR2_273(.VSS(VSS),.VDD(VDD),.Y(g6296),.A(g6247),.B(g6088));
  OR2 OR2_274(.VSS(VSS),.VDD(VDD),.Y(g6297),.A(g6248),.B(g6089));
  OR2 OR2_275(.VSS(VSS),.VDD(VDD),.Y(g6298),.A(g6255),.B(g6093));
  OR2 OR2_276(.VSS(VSS),.VDD(VDD),.Y(g6300),.A(g6253),.B(g6091));
  OR2 OR2_277(.VSS(VSS),.VDD(VDD),.Y(g6301),.A(g6254),.B(g6092));
  OR2 OR2_278(.VSS(VSS),.VDD(VDD),.Y(g6303),.A(g6258),.B(g6094));
  OR2 OR2_279(.VSS(VSS),.VDD(VDD),.Y(g6307),.A(g6262),.B(g6096));
  OR2 OR2_280(.VSS(VSS),.VDD(VDD),.Y(g6309),.A(g6265),.B(g6098));
  OR2 OR2_281(.VSS(VSS),.VDD(VDD),.Y(g6310),.A(g6269),.B(g6099));
  OR4 OR4_9(.VSS(VSS),.VDD(VDD),.Y(I8079),.A(g6194),.B(g5958),.C(g5975),.D(g5997));
  OR4 OR4_10(.VSS(VSS),.VDD(VDD),.Y(I8080),.A(g6015),.B(g6212),.C(g4950),.D(g4877));
  OR4 OR4_11(.VSS(VSS),.VDD(VDD),.Y(I8081),.A(g4894),.B(g4904),.C(g4993),.D(g4967));
  OR4 OR4_12(.VSS(VSS),.VDD(VDD),.Y(I8082),.A(g4980),.B(g4915),.C(g5025),.D(g5054));
  OR4 OR4_13(.VSS(VSS),.VDD(VDD),.Y(I8117),.A(g6194),.B(g5958),.C(g5975),.D(g5997));
  OR4 OR4_14(.VSS(VSS),.VDD(VDD),.Y(I8118),.A(g6015),.B(g6212),.C(g4950),.D(g4877));
  OR4 OR4_15(.VSS(VSS),.VDD(VDD),.Y(I8119),.A(g5202),.B(g4993),.C(g4967),.D(g4980));
  OR2 OR2_282(.VSS(VSS),.VDD(VDD),.Y(I8120),.A(g4915),.B(g5025));
  OR4 OR4_16(.VSS(VSS),.VDD(VDD),.Y(I8126),.A(g6194),.B(g5958),.C(g5975),.D(g5997));
  OR4 OR4_17(.VSS(VSS),.VDD(VDD),.Y(I8127),.A(g6015),.B(g6212),.C(g4950),.D(g4877));
  OR4 OR4_18(.VSS(VSS),.VDD(VDD),.Y(I8128),.A(g5202),.B(g4993),.C(g4967),.D(g4980));
  OR2 OR2_283(.VSS(VSS),.VDD(VDD),.Y(I8129),.A(g4915),.B(g5025));
  OR4 OR4_19(.VSS(VSS),.VDD(VDD),.Y(I8135),.A(g6194),.B(g5958),.C(g5975),.D(g5997));
  OR4 OR4_20(.VSS(VSS),.VDD(VDD),.Y(I8136),.A(g6015),.B(g6212),.C(g4950),.D(g4877));
  OR4 OR4_21(.VSS(VSS),.VDD(VDD),.Y(I8137),.A(g4894),.B(g4904),.C(g4993),.D(g4967));
  OR4 OR4_22(.VSS(VSS),.VDD(VDD),.Y(I8138),.A(g4980),.B(g4915),.C(g5025),.D(g5054));
  OR4 OR4_23(.VSS(VSS),.VDD(VDD),.Y(I8208),.A(g6194),.B(g5958),.C(g5975),.D(g5997));
  OR4 OR4_24(.VSS(VSS),.VDD(VDD),.Y(I8209),.A(g6015),.B(g6212),.C(g4950),.D(g4877));
  OR4 OR4_25(.VSS(VSS),.VDD(VDD),.Y(I8210),.A(g5202),.B(g4993),.C(g4967),.D(g4980));
  OR2 OR2_284(.VSS(VSS),.VDD(VDD),.Y(I8211),.A(g4915),.B(g5025));
  OR2 OR2_285(.VSS(VSS),.VDD(VDD),.Y(g6426),.A(g6288),.B(g6119));
  OR2 OR2_286(.VSS(VSS),.VDD(VDD),.Y(g6437),.A(g6302),.B(g6121));
  OR2 OR2_287(.VSS(VSS),.VDD(VDD),.Y(g6440),.A(g6336),.B(g5935));
  OR2 OR2_288(.VSS(VSS),.VDD(VDD),.Y(g6444),.A(g6338),.B(g5936));
  OR2 OR2_289(.VSS(VSS),.VDD(VDD),.Y(g6447),.A(g6340),.B(g5938));
  OR2 OR2_290(.VSS(VSS),.VDD(VDD),.Y(g6450),.A(g6341),.B(g5940));
  OR2 OR2_291(.VSS(VSS),.VDD(VDD),.Y(g6452),.A(g6342),.B(g5942));
  OR2 OR2_292(.VSS(VSS),.VDD(VDD),.Y(g6453),.A(g6343),.B(g5945));
  OR2 OR2_293(.VSS(VSS),.VDD(VDD),.Y(g6454),.A(g6344),.B(g5949));
  OR2 OR2_294(.VSS(VSS),.VDD(VDD),.Y(g6455),.A(g6345),.B(g5952));
  OR2 OR2_295(.VSS(VSS),.VDD(VDD),.Y(g6456),.A(g6346),.B(g5954));
  OR2 OR2_296(.VSS(VSS),.VDD(VDD),.Y(g6457),.A(g6352),.B(g6347));
  OR2 OR2_297(.VSS(VSS),.VDD(VDD),.Y(g6461),.A(g6353),.B(g6351));
  OR4 OR4_26(.VSS(VSS),.VDD(VDD),.Y(I8345),.A(g6326),.B(g6135),.C(g6140),.D(g6157));
  OR4 OR4_27(.VSS(VSS),.VDD(VDD),.Y(I8346),.A(g6159),.B(g6334),.C(g5163),.D(g5191));
  OR4 OR4_28(.VSS(VSS),.VDD(VDD),.Y(I8347),.A(g5188),.B(g5157),.C(g5154),.D(g5193));
  OR4 OR4_29(.VSS(VSS),.VDD(VDD),.Y(I8348),.A(g5229),.B(g5234),.C(g5218),.D(g5225));
  OR4 OR4_30(.VSS(VSS),.VDD(VDD),.Y(I8349),.A(I8345),.B(I8346),.C(I8347),.D(I8348));
  OR2 OR2_298(.VSS(VSS),.VDD(VDD),.Y(g6479),.A(I8349),.B(g6335));
  OR4 OR4_31(.VSS(VSS),.VDD(VDD),.Y(I8356),.A(g6311),.B(g6123),.C(g6125),.D(g6141));
  OR4 OR4_32(.VSS(VSS),.VDD(VDD),.Y(I8357),.A(g6145),.B(g6318),.C(g5171),.D(g5187));
  OR4 OR4_33(.VSS(VSS),.VDD(VDD),.Y(I8358),.A(g5192),.B(g5153),.C(g5158),.D(g5197));
  OR4 OR4_34(.VSS(VSS),.VDD(VDD),.Y(I8359),.A(g5232),.B(g5236),.C(g5216),.D(g5226));
  OR4 OR4_35(.VSS(VSS),.VDD(VDD),.Y(I8360),.A(I8356),.B(I8357),.C(I8358),.D(I8359));
  OR2 OR2_299(.VSS(VSS),.VDD(VDD),.Y(g6480),.A(I8360),.B(g6359));
  OR4 OR4_36(.VSS(VSS),.VDD(VDD),.Y(I8367),.A(g6313),.B(g6124),.C(g6127),.D(g6144));
  OR4 OR4_37(.VSS(VSS),.VDD(VDD),.Y(I8368),.A(g6148),.B(g6321),.C(g5176),.D(g5184));
  OR4 OR4_38(.VSS(VSS),.VDD(VDD),.Y(I8369),.A(g5165),.B(g5159),.C(g5233),.D(g5240));
  OR2 OR2_300(.VSS(VSS),.VDD(VDD),.Y(I8370),.A(g5214),.B(g6358));
  OR4 OR4_39(.VSS(VSS),.VDD(VDD),.Y(g6481),.A(I8367),.B(I8368),.C(I8369),.D(I8370));
  OR4 OR4_40(.VSS(VSS),.VDD(VDD),.Y(I8376),.A(g6315),.B(g6126),.C(g6129),.D(g6146));
  OR4 OR4_41(.VSS(VSS),.VDD(VDD),.Y(I8377),.A(g6150),.B(g6324),.C(g5180),.D(g5181));
  OR4 OR4_42(.VSS(VSS),.VDD(VDD),.Y(I8378),.A(g5173),.B(g5166),.C(g5235),.D(g5245));
  OR2 OR2_301(.VSS(VSS),.VDD(VDD),.Y(I8379),.A(g5212),.B(g6357));
  OR4 OR4_43(.VSS(VSS),.VDD(VDD),.Y(g6482),.A(I8376),.B(I8377),.C(I8378),.D(I8379));
  OR4 OR4_44(.VSS(VSS),.VDD(VDD),.Y(I8385),.A(g6316),.B(g6128),.C(g6131),.D(g6149));
  OR4 OR4_45(.VSS(VSS),.VDD(VDD),.Y(I8386),.A(g6152),.B(g6327),.C(g5183),.D(g5177));
  OR3 OR3_5(.VSS(VSS),.VDD(VDD),.Y(I8387),.A(g5178),.B(g5209),.C(g6281));
  OR3 OR3_6(.VSS(VSS),.VDD(VDD),.Y(g6483),.A(I8385),.B(I8386),.C(I8387));
  OR4 OR4_46(.VSS(VSS),.VDD(VDD),.Y(I8393),.A(g6317),.B(g6130),.C(g6133),.D(g6151));
  OR4 OR4_47(.VSS(VSS),.VDD(VDD),.Y(I8394),.A(g6154),.B(g6329),.C(g5186),.D(g5172));
  OR3 OR3_7(.VSS(VSS),.VDD(VDD),.Y(I8395),.A(g5182),.B(g5200),.C(g6280));
  OR3 OR3_8(.VSS(VSS),.VDD(VDD),.Y(g6485),.A(I8393),.B(I8394),.C(I8395));
  OR2 OR2_302(.VSS(VSS),.VDD(VDD),.Y(g6545),.A(g6468),.B(g4244));
  OR2 OR2_303(.VSS(VSS),.VDD(VDD),.Y(g6549),.A(g6473),.B(g4247));
  OR2 OR2_304(.VSS(VSS),.VDD(VDD),.Y(g6554),.A(g6337),.B(g6466));
  OR2 OR2_305(.VSS(VSS),.VDD(VDD),.Y(g6556),.A(g6339),.B(g6467));
  OR2 OR2_306(.VSS(VSS),.VDD(VDD),.Y(g6658),.A(g6132),.B(g6620));
  OR2 OR2_307(.VSS(VSS),.VDD(VDD),.Y(g6659),.A(g6634),.B(g6631));
  OR2 OR2_308(.VSS(VSS),.VDD(VDD),.Y(g6660),.A(g6640),.B(g6637));
  OR4 OR4_48(.VSS(VSS),.VDD(VDD),.Y(I8773),.A(g6610),.B(g6608),.C(g6606),.D(g6604));
  OR4 OR4_49(.VSS(VSS),.VDD(VDD),.Y(I8774),.A(g6655),.B(g6653),.C(g6651),.D(g6649));
  OR2 OR2_309(.VSS(VSS),.VDD(VDD),.Y(g6661),.A(I8773),.B(I8774));
  OR4 OR4_50(.VSS(VSS),.VDD(VDD),.Y(I8778),.A(g6612),.B(g6611),.C(g6609),.D(g6607));
  OR4 OR4_51(.VSS(VSS),.VDD(VDD),.Y(I8779),.A(g6605),.B(g6656),.C(g6654),.D(g6652));
  OR2 OR2_310(.VSS(VSS),.VDD(VDD),.Y(g6665),.A(I8778),.B(I8779));
  OR2 OR2_311(.VSS(VSS),.VDD(VDD),.Y(g6669),.A(g6613),.B(g4679));
  OR4 OR4_52(.VSS(VSS),.VDD(VDD),.Y(g6670),.A(g6557),.B(g6634),.C(g4410),.D(g2948));
  OR4 OR4_53(.VSS(VSS),.VDD(VDD),.Y(g6673),.A(g6559),.B(g6640),.C(g4416),.D(g2950));
  OR2 OR2_312(.VSS(VSS),.VDD(VDD),.Y(g6676),.A(g6631),.B(g6555));
  OR2 OR2_313(.VSS(VSS),.VDD(VDD),.Y(g6679),.A(g6637),.B(g6558));
  OR3 OR3_9(.VSS(VSS),.VDD(VDD),.Y(g6682),.A(g6478),.B(g6624),.C(g6623));
  OR3 OR3_10(.VSS(VSS),.VDD(VDD),.Y(g6683),.A(g6465),.B(g6622),.C(g6621));
  OR2 OR2_314(.VSS(VSS),.VDD(VDD),.Y(g6684),.A(g6250),.B(g6643));
  OR2 OR2_315(.VSS(VSS),.VDD(VDD),.Y(g6685),.A(g6256),.B(g6644));
  OR2 OR2_316(.VSS(VSS),.VDD(VDD),.Y(g6686),.A(g6259),.B(g6645));
  OR2 OR2_317(.VSS(VSS),.VDD(VDD),.Y(g6687),.A(g6260),.B(g6646));
  OR2 OR2_318(.VSS(VSS),.VDD(VDD),.Y(g6688),.A(g6263),.B(g6647));
  OR2 OR2_319(.VSS(VSS),.VDD(VDD),.Y(g6689),.A(g6266),.B(g6648));
  OR2 OR2_320(.VSS(VSS),.VDD(VDD),.Y(g6690),.A(g6270),.B(g6650));
  OR2 OR2_321(.VSS(VSS),.VDD(VDD),.Y(g6691),.A(g6275),.B(g6603));
  OR2 OR2_322(.VSS(VSS),.VDD(VDD),.Y(g6702),.A(g6659),.B(g496));
  OR2 OR2_323(.VSS(VSS),.VDD(VDD),.Y(g6703),.A(g6692),.B(g4831));
  OR2 OR2_324(.VSS(VSS),.VDD(VDD),.Y(g6704),.A(g6660),.B(g492));
  OR2 OR2_325(.VSS(VSS),.VDD(VDD),.Y(g6705),.A(g6693),.B(g4835));
  OR2 OR2_326(.VSS(VSS),.VDD(VDD),.Y(g6747),.A(g6614),.B(g6731));
  OR3 OR3_11(.VSS(VSS),.VDD(VDD),.Y(g6750),.A(g6670),.B(g6625),.C(g6736));
  OR3 OR3_12(.VSS(VSS),.VDD(VDD),.Y(g6754),.A(g6676),.B(g6625),.C(g6737));
  OR3 OR3_13(.VSS(VSS),.VDD(VDD),.Y(g6758),.A(g6673),.B(g6628),.C(g6738));
  OR3 OR3_14(.VSS(VSS),.VDD(VDD),.Y(g6762),.A(g6679),.B(g6628),.C(g6739));
  OR2 OR2_327(.VSS(VSS),.VDD(VDD),.Y(g6781),.A(g6718),.B(g6748));
  OR2 OR2_328(.VSS(VSS),.VDD(VDD),.Y(g6782),.A(g6719),.B(g6749));
  OR2 OR2_329(.VSS(VSS),.VDD(VDD),.Y(g6787),.A(g3758),.B(g6766));
  OR2 OR2_330(.VSS(VSS),.VDD(VDD),.Y(g6788),.A(g3760),.B(g6767));
  OR2 OR2_331(.VSS(VSS),.VDD(VDD),.Y(g6789),.A(g3764),.B(g6769));
  OR2 OR2_332(.VSS(VSS),.VDD(VDD),.Y(g6790),.A(g3765),.B(g6773));
  OR2 OR2_333(.VSS(VSS),.VDD(VDD),.Y(g6791),.A(g6768),.B(g3307));
  OR2 OR2_334(.VSS(VSS),.VDD(VDD),.Y(g6792),.A(g6770),.B(g3321));
  OR2 OR2_335(.VSS(VSS),.VDD(VDD),.Y(g6793),.A(g6771),.B(g3323));
  OR2 OR2_336(.VSS(VSS),.VDD(VDD),.Y(g6794),.A(g6777),.B(g3333));
  OR2 OR2_337(.VSS(VSS),.VDD(VDD),.Y(g6795),.A(g4867),.B(g6772));
  OR4 OR4_54(.VSS(VSS),.VDD(VDD),.Y(I9057),.A(g6320),.B(g6828),.C(g6830),.D(g6153));
  OR4 OR4_55(.VSS(VSS),.VDD(VDD),.Y(I9058),.A(g6156),.B(g6331),.C(g5190),.D(g5164));
  OR3 OR3_15(.VSS(VSS),.VDD(VDD),.Y(I9059),.A(g5185),.B(g5198),.C(g6279));
  OR3 OR3_16(.VSS(VSS),.VDD(VDD),.Y(g6844),.A(I9057),.B(I9058),.C(I9059));
  OR4 OR4_56(.VSS(VSS),.VDD(VDD),.Y(I9064),.A(g6323),.B(g6829),.C(g6831),.D(g6155));
  OR4 OR4_57(.VSS(VSS),.VDD(VDD),.Y(I9065),.A(g6158),.B(g6333),.C(g5152),.D(g5156));
  OR3 OR3_17(.VSS(VSS),.VDD(VDD),.Y(I9066),.A(g5189),.B(g5269),.C(g6400));
  OR3 OR3_18(.VSS(VSS),.VDD(VDD),.Y(g6845),.A(I9064),.B(I9065),.C(I9066));
  OR2 OR2_338(.VSS(VSS),.VDD(VDD),.Y(g6846),.A(g5860),.B(g6834));
  OR2 OR2_339(.VSS(VSS),.VDD(VDD),.Y(g6847),.A(g5861),.B(g6837));
  OR2 OR2_340(.VSS(VSS),.VDD(VDD),.Y(g6855),.A(g6851),.B(g2085));
  OR2 OR2_341(.VSS(VSS),.VDD(VDD),.Y(g6864),.A(g6852),.B(g2089));
  OR2 OR2_342(.VSS(VSS),.VDD(VDD),.Y(g6907),.A(g6874),.B(g3358));
  OR2 OR2_343(.VSS(VSS),.VDD(VDD),.Y(g6917),.A(g6909),.B(g6910));
  OR2 OR2_344(.VSS(VSS),.VDD(VDD),.Y(g6918),.A(g6911),.B(g6913));
  OR2 OR2_345(.VSS(VSS),.VDD(VDD),.Y(g6919),.A(g6912),.B(g6914));
  OR2 OR2_346(.VSS(VSS),.VDD(VDD),.Y(g6920),.A(g6915),.B(g6916));
  OR2 OR2_347(.VSS(VSS),.VDD(VDD),.Y(g6921),.A(g6908),.B(g6816));
  OR2 OR2_348(.VSS(VSS),.VDD(VDD),.Y(g6926),.A(g6798),.B(g6923));
  OR2 OR2_349(.VSS(VSS),.VDD(VDD),.Y(g6927),.A(g6799),.B(g6924));
  OR2 OR2_350(.VSS(VSS),.VDD(VDD),.Y(g6930),.A(g6740),.B(g6928));
  OR2 OR2_351(.VSS(VSS),.VDD(VDD),.Y(g6931),.A(g6741),.B(g6929));
  OR2 OR2_352(.VSS(VSS),.VDD(VDD),.Y(g6936),.A(g5438),.B(g6935));
  OR2 OR2_353(.VSS(VSS),.VDD(VDD),.Y(g6937),.A(g4616),.B(g6934));
//
  NAND2 NAND2_0(.VSS(VSS),.VDD(VDD),.Y(g901),.A(g314),.B(g310));
  NAND2 NAND2_1(.VSS(VSS),.VDD(VDD),.Y(g905),.A(g301),.B(g319));
  NAND2 NAND2_2(.VSS(VSS),.VDD(VDD),.Y(I1951),.A(g524),.B(g248));
  NAND2 NAND2_3(.VSS(VSS),.VDD(VDD),.Y(I1952),.A(g524),.B(I1951));
  NAND2 NAND2_4(.VSS(VSS),.VDD(VDD),.Y(I1953),.A(g248),.B(I1951));
  NAND2 NAND2_5(.VSS(VSS),.VDD(VDD),.Y(g926),.A(I1952),.B(I1953));
  NAND2 NAND2_6(.VSS(VSS),.VDD(VDD),.Y(I1961),.A(g520),.B(g242));
  NAND2 NAND2_7(.VSS(VSS),.VDD(VDD),.Y(I1962),.A(g520),.B(I1961));
  NAND2 NAND2_8(.VSS(VSS),.VDD(VDD),.Y(I1963),.A(g242),.B(I1961));
  NAND2 NAND2_9(.VSS(VSS),.VDD(VDD),.Y(g928),.A(I1962),.B(I1963));
  NAND2 NAND2_10(.VSS(VSS),.VDD(VDD),.Y(I1969),.A(g516),.B(g236));
  NAND2 NAND2_11(.VSS(VSS),.VDD(VDD),.Y(I1970),.A(g516),.B(I1969));
  NAND2 NAND2_12(.VSS(VSS),.VDD(VDD),.Y(I1971),.A(g236),.B(I1969));
  NAND2 NAND2_13(.VSS(VSS),.VDD(VDD),.Y(g930),.A(I1970),.B(I1971));
  NAND2 NAND2_14(.VSS(VSS),.VDD(VDD),.Y(I1978),.A(g512),.B(g230));
  NAND2 NAND2_15(.VSS(VSS),.VDD(VDD),.Y(I1979),.A(g512),.B(I1978));
  NAND2 NAND2_16(.VSS(VSS),.VDD(VDD),.Y(I1980),.A(g230),.B(I1978));
  NAND2 NAND2_17(.VSS(VSS),.VDD(VDD),.Y(g937),.A(I1979),.B(I1980));
  NAND2 NAND2_18(.VSS(VSS),.VDD(VDD),.Y(I1986),.A(g508),.B(g224));
  NAND2 NAND2_19(.VSS(VSS),.VDD(VDD),.Y(I1987),.A(g508),.B(I1986));
  NAND2 NAND2_20(.VSS(VSS),.VDD(VDD),.Y(I1988),.A(g224),.B(I1986));
  NAND2 NAND2_21(.VSS(VSS),.VDD(VDD),.Y(g939),.A(I1987),.B(I1988));
  NAND2 NAND2_22(.VSS(VSS),.VDD(VDD),.Y(I1994),.A(g504),.B(g218));
  NAND2 NAND2_23(.VSS(VSS),.VDD(VDD),.Y(I1995),.A(g504),.B(I1994));
  NAND2 NAND2_24(.VSS(VSS),.VDD(VDD),.Y(I1996),.A(g218),.B(I1994));
  NAND2 NAND2_25(.VSS(VSS),.VDD(VDD),.Y(g941),.A(I1995),.B(I1996));
  NAND2 NAND2_26(.VSS(VSS),.VDD(VDD),.Y(I2003),.A(g500),.B(g212));
  NAND2 NAND2_27(.VSS(VSS),.VDD(VDD),.Y(I2004),.A(g500),.B(I2003));
  NAND2 NAND2_28(.VSS(VSS),.VDD(VDD),.Y(I2005),.A(g212),.B(I2003));
  NAND2 NAND2_29(.VSS(VSS),.VDD(VDD),.Y(g944),.A(I2004),.B(I2005));
  NAND2 NAND2_30(.VSS(VSS),.VDD(VDD),.Y(I2013),.A(g532),.B(g260));
  NAND2 NAND2_31(.VSS(VSS),.VDD(VDD),.Y(I2014),.A(g532),.B(I2013));
  NAND2 NAND2_32(.VSS(VSS),.VDD(VDD),.Y(I2015),.A(g260),.B(I2013));
  NAND2 NAND2_33(.VSS(VSS),.VDD(VDD),.Y(g948),.A(I2014),.B(I2015));
  NAND2 NAND2_34(.VSS(VSS),.VDD(VDD),.Y(I2021),.A(g528),.B(g254));
  NAND2 NAND2_35(.VSS(VSS),.VDD(VDD),.Y(I2022),.A(g528),.B(I2021));
  NAND2 NAND2_36(.VSS(VSS),.VDD(VDD),.Y(I2023),.A(g254),.B(I2021));
  NAND2 NAND2_37(.VSS(VSS),.VDD(VDD),.Y(g950),.A(I2022),.B(I2023));
  NAND2 NAND2_38(.VSS(VSS),.VDD(VDD),.Y(I2060),.A(g7),.B(g3));
  NAND2 NAND2_39(.VSS(VSS),.VDD(VDD),.Y(I2061),.A(g7),.B(I2060));
  NAND2 NAND2_40(.VSS(VSS),.VDD(VDD),.Y(I2062),.A(g3),.B(I2060));
  NAND2 NAND2_41(.VSS(VSS),.VDD(VDD),.Y(g1036),.A(I2061),.B(I2062));
  NAND2 NAND2_42(.VSS(VSS),.VDD(VDD),.Y(I2072),.A(g15),.B(g11));
  NAND2 NAND2_43(.VSS(VSS),.VDD(VDD),.Y(I2073),.A(g15),.B(I2072));
  NAND2 NAND2_44(.VSS(VSS),.VDD(VDD),.Y(I2074),.A(g11),.B(I2072));
  NAND2 NAND2_45(.VSS(VSS),.VDD(VDD),.Y(g1042),.A(I2073),.B(I2074));
  NAND2 NAND2_46(.VSS(VSS),.VDD(VDD),.Y(I2080),.A(g25),.B(g19));
  NAND2 NAND2_47(.VSS(VSS),.VDD(VDD),.Y(I2081),.A(g25),.B(I2080));
  NAND2 NAND2_48(.VSS(VSS),.VDD(VDD),.Y(I2082),.A(g19),.B(I2080));
  NAND2 NAND2_49(.VSS(VSS),.VDD(VDD),.Y(g1044),.A(I2081),.B(I2082));
  NAND2 NAND2_50(.VSS(VSS),.VDD(VDD),.Y(I2089),.A(g33),.B(g29));
  NAND2 NAND2_51(.VSS(VSS),.VDD(VDD),.Y(I2090),.A(g33),.B(I2089));
  NAND2 NAND2_52(.VSS(VSS),.VDD(VDD),.Y(I2091),.A(g29),.B(I2089));
  NAND2 NAND2_53(.VSS(VSS),.VDD(VDD),.Y(g1047),.A(I2090),.B(I2091));
  NAND2 NAND2_54(.VSS(VSS),.VDD(VDD),.Y(I2108),.A(g602),.B(g610));
  NAND2 NAND2_55(.VSS(VSS),.VDD(VDD),.Y(I2109),.A(g602),.B(I2108));
  NAND2 NAND2_56(.VSS(VSS),.VDD(VDD),.Y(I2110),.A(g610),.B(I2108));
  NAND2 NAND2_57(.VSS(VSS),.VDD(VDD),.Y(g1075),.A(I2109),.B(I2110));
  NAND2 NAND2_58(.VSS(VSS),.VDD(VDD),.Y(g1138),.A(g102),.B(g98));
  NAND2 NAND2_59(.VSS(VSS),.VDD(VDD),.Y(g1157),.A(g89),.B(g107));
  NAND2 NAND2_60(.VSS(VSS),.VDD(VDD),.Y(I2244),.A(g567),.B(g598));
  NAND2 NAND2_61(.VSS(VSS),.VDD(VDD),.Y(I2245),.A(g567),.B(I2244));
  NAND2 NAND2_62(.VSS(VSS),.VDD(VDD),.Y(I2246),.A(g598),.B(I2244));
  NAND2 NAND2_63(.VSS(VSS),.VDD(VDD),.Y(g1253),.A(I2245),.B(I2246));
  NAND2 NAND2_64(.VSS(VSS),.VDD(VDD),.Y(I2299),.A(g830),.B(g341));
  NAND2 NAND2_65(.VSS(VSS),.VDD(VDD),.Y(I2300),.A(g830),.B(I2299));
  NAND2 NAND2_66(.VSS(VSS),.VDD(VDD),.Y(I2301),.A(g341),.B(I2299));
  NAND2 NAND2_67(.VSS(VSS),.VDD(VDD),.Y(g1316),.A(I2300),.B(I2301));
  NAND2 NAND2_68(.VSS(VSS),.VDD(VDD),.Y(g1359),.A(g866),.B(g306));
  NAND3 NAND3_0(.VSS(VSS),.VDD(VDD),.Y(g1387),.A(g862),.B(g314),.C(g301));
  NAND2 NAND2_69(.VSS(VSS),.VDD(VDD),.Y(g1398),.A(g306),.B(g889));
  NAND3 NAND3_1(.VSS(VSS),.VDD(VDD),.Y(g1402),.A(g310),.B(g866),.C(g873));
  NAND2 NAND2_70(.VSS(VSS),.VDD(VDD),.Y(g1411),.A(g314),.B(g873));
  NAND2 NAND2_71(.VSS(VSS),.VDD(VDD),.Y(g1417),.A(g873),.B(g889));
  NAND2 NAND2_72(.VSS(VSS),.VDD(VDD),.Y(I2497),.A(g1042),.B(g1036));
  NAND2 NAND2_73(.VSS(VSS),.VDD(VDD),.Y(I2498),.A(g1042),.B(I2497));
  NAND2 NAND2_74(.VSS(VSS),.VDD(VDD),.Y(I2499),.A(g1036),.B(I2497));
  NAND2 NAND2_75(.VSS(VSS),.VDD(VDD),.Y(g1534),.A(I2498),.B(I2499));
  NAND2 NAND2_76(.VSS(VSS),.VDD(VDD),.Y(I2506),.A(g1047),.B(g1044));
  NAND2 NAND2_77(.VSS(VSS),.VDD(VDD),.Y(I2507),.A(g1047),.B(I2506));
  NAND2 NAND2_78(.VSS(VSS),.VDD(VDD),.Y(I2508),.A(g1044),.B(I2506));
  NAND2 NAND2_79(.VSS(VSS),.VDD(VDD),.Y(g1540),.A(I2507),.B(I2508));
  NAND2 NAND2_80(.VSS(VSS),.VDD(VDD),.Y(I2526),.A(g766),.B(g719));
  NAND2 NAND2_81(.VSS(VSS),.VDD(VDD),.Y(I2527),.A(g766),.B(I2526));
  NAND2 NAND2_82(.VSS(VSS),.VDD(VDD),.Y(I2528),.A(g719),.B(I2526));
  NAND2 NAND2_83(.VSS(VSS),.VDD(VDD),.Y(g1558),.A(I2527),.B(I2528));
  NAND3 NAND3_2(.VSS(VSS),.VDD(VDD),.Y(g1573),.A(g729),.B(g719),.C(g766));
  NAND2 NAND2_84(.VSS(VSS),.VDD(VDD),.Y(I2542),.A(g821),.B(g774));
  NAND2 NAND2_85(.VSS(VSS),.VDD(VDD),.Y(I2543),.A(g821),.B(I2542));
  NAND2 NAND2_86(.VSS(VSS),.VDD(VDD),.Y(I2544),.A(g774),.B(I2542));
  NAND2 NAND2_87(.VSS(VSS),.VDD(VDD),.Y(g1574),.A(I2543),.B(I2544));
  NAND3 NAND3_3(.VSS(VSS),.VDD(VDD),.Y(g1582),.A(g784),.B(g774),.C(g821));
  NAND2 NAND2_88(.VSS(VSS),.VDD(VDD),.Y(I2674),.A(g710),.B(g131));
  NAND2 NAND2_89(.VSS(VSS),.VDD(VDD),.Y(I2675),.A(g710),.B(I2674));
  NAND2 NAND2_90(.VSS(VSS),.VDD(VDD),.Y(I2676),.A(g131),.B(I2674));
  NAND2 NAND2_91(.VSS(VSS),.VDD(VDD),.Y(g1686),.A(I2675),.B(I2676));
  NAND2 NAND2_92(.VSS(VSS),.VDD(VDD),.Y(I2681),.A(g918),.B(g613));
  NAND2 NAND2_93(.VSS(VSS),.VDD(VDD),.Y(I2682),.A(g918),.B(I2681));
  NAND2 NAND2_94(.VSS(VSS),.VDD(VDD),.Y(I2683),.A(g613),.B(I2681));
  NAND2 NAND2_95(.VSS(VSS),.VDD(VDD),.Y(g1687),.A(I2682),.B(I2683));
  NAND2 NAND2_96(.VSS(VSS),.VDD(VDD),.Y(g1743),.A(g1064),.B(g94));
  NAND2 NAND2_97(.VSS(VSS),.VDD(VDD),.Y(I2766),.A(g749),.B(g743));
  NAND2 NAND2_98(.VSS(VSS),.VDD(VDD),.Y(I2767),.A(g749),.B(I2766));
  NAND2 NAND2_99(.VSS(VSS),.VDD(VDD),.Y(I2768),.A(g743),.B(I2766));
  NAND2 NAND2_100(.VSS(VSS),.VDD(VDD),.Y(g1749),.A(I2767),.B(I2768));
  NAND2 NAND2_101(.VSS(VSS),.VDD(VDD),.Y(I2795),.A(g804),.B(g798));
  NAND2 NAND2_102(.VSS(VSS),.VDD(VDD),.Y(I2796),.A(g804),.B(I2795));
  NAND2 NAND2_103(.VSS(VSS),.VDD(VDD),.Y(I2797),.A(g798),.B(I2795));
  NAND2 NAND2_104(.VSS(VSS),.VDD(VDD),.Y(g1764),.A(I2796),.B(I2797));
  NAND3 NAND3_4(.VSS(VSS),.VDD(VDD),.Y(g1777),.A(g1060),.B(g102),.C(g89));
  NAND2 NAND2_105(.VSS(VSS),.VDD(VDD),.Y(g1793),.A(g94),.B(g1084));
  NAND3 NAND3_5(.VSS(VSS),.VDD(VDD),.Y(g1797),.A(g98),.B(g1064),.C(g1070));
  NAND2 NAND2_106(.VSS(VSS),.VDD(VDD),.Y(g1815),.A(g102),.B(g1070));
  NAND2 NAND2_107(.VSS(VSS),.VDD(VDD),.Y(g1822),.A(g1070),.B(g1084));
  NAND2 NAND2_108(.VSS(VSS),.VDD(VDD),.Y(I2897),.A(g1027),.B(g634));
  NAND2 NAND2_109(.VSS(VSS),.VDD(VDD),.Y(I2898),.A(g1027),.B(I2897));
  NAND2 NAND2_110(.VSS(VSS),.VDD(VDD),.Y(I2899),.A(g634),.B(I2897));
  NAND2 NAND2_111(.VSS(VSS),.VDD(VDD),.Y(g1829),.A(I2898),.B(I2899));
  NAND2 NAND2_112(.VSS(VSS),.VDD(VDD),.Y(I2933),.A(g1436),.B(g345));
  NAND2 NAND2_113(.VSS(VSS),.VDD(VDD),.Y(I2934),.A(g1436),.B(I2933));
  NAND2 NAND2_114(.VSS(VSS),.VDD(VDD),.Y(I2935),.A(g345),.B(I2933));
  NAND2 NAND2_115(.VSS(VSS),.VDD(VDD),.Y(g1845),.A(I2934),.B(I2935));
  NAND3 NAND3_6(.VSS(VSS),.VDD(VDD),.Y(g2008),.A(g866),.B(g873),.C(g1784));
  NAND3 NAND3_7(.VSS(VSS),.VDD(VDD),.Y(g2009),.A(g901),.B(g1387),.C(g905));
  NAND3 NAND3_8(.VSS(VSS),.VDD(VDD),.Y(g2010),.A(g1473),.B(g1470),.C(g1459));
  NAND2 NAND2_116(.VSS(VSS),.VDD(VDD),.Y(I3125),.A(g1279),.B(g1276));
  NAND2 NAND2_117(.VSS(VSS),.VDD(VDD),.Y(I3126),.A(g1279),.B(I3125));
  NAND2 NAND2_118(.VSS(VSS),.VDD(VDD),.Y(I3127),.A(g1276),.B(I3125));
  NAND2 NAND2_119(.VSS(VSS),.VDD(VDD),.Y(g2024),.A(I3126),.B(I3127));
  NAND2 NAND2_120(.VSS(VSS),.VDD(VDD),.Y(I3168),.A(g1540),.B(g1534));
  NAND2 NAND2_121(.VSS(VSS),.VDD(VDD),.Y(I3169),.A(g1540),.B(I3168));
  NAND2 NAND2_122(.VSS(VSS),.VDD(VDD),.Y(I3170),.A(g1534),.B(I3168));
  NAND2 NAND2_123(.VSS(VSS),.VDD(VDD),.Y(g2061),.A(I3169),.B(I3170));
  NAND2 NAND2_124(.VSS(VSS),.VDD(VDD),.Y(I3177),.A(g1706),.B(g736));
  NAND2 NAND2_125(.VSS(VSS),.VDD(VDD),.Y(I3178),.A(g1706),.B(I3177));
  NAND2 NAND2_126(.VSS(VSS),.VDD(VDD),.Y(I3179),.A(g736),.B(I3177));
  NAND2 NAND2_127(.VSS(VSS),.VDD(VDD),.Y(g2067),.A(I3178),.B(I3179));
  NAND2 NAND2_128(.VSS(VSS),.VDD(VDD),.Y(I3188),.A(g1716),.B(g791));
  NAND2 NAND2_129(.VSS(VSS),.VDD(VDD),.Y(I3189),.A(g1716),.B(I3188));
  NAND2 NAND2_130(.VSS(VSS),.VDD(VDD),.Y(I3190),.A(g791),.B(I3188));
  NAND2 NAND2_131(.VSS(VSS),.VDD(VDD),.Y(g2080),.A(I3189),.B(I3190));
  NAND3 NAND3_9(.VSS(VSS),.VDD(VDD),.Y(g2095),.A(g1584),.B(g749),.C(g736));
  NAND3 NAND3_10(.VSS(VSS),.VDD(VDD),.Y(g2100),.A(g1588),.B(g804),.C(g791));
  NAND2 NAND2_132(.VSS(VSS),.VDD(VDD),.Y(I3398),.A(g1826),.B(g135));
  NAND2 NAND2_133(.VSS(VSS),.VDD(VDD),.Y(I3399),.A(g1826),.B(I3398));
  NAND2 NAND2_134(.VSS(VSS),.VDD(VDD),.Y(I3400),.A(g135),.B(I3398));
  NAND2 NAND2_135(.VSS(VSS),.VDD(VDD),.Y(g2263),.A(I3399),.B(I3400));
  NAND2 NAND2_136(.VSS(VSS),.VDD(VDD),.Y(I3411),.A(g1419),.B(g616));
  NAND2 NAND2_137(.VSS(VSS),.VDD(VDD),.Y(I3412),.A(g1419),.B(I3411));
  NAND2 NAND2_138(.VSS(VSS),.VDD(VDD),.Y(I3413),.A(g616),.B(I3411));
  NAND2 NAND2_139(.VSS(VSS),.VDD(VDD),.Y(g2266),.A(I3412),.B(I3413));
  NAND2 NAND2_140(.VSS(VSS),.VDD(VDD),.Y(I3445),.A(g1689),.B(g729));
  NAND2 NAND2_141(.VSS(VSS),.VDD(VDD),.Y(I3446),.A(g1689),.B(I3445));
  NAND2 NAND2_142(.VSS(VSS),.VDD(VDD),.Y(I3447),.A(g729),.B(I3445));
  NAND2 NAND2_143(.VSS(VSS),.VDD(VDD),.Y(g2307),.A(I3446),.B(I3447));
  NAND2 NAND2_144(.VSS(VSS),.VDD(VDD),.Y(I3455),.A(g1691),.B(g784));
  NAND2 NAND2_145(.VSS(VSS),.VDD(VDD),.Y(I3456),.A(g1691),.B(I3455));
  NAND2 NAND2_146(.VSS(VSS),.VDD(VDD),.Y(I3457),.A(g784),.B(I3455));
  NAND2 NAND2_147(.VSS(VSS),.VDD(VDD),.Y(g2311),.A(I3456),.B(I3457));
  NAND3 NAND3_11(.VSS(VSS),.VDD(VDD),.Y(g2434),.A(g1064),.B(g1070),.C(g1620));
  NAND3 NAND3_12(.VSS(VSS),.VDD(VDD),.Y(g2435),.A(g1138),.B(g1777),.C(g1157));
  NAND2 NAND2_148(.VSS(VSS),.VDD(VDD),.Y(I3697),.A(g1570),.B(g642));
  NAND2 NAND2_149(.VSS(VSS),.VDD(VDD),.Y(I3698),.A(g1570),.B(I3697));
  NAND2 NAND2_150(.VSS(VSS),.VDD(VDD),.Y(I3699),.A(g642),.B(I3697));
  NAND2 NAND2_151(.VSS(VSS),.VDD(VDD),.Y(g2582),.A(I3698),.B(I3699));
  NAND2 NAND2_152(.VSS(VSS),.VDD(VDD),.Y(I3739),.A(g2021),.B(g349));
  NAND2 NAND2_153(.VSS(VSS),.VDD(VDD),.Y(I3740),.A(g2021),.B(I3739));
  NAND2 NAND2_154(.VSS(VSS),.VDD(VDD),.Y(I3741),.A(g349),.B(I3739));
  NAND2 NAND2_155(.VSS(VSS),.VDD(VDD),.Y(g2607),.A(I3740),.B(I3741));
  NAND2 NAND2_156(.VSS(VSS),.VDD(VDD),.Y(I3846),.A(g284),.B(g2370));
  NAND2 NAND2_157(.VSS(VSS),.VDD(VDD),.Y(I3847),.A(g284),.B(I3846));
  NAND2 NAND2_158(.VSS(VSS),.VDD(VDD),.Y(I3848),.A(g2370),.B(I3846));
  NAND2 NAND2_159(.VSS(VSS),.VDD(VDD),.Y(g2698),.A(I3847),.B(I3848));
  NAND2 NAND2_160(.VSS(VSS),.VDD(VDD),.Y(I3874),.A(g285),.B(g2397));
  NAND2 NAND2_161(.VSS(VSS),.VDD(VDD),.Y(I3875),.A(g285),.B(I3874));
  NAND2 NAND2_162(.VSS(VSS),.VDD(VDD),.Y(I3876),.A(g2397),.B(I3874));
  NAND2 NAND2_163(.VSS(VSS),.VDD(VDD),.Y(g2719),.A(I3875),.B(I3876));
  NAND2 NAND2_164(.VSS(VSS),.VDD(VDD),.Y(I3893),.A(g286),.B(g2422));
  NAND2 NAND2_165(.VSS(VSS),.VDD(VDD),.Y(I3894),.A(g286),.B(I3893));
  NAND2 NAND2_166(.VSS(VSS),.VDD(VDD),.Y(I3895),.A(g2422),.B(I3893));
  NAND2 NAND2_167(.VSS(VSS),.VDD(VDD),.Y(g2731),.A(I3894),.B(I3895));
  NAND2 NAND2_168(.VSS(VSS),.VDD(VDD),.Y(I3914),.A(g287),.B(g2449));
  NAND2 NAND2_169(.VSS(VSS),.VDD(VDD),.Y(I3915),.A(g287),.B(I3914));
  NAND2 NAND2_170(.VSS(VSS),.VDD(VDD),.Y(I3916),.A(g2449),.B(I3914));
  NAND2 NAND2_171(.VSS(VSS),.VDD(VDD),.Y(g2745),.A(I3915),.B(I3916));
  NAND2 NAND2_172(.VSS(VSS),.VDD(VDD),.Y(I3933),.A(g288),.B(g2473));
  NAND2 NAND2_173(.VSS(VSS),.VDD(VDD),.Y(I3934),.A(g288),.B(I3933));
  NAND2 NAND2_174(.VSS(VSS),.VDD(VDD),.Y(I3935),.A(g2473),.B(I3933));
  NAND2 NAND2_175(.VSS(VSS),.VDD(VDD),.Y(g2757),.A(I3934),.B(I3935));
  NAND2 NAND2_176(.VSS(VSS),.VDD(VDD),.Y(I3952),.A(g289),.B(g2497));
  NAND2 NAND2_177(.VSS(VSS),.VDD(VDD),.Y(I3953),.A(g289),.B(I3952));
  NAND2 NAND2_178(.VSS(VSS),.VDD(VDD),.Y(I3954),.A(g2497),.B(I3952));
  NAND2 NAND2_179(.VSS(VSS),.VDD(VDD),.Y(g2769),.A(I3953),.B(I3954));
  NAND2 NAND2_180(.VSS(VSS),.VDD(VDD),.Y(I3970),.A(g290),.B(g2518));
  NAND2 NAND2_181(.VSS(VSS),.VDD(VDD),.Y(I3971),.A(g290),.B(I3970));
  NAND2 NAND2_182(.VSS(VSS),.VDD(VDD),.Y(I3972),.A(g2518),.B(I3970));
  NAND2 NAND2_183(.VSS(VSS),.VDD(VDD),.Y(g2780),.A(I3971),.B(I3972));
  NAND2 NAND2_184(.VSS(VSS),.VDD(VDD),.Y(I3988),.A(g291),.B(g2544));
  NAND2 NAND2_185(.VSS(VSS),.VDD(VDD),.Y(I3989),.A(g291),.B(I3988));
  NAND2 NAND2_186(.VSS(VSS),.VDD(VDD),.Y(I3990),.A(g2544),.B(I3988));
  NAND2 NAND2_187(.VSS(VSS),.VDD(VDD),.Y(g2791),.A(I3989),.B(I3990));
  NAND2 NAND2_188(.VSS(VSS),.VDD(VDD),.Y(g2795),.A(g1997),.B(g866));
  NAND2 NAND2_189(.VSS(VSS),.VDD(VDD),.Y(I4008),.A(g292),.B(g2568));
  NAND2 NAND2_190(.VSS(VSS),.VDD(VDD),.Y(I4009),.A(g292),.B(I4008));
  NAND2 NAND2_191(.VSS(VSS),.VDD(VDD),.Y(I4010),.A(g2568),.B(I4008));
  NAND2 NAND2_192(.VSS(VSS),.VDD(VDD),.Y(g2804),.A(I4009),.B(I4010));
  NAND3 NAND3_13(.VSS(VSS),.VDD(VDD),.Y(g2831),.A(g2007),.B(g862),.C(g1784));
  NAND2 NAND2_193(.VSS(VSS),.VDD(VDD),.Y(g2858),.A(g1815),.B(g2577));
  NAND2 NAND2_194(.VSS(VSS),.VDD(VDD),.Y(g2940),.A(g197),.B(g2381));
  NAND2 NAND2_195(.VSS(VSS),.VDD(VDD),.Y(g2944),.A(g269),.B(g2381));
  NAND2 NAND2_196(.VSS(VSS),.VDD(VDD),.Y(g2947),.A(g1411),.B(g2026));
  NAND2 NAND2_197(.VSS(VSS),.VDD(VDD),.Y(g2951),.A(g2142),.B(g1797));
  NAND2 NAND2_198(.VSS(VSS),.VDD(VDD),.Y(I4150),.A(g2551),.B(g139));
  NAND2 NAND2_199(.VSS(VSS),.VDD(VDD),.Y(I4151),.A(g2551),.B(I4150));
  NAND2 NAND2_200(.VSS(VSS),.VDD(VDD),.Y(I4152),.A(g139),.B(I4150));
  NAND2 NAND2_201(.VSS(VSS),.VDD(VDD),.Y(g2960),.A(I4151),.B(I4152));
  NAND2 NAND2_202(.VSS(VSS),.VDD(VDD),.Y(I4159),.A(g2015),.B(g619));
  NAND2 NAND2_203(.VSS(VSS),.VDD(VDD),.Y(I4160),.A(g2015),.B(I4159));
  NAND2 NAND2_204(.VSS(VSS),.VDD(VDD),.Y(I4161),.A(g619),.B(I4159));
  NAND2 NAND2_205(.VSS(VSS),.VDD(VDD),.Y(g2966),.A(I4160),.B(I4161));
  NAND2 NAND2_206(.VSS(VSS),.VDD(VDD),.Y(I4182),.A(g2292),.B(g749));
  NAND2 NAND2_207(.VSS(VSS),.VDD(VDD),.Y(I4183),.A(g2292),.B(I4182));
  NAND2 NAND2_208(.VSS(VSS),.VDD(VDD),.Y(I4184),.A(g749),.B(I4182));
  NAND2 NAND2_209(.VSS(VSS),.VDD(VDD),.Y(g2995),.A(I4183),.B(I4184));
  NAND2 NAND2_210(.VSS(VSS),.VDD(VDD),.Y(I4203),.A(g2255),.B(g743));
  NAND2 NAND2_211(.VSS(VSS),.VDD(VDD),.Y(I4204),.A(g2255),.B(I4203));
  NAND2 NAND2_212(.VSS(VSS),.VDD(VDD),.Y(I4205),.A(g743),.B(I4203));
  NAND2 NAND2_213(.VSS(VSS),.VDD(VDD),.Y(g3012),.A(I4204),.B(I4205));
  NAND2 NAND2_214(.VSS(VSS),.VDD(VDD),.Y(I4210),.A(g2294),.B(g804));
  NAND2 NAND2_215(.VSS(VSS),.VDD(VDD),.Y(I4211),.A(g2294),.B(I4210));
  NAND2 NAND2_216(.VSS(VSS),.VDD(VDD),.Y(I4212),.A(g804),.B(I4210));
  NAND2 NAND2_217(.VSS(VSS),.VDD(VDD),.Y(g3013),.A(I4211),.B(I4212));
  NAND2 NAND2_218(.VSS(VSS),.VDD(VDD),.Y(I4233),.A(g2267),.B(g798));
  NAND2 NAND2_219(.VSS(VSS),.VDD(VDD),.Y(I4234),.A(g2267),.B(I4233));
  NAND2 NAND2_220(.VSS(VSS),.VDD(VDD),.Y(I4235),.A(g798),.B(I4233));
  NAND2 NAND2_221(.VSS(VSS),.VDD(VDD),.Y(g3028),.A(I4234),.B(I4235));
  NAND2 NAND2_222(.VSS(VSS),.VDD(VDD),.Y(g3109),.A(g2360),.B(g1064));
  NAND3 NAND3_14(.VSS(VSS),.VDD(VDD),.Y(g3140),.A(g2409),.B(g1060),.C(g1620));
  NAND2 NAND2_223(.VSS(VSS),.VDD(VDD),.Y(I4444),.A(g2092),.B(g606));
  NAND2 NAND2_224(.VSS(VSS),.VDD(VDD),.Y(I4445),.A(g2092),.B(I4444));
  NAND2 NAND2_225(.VSS(VSS),.VDD(VDD),.Y(I4446),.A(g606),.B(I4444));
  NAND2 NAND2_226(.VSS(VSS),.VDD(VDD),.Y(g3207),.A(I4445),.B(I4446));
  NAND2 NAND2_227(.VSS(VSS),.VDD(VDD),.Y(g3215),.A(g2340),.B(g1402));
  NAND2 NAND2_228(.VSS(VSS),.VDD(VDD),.Y(I4526),.A(g2909),.B(g646));
  NAND2 NAND2_229(.VSS(VSS),.VDD(VDD),.Y(I4527),.A(g2909),.B(I4526));
  NAND2 NAND2_230(.VSS(VSS),.VDD(VDD),.Y(I4528),.A(g646),.B(I4526));
  NAND2 NAND2_231(.VSS(VSS),.VDD(VDD),.Y(g3246),.A(I4527),.B(I4528));
  NAND2 NAND2_232(.VSS(VSS),.VDD(VDD),.Y(I4545),.A(g2853),.B(g353));
  NAND2 NAND2_233(.VSS(VSS),.VDD(VDD),.Y(I4546),.A(g2853),.B(I4545));
  NAND2 NAND2_234(.VSS(VSS),.VDD(VDD),.Y(I4547),.A(g353),.B(I4545));
  NAND2 NAND2_235(.VSS(VSS),.VDD(VDD),.Y(g3276),.A(I4546),.B(I4547));
  NAND3 NAND3_15(.VSS(VSS),.VDD(VDD),.Y(g3330),.A(g1815),.B(g1797),.C(g3109));
  NAND3 NAND3_16(.VSS(VSS),.VDD(VDD),.Y(g3502),.A(g1411),.B(g1402),.C(g2795));
  NAND4 NAND4_0(.VSS(VSS),.VDD(VDD),.Y(g3511),.A(g3158),.B(g3002),.C(g2976),.D(g2968));
  NAND4 NAND4_1(.VSS(VSS),.VDD(VDD),.Y(g3517),.A(g3173),.B(g3002),.C(g2976),.D(g2179));
  NAND4 NAND4_2(.VSS(VSS),.VDD(VDD),.Y(g3518),.A(g3177),.B(g3023),.C(g3007),.D(g2981));
  NAND4 NAND4_3(.VSS(VSS),.VDD(VDD),.Y(g3520),.A(g3183),.B(g3002),.C(g2197),.D(g2968));
  NAND4 NAND4_4(.VSS(VSS),.VDD(VDD),.Y(g3521),.A(g3187),.B(g3023),.C(g3007),.D(g2179));
  NAND4 NAND4_5(.VSS(VSS),.VDD(VDD),.Y(g3525),.A(g3192),.B(g3002),.C(g2197),.D(g2179));
  NAND4 NAND4_6(.VSS(VSS),.VDD(VDD),.Y(g3526),.A(g3196),.B(g3023),.C(g2197),.D(g2981));
  NAND4 NAND4_7(.VSS(VSS),.VDD(VDD),.Y(g3529),.A(g3200),.B(g2215),.C(g2976),.D(g2968));
  NAND4 NAND4_8(.VSS(VSS),.VDD(VDD),.Y(g3530),.A(g3204),.B(g3023),.C(g2197),.D(g2179));
  NAND4 NAND4_9(.VSS(VSS),.VDD(VDD),.Y(g3531),.A(g3209),.B(g2215),.C(g2976),.D(g2179));
  NAND4 NAND4_10(.VSS(VSS),.VDD(VDD),.Y(g3532),.A(g3212),.B(g2215),.C(g3007),.D(g2981));
  NAND4 NAND4_11(.VSS(VSS),.VDD(VDD),.Y(g3535),.A(g3216),.B(g2215),.C(g2197),.D(g2968));
  NAND4 NAND4_12(.VSS(VSS),.VDD(VDD),.Y(g3536),.A(g3219),.B(g2215),.C(g3007),.D(g2179));
  NAND4 NAND4_13(.VSS(VSS),.VDD(VDD),.Y(g3538),.A(g2588),.B(g2215),.C(g2197),.D(g2179));
  NAND4 NAND4_14(.VSS(VSS),.VDD(VDD),.Y(g3539),.A(g2591),.B(g2215),.C(g2197),.D(g2981));
  NAND4 NAND4_15(.VSS(VSS),.VDD(VDD),.Y(g3544),.A(g2594),.B(g2215),.C(g2197),.D(g2179));
  NAND2 NAND2_236(.VSS(VSS),.VDD(VDD),.Y(I4782),.A(g2846),.B(g622));
  NAND2 NAND2_237(.VSS(VSS),.VDD(VDD),.Y(I4783),.A(g2846),.B(I4782));
  NAND2 NAND2_238(.VSS(VSS),.VDD(VDD),.Y(I4784),.A(g622),.B(I4782));
  NAND2 NAND2_239(.VSS(VSS),.VDD(VDD),.Y(g3597),.A(I4783),.B(I4784));
  NAND3 NAND3_17(.VSS(VSS),.VDD(VDD),.Y(g3741),.A(g901),.B(g3433),.C(g2340));
  NAND2 NAND2_240(.VSS(VSS),.VDD(VDD),.Y(I4919),.A(g3522),.B(g650));
  NAND2 NAND2_241(.VSS(VSS),.VDD(VDD),.Y(I4920),.A(g3522),.B(I4919));
  NAND2 NAND2_242(.VSS(VSS),.VDD(VDD),.Y(I4921),.A(g650),.B(I4919));
  NAND2 NAND2_243(.VSS(VSS),.VDD(VDD),.Y(g3742),.A(I4920),.B(I4921));
  NAND2 NAND2_244(.VSS(VSS),.VDD(VDD),.Y(I4939),.A(g3437),.B(g357));
  NAND2 NAND2_245(.VSS(VSS),.VDD(VDD),.Y(I4940),.A(g3437),.B(I4939));
  NAND2 NAND2_246(.VSS(VSS),.VDD(VDD),.Y(I4941),.A(g357),.B(I4939));
  NAND2 NAND2_247(.VSS(VSS),.VDD(VDD),.Y(g3756),.A(I4940),.B(I4941));
  NAND3 NAND3_18(.VSS(VSS),.VDD(VDD),.Y(g3893),.A(g3664),.B(g3656),.C(g3647));
  NAND2 NAND2_248(.VSS(VSS),.VDD(VDD),.Y(I5187),.A(g3589),.B(g3593));
  NAND2 NAND2_249(.VSS(VSS),.VDD(VDD),.Y(I5188),.A(g3589),.B(I5187));
  NAND2 NAND2_250(.VSS(VSS),.VDD(VDD),.Y(I5189),.A(g3593),.B(I5187));
  NAND2 NAND2_251(.VSS(VSS),.VDD(VDD),.Y(g3955),.A(I5188),.B(I5189));
  NAND2 NAND2_252(.VSS(VSS),.VDD(VDD),.Y(I5195),.A(g3567),.B(g3571));
  NAND2 NAND2_253(.VSS(VSS),.VDD(VDD),.Y(I5196),.A(g3567),.B(I5195));
  NAND2 NAND2_254(.VSS(VSS),.VDD(VDD),.Y(I5197),.A(g3571),.B(I5195));
  NAND2 NAND2_255(.VSS(VSS),.VDD(VDD),.Y(g3957),.A(I5196),.B(I5197));
  NAND2 NAND2_256(.VSS(VSS),.VDD(VDD),.Y(I5207),.A(g3267),.B(g3271));
  NAND2 NAND2_257(.VSS(VSS),.VDD(VDD),.Y(I5208),.A(g3267),.B(I5207));
  NAND2 NAND2_258(.VSS(VSS),.VDD(VDD),.Y(I5209),.A(g3271),.B(I5207));
  NAND2 NAND2_259(.VSS(VSS),.VDD(VDD),.Y(g3961),.A(I5208),.B(I5209));
  NAND2 NAND2_260(.VSS(VSS),.VDD(VDD),.Y(I5226),.A(g3259),.B(g3263));
  NAND2 NAND2_261(.VSS(VSS),.VDD(VDD),.Y(I5227),.A(g3259),.B(I5226));
  NAND2 NAND2_262(.VSS(VSS),.VDD(VDD),.Y(I5228),.A(g3263),.B(I5226));
  NAND2 NAND2_263(.VSS(VSS),.VDD(VDD),.Y(g3968),.A(I5227),.B(I5228));
  NAND2 NAND2_264(.VSS(VSS),.VDD(VDD),.Y(I5242),.A(g3242),.B(g3247));
  NAND2 NAND2_265(.VSS(VSS),.VDD(VDD),.Y(I5243),.A(g3242),.B(I5242));
  NAND2 NAND2_266(.VSS(VSS),.VDD(VDD),.Y(I5244),.A(g3247),.B(I5242));
  NAND2 NAND2_267(.VSS(VSS),.VDD(VDD),.Y(g3974),.A(I5243),.B(I5244));
  NAND2 NAND2_268(.VSS(VSS),.VDD(VDD),.Y(I5257),.A(g3714),.B(g3719));
  NAND2 NAND2_269(.VSS(VSS),.VDD(VDD),.Y(I5258),.A(g3714),.B(I5257));
  NAND2 NAND2_270(.VSS(VSS),.VDD(VDD),.Y(I5259),.A(g3719),.B(I5257));
  NAND2 NAND2_271(.VSS(VSS),.VDD(VDD),.Y(g3979),.A(I5258),.B(I5259));
  NAND2 NAND2_272(.VSS(VSS),.VDD(VDD),.Y(I5269),.A(g3705),.B(g3710));
  NAND2 NAND2_273(.VSS(VSS),.VDD(VDD),.Y(I5270),.A(g3705),.B(I5269));
  NAND2 NAND2_274(.VSS(VSS),.VDD(VDD),.Y(I5271),.A(g3710),.B(I5269));
  NAND2 NAND2_275(.VSS(VSS),.VDD(VDD),.Y(g3983),.A(I5270),.B(I5271));
  NAND3 NAND3_19(.VSS(VSS),.VDD(VDD),.Y(g3985),.A(g1138),.B(g3718),.C(g2142));
  NAND2 NAND2_276(.VSS(VSS),.VDD(VDD),.Y(I5292),.A(g3421),.B(g625));
  NAND2 NAND2_277(.VSS(VSS),.VDD(VDD),.Y(I5293),.A(g3421),.B(I5292));
  NAND2 NAND2_278(.VSS(VSS),.VDD(VDD),.Y(I5294),.A(g625),.B(I5292));
  NAND2 NAND2_279(.VSS(VSS),.VDD(VDD),.Y(g4002),.A(I5293),.B(I5294));
  NAND2 NAND2_280(.VSS(VSS),.VDD(VDD),.Y(I5300),.A(g471),.B(g3505));
  NAND2 NAND2_281(.VSS(VSS),.VDD(VDD),.Y(I5301),.A(g471),.B(I5300));
  NAND2 NAND2_282(.VSS(VSS),.VDD(VDD),.Y(I5302),.A(g3505),.B(I5300));
  NAND2 NAND2_283(.VSS(VSS),.VDD(VDD),.Y(g4004),.A(I5301),.B(I5302));
  NAND2 NAND2_284(.VSS(VSS),.VDD(VDD),.Y(I5307),.A(g478),.B(g3512));
  NAND2 NAND2_285(.VSS(VSS),.VDD(VDD),.Y(I5308),.A(g478),.B(I5307));
  NAND2 NAND2_286(.VSS(VSS),.VDD(VDD),.Y(I5309),.A(g3512),.B(I5307));
  NAND2 NAND2_287(.VSS(VSS),.VDD(VDD),.Y(g4007),.A(I5308),.B(I5309));
  NAND2 NAND2_288(.VSS(VSS),.VDD(VDD),.Y(g4017),.A(g107),.B(g3425));
  NAND2 NAND2_289(.VSS(VSS),.VDD(VDD),.Y(g4049),.A(g3677),.B(g3425));
  NAND2 NAND2_290(.VSS(VSS),.VDD(VDD),.Y(I5535),.A(g3907),.B(g654));
  NAND2 NAND2_291(.VSS(VSS),.VDD(VDD),.Y(I5536),.A(g3907),.B(I5535));
  NAND2 NAND2_292(.VSS(VSS),.VDD(VDD),.Y(I5537),.A(g654),.B(I5535));
  NAND2 NAND2_293(.VSS(VSS),.VDD(VDD),.Y(g4151),.A(I5536),.B(I5537));
  NAND2 NAND2_294(.VSS(VSS),.VDD(VDD),.Y(I5647),.A(g3974),.B(g3968));
  NAND2 NAND2_295(.VSS(VSS),.VDD(VDD),.Y(I5648),.A(g3974),.B(I5647));
  NAND2 NAND2_296(.VSS(VSS),.VDD(VDD),.Y(I5649),.A(g3968),.B(I5647));
  NAND2 NAND2_297(.VSS(VSS),.VDD(VDD),.Y(g4221),.A(I5648),.B(I5649));
  NAND2 NAND2_298(.VSS(VSS),.VDD(VDD),.Y(I5657),.A(g3983),.B(g3979));
  NAND2 NAND2_299(.VSS(VSS),.VDD(VDD),.Y(I5658),.A(g3983),.B(I5657));
  NAND2 NAND2_300(.VSS(VSS),.VDD(VDD),.Y(I5659),.A(g3979),.B(I5657));
  NAND2 NAND2_301(.VSS(VSS),.VDD(VDD),.Y(g4223),.A(I5658),.B(I5659));
  NAND2 NAND2_302(.VSS(VSS),.VDD(VDD),.Y(g4237),.A(g4049),.B(g4017));
  NAND2 NAND2_303(.VSS(VSS),.VDD(VDD),.Y(I5759),.A(g3836),.B(g3503));
  NAND2 NAND2_304(.VSS(VSS),.VDD(VDD),.Y(I5760),.A(g3836),.B(I5759));
  NAND2 NAND2_305(.VSS(VSS),.VDD(VDD),.Y(I5761),.A(g3503),.B(I5759));
  NAND2 NAND2_306(.VSS(VSS),.VDD(VDD),.Y(g4300),.A(I5760),.B(I5761));
  NAND2 NAND2_307(.VSS(VSS),.VDD(VDD),.Y(I5766),.A(g3961),.B(g3957));
  NAND2 NAND2_308(.VSS(VSS),.VDD(VDD),.Y(I5767),.A(g3961),.B(I5766));
  NAND2 NAND2_309(.VSS(VSS),.VDD(VDD),.Y(I5768),.A(g3957),.B(I5766));
  NAND2 NAND2_310(.VSS(VSS),.VDD(VDD),.Y(g4301),.A(I5767),.B(I5768));
  NAND2 NAND2_311(.VSS(VSS),.VDD(VDD),.Y(I5782),.A(g3810),.B(g628));
  NAND2 NAND2_312(.VSS(VSS),.VDD(VDD),.Y(I5783),.A(g3810),.B(I5782));
  NAND2 NAND2_313(.VSS(VSS),.VDD(VDD),.Y(I5784),.A(g628),.B(I5782));
  NAND2 NAND2_314(.VSS(VSS),.VDD(VDD),.Y(g4319),.A(I5783),.B(I5784));
  NAND2 NAND2_315(.VSS(VSS),.VDD(VDD),.Y(g4465),.A(g319),.B(g4253));
  NAND2 NAND2_316(.VSS(VSS),.VDD(VDD),.Y(g4472),.A(g3380),.B(g4253));
  NAND2 NAND2_317(.VSS(VSS),.VDD(VDD),.Y(I6026),.A(g4223),.B(g4221));
  NAND2 NAND2_318(.VSS(VSS),.VDD(VDD),.Y(I6027),.A(g4223),.B(I6026));
  NAND2 NAND2_319(.VSS(VSS),.VDD(VDD),.Y(I6028),.A(g4221),.B(I6026));
  NAND2 NAND2_320(.VSS(VSS),.VDD(VDD),.Y(g4504),.A(I6027),.B(I6028));
  NAND2 NAND2_321(.VSS(VSS),.VDD(VDD),.Y(I6175),.A(g4236),.B(g571));
  NAND2 NAND2_322(.VSS(VSS),.VDD(VDD),.Y(I6176),.A(g4236),.B(I6175));
  NAND2 NAND2_323(.VSS(VSS),.VDD(VDD),.Y(I6177),.A(g571),.B(I6175));
  NAND2 NAND2_324(.VSS(VSS),.VDD(VDD),.Y(g4608),.A(I6176),.B(I6177));
  NAND2 NAND2_325(.VSS(VSS),.VDD(VDD),.Y(I6185),.A(g4301),.B(g3955));
  NAND2 NAND2_326(.VSS(VSS),.VDD(VDD),.Y(I6186),.A(g4301),.B(I6185));
  NAND2 NAND2_327(.VSS(VSS),.VDD(VDD),.Y(I6187),.A(g3955),.B(I6185));
  NAND2 NAND2_328(.VSS(VSS),.VDD(VDD),.Y(g4610),.A(I6186),.B(I6187));
  NAND2 NAND2_329(.VSS(VSS),.VDD(VDD),.Y(I6194),.A(g4199),.B(g631));
  NAND2 NAND2_330(.VSS(VSS),.VDD(VDD),.Y(I6195),.A(g4199),.B(I6194));
  NAND2 NAND2_331(.VSS(VSS),.VDD(VDD),.Y(I6196),.A(g631),.B(I6194));
  NAND2 NAND2_332(.VSS(VSS),.VDD(VDD),.Y(g4613),.A(I6195),.B(I6196));
  NAND2 NAND2_333(.VSS(VSS),.VDD(VDD),.Y(g4640),.A(g4402),.B(g1056));
  NAND4 NAND4_16(.VSS(VSS),.VDD(VDD),.Y(g4669),.A(g4550),.B(g1017),.C(g1680),.D(g2897));
  NAND2 NAND2_334(.VSS(VSS),.VDD(VDD),.Y(g4670),.A(g4611),.B(g3528));
  NAND4 NAND4_17(.VSS(VSS),.VDD(VDD),.Y(g4674),.A(g4550),.B(g1514),.C(g2107),.D(g2897));
  NAND4 NAND4_18(.VSS(VSS),.VDD(VDD),.Y(g4678),.A(g2897),.B(g2101),.C(g1514),.D(g4550));
  NAND4 NAND4_19(.VSS(VSS),.VDD(VDD),.Y(g4680),.A(g4550),.B(g1514),.C(g1006),.D(g2897));
  NAND2 NAND2_335(.VSS(VSS),.VDD(VDD),.Y(I6390),.A(g4504),.B(g4610));
  NAND2 NAND2_336(.VSS(VSS),.VDD(VDD),.Y(I6391),.A(g4504),.B(I6390));
  NAND2 NAND2_337(.VSS(VSS),.VDD(VDD),.Y(I6392),.A(g4610),.B(I6390));
  NAND2 NAND2_338(.VSS(VSS),.VDD(VDD),.Y(g4762),.A(I6391),.B(I6392));
  NAND2 NAND2_339(.VSS(VSS),.VDD(VDD),.Y(I6473),.A(g4541),.B(g578));
  NAND2 NAND2_340(.VSS(VSS),.VDD(VDD),.Y(I6474),.A(g4541),.B(I6473));
  NAND2 NAND2_341(.VSS(VSS),.VDD(VDD),.Y(I6475),.A(g578),.B(I6473));
  NAND2 NAND2_342(.VSS(VSS),.VDD(VDD),.Y(g4803),.A(I6474),.B(I6475));
  NAND4 NAND4_20(.VSS(VSS),.VDD(VDD),.Y(g4812),.A(g4550),.B(g1560),.C(g1559),.D(g2073));
  NAND4 NAND4_21(.VSS(VSS),.VDD(VDD),.Y(g4813),.A(g4550),.B(g965),.C(g1560),.D(g2073));
  NAND4 NAND4_22(.VSS(VSS),.VDD(VDD),.Y(g4814),.A(g4550),.B(g1575),.C(g1550),.D(g2073));
  NAND4 NAND4_23(.VSS(VSS),.VDD(VDD),.Y(g4816),.A(g996),.B(g4550),.C(g1518),.D(g2073));
  NAND2 NAND2_343(.VSS(VSS),.VDD(VDD),.Y(I6499),.A(g4504),.B(g3541));
  NAND2 NAND2_344(.VSS(VSS),.VDD(VDD),.Y(I6500),.A(g4504),.B(I6499));
  NAND2 NAND2_345(.VSS(VSS),.VDD(VDD),.Y(I6501),.A(g3541),.B(I6499));
  NAND2 NAND2_346(.VSS(VSS),.VDD(VDD),.Y(g4819),.A(I6500),.B(I6501));
  NAND2 NAND2_347(.VSS(VSS),.VDD(VDD),.Y(g4825),.A(g4472),.B(g4465));
  NAND2 NAND2_348(.VSS(VSS),.VDD(VDD),.Y(g4903),.A(g4717),.B(g858));
  NAND2 NAND2_349(.VSS(VSS),.VDD(VDD),.Y(I6659),.A(g4762),.B(g3541));
  NAND2 NAND2_350(.VSS(VSS),.VDD(VDD),.Y(I6660),.A(g4762),.B(I6659));
  NAND2 NAND2_351(.VSS(VSS),.VDD(VDD),.Y(I6661),.A(g3541),.B(I6659));
  NAND2 NAND2_352(.VSS(VSS),.VDD(VDD),.Y(g5019),.A(I6660),.B(I6661));
  NAND2 NAND2_353(.VSS(VSS),.VDD(VDD),.Y(I6743),.A(g4708),.B(g582));
  NAND2 NAND2_354(.VSS(VSS),.VDD(VDD),.Y(I6744),.A(g4708),.B(I6743));
  NAND2 NAND2_355(.VSS(VSS),.VDD(VDD),.Y(I6745),.A(g582),.B(I6743));
  NAND2 NAND2_356(.VSS(VSS),.VDD(VDD),.Y(g5111),.A(I6744),.B(I6745));
  NAND2 NAND2_357(.VSS(VSS),.VDD(VDD),.Y(I6962),.A(g4874),.B(g586));
  NAND2 NAND2_358(.VSS(VSS),.VDD(VDD),.Y(I6963),.A(g4874),.B(I6962));
  NAND2 NAND2_359(.VSS(VSS),.VDD(VDD),.Y(I6964),.A(g586),.B(I6962));
  NAND2 NAND2_360(.VSS(VSS),.VDD(VDD),.Y(g5308),.A(I6963),.B(I6964));
  NAND2 NAND2_361(.VSS(VSS),.VDD(VDD),.Y(g5318),.A(g676),.B(g5060));
  NAND2 NAND2_362(.VSS(VSS),.VDD(VDD),.Y(I7097),.A(g5194),.B(g574));
  NAND2 NAND2_363(.VSS(VSS),.VDD(VDD),.Y(I7098),.A(g5194),.B(I7097));
  NAND2 NAND2_364(.VSS(VSS),.VDD(VDD),.Y(I7099),.A(g574),.B(I7097));
  NAND2 NAND2_365(.VSS(VSS),.VDD(VDD),.Y(g5431),.A(I7098),.B(I7099));
  NAND2 NAND2_366(.VSS(VSS),.VDD(VDD),.Y(g5455),.A(g2330),.B(g5311));
  NAND2 NAND2_367(.VSS(VSS),.VDD(VDD),.Y(I7208),.A(g143),.B(g5367));
  NAND2 NAND2_368(.VSS(VSS),.VDD(VDD),.Y(I7209),.A(g143),.B(I7208));
  NAND2 NAND2_369(.VSS(VSS),.VDD(VDD),.Y(I7210),.A(g5367),.B(I7208));
  NAND2 NAND2_370(.VSS(VSS),.VDD(VDD),.Y(g5502),.A(I7209),.B(I7210));
  NAND2 NAND2_371(.VSS(VSS),.VDD(VDD),.Y(I7216),.A(g152),.B(g5368));
  NAND2 NAND2_372(.VSS(VSS),.VDD(VDD),.Y(I7217),.A(g152),.B(I7216));
  NAND2 NAND2_373(.VSS(VSS),.VDD(VDD),.Y(I7218),.A(g5368),.B(I7216));
  NAND2 NAND2_374(.VSS(VSS),.VDD(VDD),.Y(g5504),.A(I7217),.B(I7218));
  NAND2 NAND2_375(.VSS(VSS),.VDD(VDD),.Y(I7223),.A(g161),.B(g5370));
  NAND2 NAND2_376(.VSS(VSS),.VDD(VDD),.Y(I7224),.A(g161),.B(I7223));
  NAND2 NAND2_377(.VSS(VSS),.VDD(VDD),.Y(I7225),.A(g5370),.B(I7223));
  NAND2 NAND2_378(.VSS(VSS),.VDD(VDD),.Y(g5505),.A(I7224),.B(I7225));
  NAND2 NAND2_379(.VSS(VSS),.VDD(VDD),.Y(I7230),.A(g170),.B(g5372));
  NAND2 NAND2_380(.VSS(VSS),.VDD(VDD),.Y(I7231),.A(g170),.B(I7230));
  NAND2 NAND2_381(.VSS(VSS),.VDD(VDD),.Y(I7232),.A(g5372),.B(I7230));
  NAND2 NAND2_382(.VSS(VSS),.VDD(VDD),.Y(g5506),.A(I7231),.B(I7232));
  NAND2 NAND2_383(.VSS(VSS),.VDD(VDD),.Y(I7237),.A(g179),.B(g5374));
  NAND2 NAND2_384(.VSS(VSS),.VDD(VDD),.Y(I7238),.A(g179),.B(I7237));
  NAND2 NAND2_385(.VSS(VSS),.VDD(VDD),.Y(I7239),.A(g5374),.B(I7237));
  NAND2 NAND2_386(.VSS(VSS),.VDD(VDD),.Y(g5507),.A(I7238),.B(I7239));
  NAND2 NAND2_387(.VSS(VSS),.VDD(VDD),.Y(I7244),.A(g188),.B(g5377));
  NAND2 NAND2_388(.VSS(VSS),.VDD(VDD),.Y(I7245),.A(g188),.B(I7244));
  NAND2 NAND2_389(.VSS(VSS),.VDD(VDD),.Y(I7246),.A(g5377),.B(I7244));
  NAND2 NAND2_390(.VSS(VSS),.VDD(VDD),.Y(g5508),.A(I7245),.B(I7246));
  NAND2 NAND2_391(.VSS(VSS),.VDD(VDD),.Y(I7311),.A(g5364),.B(g590));
  NAND2 NAND2_392(.VSS(VSS),.VDD(VDD),.Y(I7312),.A(g5364),.B(I7311));
  NAND2 NAND2_393(.VSS(VSS),.VDD(VDD),.Y(I7313),.A(g590),.B(I7311));
  NAND2 NAND2_394(.VSS(VSS),.VDD(VDD),.Y(g5565),.A(I7312),.B(I7313));
  NAND2 NAND2_395(.VSS(VSS),.VDD(VDD),.Y(g5634),.A(g5563),.B(g4767));
  NAND2 NAND2_396(.VSS(VSS),.VDD(VDD),.Y(g5636),.A(g5564),.B(g4769));
  NAND2 NAND2_397(.VSS(VSS),.VDD(VDD),.Y(I7432),.A(g111),.B(g5554));
  NAND2 NAND2_398(.VSS(VSS),.VDD(VDD),.Y(I7433),.A(g111),.B(I7432));
  NAND2 NAND2_399(.VSS(VSS),.VDD(VDD),.Y(I7434),.A(g5554),.B(I7432));
  NAND2 NAND2_400(.VSS(VSS),.VDD(VDD),.Y(g5683),.A(I7433),.B(I7434));
  NAND2 NAND2_401(.VSS(VSS),.VDD(VDD),.Y(I7439),.A(g5515),.B(g594));
  NAND2 NAND2_402(.VSS(VSS),.VDD(VDD),.Y(I7440),.A(g5515),.B(I7439));
  NAND2 NAND2_403(.VSS(VSS),.VDD(VDD),.Y(I7441),.A(g594),.B(I7439));
  NAND2 NAND2_404(.VSS(VSS),.VDD(VDD),.Y(g5684),.A(I7440),.B(I7441));
  NAND4 NAND4_24(.VSS(VSS),.VDD(VDD),.Y(g5686),.A(g5546),.B(g1017),.C(g1551),.D(g2916));
  NAND4 NAND4_25(.VSS(VSS),.VDD(VDD),.Y(g5688),.A(g5546),.B(g1585),.C(g2084),.D(g2916));
  NAND2 NAND2_405(.VSS(VSS),.VDD(VDD),.Y(I7520),.A(g361),.B(g5659));
  NAND2 NAND2_406(.VSS(VSS),.VDD(VDD),.Y(I7521),.A(g361),.B(I7520));
  NAND2 NAND2_407(.VSS(VSS),.VDD(VDD),.Y(I7522),.A(g5659),.B(I7520));
  NAND2 NAND2_408(.VSS(VSS),.VDD(VDD),.Y(g5775),.A(I7521),.B(I7522));
  NAND2 NAND2_409(.VSS(VSS),.VDD(VDD),.Y(I7527),.A(g49),.B(g5662));
  NAND2 NAND2_410(.VSS(VSS),.VDD(VDD),.Y(I7528),.A(g49),.B(I7527));
  NAND2 NAND2_411(.VSS(VSS),.VDD(VDD),.Y(I7529),.A(g5662),.B(I7527));
  NAND2 NAND2_412(.VSS(VSS),.VDD(VDD),.Y(g5776),.A(I7528),.B(I7529));
  NAND2 NAND2_413(.VSS(VSS),.VDD(VDD),.Y(I7534),.A(g54),.B(g5666));
  NAND2 NAND2_414(.VSS(VSS),.VDD(VDD),.Y(I7535),.A(g54),.B(I7534));
  NAND2 NAND2_415(.VSS(VSS),.VDD(VDD),.Y(I7536),.A(g5666),.B(I7534));
  NAND2 NAND2_416(.VSS(VSS),.VDD(VDD),.Y(g5777),.A(I7535),.B(I7536));
  NAND2 NAND2_417(.VSS(VSS),.VDD(VDD),.Y(I7541),.A(g59),.B(g5669));
  NAND2 NAND2_418(.VSS(VSS),.VDD(VDD),.Y(I7542),.A(g59),.B(I7541));
  NAND2 NAND2_419(.VSS(VSS),.VDD(VDD),.Y(I7543),.A(g5669),.B(I7541));
  NAND2 NAND2_420(.VSS(VSS),.VDD(VDD),.Y(g5778),.A(I7542),.B(I7543));
  NAND2 NAND2_421(.VSS(VSS),.VDD(VDD),.Y(I7548),.A(g64),.B(g5672));
  NAND2 NAND2_422(.VSS(VSS),.VDD(VDD),.Y(I7549),.A(g64),.B(I7548));
  NAND2 NAND2_423(.VSS(VSS),.VDD(VDD),.Y(I7550),.A(g5672),.B(I7548));
  NAND2 NAND2_424(.VSS(VSS),.VDD(VDD),.Y(g5779),.A(I7549),.B(I7550));
  NAND2 NAND2_425(.VSS(VSS),.VDD(VDD),.Y(I7555),.A(g69),.B(g5674));
  NAND2 NAND2_426(.VSS(VSS),.VDD(VDD),.Y(I7556),.A(g69),.B(I7555));
  NAND2 NAND2_427(.VSS(VSS),.VDD(VDD),.Y(I7557),.A(g5674),.B(I7555));
  NAND2 NAND2_428(.VSS(VSS),.VDD(VDD),.Y(g5780),.A(I7556),.B(I7557));
  NAND2 NAND2_429(.VSS(VSS),.VDD(VDD),.Y(I7562),.A(g74),.B(g5676));
  NAND2 NAND2_430(.VSS(VSS),.VDD(VDD),.Y(I7563),.A(g74),.B(I7562));
  NAND2 NAND2_431(.VSS(VSS),.VDD(VDD),.Y(I7564),.A(g5676),.B(I7562));
  NAND2 NAND2_432(.VSS(VSS),.VDD(VDD),.Y(g5781),.A(I7563),.B(I7564));
  NAND2 NAND2_433(.VSS(VSS),.VDD(VDD),.Y(I7569),.A(g79),.B(g5678));
  NAND2 NAND2_434(.VSS(VSS),.VDD(VDD),.Y(I7570),.A(g79),.B(I7569));
  NAND2 NAND2_435(.VSS(VSS),.VDD(VDD),.Y(I7571),.A(g5678),.B(I7569));
  NAND2 NAND2_436(.VSS(VSS),.VDD(VDD),.Y(g5782),.A(I7570),.B(I7571));
  NAND2 NAND2_437(.VSS(VSS),.VDD(VDD),.Y(I7576),.A(g84),.B(g5680));
  NAND2 NAND2_438(.VSS(VSS),.VDD(VDD),.Y(I7577),.A(g84),.B(I7576));
  NAND2 NAND2_439(.VSS(VSS),.VDD(VDD),.Y(I7578),.A(g5680),.B(I7576));
  NAND2 NAND2_440(.VSS(VSS),.VDD(VDD),.Y(g5783),.A(I7577),.B(I7578));
  NAND4 NAND4_26(.VSS(VSS),.VDD(VDD),.Y(g5818),.A(g5638),.B(g2056),.C(g1666),.D(g1661));
  NAND4 NAND4_27(.VSS(VSS),.VDD(VDD),.Y(g5821),.A(g5638),.B(g2056),.C(g1076),.D(g1666));
  NAND3 NAND3_20(.VSS(VSS),.VDD(VDD),.Y(g5852),.A(g5638),.B(g2053),.C(g1661));
  NAND3 NAND3_21(.VSS(VSS),.VDD(VDD),.Y(g5853),.A(g5638),.B(g2053),.C(g1076));
  NAND4 NAND4_28(.VSS(VSS),.VDD(VDD),.Y(g5854),.A(g5638),.B(g1683),.C(g1552),.D(g2062));
  NAND4 NAND4_29(.VSS(VSS),.VDD(VDD),.Y(g5857),.A(g5638),.B(g1552),.C(g1017),.D(g2062));
  NAND4 NAND4_30(.VSS(VSS),.VDD(VDD),.Y(g5862),.A(g5649),.B(g1529),.C(g1535),.D(g2068));
  NAND4 NAND4_31(.VSS(VSS),.VDD(VDD),.Y(g5863),.A(g5649),.B(g1076),.C(g1535),.D(g2068));
  NAND4 NAND4_32(.VSS(VSS),.VDD(VDD),.Y(g5864),.A(g5649),.B(g1529),.C(g1088),.D(g2068));
  NAND4 NAND4_33(.VSS(VSS),.VDD(VDD),.Y(g5865),.A(g5649),.B(g1088),.C(g1076),.D(g2068));
  NAND3 NAND3_22(.VSS(VSS),.VDD(VDD),.Y(g5866),.A(g5649),.B(g1529),.C(g2081));
  NAND3 NAND3_23(.VSS(VSS),.VDD(VDD),.Y(g5869),.A(g5649),.B(g1076),.C(g2081));
  NAND4 NAND4_34(.VSS(VSS),.VDD(VDD),.Y(g5872),.A(g5649),.B(g1557),.C(g1564),.D(g2113));
  NAND4 NAND4_35(.VSS(VSS),.VDD(VDD),.Y(g5873),.A(g5649),.B(g1017),.C(g1564),.D(g2113));
  NAND2 NAND2_441(.VSS(VSS),.VDD(VDD),.Y(g5926),.A(g5741),.B(g639));
  NAND2 NAND2_442(.VSS(VSS),.VDD(VDD),.Y(g5943),.A(g5818),.B(g2940));
  NAND2 NAND2_443(.VSS(VSS),.VDD(VDD),.Y(g5947),.A(g5821),.B(g2944));
  NAND2 NAND2_444(.VSS(VSS),.VDD(VDD),.Y(g6095),.A(g2952),.B(g5854));
  NAND2 NAND2_445(.VSS(VSS),.VDD(VDD),.Y(g6097),.A(g2954),.B(g5857));
  NAND2 NAND2_446(.VSS(VSS),.VDD(VDD),.Y(I8194),.A(g471),.B(g6188));
  NAND2 NAND2_447(.VSS(VSS),.VDD(VDD),.Y(I8195),.A(g471),.B(I8194));
  NAND2 NAND2_448(.VSS(VSS),.VDD(VDD),.Y(I8196),.A(g6188),.B(I8194));
  NAND2 NAND2_449(.VSS(VSS),.VDD(VDD),.Y(g6394),.A(I8195),.B(I8196));
  NAND2 NAND2_450(.VSS(VSS),.VDD(VDD),.Y(I8201),.A(g478),.B(g6192));
  NAND2 NAND2_451(.VSS(VSS),.VDD(VDD),.Y(I8202),.A(g478),.B(I8201));
  NAND2 NAND2_452(.VSS(VSS),.VDD(VDD),.Y(I8203),.A(g6192),.B(I8201));
  NAND2 NAND2_453(.VSS(VSS),.VDD(VDD),.Y(g6397),.A(I8202),.B(I8203));
  NAND3 NAND3_24(.VSS(VSS),.VDD(VDD),.Y(g6717),.A(g6669),.B(g5065),.C(g5062));
  NAND3 NAND3_25(.VSS(VSS),.VDD(VDD),.Y(g6740),.A(g6703),.B(g6457),.C(g4936));
  NAND3 NAND3_26(.VSS(VSS),.VDD(VDD),.Y(g6741),.A(g6705),.B(g6461),.C(g4941));
  NAND3 NAND3_27(.VSS(VSS),.VDD(VDD),.Y(g6742),.A(g6683),.B(g932),.C(g6716));
  NAND2 NAND2_454(.VSS(VSS),.VDD(VDD),.Y(g6774),.A(g6754),.B(g6750));
  NAND2 NAND2_455(.VSS(VSS),.VDD(VDD),.Y(g6778),.A(g6762),.B(g6758));
  NAND3 NAND3_28(.VSS(VSS),.VDD(VDD),.Y(g6783),.A(g6747),.B(g5068),.C(g5066));
  NAND2 NAND2_456(.VSS(VSS),.VDD(VDD),.Y(I9050),.A(g6832),.B(g3598));
  NAND2 NAND2_457(.VSS(VSS),.VDD(VDD),.Y(I9051),.A(g6832),.B(I9050));
  NAND2 NAND2_458(.VSS(VSS),.VDD(VDD),.Y(I9052),.A(g3598),.B(I9050));
  NAND2 NAND2_459(.VSS(VSS),.VDD(VDD),.Y(g6843),.A(I9051),.B(I9052));
  NAND2 NAND2_460(.VSS(VSS),.VDD(VDD),.Y(g6873),.A(g6848),.B(g3621));
  NAND2 NAND2_461(.VSS(VSS),.VDD(VDD),.Y(g6928),.A(g4532),.B(g6926));
  NAND2 NAND2_462(.VSS(VSS),.VDD(VDD),.Y(g6929),.A(g4536),.B(g6927));
//
  NOR2 NOR2_0(.VSS(VSS),.VDD(VDD),.Y(g1418),.A(g486),.B(g943));
  NOR2 NOR2_1(.VSS(VSS),.VDD(VDD),.Y(g1422),.A(g1039),.B(g913));
  NOR2 NOR2_2(.VSS(VSS),.VDD(VDD),.Y(g1449),.A(g489),.B(g1048));
  NOR3 NOR3_0(.VSS(VSS),.VDD(VDD),.Y(g1459),.A(g926),.B(g950),.C(g948));
  NOR3 NOR3_1(.VSS(VSS),.VDD(VDD),.Y(g1470),.A(g937),.B(g930),.C(g928));
  NOR3 NOR3_2(.VSS(VSS),.VDD(VDD),.Y(g1473),.A(g944),.B(g941),.C(g939));
  NOR2 NOR2_3(.VSS(VSS),.VDD(VDD),.Y(g1474),.A(g760),.B(g754));
  NOR2 NOR2_4(.VSS(VSS),.VDD(VDD),.Y(g1481),.A(g815),.B(g809));
  NOR2 NOR2_5(.VSS(VSS),.VDD(VDD),.Y(g1518),.A(g980),.B(g965));
  NOR2 NOR2_6(.VSS(VSS),.VDD(VDD),.Y(g1560),.A(g996),.B(g980));
  NOR2 NOR2_7(.VSS(VSS),.VDD(VDD),.Y(g1603),.A(g1039),.B(g658));
  NOR2 NOR2_8(.VSS(VSS),.VDD(VDD),.Y(g1879),.A(g1603),.B(g1416));
  NOR2 NOR2_9(.VSS(VSS),.VDD(VDD),.Y(g2433),.A(g1418),.B(g1449));
  NOR3 NOR3_3(.VSS(VSS),.VDD(VDD),.Y(g2908),.A(g536),.B(g2010),.C(g541));
  NOR2 NOR2_10(.VSS(VSS),.VDD(VDD),.Y(g3528),.A(g1802),.B(g3167));
  NOR2 NOR2_11(.VSS(VSS),.VDD(VDD),.Y(g3621),.A(g1407),.B(g2842));
  NOR3 NOR3_4(.VSS(VSS),.VDD(VDD),.Y(g3647),.A(g2731),.B(g2719),.C(g2698));
  NOR3 NOR3_5(.VSS(VSS),.VDD(VDD),.Y(g3656),.A(g2769),.B(g2757),.C(g2745));
  NOR3 NOR3_6(.VSS(VSS),.VDD(VDD),.Y(g3664),.A(g2804),.B(g2791),.C(g2780));
  NOR2 NOR2_12(.VSS(VSS),.VDD(VDD),.Y(g3903),.A(g3505),.B(g471));
  NOR2 NOR2_13(.VSS(VSS),.VDD(VDD),.Y(g3905),.A(g3512),.B(g478));
  NOR2 NOR2_14(.VSS(VSS),.VDD(VDD),.Y(g3923),.A(g3378),.B(g3381));
  NOR2 NOR2_15(.VSS(VSS),.VDD(VDD),.Y(g3925),.A(g3303),.B(g3315));
  NOR2 NOR2_16(.VSS(VSS),.VDD(VDD),.Y(g3926),.A(g3338),.B(g3350));
  NOR2 NOR2_17(.VSS(VSS),.VDD(VDD),.Y(g3927),.A(g3382),.B(g3383));
  NOR2 NOR2_18(.VSS(VSS),.VDD(VDD),.Y(g3929),.A(g3373),.B(g3376));
  NOR2 NOR2_19(.VSS(VSS),.VDD(VDD),.Y(g3930),.A(g3317),.B(g3328));
  NOR2 NOR2_20(.VSS(VSS),.VDD(VDD),.Y(g3931),.A(g3353),.B(g3361));
  NOR2 NOR2_21(.VSS(VSS),.VDD(VDD),.Y(g3933),.A(g3327),.B(g3336));
  NOR2 NOR2_22(.VSS(VSS),.VDD(VDD),.Y(g3934),.A(g3377),.B(g3379));
  NOR2 NOR2_23(.VSS(VSS),.VDD(VDD),.Y(g3939),.A(g3340),.B(g3351));
  NOR2 NOR2_24(.VSS(VSS),.VDD(VDD),.Y(g3956),.A(g3337),.B(g3349));
  NOR2 NOR2_25(.VSS(VSS),.VDD(VDD),.Y(g3958),.A(g3316),.B(g3326));
  NOR2 NOR2_26(.VSS(VSS),.VDD(VDD),.Y(g3959),.A(g3352),.B(g3360));
  NOR2 NOR2_27(.VSS(VSS),.VDD(VDD),.Y(g3965),.A(g3359),.B(g3367));
  NOR2 NOR2_28(.VSS(VSS),.VDD(VDD),.Y(g3966),.A(g3329),.B(g3339));
  NOR2 NOR2_29(.VSS(VSS),.VDD(VDD),.Y(g3973),.A(g3368),.B(g3374));
  NOR2 NOR2_30(.VSS(VSS),.VDD(VDD),.Y(g4000),.A(g1250),.B(g3425));
  NOR2 NOR2_31(.VSS(VSS),.VDD(VDD),.Y(g4235),.A(g3780),.B(g3362));
  NOR2 NOR2_32(.VSS(VSS),.VDD(VDD),.Y(g4238),.A(g3755),.B(g3279));
  NOR2 NOR2_33(.VSS(VSS),.VDD(VDD),.Y(g4239),.A(g3763),.B(g3296));
  NOR3 NOR3_7(.VSS(VSS),.VDD(VDD),.Y(g4240),.A(g1589),.B(g1879),.C(g3793));
  NOR2 NOR2_34(.VSS(VSS),.VDD(VDD),.Y(g4241),.A(g3774),.B(g3341));
  NOR2 NOR2_35(.VSS(VSS),.VDD(VDD),.Y(g4245),.A(g3759),.B(g3288));
  NOR2 NOR2_36(.VSS(VSS),.VDD(VDD),.Y(g4261),.A(g3762),.B(g3295));
  NOR2 NOR2_37(.VSS(VSS),.VDD(VDD),.Y(g4266),.A(g3757),.B(g3283));
  NOR2 NOR2_38(.VSS(VSS),.VDD(VDD),.Y(g4272),.A(g3767),.B(g3319));
  NOR2 NOR2_39(.VSS(VSS),.VDD(VDD),.Y(g4432),.A(g923),.B(g4253));
  NOR2 NOR2_40(.VSS(VSS),.VDD(VDD),.Y(g4568),.A(g4233),.B(g3924));
  NOR2 NOR2_41(.VSS(VSS),.VDD(VDD),.Y(g4578),.A(g4234),.B(g3928));
  NOR2 NOR2_42(.VSS(VSS),.VDD(VDD),.Y(g4581),.A(g4156),.B(g4160));
  NOR2 NOR2_43(.VSS(VSS),.VDD(VDD),.Y(g4584),.A(g4164),.B(g4168));
  NOR2 NOR2_44(.VSS(VSS),.VDD(VDD),.Y(g4585),.A(g4171),.B(g4177));
  NOR2 NOR2_45(.VSS(VSS),.VDD(VDD),.Y(g4586),.A(g4161),.B(g4165));
  NOR2 NOR2_46(.VSS(VSS),.VDD(VDD),.Y(g4589),.A(g4180),.B(g4183));
  NOR2 NOR2_47(.VSS(VSS),.VDD(VDD),.Y(g4590),.A(g4169),.B(g4172));
  NOR2 NOR2_48(.VSS(VSS),.VDD(VDD),.Y(g4591),.A(g4178),.B(g4181));
  NOR2 NOR2_49(.VSS(VSS),.VDD(VDD),.Y(g4596),.A(g4184),.B(g4186));
  NOR2 NOR2_50(.VSS(VSS),.VDD(VDD),.Y(g4774),.A(g4442),.B(g4445));
  NOR2 NOR2_51(.VSS(VSS),.VDD(VDD),.Y(g4776),.A(g4449),.B(g4453));
  NOR2 NOR2_52(.VSS(VSS),.VDD(VDD),.Y(g4777),.A(g4457),.B(g4459));
  NOR2 NOR2_53(.VSS(VSS),.VDD(VDD),.Y(g4779),.A(g4461),.B(g4464));
  NOR2 NOR2_54(.VSS(VSS),.VDD(VDD),.Y(g4877),.A(g952),.B(g4680));
  NOR2 NOR2_55(.VSS(VSS),.VDD(VDD),.Y(g4950),.A(g1472),.B(g4680));
  NOR2 NOR2_56(.VSS(VSS),.VDD(VDD),.Y(g4967),.A(g4674),.B(g952));
  NOR2 NOR2_57(.VSS(VSS),.VDD(VDD),.Y(g4993),.A(g4674),.B(g1477));
  NOR3 NOR3_8(.VSS(VSS),.VDD(VDD),.Y(g5048),.A(g4819),.B(g3491),.C(g3559));
  NOR2 NOR2_58(.VSS(VSS),.VDD(VDD),.Y(g5088),.A(g4691),.B(g4697));
  NOR2 NOR2_59(.VSS(VSS),.VDD(VDD),.Y(g5091),.A(g4698),.B(g4701));
  NOR2 NOR2_60(.VSS(VSS),.VDD(VDD),.Y(g5093),.A(g4683),.B(g4684));
  NOR2 NOR2_61(.VSS(VSS),.VDD(VDD),.Y(g5094),.A(g4685),.B(g4686));
  NOR2 NOR2_62(.VSS(VSS),.VDD(VDD),.Y(g5227),.A(g5019),.B(g3559));
  NOR2 NOR2_63(.VSS(VSS),.VDD(VDD),.Y(g5249),.A(g4868),.B(g4870));
  NOR2 NOR2_64(.VSS(VSS),.VDD(VDD),.Y(g5265),.A(g4863),.B(g4865));
  NOR3 NOR3_9(.VSS(VSS),.VDD(VDD),.Y(g5324),.A(g5069),.B(g4410),.C(g766));
  NOR3 NOR3_10(.VSS(VSS),.VDD(VDD),.Y(g5325),.A(g5077),.B(g4416),.C(g821));
  NOR2 NOR2_65(.VSS(VSS),.VDD(VDD),.Y(g5418),.A(g5162),.B(g5169));
  NOR2 NOR2_66(.VSS(VSS),.VDD(VDD),.Y(g5423),.A(g5170),.B(g5175));
  NOR2 NOR2_67(.VSS(VSS),.VDD(VDD),.Y(g5541),.A(g5388),.B(g1880));
  NOR2 NOR2_68(.VSS(VSS),.VDD(VDD),.Y(g5552),.A(g5354),.B(g5356));
  NOR4 NOR4_0(.VSS(VSS),.VDD(VDD),.Y(g5561),.A(g5391),.B(g1589),.C(g3793),.D(g1880));
  NOR2 NOR2_69(.VSS(VSS),.VDD(VDD),.Y(g5731),.A(g952),.B(g5688));
  NOR2 NOR2_70(.VSS(VSS),.VDD(VDD),.Y(g5753),.A(g1477),.B(g5688));
  NOR2 NOR2_71(.VSS(VSS),.VDD(VDD),.Y(g6073),.A(g197),.B(g5862));
  NOR2 NOR2_72(.VSS(VSS),.VDD(VDD),.Y(g6075),.A(g269),.B(g5863));
  NOR4 NOR4_1(.VSS(VSS),.VDD(VDD),.Y(g6279),.A(I7969),.B(I7970),.C(I7971),.D(I7972));
  NOR4 NOR4_2(.VSS(VSS),.VDD(VDD),.Y(g6280),.A(I7978),.B(I7979),.C(I7980),.D(I7981));
  NOR4 NOR4_3(.VSS(VSS),.VDD(VDD),.Y(g6281),.A(I7987),.B(I7988),.C(I7989),.D(I7990));
  NOR4 NOR4_4(.VSS(VSS),.VDD(VDD),.Y(g6335),.A(I8079),.B(I8080),.C(I8081),.D(I8082));
  NOR4 NOR4_5(.VSS(VSS),.VDD(VDD),.Y(g6357),.A(I8117),.B(I8118),.C(I8119),.D(I8120));
  NOR4 NOR4_6(.VSS(VSS),.VDD(VDD),.Y(g6358),.A(I8126),.B(I8127),.C(I8128),.D(I8129));
  NOR4 NOR4_7(.VSS(VSS),.VDD(VDD),.Y(g6359),.A(I8135),.B(I8136),.C(I8137),.D(I8138));
  NOR4 NOR4_8(.VSS(VSS),.VDD(VDD),.Y(g6400),.A(I8208),.B(I8209),.C(I8210),.D(I8211));
  NOR4 NOR4_9(.VSS(VSS),.VDD(VDD),.Y(g6427),.A(g6376),.B(g4086),.C(g4074),.D(g4068));
  NOR4 NOR4_10(.VSS(VSS),.VDD(VDD),.Y(g6429),.A(g6376),.B(g4086),.C(g4074),.D(g4302));
  NOR4 NOR4_11(.VSS(VSS),.VDD(VDD),.Y(g6430),.A(g6385),.B(g3733),.C(g4092),.D(g4080));
  NOR4 NOR4_12(.VSS(VSS),.VDD(VDD),.Y(g6432),.A(g6376),.B(g4086),.C(g4309),.D(g4068));
  NOR4 NOR4_13(.VSS(VSS),.VDD(VDD),.Y(g6433),.A(g6385),.B(g3733),.C(g4092),.D(g4314));
  NOR4 NOR4_14(.VSS(VSS),.VDD(VDD),.Y(g6435),.A(g6376),.B(g4086),.C(g4309),.D(g4302));
  NOR4 NOR4_15(.VSS(VSS),.VDD(VDD),.Y(g6436),.A(g6385),.B(g3733),.C(g4328),.D(g4080));
  NOR4 NOR4_16(.VSS(VSS),.VDD(VDD),.Y(g6438),.A(g6376),.B(g4323),.C(g4074),.D(g4068));
  NOR4 NOR4_17(.VSS(VSS),.VDD(VDD),.Y(g6439),.A(g6385),.B(g3733),.C(g4328),.D(g4314));
  NOR4 NOR4_18(.VSS(VSS),.VDD(VDD),.Y(g6442),.A(g6376),.B(g4323),.C(g4074),.D(g4302));
  NOR4 NOR4_19(.VSS(VSS),.VDD(VDD),.Y(g6443),.A(g6385),.B(g4334),.C(g4092),.D(g4080));
  NOR4 NOR4_20(.VSS(VSS),.VDD(VDD),.Y(g6445),.A(g6376),.B(g4323),.C(g4309),.D(g4068));
  NOR4 NOR4_21(.VSS(VSS),.VDD(VDD),.Y(g6446),.A(g6385),.B(g4334),.C(g4092),.D(g4314));
  NOR4 NOR4_22(.VSS(VSS),.VDD(VDD),.Y(g6448),.A(g6376),.B(g4323),.C(g4309),.D(g4302));
  NOR4 NOR4_23(.VSS(VSS),.VDD(VDD),.Y(g6449),.A(g6385),.B(g4334),.C(g4328),.D(g4080));
  NOR4 NOR4_24(.VSS(VSS),.VDD(VDD),.Y(g6451),.A(g6385),.B(g4334),.C(g4328),.D(g4314));
  NOR2 NOR2_73(.VSS(VSS),.VDD(VDD),.Y(g6492),.A(g6348),.B(g1734));
  NOR2 NOR2_74(.VSS(VSS),.VDD(VDD),.Y(g6494),.A(g952),.B(g6348));
  NOR2 NOR2_75(.VSS(VSS),.VDD(VDD),.Y(g6495),.A(g6354),.B(g1775));
  NOR2 NOR2_76(.VSS(VSS),.VDD(VDD),.Y(g6496),.A(g952),.B(g6354));

endmodule