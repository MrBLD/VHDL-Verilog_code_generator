module s298w(G117,G132,G133,G0,G118,CLOCK,G66,VDD,G1,VSS,G2,G67);
input G0,CLOCK,VDD,G1,VSS,G2;
output G117,G132,G133,G118,G66,G67;

  wire G131,G90,G102,G93,G114,G53,G75,G55,G98,G14,G47,G26,G127,G121,G25,I235,G130,G28,G54,G74,G80,G59,G32,G86,G79,G116,I221,G128,G29,G42,G52,G61,G91,G20,G110,G41,G122,G62,G23,G35,G111,G18,G78,G60,G70,G77,G10,G104,G21,G30,G50,G73,G85,G115,G101,G100,G119,G109,I238,G13,I210,I158,G83,G24,G40,G37,G125,G124,G68,G94,G106,G27,G48,G71,G58,G64,G112,G105,G36,I155,G92,G84,G97,G17,G15,G129,G69,G43,G31,G16,G12,G87,G33,G88,G49,G38,G56,G22,G39,G82,I232,G99,G19,G89,G46,G11,G126,G65,G45,G96,G113,G81,G72,I213,G34,G76,G51,G95,G103,G44,G107,G123,G63,G120,I229,G108,G57;
//# 3 inputs
//# 6 outputs
//# 14 D-type flipflops
//# 44 inverters
//# 75 gates (31 ANDs + 9 NANDs + 16 ORs + 19 NORs)
//
//
//
  MSFF DFF_0(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G10),.DATA(G29));
  MSFF DFF_1(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G11),.DATA(G30));
  MSFF DFF_2(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G12),.DATA(G34));
  MSFF DFF_3(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G13),.DATA(G39));
  MSFF DFF_4(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G14),.DATA(G44));
  MSFF DFF_5(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G15),.DATA(G56));
  MSFF DFF_6(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G16),.DATA(G86));
  MSFF DFF_7(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G17),.DATA(G92));
  MSFF DFF_8(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G18),.DATA(G98));
  MSFF DFF_9(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G19),.DATA(G102));
  MSFF DFF_10(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G20),.DATA(G107));
  MSFF DFF_11(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G21),.DATA(G113));
  MSFF DFF_12(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G22),.DATA(G119));
  MSFF DFF_13(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G23),.DATA(G125));
//
  NOT NOT1_0(.VSS(VSS),.VDD(VDD),.Y(G28),.A(G130));
  NOT NOT1_1(.VSS(VSS),.VDD(VDD),.Y(G38),.A(G10));
  NOT NOT1_2(.VSS(VSS),.VDD(VDD),.Y(G40),.A(G13));
  NOT NOT1_3(.VSS(VSS),.VDD(VDD),.Y(G45),.A(G12));
  NOT NOT1_4(.VSS(VSS),.VDD(VDD),.Y(G46),.A(G11));
  NOT NOT1_5(.VSS(VSS),.VDD(VDD),.Y(G50),.A(G14));
  NOT NOT1_6(.VSS(VSS),.VDD(VDD),.Y(G51),.A(G23));
  NOT NOT1_7(.VSS(VSS),.VDD(VDD),.Y(G54),.A(G11));
  NOT NOT1_8(.VSS(VSS),.VDD(VDD),.Y(G55),.A(G13));
  NOT NOT1_9(.VSS(VSS),.VDD(VDD),.Y(G59),.A(G12));
  NOT NOT1_10(.VSS(VSS),.VDD(VDD),.Y(G60),.A(G22));
  NOT NOT1_11(.VSS(VSS),.VDD(VDD),.Y(G64),.A(G15));
  NOT NOT1_12(.VSS(VSS),.VDD(VDD),.Y(I155),.A(G16));
  NOT NOT1_13(.VSS(VSS),.VDD(VDD),.Y(G66),.A(I155));
  NOT NOT1_14(.VSS(VSS),.VDD(VDD),.Y(I158),.A(G17));
  NOT NOT1_15(.VSS(VSS),.VDD(VDD),.Y(G67),.A(I158));
  NOT NOT1_16(.VSS(VSS),.VDD(VDD),.Y(G76),.A(G10));
  NOT NOT1_17(.VSS(VSS),.VDD(VDD),.Y(G82),.A(G11));
  NOT NOT1_18(.VSS(VSS),.VDD(VDD),.Y(G87),.A(G16));
  NOT NOT1_19(.VSS(VSS),.VDD(VDD),.Y(G91),.A(G12));
  NOT NOT1_20(.VSS(VSS),.VDD(VDD),.Y(G93),.A(G17));
  NOT NOT1_21(.VSS(VSS),.VDD(VDD),.Y(G96),.A(G14));
  NOT NOT1_22(.VSS(VSS),.VDD(VDD),.Y(G99),.A(G18));
  NOT NOT1_23(.VSS(VSS),.VDD(VDD),.Y(G103),.A(G13));
  NOT NOT1_24(.VSS(VSS),.VDD(VDD),.Y(G108),.A(G112));
  NOT NOT1_25(.VSS(VSS),.VDD(VDD),.Y(G114),.A(G21));
  NOT NOT1_26(.VSS(VSS),.VDD(VDD),.Y(I210),.A(G18));
  NOT NOT1_27(.VSS(VSS),.VDD(VDD),.Y(G117),.A(I210));
  NOT NOT1_28(.VSS(VSS),.VDD(VDD),.Y(I213),.A(G19));
  NOT NOT1_29(.VSS(VSS),.VDD(VDD),.Y(G118),.A(I213));
  NOT NOT1_30(.VSS(VSS),.VDD(VDD),.Y(G120),.A(G124));
  NOT NOT1_31(.VSS(VSS),.VDD(VDD),.Y(G121),.A(G22));
  NOT NOT1_32(.VSS(VSS),.VDD(VDD),.Y(I221),.A(G2));
  NOT NOT1_33(.VSS(VSS),.VDD(VDD),.Y(G124),.A(I221));
  NOT NOT1_34(.VSS(VSS),.VDD(VDD),.Y(G126),.A(G131));
  NOT NOT1_35(.VSS(VSS),.VDD(VDD),.Y(G127),.A(G23));
  NOT NOT1_36(.VSS(VSS),.VDD(VDD),.Y(I229),.A(G0));
  NOT NOT1_37(.VSS(VSS),.VDD(VDD),.Y(G130),.A(I229));
  NOT NOT1_38(.VSS(VSS),.VDD(VDD),.Y(I232),.A(G1));
  NOT NOT1_39(.VSS(VSS),.VDD(VDD),.Y(G131),.A(I232));
  NOT NOT1_40(.VSS(VSS),.VDD(VDD),.Y(I235),.A(G20));
  NOT NOT1_41(.VSS(VSS),.VDD(VDD),.Y(G132),.A(I235));
  NOT NOT1_42(.VSS(VSS),.VDD(VDD),.Y(I238),.A(G21));
  NOT NOT1_43(.VSS(VSS),.VDD(VDD),.Y(G133),.A(I238));
//
  AND2 AND2_0(.VSS(VSS),.VDD(VDD),.Y(G26),.A(G28),.B(G50));
  AND2 AND2_1(.VSS(VSS),.VDD(VDD),.Y(G27),.A(G51),.B(G28));
  AND3 AND3_0(.VSS(VSS),.VDD(VDD),.Y(G31),.A(G10),.B(G45),.C(G13));
  AND2 AND2_2(.VSS(VSS),.VDD(VDD),.Y(G32),.A(G10),.B(G11));
  AND2 AND2_3(.VSS(VSS),.VDD(VDD),.Y(G33),.A(G38),.B(G46));
  AND3 AND3_1(.VSS(VSS),.VDD(VDD),.Y(G35),.A(G10),.B(G11),.C(G12));
  AND2 AND2_4(.VSS(VSS),.VDD(VDD),.Y(G36),.A(G38),.B(G45));
  AND2 AND2_5(.VSS(VSS),.VDD(VDD),.Y(G37),.A(G46),.B(G45));
  AND2 AND2_6(.VSS(VSS),.VDD(VDD),.Y(G42),.A(G40),.B(G41));
  AND4 AND4_0(.VSS(VSS),.VDD(VDD),.Y(G48),.A(G45),.B(G46),.C(G10),.D(G47));
  AND3 AND3_2(.VSS(VSS),.VDD(VDD),.Y(G49),.A(G50),.B(G51),.C(G52));
  AND4 AND4_1(.VSS(VSS),.VDD(VDD),.Y(G57),.A(G59),.B(G11),.C(G60),.D(G61));
  AND2 AND2_7(.VSS(VSS),.VDD(VDD),.Y(G58),.A(G64),.B(G65));
  AND4 AND4_2(.VSS(VSS),.VDD(VDD),.Y(G62),.A(G59),.B(G11),.C(G60),.D(G61));
  AND2 AND2_8(.VSS(VSS),.VDD(VDD),.Y(G63),.A(G64),.B(G65));
  AND3 AND3_3(.VSS(VSS),.VDD(VDD),.Y(G74),.A(G12),.B(G14),.C(G19));
  AND3 AND3_4(.VSS(VSS),.VDD(VDD),.Y(G75),.A(G82),.B(G91),.C(G14));
  AND2 AND2_9(.VSS(VSS),.VDD(VDD),.Y(G88),.A(G14),.B(G87));
  AND2 AND2_10(.VSS(VSS),.VDD(VDD),.Y(G89),.A(G103),.B(G96));
  AND2 AND2_11(.VSS(VSS),.VDD(VDD),.Y(G90),.A(G91),.B(G103));
  AND2 AND2_12(.VSS(VSS),.VDD(VDD),.Y(G94),.A(G93),.B(G13));
  AND2 AND2_13(.VSS(VSS),.VDD(VDD),.Y(G95),.A(G96),.B(G13));
  AND3 AND3_5(.VSS(VSS),.VDD(VDD),.Y(G100),.A(G99),.B(G14),.C(G12));
  AND3 AND3_6(.VSS(VSS),.VDD(VDD),.Y(G105),.A(G103),.B(G108),.C(G104));
  AND2 AND2_14(.VSS(VSS),.VDD(VDD),.Y(G110),.A(G108),.B(G109));
  AND2 AND2_15(.VSS(VSS),.VDD(VDD),.Y(G111),.A(G10),.B(G112));
  AND2 AND2_16(.VSS(VSS),.VDD(VDD),.Y(G115),.A(G114),.B(G14));
  AND2 AND2_17(.VSS(VSS),.VDD(VDD),.Y(G122),.A(G120),.B(G121));
  AND2 AND2_18(.VSS(VSS),.VDD(VDD),.Y(G123),.A(G124),.B(G22));
  AND2 AND2_19(.VSS(VSS),.VDD(VDD),.Y(G128),.A(G126),.B(G127));
  AND2 AND2_20(.VSS(VSS),.VDD(VDD),.Y(G129),.A(G131),.B(G23));
//
  OR4 OR4_0(.VSS(VSS),.VDD(VDD),.Y(G24),.A(G38),.B(G46),.C(G45),.D(G40));
  OR3 OR3_0(.VSS(VSS),.VDD(VDD),.Y(G25),.A(G38),.B(G11),.C(G12));
  OR4 OR4_1(.VSS(VSS),.VDD(VDD),.Y(G68),.A(G11),.B(G12),.C(G13),.D(G96));
  OR2 OR2_0(.VSS(VSS),.VDD(VDD),.Y(G69),.A(G103),.B(G18));
  OR2 OR2_1(.VSS(VSS),.VDD(VDD),.Y(G70),.A(G103),.B(G14));
  OR3 OR3_1(.VSS(VSS),.VDD(VDD),.Y(G71),.A(G82),.B(G12),.C(G13));
  OR2 OR2_2(.VSS(VSS),.VDD(VDD),.Y(G72),.A(G91),.B(G20));
  OR2 OR2_3(.VSS(VSS),.VDD(VDD),.Y(G73),.A(G103),.B(G20));
  OR4 OR4_2(.VSS(VSS),.VDD(VDD),.Y(G77),.A(G112),.B(G103),.C(G96),.D(G19));
  OR2 OR2_4(.VSS(VSS),.VDD(VDD),.Y(G78),.A(G108),.B(G76));
  OR2 OR2_5(.VSS(VSS),.VDD(VDD),.Y(G79),.A(G103),.B(G14));
  OR2 OR2_6(.VSS(VSS),.VDD(VDD),.Y(G80),.A(G11),.B(G14));
  OR2 OR2_7(.VSS(VSS),.VDD(VDD),.Y(G81),.A(G12),.B(G13));
  OR4 OR4_3(.VSS(VSS),.VDD(VDD),.Y(G83),.A(G11),.B(G12),.C(G13),.D(G96));
  OR3 OR3_2(.VSS(VSS),.VDD(VDD),.Y(G84),.A(G82),.B(G91),.C(G14));
  OR3 OR3_3(.VSS(VSS),.VDD(VDD),.Y(G85),.A(G91),.B(G96),.C(G17));
//
  NAND3 NAND3_0(.VSS(VSS),.VDD(VDD),.Y(G41),.A(G12),.B(G11),.C(G10));
  NAND3 NAND3_1(.VSS(VSS),.VDD(VDD),.Y(G43),.A(G24),.B(G25),.C(G28));
  NAND4 NAND4_0(.VSS(VSS),.VDD(VDD),.Y(G52),.A(G13),.B(G45),.C(G46),.D(G10));
  NAND4 NAND4_1(.VSS(VSS),.VDD(VDD),.Y(G65),.A(G59),.B(G54),.C(G22),.D(G61));
  NAND4 NAND4_2(.VSS(VSS),.VDD(VDD),.Y(G97),.A(G83),.B(G84),.C(G85),.D(G108));
  NAND4 NAND4_3(.VSS(VSS),.VDD(VDD),.Y(G101),.A(G68),.B(G69),.C(G70),.D(G108));
  NAND2 NAND2_0(.VSS(VSS),.VDD(VDD),.Y(G106),.A(G77),.B(G78));
  NAND4 NAND4_4(.VSS(VSS),.VDD(VDD),.Y(G109),.A(G71),.B(G72),.C(G73),.D(G14));
  NAND4 NAND4_5(.VSS(VSS),.VDD(VDD),.Y(G116),.A(G79),.B(G80),.C(G81),.D(G108));
//
  NOR2 NOR2_0(.VSS(VSS),.VDD(VDD),.Y(G29),.A(G10),.B(G130));
  NOR4 NOR4_0(.VSS(VSS),.VDD(VDD),.Y(G30),.A(G31),.B(G32),.C(G33),.D(G130));
  NOR4 NOR4_1(.VSS(VSS),.VDD(VDD),.Y(G34),.A(G35),.B(G36),.C(G37),.D(G130));
  NOR2 NOR2_1(.VSS(VSS),.VDD(VDD),.Y(G39),.A(G42),.B(G43));
  NOR3 NOR3_0(.VSS(VSS),.VDD(VDD),.Y(G44),.A(G48),.B(G49),.C(G53));
  NOR2 NOR2_2(.VSS(VSS),.VDD(VDD),.Y(G47),.A(G50),.B(G40));
  NOR2 NOR2_3(.VSS(VSS),.VDD(VDD),.Y(G53),.A(G26),.B(G27));
  NOR3 NOR3_1(.VSS(VSS),.VDD(VDD),.Y(G56),.A(G57),.B(G58),.C(G130));
  NOR2 NOR2_4(.VSS(VSS),.VDD(VDD),.Y(G61),.A(G14),.B(G55));
  NOR4 NOR4_2(.VSS(VSS),.VDD(VDD),.Y(G86),.A(G88),.B(G89),.C(G90),.D(G112));
  NOR3 NOR3_2(.VSS(VSS),.VDD(VDD),.Y(G92),.A(G94),.B(G95),.C(G97));
  NOR2 NOR2_5(.VSS(VSS),.VDD(VDD),.Y(G98),.A(G100),.B(G101));
  NOR2 NOR2_6(.VSS(VSS),.VDD(VDD),.Y(G102),.A(G105),.B(G106));
  NOR2 NOR2_7(.VSS(VSS),.VDD(VDD),.Y(G104),.A(G74),.B(G75));
  NOR2 NOR2_8(.VSS(VSS),.VDD(VDD),.Y(G107),.A(G110),.B(G111));
  NOR2 NOR2_9(.VSS(VSS),.VDD(VDD),.Y(G112),.A(G62),.B(G63));
  NOR2 NOR2_10(.VSS(VSS),.VDD(VDD),.Y(G113),.A(G115),.B(G116));
  NOR3 NOR3_3(.VSS(VSS),.VDD(VDD),.Y(G119),.A(G122),.B(G123),.C(G130));
  NOR3 NOR3_4(.VSS(VSS),.VDD(VDD),.Y(G125),.A(G128),.B(G129),.C(G130));
//

endmodule