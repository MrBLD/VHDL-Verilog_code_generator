module s444w(G118,G2,G108,G119,G167,G168,VDD,G0,CLOCK,G1,G107,VSS);
input G2,VDD,G0,CLOCK,G1,VSS;
output G118,G108,G119,G167,G168,G107;

  wire G125,G146,G144,I272,G23,G113,G67,G31,G111,I181,I191,G36,G17,I212,G72,G155,G121,I236,G73,G70,I392,G139,G33,G128,G127,G22,G37,G48,I292,G76,G40,G74,I257,G130,G53,G43,G82,I200,G148,G30,G138,I256,I303,I226,G12,G96,G20,G59,G116,G19,G97,G65,G88,G42,G164,G54,G159,G145,G133,I190,I227,G38,G63,G149,G18,G102,G34,G115,G80,G78,G11,G162BF,G143,G24,G105,G58,I211,I282,G47,G120,G151,G85,I210,I201,G136,G92,G135,G71,G147,G87,G93,G55,G165,G14,G142,G161,G131,G50,I304,G103,G61,G21,G25,G62,G160,I105,G122,I225,G32,G106,G90,G15,G163,G81,G27,G132,G129,G79,G86,I246,I283,I291,G35,G52,G83,G68,G60,G91,G154,G57,G158,I302,I382,G101,G41,G16,G150,I192,I255,I293,G94,G134,I271,G166,I245,G56,G29,G51,G140,G66,G46,I182,G89,G98,I202,G13,G95,G137,G104,G110,G114,G49,G26,G100,G45,G162,G99,G69,I237,G64,I324,G156,G28,I273,I321,I235,G157,G44,I372,G141,G152,G126,G117,G109,G124,G84,G112,G123,G153,I180,I281,I247,G75,I336,I318,G77;
//# 3 inputs
//# 6 outputs
//# 21 D-type flipflops
//# 62 inverters
//# 119 gates (13 ANDs + 58 NANDs + 14 ORs + 34 NORs)
//
//
//
  MSFF DFF_0(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G11),.DATA(G37));
  MSFF DFF_1(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G12),.DATA(G41));
  MSFF DFF_2(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G13),.DATA(G45));
  MSFF DFF_3(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G14),.DATA(G49));
  MSFF DFF_4(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G15),.DATA(G58));
  MSFF DFF_5(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G16),.DATA(G62));
  MSFF DFF_6(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G17),.DATA(G66));
  MSFF DFF_7(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G18),.DATA(G70));
  MSFF DFF_8(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G19),.DATA(G80));
  MSFF DFF_9(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G20),.DATA(G84));
  MSFF DFF_10(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G21),.DATA(G88));
  MSFF DFF_11(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G22),.DATA(G92));
  MSFF DFF_12(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G23),.DATA(G101));
  MSFF DFF_13(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G24),.DATA(G162BF));
  MSFF DFF_14(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G25),.DATA(G109));
  MSFF DFF_15(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G26),.DATA(G110));
  MSFF DFF_16(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G27),.DATA(G111));
  MSFF DFF_17(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G28),.DATA(G112));
  MSFF DFF_18(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G29),.DATA(G113));
  MSFF DFF_19(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G30),.DATA(G114));
  MSFF DFF_20(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(G31),.DATA(G155));
//
  NOT NOT1_0(.VSS(VSS),.VDD(VDD),.Y(I372),.A(G0));
  NOT NOT1_1(.VSS(VSS),.VDD(VDD),.Y(I382),.A(G1));
  NOT NOT1_2(.VSS(VSS),.VDD(VDD),.Y(I318),.A(G2));
  NOT NOT1_3(.VSS(VSS),.VDD(VDD),.Y(G34),.A(G11));
  NOT NOT1_4(.VSS(VSS),.VDD(VDD),.Y(I180),.A(G11));
  NOT NOT1_5(.VSS(VSS),.VDD(VDD),.Y(G35),.A(G12));
  NOT NOT1_6(.VSS(VSS),.VDD(VDD),.Y(G77),.A(G20));
  NOT NOT1_7(.VSS(VSS),.VDD(VDD),.Y(G135),.A(G20));
  NOT NOT1_8(.VSS(VSS),.VDD(VDD),.Y(G36),.A(G13));
  NOT NOT1_9(.VSS(VSS),.VDD(VDD),.Y(G78),.A(G21));
  NOT NOT1_10(.VSS(VSS),.VDD(VDD),.Y(G144),.A(G21));
  NOT NOT1_11(.VSS(VSS),.VDD(VDD),.Y(G32),.A(G14));
  NOT NOT1_12(.VSS(VSS),.VDD(VDD),.Y(G74),.A(G22));
  NOT NOT1_13(.VSS(VSS),.VDD(VDD),.Y(G142),.A(G22));
  NOT NOT1_14(.VSS(VSS),.VDD(VDD),.Y(I392),.A(G30));
  NOT NOT1_15(.VSS(VSS),.VDD(VDD),.Y(G55),.A(G15));
  NOT NOT1_16(.VSS(VSS),.VDD(VDD),.Y(G102),.A(G23));
  NOT NOT1_17(.VSS(VSS),.VDD(VDD),.Y(G136),.A(G23));
  NOT NOT1_18(.VSS(VSS),.VDD(VDD),.Y(G156),.A(G31));
  NOT NOT1_19(.VSS(VSS),.VDD(VDD),.Y(G56),.A(G16));
  NOT NOT1_20(.VSS(VSS),.VDD(VDD),.Y(G143),.A(G24));
  NOT NOT1_21(.VSS(VSS),.VDD(VDD),.Y(G161),.A(G17));
  NOT NOT1_22(.VSS(VSS),.VDD(VDD),.Y(I321),.A(G25));
  NOT NOT1_23(.VSS(VSS),.VDD(VDD),.Y(G53),.A(G18));
  NOT NOT1_24(.VSS(VSS),.VDD(VDD),.Y(I324),.A(G26));
  NOT NOT1_25(.VSS(VSS),.VDD(VDD),.Y(G76),.A(G19));
  NOT NOT1_26(.VSS(VSS),.VDD(VDD),.Y(G150),.A(G19));
  NOT NOT1_27(.VSS(VSS),.VDD(VDD),.Y(I336),.A(G27));
  NOT NOT1_28(.VSS(VSS),.VDD(VDD),.Y(G119),.A(G28));
  NOT NOT1_29(.VSS(VSS),.VDD(VDD),.Y(G167),.A(G29));
  NOT NOT1_30(.VSS(VSS),.VDD(VDD),.Y(G152),.A(I372));
  NOT NOT1_31(.VSS(VSS),.VDD(VDD),.Y(G160),.A(I382));
  NOT NOT1_32(.VSS(VSS),.VDD(VDD),.Y(G106),.A(I318));
  NOT NOT1_33(.VSS(VSS),.VDD(VDD),.Y(G43),.A(G34));
  NOT NOT1_34(.VSS(VSS),.VDD(VDD),.Y(I182),.A(I180));
  NOT NOT1_35(.VSS(VSS),.VDD(VDD),.Y(G168),.A(I392));
  NOT NOT1_36(.VSS(VSS),.VDD(VDD),.Y(G107),.A(I321));
  NOT NOT1_37(.VSS(VSS),.VDD(VDD),.Y(G108),.A(I324));
  NOT NOT1_38(.VSS(VSS),.VDD(VDD),.Y(G118),.A(I336));
  NOT NOT1_39(.VSS(VSS),.VDD(VDD),.Y(G99),.A(G152));
  NOT NOT1_40(.VSS(VSS),.VDD(VDD),.Y(G139),.A(G152));
  NOT NOT1_41(.VSS(VSS),.VDD(VDD),.Y(G153),.A(G152));
  NOT NOT1_42(.VSS(VSS),.VDD(VDD),.Y(G157),.A(G160));
  NOT NOT1_43(.VSS(VSS),.VDD(VDD),.Y(G103),.A(G106));
  NOT NOT1_44(.VSS(VSS),.VDD(VDD),.Y(G38),.A(G40));
  NOT NOT1_45(.VSS(VSS),.VDD(VDD),.Y(G60),.A(G57));
  NOT NOT1_46(.VSS(VSS),.VDD(VDD),.Y(G79),.A(G97));
  NOT NOT1_47(.VSS(VSS),.VDD(VDD),.Y(G42),.A(G44));
  NOT NOT1_48(.VSS(VSS),.VDD(VDD),.Y(G46),.A(G48));
  NOT NOT1_49(.VSS(VSS),.VDD(VDD),.Y(I105),.A(G162));
  NOT NOT1_50(.VSS(VSS),.VDD(VDD),.Y(G166),.A(G162));
  NOT NOT1_51(.VSS(VSS),.VDD(VDD),.Y(G50),.A(G52));
  NOT NOT1_52(.VSS(VSS),.VDD(VDD),.Y(G82),.A(G79));
  NOT NOT1_53(.VSS(VSS),.VDD(VDD),.Y(G162BF),.A(I105));
  NOT NOT1_54(.VSS(VSS),.VDD(VDD),.Y(G59),.A(G61));
  NOT NOT1_55(.VSS(VSS),.VDD(VDD),.Y(G63),.A(G65));
  NOT NOT1_56(.VSS(VSS),.VDD(VDD),.Y(G67),.A(G69));
  NOT NOT1_57(.VSS(VSS),.VDD(VDD),.Y(G71),.A(G73));
  NOT NOT1_58(.VSS(VSS),.VDD(VDD),.Y(G81),.A(G83));
  NOT NOT1_59(.VSS(VSS),.VDD(VDD),.Y(G85),.A(G87));
  NOT NOT1_60(.VSS(VSS),.VDD(VDD),.Y(G89),.A(G91));
  NOT NOT1_61(.VSS(VSS),.VDD(VDD),.Y(G94),.A(G96));
//
  AND2 AND2_0(.VSS(VSS),.VDD(VDD),.Y(G122),.A(G24),.B(G121));
  AND3 AND3_0(.VSS(VSS),.VDD(VDD),.Y(G124),.A(G139),.B(G22),.C(G150));
  AND3 AND3_1(.VSS(VSS),.VDD(VDD),.Y(G125),.A(G139),.B(G20),.C(G19));
  AND2 AND2_1(.VSS(VSS),.VDD(VDD),.Y(G126),.A(G139),.B(G21));
  AND2 AND2_2(.VSS(VSS),.VDD(VDD),.Y(G127),.A(G139),.B(G24));
  AND2 AND2_3(.VSS(VSS),.VDD(VDD),.Y(G154),.A(G158),.B(G159));
  AND2 AND2_4(.VSS(VSS),.VDD(VDD),.Y(G100),.A(G104),.B(G105));
  AND2 AND2_5(.VSS(VSS),.VDD(VDD),.Y(G155),.A(G154),.B(G153));
  AND2 AND2_6(.VSS(VSS),.VDD(VDD),.Y(G101),.A(G100),.B(G99));
  AND3 AND3_2(.VSS(VSS),.VDD(VDD),.Y(G115),.A(G161),.B(G117),.C(G162));
  AND3 AND3_3(.VSS(VSS),.VDD(VDD),.Y(G163),.A(G161),.B(G165),.C(G162));
  AND2 AND2_7(.VSS(VSS),.VDD(VDD),.Y(G116),.A(G117),.B(G166));
  AND2 AND2_8(.VSS(VSS),.VDD(VDD),.Y(G164),.A(G165),.B(G166));
//
  OR3 OR3_0(.VSS(VSS),.VDD(VDD),.Y(G141),.A(G24),.B(G22),.C(G21));
  OR3 OR3_1(.VSS(VSS),.VDD(VDD),.Y(G137),.A(G136),.B(G20),.C(G19));
  OR2 OR2_0(.VSS(VSS),.VDD(VDD),.Y(G138),.A(G136),.B(G142));
  OR4 OR4_0(.VSS(VSS),.VDD(VDD),.Y(G140),.A(G24),.B(G21),.C(G20),.D(G150));
  OR4 OR4_1(.VSS(VSS),.VDD(VDD),.Y(G133),.A(G152),.B(G136),.C(G22),.D(G144));
  OR3 OR3_2(.VSS(VSS),.VDD(VDD),.Y(G134),.A(G152),.B(G142),.C(G21));
  OR4 OR4_2(.VSS(VSS),.VDD(VDD),.Y(G145),.A(G152),.B(G142),.C(G20),.D(G19));
  OR2 OR2_1(.VSS(VSS),.VDD(VDD),.Y(G146),.A(G152),.B(G143));
  OR2 OR2_2(.VSS(VSS),.VDD(VDD),.Y(G147),.A(G152),.B(G144));
  OR2 OR2_3(.VSS(VSS),.VDD(VDD),.Y(G158),.A(G31),.B(G160));
  OR2 OR2_4(.VSS(VSS),.VDD(VDD),.Y(G104),.A(G23),.B(G106));
  OR4 OR4_3(.VSS(VSS),.VDD(VDD),.Y(G131),.A(G144),.B(G22),.C(G23),.D(G129));
  OR2 OR2_5(.VSS(VSS),.VDD(VDD),.Y(G159),.A(G156),.B(G157));
  OR2 OR2_6(.VSS(VSS),.VDD(VDD),.Y(G105),.A(G102),.B(G103));
//
  NAND2 NAND2_0(.VSS(VSS),.VDD(VDD),.Y(I181),.A(G11),.B(I180));
  NAND2 NAND2_1(.VSS(VSS),.VDD(VDD),.Y(G129),.A(G19),.B(G135));
  NAND4 NAND4_0(.VSS(VSS),.VDD(VDD),.Y(G121),.A(G19),.B(G135),.C(G142),.D(G136));
  NAND2 NAND2_2(.VSS(VSS),.VDD(VDD),.Y(I190),.A(G12),.B(G43));
  NAND2 NAND2_3(.VSS(VSS),.VDD(VDD),.Y(G40),.A(I181),.B(I182));
  NAND2 NAND2_4(.VSS(VSS),.VDD(VDD),.Y(I200),.A(G13),.B(G47));
  NAND2 NAND2_5(.VSS(VSS),.VDD(VDD),.Y(I210),.A(G14),.B(G51));
  NAND2 NAND2_6(.VSS(VSS),.VDD(VDD),.Y(G120),.A(G150),.B(G128));
  NAND2 NAND2_7(.VSS(VSS),.VDD(VDD),.Y(G132),.A(G133),.B(G134));
  NAND3 NAND3_0(.VSS(VSS),.VDD(VDD),.Y(G111),.A(G140),.B(G141),.C(G139));
  NAND4 NAND4_1(.VSS(VSS),.VDD(VDD),.Y(G123),.A(G137),.B(G138),.C(G21),.D(G139));
  NAND4 NAND4_2(.VSS(VSS),.VDD(VDD),.Y(G151),.A(G20),.B(G144),.C(G143),.D(G139));
  NAND3 NAND3_1(.VSS(VSS),.VDD(VDD),.Y(G117),.A(G145),.B(G146),.C(G147));
  NAND2 NAND2_8(.VSS(VSS),.VDD(VDD),.Y(I191),.A(G12),.B(I190));
  NAND2 NAND2_9(.VSS(VSS),.VDD(VDD),.Y(I192),.A(G43),.B(I190));
  NAND2 NAND2_10(.VSS(VSS),.VDD(VDD),.Y(I201),.A(G13),.B(I200));
  NAND2 NAND2_11(.VSS(VSS),.VDD(VDD),.Y(I202),.A(G47),.B(I200));
  NAND2 NAND2_12(.VSS(VSS),.VDD(VDD),.Y(G149),.A(G131),.B(G130));
  NAND2 NAND2_13(.VSS(VSS),.VDD(VDD),.Y(I211),.A(G14),.B(I210));
  NAND2 NAND2_14(.VSS(VSS),.VDD(VDD),.Y(I212),.A(G51),.B(I210));
  NAND3 NAND3_2(.VSS(VSS),.VDD(VDD),.Y(G148),.A(G150),.B(G135),.C(G132));
  NAND2 NAND2_15(.VSS(VSS),.VDD(VDD),.Y(G44),.A(I191),.B(I192));
  NAND2 NAND2_16(.VSS(VSS),.VDD(VDD),.Y(G48),.A(I201),.B(I202));
  NAND2 NAND2_17(.VSS(VSS),.VDD(VDD),.Y(G162),.A(G120),.B(G149));
  NAND2 NAND2_18(.VSS(VSS),.VDD(VDD),.Y(G52),.A(I211),.B(I212));
  NAND2 NAND2_19(.VSS(VSS),.VDD(VDD),.Y(I225),.A(G15),.B(G60));
  NAND2 NAND2_20(.VSS(VSS),.VDD(VDD),.Y(I235),.A(G16),.B(G64));
  NAND2 NAND2_21(.VSS(VSS),.VDD(VDD),.Y(I245),.A(G17),.B(G68));
  NAND2 NAND2_22(.VSS(VSS),.VDD(VDD),.Y(I255),.A(G18),.B(G72));
  NAND2 NAND2_23(.VSS(VSS),.VDD(VDD),.Y(G165),.A(G148),.B(G149));
  NAND2 NAND2_24(.VSS(VSS),.VDD(VDD),.Y(I226),.A(G15),.B(I225));
  NAND2 NAND2_25(.VSS(VSS),.VDD(VDD),.Y(I227),.A(G60),.B(I225));
  NAND2 NAND2_26(.VSS(VSS),.VDD(VDD),.Y(I236),.A(G16),.B(I235));
  NAND2 NAND2_27(.VSS(VSS),.VDD(VDD),.Y(I237),.A(G64),.B(I235));
  NAND2 NAND2_28(.VSS(VSS),.VDD(VDD),.Y(I246),.A(G17),.B(I245));
  NAND2 NAND2_29(.VSS(VSS),.VDD(VDD),.Y(I247),.A(G68),.B(I245));
  NAND2 NAND2_30(.VSS(VSS),.VDD(VDD),.Y(I256),.A(G18),.B(I255));
  NAND2 NAND2_31(.VSS(VSS),.VDD(VDD),.Y(I257),.A(G72),.B(I255));
  NAND2 NAND2_32(.VSS(VSS),.VDD(VDD),.Y(G61),.A(I226),.B(I227));
  NAND2 NAND2_33(.VSS(VSS),.VDD(VDD),.Y(G65),.A(I236),.B(I237));
  NAND2 NAND2_34(.VSS(VSS),.VDD(VDD),.Y(G69),.A(I246),.B(I247));
  NAND2 NAND2_35(.VSS(VSS),.VDD(VDD),.Y(G73),.A(I256),.B(I257));
  NAND2 NAND2_36(.VSS(VSS),.VDD(VDD),.Y(I271),.A(G19),.B(G82));
  NAND2 NAND2_37(.VSS(VSS),.VDD(VDD),.Y(I281),.A(G20),.B(G86));
  NAND2 NAND2_38(.VSS(VSS),.VDD(VDD),.Y(I291),.A(G21),.B(G90));
  NAND2 NAND2_39(.VSS(VSS),.VDD(VDD),.Y(I302),.A(G22),.B(G95));
  NAND2 NAND2_40(.VSS(VSS),.VDD(VDD),.Y(I272),.A(G19),.B(I271));
  NAND2 NAND2_41(.VSS(VSS),.VDD(VDD),.Y(I273),.A(G82),.B(I271));
  NAND2 NAND2_42(.VSS(VSS),.VDD(VDD),.Y(I282),.A(G20),.B(I281));
  NAND2 NAND2_43(.VSS(VSS),.VDD(VDD),.Y(I283),.A(G86),.B(I281));
  NAND2 NAND2_44(.VSS(VSS),.VDD(VDD),.Y(I292),.A(G21),.B(I291));
  NAND2 NAND2_45(.VSS(VSS),.VDD(VDD),.Y(I293),.A(G90),.B(I291));
  NAND2 NAND2_46(.VSS(VSS),.VDD(VDD),.Y(I303),.A(G22),.B(I302));
  NAND2 NAND2_47(.VSS(VSS),.VDD(VDD),.Y(I304),.A(G95),.B(I302));
  NAND2 NAND2_48(.VSS(VSS),.VDD(VDD),.Y(G83),.A(I272),.B(I273));
  NAND2 NAND2_49(.VSS(VSS),.VDD(VDD),.Y(G87),.A(I282),.B(I283));
  NAND2 NAND2_50(.VSS(VSS),.VDD(VDD),.Y(G91),.A(I292),.B(I293));
  NAND2 NAND2_51(.VSS(VSS),.VDD(VDD),.Y(G96),.A(I303),.B(I304));
//
  NOR3 NOR3_0(.VSS(VSS),.VDD(VDD),.Y(G33),.A(G11),.B(G12),.C(G13));
  NOR3 NOR3_1(.VSS(VSS),.VDD(VDD),.Y(G54),.A(G15),.B(G16),.C(G17));
  NOR3 NOR3_2(.VSS(VSS),.VDD(VDD),.Y(G75),.A(G19),.B(G20),.C(G21));
  NOR2 NOR2_0(.VSS(VSS),.VDD(VDD),.Y(G47),.A(G34),.B(G35));
  NOR3 NOR3_3(.VSS(VSS),.VDD(VDD),.Y(G51),.A(G34),.B(G35),.C(G36));
  NOR2 NOR2_1(.VSS(VSS),.VDD(VDD),.Y(G98),.A(G32),.B(G33));
  NOR4 NOR4_0(.VSS(VSS),.VDD(VDD),.Y(G128),.A(G20),.B(G144),.C(G136),.D(G152));
  NOR2 NOR2_2(.VSS(VSS),.VDD(VDD),.Y(G130),.A(G143),.B(G152));
  NOR2 NOR2_3(.VSS(VSS),.VDD(VDD),.Y(G57),.A(G31),.B(G98));
  NOR2 NOR2_4(.VSS(VSS),.VDD(VDD),.Y(G64),.A(G55),.B(G57));
  NOR3 NOR3_4(.VSS(VSS),.VDD(VDD),.Y(G68),.A(G55),.B(G56),.C(G57));
  NOR4 NOR4_1(.VSS(VSS),.VDD(VDD),.Y(G72),.A(G55),.B(G56),.C(G161),.D(G57));
  NOR3 NOR3_5(.VSS(VSS),.VDD(VDD),.Y(G97),.A(G53),.B(G57),.C(G54));
  NOR2 NOR2_5(.VSS(VSS),.VDD(VDD),.Y(G109),.A(G122),.B(G123));
  NOR4 NOR4_2(.VSS(VSS),.VDD(VDD),.Y(G110),.A(G124),.B(G125),.C(G126),.D(G127));
  NOR2 NOR2_6(.VSS(VSS),.VDD(VDD),.Y(G114),.A(G150),.B(G151));
  NOR3 NOR3_6(.VSS(VSS),.VDD(VDD),.Y(G37),.A(G98),.B(G38),.C(G152));
  NOR2 NOR2_7(.VSS(VSS),.VDD(VDD),.Y(G86),.A(G76),.B(G79));
  NOR3 NOR3_7(.VSS(VSS),.VDD(VDD),.Y(G90),.A(G76),.B(G77),.C(G79));
  NOR3 NOR3_8(.VSS(VSS),.VDD(VDD),.Y(G93),.A(G74),.B(G79),.C(G75));
  NOR4 NOR4_3(.VSS(VSS),.VDD(VDD),.Y(G95),.A(G76),.B(G77),.C(G78),.D(G79));
  NOR3 NOR3_9(.VSS(VSS),.VDD(VDD),.Y(G41),.A(G98),.B(G42),.C(G152));
  NOR3 NOR3_10(.VSS(VSS),.VDD(VDD),.Y(G45),.A(G98),.B(G46),.C(G152));
  NOR3 NOR3_11(.VSS(VSS),.VDD(VDD),.Y(G49),.A(G98),.B(G50),.C(G152));
  NOR2 NOR2_8(.VSS(VSS),.VDD(VDD),.Y(G112),.A(G115),.B(G116));
  NOR2 NOR2_9(.VSS(VSS),.VDD(VDD),.Y(G113),.A(G163),.B(G164));
  NOR3 NOR3_12(.VSS(VSS),.VDD(VDD),.Y(G58),.A(G97),.B(G59),.C(G152));
  NOR3 NOR3_13(.VSS(VSS),.VDD(VDD),.Y(G62),.A(G97),.B(G63),.C(G152));
  NOR3 NOR3_14(.VSS(VSS),.VDD(VDD),.Y(G66),.A(G97),.B(G67),.C(G152));
  NOR3 NOR3_15(.VSS(VSS),.VDD(VDD),.Y(G70),.A(G97),.B(G71),.C(G152));
  NOR3 NOR3_16(.VSS(VSS),.VDD(VDD),.Y(G80),.A(G93),.B(G81),.C(G152));
  NOR3 NOR3_17(.VSS(VSS),.VDD(VDD),.Y(G84),.A(G93),.B(G85),.C(G152));
  NOR3 NOR3_18(.VSS(VSS),.VDD(VDD),.Y(G88),.A(G93),.B(G89),.C(G152));
  NOR3 NOR3_19(.VSS(VSS),.VDD(VDD),.Y(G92),.A(G93),.B(G94),.C(G152));
//

endmodule