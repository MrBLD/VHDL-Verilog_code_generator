module s386w(v13_D_12,v13_D_10,v13_D_6,v2,v13_D_9,v13_D_7,v1,v4,v0,v5,v13_D_11,CLOCK,VDD,VSS,v13_D_8,v3,v6);
input v2,v1,v4,v0,v5,CLOCK,VDD,VSS,v3,v6;
output v13_D_10,v13_D_6,v13_D_9,v13_D_7,v13_D_11,v13_D_8,v13_D_12;

  wire B35B,B30B,I228,I43,I109,B38B,B39B,v13_D_2,I234,v7,Lv13_D_7,I69,Lv13_D_4,v7bar,I76,v8,v5bar,I25,I124,I89,v11,I198,I87,I207,v13_D_1,I84,I63,B43B,B15B,B26B,I204,Lv13_D_5,I65,I108,Lv13_D_0,I104,I167,B44B,I114,I22,B17B,I60,I106,I30,v9bar,I71,Lv13_D_10,v6bar,I50,I77,v13_D_3,B21B,B40B,I103,v11bar,I17,I91,I93,I53,B19B,I216,I27,v3bar,II98,v13_D_5,v8bar,B34B,v9,I210,Lv13_D_6,I79,I90,I102,I158,v12bar,I74,I39,I94,I231,I186,v12,Lv13_D_1,I225,Lv13_D_9,I28,B32B,I47,B14B,I56,I175,I192,B20B,B24B,B25B,B14Bbar,B35Bbar,B31B,II65,B28B,I73,I48,I35,I201,B45B,v1bar,v13_D_0,Lv13_D_8,I51,I44,Lv13_D_12,B16B,I222,v10,I54,I66,I18,Lv13_D_3,B23B,I40,B29B,I96,I36,I57,I171,B33B,B41B,I100,I148,Lv13_D_11,I31,I113,I98,I64,v4bar,B42B,I195,v0bar,B22B,I111,B37B,B27B,I85,I62,v13_D_4,I213,Lv13_D_2,B34Bbar,I41,v10bar,B18B,B36B,I164,I24,I59,I219,I105,I97,I21;
//# 7 inputs
//# 7 outputs
//# 6 D-type flipflops
//# 41 inverters
//# 118 gates (83 ANDs + 0 NANDs + 35 ORs + 0 NORs)
//
//
//
  MSFF DFF_0(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(v12),.DATA(v13_D_5));
  MSFF DFF_1(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(v11),.DATA(v13_D_4));
  MSFF DFF_2(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(v10),.DATA(v13_D_3));
  MSFF DFF_3(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(v9),.DATA(v13_D_2));
  MSFF DFF_4(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(v8),.DATA(v13_D_1));
  MSFF DFF_5(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(v7),.DATA(v13_D_0));
//
  NOT NOT1_0(.VSS(VSS),.VDD(VDD),.Y(v3bar),.A(v3));
  NOT NOT1_1(.VSS(VSS),.VDD(VDD),.Y(v6bar),.A(v6));
  NOT NOT1_2(.VSS(VSS),.VDD(VDD),.Y(v5bar),.A(v5));
  NOT NOT1_3(.VSS(VSS),.VDD(VDD),.Y(B35Bbar),.A(B35B));
  NOT NOT1_4(.VSS(VSS),.VDD(VDD),.Y(B14Bbar),.A(B14B));
  NOT NOT1_5(.VSS(VSS),.VDD(VDD),.Y(B34Bbar),.A(B34B));
  NOT NOT1_6(.VSS(VSS),.VDD(VDD),.Y(v4bar),.A(v4));
  NOT NOT1_7(.VSS(VSS),.VDD(VDD),.Y(v11bar),.A(v11));
  NOT NOT1_8(.VSS(VSS),.VDD(VDD),.Y(v8bar),.A(v8));
  NOT NOT1_9(.VSS(VSS),.VDD(VDD),.Y(v7bar),.A(v7));
  NOT NOT1_10(.VSS(VSS),.VDD(VDD),.Y(v12bar),.A(v12));
  NOT NOT1_11(.VSS(VSS),.VDD(VDD),.Y(v0bar),.A(v0));
  NOT NOT1_12(.VSS(VSS),.VDD(VDD),.Y(v10bar),.A(v10));
  NOT NOT1_13(.VSS(VSS),.VDD(VDD),.Y(v9bar),.A(v9));
  NOT NOT1_14(.VSS(VSS),.VDD(VDD),.Y(v1bar),.A(v1));
  NOT NOT1_15(.VSS(VSS),.VDD(VDD),.Y(I198),.A(Lv13_D_12));
  NOT NOT1_16(.VSS(VSS),.VDD(VDD),.Y(v13_D_12),.A(I198));
  NOT NOT1_17(.VSS(VSS),.VDD(VDD),.Y(I201),.A(Lv13_D_11));
  NOT NOT1_18(.VSS(VSS),.VDD(VDD),.Y(v13_D_11),.A(I201));
  NOT NOT1_19(.VSS(VSS),.VDD(VDD),.Y(I204),.A(Lv13_D_10));
  NOT NOT1_20(.VSS(VSS),.VDD(VDD),.Y(v13_D_10),.A(I204));
  NOT NOT1_21(.VSS(VSS),.VDD(VDD),.Y(I207),.A(Lv13_D_9));
  NOT NOT1_22(.VSS(VSS),.VDD(VDD),.Y(v13_D_9),.A(I207));
  NOT NOT1_23(.VSS(VSS),.VDD(VDD),.Y(I210),.A(Lv13_D_8));
  NOT NOT1_24(.VSS(VSS),.VDD(VDD),.Y(v13_D_8),.A(I210));
  NOT NOT1_25(.VSS(VSS),.VDD(VDD),.Y(I213),.A(Lv13_D_7));
  NOT NOT1_26(.VSS(VSS),.VDD(VDD),.Y(v13_D_7),.A(I213));
  NOT NOT1_27(.VSS(VSS),.VDD(VDD),.Y(I216),.A(Lv13_D_6));
  NOT NOT1_28(.VSS(VSS),.VDD(VDD),.Y(v13_D_6),.A(I216));
  NOT NOT1_29(.VSS(VSS),.VDD(VDD),.Y(I219),.A(Lv13_D_5));
  NOT NOT1_30(.VSS(VSS),.VDD(VDD),.Y(v13_D_5),.A(I219));
  NOT NOT1_31(.VSS(VSS),.VDD(VDD),.Y(I222),.A(Lv13_D_4));
  NOT NOT1_32(.VSS(VSS),.VDD(VDD),.Y(v13_D_4),.A(I222));
  NOT NOT1_33(.VSS(VSS),.VDD(VDD),.Y(I225),.A(Lv13_D_3));
  NOT NOT1_34(.VSS(VSS),.VDD(VDD),.Y(v13_D_3),.A(I225));
  NOT NOT1_35(.VSS(VSS),.VDD(VDD),.Y(I228),.A(Lv13_D_2));
  NOT NOT1_36(.VSS(VSS),.VDD(VDD),.Y(v13_D_2),.A(I228));
  NOT NOT1_37(.VSS(VSS),.VDD(VDD),.Y(I231),.A(Lv13_D_1));
  NOT NOT1_38(.VSS(VSS),.VDD(VDD),.Y(v13_D_1),.A(I231));
  NOT NOT1_39(.VSS(VSS),.VDD(VDD),.Y(I234),.A(Lv13_D_0));
  NOT NOT1_40(.VSS(VSS),.VDD(VDD),.Y(v13_D_0),.A(I234));
//
  AND4 AND4_0(.VSS(VSS),.VDD(VDD),.Y(I64),.A(v0bar),.B(v5),.C(v7bar),.D(v8bar));
  AND4 AND4_1(.VSS(VSS),.VDD(VDD),.Y(I65),.A(v9),.B(v10),.C(v11bar),.D(v12bar));
  AND2 AND2_0(.VSS(VSS),.VDD(VDD),.Y(Lv13_D_12),.A(I64),.B(I65));
  AND2 AND2_1(.VSS(VSS),.VDD(VDD),.Y(I114),.A(v9bar),.B(v12bar));
  AND2 AND2_2(.VSS(VSS),.VDD(VDD),.Y(I113),.A(v7bar),.B(v8bar));
  AND2 AND2_3(.VSS(VSS),.VDD(VDD),.Y(I111),.A(v7bar),.B(v8bar));
  AND3 AND3_0(.VSS(VSS),.VDD(VDD),.Y(I109),.A(v3bar),.B(v4bar),.C(v11bar));
  AND2 AND2_4(.VSS(VSS),.VDD(VDD),.Y(I108),.A(v7),.B(v11));
  AND4 AND4_2(.VSS(VSS),.VDD(VDD),.Y(I106),.A(v5bar),.B(v7bar),.C(v11),.D(v12));
  AND3 AND3_1(.VSS(VSS),.VDD(VDD),.Y(I105),.A(v2),.B(v11bar),.C(v12bar));
  AND3 AND3_2(.VSS(VSS),.VDD(VDD),.Y(I103),.A(v8),.B(v11),.C(v12bar));
  AND3 AND3_3(.VSS(VSS),.VDD(VDD),.Y(I102),.A(v8bar),.B(v11bar),.C(v12));
  AND2 AND2_5(.VSS(VSS),.VDD(VDD),.Y(I100),.A(v2),.B(v8bar));
  AND2 AND2_6(.VSS(VSS),.VDD(VDD),.Y(II98),.A(v0),.B(v5));
  AND2 AND2_7(.VSS(VSS),.VDD(VDD),.Y(I96),.A(v1),.B(v9bar));
  AND3 AND3_4(.VSS(VSS),.VDD(VDD),.Y(I89),.A(v5bar),.B(v7bar),.C(v8bar));
  AND3 AND3_5(.VSS(VSS),.VDD(VDD),.Y(I94),.A(v10),.B(v11bar),.C(I89));
  AND2 AND2_8(.VSS(VSS),.VDD(VDD),.Y(I93),.A(v9bar),.B(v10bar));
  AND3 AND3_6(.VSS(VSS),.VDD(VDD),.Y(I91),.A(v0),.B(v11bar),.C(v12bar));
  AND2 AND2_9(.VSS(VSS),.VDD(VDD),.Y(I90),.A(v9bar),.B(v10bar));
  AND4 AND4_3(.VSS(VSS),.VDD(VDD),.Y(I97),.A(v0),.B(v6bar),.C(v7bar),.D(v8bar));
  AND4 AND4_4(.VSS(VSS),.VDD(VDD),.Y(I98),.A(v9bar),.B(v10),.C(v11bar),.D(v12bar));
  AND2 AND2_10(.VSS(VSS),.VDD(VDD),.Y(Lv13_D_8),.A(I97),.B(I98));
  AND4 AND4_5(.VSS(VSS),.VDD(VDD),.Y(I87),.A(v5bar),.B(v9),.C(v11bar),.D(v12bar));
  AND3 AND3_7(.VSS(VSS),.VDD(VDD),.Y(I104),.A(v2),.B(v3),.C(v8));
  AND3 AND3_8(.VSS(VSS),.VDD(VDD),.Y(I85),.A(v11bar),.B(v12bar),.C(I104));
  AND3 AND3_9(.VSS(VSS),.VDD(VDD),.Y(I84),.A(v8bar),.B(v11),.C(v12));
  AND2 AND2_11(.VSS(VSS),.VDD(VDD),.Y(I79),.A(v11bar),.B(v12bar));
  AND3 AND3_10(.VSS(VSS),.VDD(VDD),.Y(I77),.A(v0),.B(v8bar),.C(v10));
  AND4 AND4_6(.VSS(VSS),.VDD(VDD),.Y(I76),.A(v1bar),.B(v4),.C(v10bar),.D(B34Bbar));
  AND3 AND3_11(.VSS(VSS),.VDD(VDD),.Y(I74),.A(v7),.B(v8bar),.C(v11));
  AND3 AND3_12(.VSS(VSS),.VDD(VDD),.Y(I73),.A(v4bar),.B(v11bar),.C(B34Bbar));
  AND3 AND3_13(.VSS(VSS),.VDD(VDD),.Y(I71),.A(v4bar),.B(v11bar),.C(B34Bbar));
  AND2 AND2_12(.VSS(VSS),.VDD(VDD),.Y(I69),.A(v7),.B(v11bar));
  AND4 AND4_7(.VSS(VSS),.VDD(VDD),.Y(I124),.A(B40B),.B(v1),.C(v7bar),.D(v8bar));
  AND4 AND4_8(.VSS(VSS),.VDD(VDD),.Y(Lv13_D_10),.A(v9),.B(v11bar),.C(v12bar),.D(I124));
  AND2 AND2_13(.VSS(VSS),.VDD(VDD),.Y(I66),.A(v4),.B(v7));
  AND2 AND2_14(.VSS(VSS),.VDD(VDD),.Y(II65),.A(B35B),.B(B34B));
  AND3 AND3_14(.VSS(VSS),.VDD(VDD),.Y(I63),.A(v9bar),.B(v10bar),.C(v12bar));
  AND3 AND3_15(.VSS(VSS),.VDD(VDD),.Y(I62),.A(B23B),.B(v7bar),.C(v8bar));
  AND2 AND2_15(.VSS(VSS),.VDD(VDD),.Y(I60),.A(v1),.B(B42B));
  AND3 AND3_16(.VSS(VSS),.VDD(VDD),.Y(I59),.A(B43B),.B(v8),.C(v12bar));
  AND2 AND2_16(.VSS(VSS),.VDD(VDD),.Y(I57),.A(B32B),.B(v7bar));
  AND3 AND3_17(.VSS(VSS),.VDD(VDD),.Y(I56),.A(v11),.B(v12bar),.C(B14Bbar));
  AND3 AND3_18(.VSS(VSS),.VDD(VDD),.Y(I54),.A(v0bar),.B(v9bar),.C(v10bar));
  AND2 AND2_17(.VSS(VSS),.VDD(VDD),.Y(I53),.A(B27B),.B(v1));
  AND3 AND3_19(.VSS(VSS),.VDD(VDD),.Y(I51),.A(v9bar),.B(v10bar),.C(v12bar));
  AND3 AND3_20(.VSS(VSS),.VDD(VDD),.Y(I50),.A(B21B),.B(v7bar),.C(v8bar));
  AND2 AND2_18(.VSS(VSS),.VDD(VDD),.Y(I48),.A(B14B),.B(v11));
  AND3 AND3_21(.VSS(VSS),.VDD(VDD),.Y(I47),.A(v4bar),.B(v11bar),.C(B34Bbar));
  AND3 AND3_22(.VSS(VSS),.VDD(VDD),.Y(I148),.A(B38B),.B(v0),.C(v1bar));
  AND4 AND4_9(.VSS(VSS),.VDD(VDD),.Y(Lv13_D_7),.A(v9bar),.B(v10bar),.C(v12bar),.D(I148));
  AND2 AND2_19(.VSS(VSS),.VDD(VDD),.Y(I44),.A(v8bar),.B(B29B));
  AND2 AND2_20(.VSS(VSS),.VDD(VDD),.Y(I43),.A(B30B),.B(v12bar));
  AND3 AND3_23(.VSS(VSS),.VDD(VDD),.Y(I41),.A(v4),.B(v11bar),.C(B17B));
  AND3 AND3_24(.VSS(VSS),.VDD(VDD),.Y(I40),.A(v3),.B(v8),.C(B16B));
  AND4 AND4_10(.VSS(VSS),.VDD(VDD),.Y(I39),.A(v5),.B(v7),.C(v8bar),.D(v11));
  AND3 AND3_25(.VSS(VSS),.VDD(VDD),.Y(I158),.A(B39B),.B(v7bar),.C(v9bar));
  AND3 AND3_26(.VSS(VSS),.VDD(VDD),.Y(Lv13_D_9),.A(v11bar),.B(v12bar),.C(I158));
  AND4 AND4_11(.VSS(VSS),.VDD(VDD),.Y(I36),.A(v7bar),.B(v8bar),.C(B25B),.D(B26B));
  AND2 AND2_21(.VSS(VSS),.VDD(VDD),.Y(I35),.A(B28B),.B(v12bar));
  AND3 AND3_27(.VSS(VSS),.VDD(VDD),.Y(I164),.A(B15B),.B(v0),.C(v1bar));
  AND4 AND4_12(.VSS(VSS),.VDD(VDD),.Y(Lv13_D_0),.A(v9bar),.B(v10bar),.C(v12bar),.D(I164));
  AND3 AND3_28(.VSS(VSS),.VDD(VDD),.Y(I167),.A(B33B),.B(v0),.C(v1bar));
  AND3 AND3_29(.VSS(VSS),.VDD(VDD),.Y(Lv13_D_5),.A(v9bar),.B(v10bar),.C(I167));
  AND3 AND3_30(.VSS(VSS),.VDD(VDD),.Y(I31),.A(B36B),.B(v11bar),.C(v12bar));
  AND3 AND3_31(.VSS(VSS),.VDD(VDD),.Y(I171),.A(v5),.B(v7bar),.C(v8bar));
  AND3 AND3_32(.VSS(VSS),.VDD(VDD),.Y(I30),.A(v11),.B(v12),.C(I171));
  AND3 AND3_33(.VSS(VSS),.VDD(VDD),.Y(I175),.A(v0),.B(v7bar),.C(v8bar));
  AND4 AND4_13(.VSS(VSS),.VDD(VDD),.Y(I28),.A(v10),.B(v11bar),.C(v12bar),.D(I175));
  AND2 AND2_22(.VSS(VSS),.VDD(VDD),.Y(I27),.A(B44B),.B(v10bar));
  AND2 AND2_23(.VSS(VSS),.VDD(VDD),.Y(I25),.A(v0bar),.B(B22B));
  AND2 AND2_24(.VSS(VSS),.VDD(VDD),.Y(I24),.A(B24B),.B(v1));
  AND2 AND2_25(.VSS(VSS),.VDD(VDD),.Y(I22),.A(v7bar),.B(B18B));
  AND2 AND2_26(.VSS(VSS),.VDD(VDD),.Y(I21),.A(B19B),.B(v12bar));
  AND3 AND3_34(.VSS(VSS),.VDD(VDD),.Y(I186),.A(B31B),.B(v0),.C(v1bar));
  AND3 AND3_35(.VSS(VSS),.VDD(VDD),.Y(Lv13_D_4),.A(v9bar),.B(v10bar),.C(I186));
  AND3 AND3_36(.VSS(VSS),.VDD(VDD),.Y(I18),.A(v0bar),.B(v10bar),.C(B41B));
  AND2 AND2_27(.VSS(VSS),.VDD(VDD),.Y(I17),.A(B45B),.B(v9bar));
  AND3 AND3_37(.VSS(VSS),.VDD(VDD),.Y(I192),.A(B37B),.B(v0),.C(v1bar));
  AND3 AND3_38(.VSS(VSS),.VDD(VDD),.Y(Lv13_D_6),.A(v9bar),.B(v10bar),.C(I192));
  AND3 AND3_39(.VSS(VSS),.VDD(VDD),.Y(I195),.A(B20B),.B(v0),.C(v1bar));
  AND3 AND3_40(.VSS(VSS),.VDD(VDD),.Y(Lv13_D_1),.A(v9bar),.B(v10bar),.C(I195));
//
  OR2 OR2_0(.VSS(VSS),.VDD(VDD),.Y(B41B),.A(I113),.B(I114));
  OR2 OR2_1(.VSS(VSS),.VDD(VDD),.Y(B42B),.A(I111),.B(v12bar));
  OR2 OR2_2(.VSS(VSS),.VDD(VDD),.Y(B43B),.A(I108),.B(I109));
  OR2 OR2_3(.VSS(VSS),.VDD(VDD),.Y(B29B),.A(I105),.B(I106));
  OR2 OR2_4(.VSS(VSS),.VDD(VDD),.Y(B18B),.A(I102),.B(I103));
  OR2 OR2_5(.VSS(VSS),.VDD(VDD),.Y(B17B),.A(v7),.B(I100));
  OR2 OR2_6(.VSS(VSS),.VDD(VDD),.Y(B40B),.A(II98),.B(v10bar));
  OR2 OR2_7(.VSS(VSS),.VDD(VDD),.Y(B26B),.A(v0bar),.B(I96));
  OR2 OR2_8(.VSS(VSS),.VDD(VDD),.Y(B27B),.A(I93),.B(I94));
  OR2 OR2_9(.VSS(VSS),.VDD(VDD),.Y(B23B),.A(I90),.B(I91));
  OR2 OR2_10(.VSS(VSS),.VDD(VDD),.Y(B21B),.A(v10bar),.B(I87));
  OR2 OR2_11(.VSS(VSS),.VDD(VDD),.Y(B32B),.A(I84),.B(I85));
  OR2 OR2_12(.VSS(VSS),.VDD(VDD),.Y(B34B),.A(v8bar),.B(v3));
  OR2 OR2_13(.VSS(VSS),.VDD(VDD),.Y(B14B),.A(v7bar),.B(v8bar));
  OR2 OR2_14(.VSS(VSS),.VDD(VDD),.Y(B35B),.A(v2),.B(v7));
  OR2 OR2_15(.VSS(VSS),.VDD(VDD),.Y(B25B),.A(v10bar),.B(I79));
  OR2 OR2_16(.VSS(VSS),.VDD(VDD),.Y(B39B),.A(I76),.B(I77));
  OR2 OR2_17(.VSS(VSS),.VDD(VDD),.Y(B38B),.A(I73),.B(I74));
  OR2 OR2_18(.VSS(VSS),.VDD(VDD),.Y(B30B),.A(I71),.B(v7));
  OR2 OR2_19(.VSS(VSS),.VDD(VDD),.Y(B16B),.A(B35Bbar),.B(I69));
  OR2 OR2_20(.VSS(VSS),.VDD(VDD),.Y(B36B),.A(II65),.B(I66));
  OR2 OR2_21(.VSS(VSS),.VDD(VDD),.Y(B24B),.A(I62),.B(I63));
  OR2 OR2_22(.VSS(VSS),.VDD(VDD),.Y(B44B),.A(I59),.B(I60));
  OR2 OR2_23(.VSS(VSS),.VDD(VDD),.Y(B33B),.A(I56),.B(I57));
  OR2 OR2_24(.VSS(VSS),.VDD(VDD),.Y(B28B),.A(I53),.B(I54));
  OR2 OR2_25(.VSS(VSS),.VDD(VDD),.Y(B22B),.A(I50),.B(I51));
  OR2 OR2_26(.VSS(VSS),.VDD(VDD),.Y(B15B),.A(I47),.B(I48));
  OR2 OR2_27(.VSS(VSS),.VDD(VDD),.Y(B31B),.A(I43),.B(I44));
  OR3 OR3_0(.VSS(VSS),.VDD(VDD),.Y(B19B),.A(I39),.B(I40),.C(I41));
  OR2 OR2_28(.VSS(VSS),.VDD(VDD),.Y(Lv13_D_3),.A(I35),.B(I36));
  OR2 OR2_29(.VSS(VSS),.VDD(VDD),.Y(B37B),.A(I30),.B(I31));
  OR2 OR2_30(.VSS(VSS),.VDD(VDD),.Y(B45B),.A(I27),.B(I28));
  OR2 OR2_31(.VSS(VSS),.VDD(VDD),.Y(Lv13_D_2),.A(I24),.B(I25));
  OR2 OR2_32(.VSS(VSS),.VDD(VDD),.Y(B20B),.A(I21),.B(I22));
  OR2 OR2_33(.VSS(VSS),.VDD(VDD),.Y(Lv13_D_11),.A(I17),.B(I18));
//

endmodule