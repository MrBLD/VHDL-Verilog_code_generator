module s3841(g3233,g16355,g5695,g16437,g3218,g8263,g4590,g8268,g6225,g8262,g6712,g7425,g5637,g24734,g3993,g7961,g6979,VDD,g3213,g16297,g8175,g3219,g8082,g5648,g7052,g26135,g7357,g6677,g6442,g8270,g7084,g7229,g6750,g6944,g3221,g7334,g26149,g5549,g3224,g3230,g7264,g8030,g27380,g3212,g51,g4450,g3217,g8012,g4088,g5437,g3222,g3234,g16496,g8007,g8258,g7956,g8251,g4321,g8265,g8023,g8106,g5472,g4200,g8087,g25489,g8167,g5595,g7014,g6895,g8274,g6447,g25420,g6313,g8275,g3226,g25442,g8096,g3223,g7302,g3228,g3227,g8261,g3225,g26104,g6642,g8259,g8272,g6368,g3220,g563,g3216,g5738,g7194,g5555,g6782,g1249,g5612,g5511,g16399,g6573,g3214,g7161,g5686,g8267,g8266,g8273,g8271,g5747,g1943,g5629,g7909,g3215,g3232,g5796,g4323,g6518,g7487,g8264,g4090,g8269,g6231,g3231,g6837,g7390,g3229,g7519,VSS,g6485,g8249,g8021,CLOCK,g5657,g6911,g25435,g8260,g2637,g5388);
input g3233,g3221,g1249,g3224,g3214,g3230,g3218,g3212,g51,g1943,g3217,g3215,g3226,g3232,g3223,g3222,g3228,g3227,VDD,g3213,g3225,g3231,g3234,g3229,g3219,g3220,g563,VSS,g3216,CLOCK,g2637;
output g16355,g5695,g16437,g8263,g4590,g8268,g8262,g6712,g7425,g5637,g24734,g3993,g7961,g6979,g16297,g8175,g25435,g8082,g5648,g7052,g26135,g7357,g6677,g6442,g8270,g7084,g7229,g6750,g6944,g7334,g26149,g5549,g7264,g8030,g27380,g4450,g8012,g4088,g5437,g16496,g8007,g8258,g7956,g8251,g4321,g8265,g8023,g8106,g5472,g4200,g8087,g25489,g8167,g5595,g7014,g6895,g8274,g6447,g25420,g6313,g8275,g25442,g8096,g7302,g8261,g26104,g6642,g8259,g8272,g6368,g5738,g7194,g5555,g6782,g5612,g5511,g16399,g6573,g7161,g5686,g8267,g8266,g8273,g8271,g5747,g5629,g7909,g5796,g4323,g6518,g7487,g8264,g4090,g8269,g6231,g6837,g7390,g7519,g6485,g8249,g8021,g5657,g6911,g6225,g5388,g8260;

  wire I39779,g383,g10200,g26388,I29694,I32368,g7535,I30704,g2896,g27306,I39273,g9113,g19174,g12950,g3462,g7153,g10461,g28343,g8464,g30003,I39460,g8812,g27416,I35476,g22176,g24112,g8408,I23258,g4746,I24061,g26591,g4313,g7593,g24843,g26458,I37035,g28295,g19479,g16164,I29291,g22519,I32616,g712,g4392,I37062,g2652,g21187,g30773,I40245,I39782,g18325,I19727,g15432,I39976,g29865,g22421,g10390,I31171,g30921,g10449,g17167,I30197,g14143,g16394,g5550,g26465,g26784,g22078,g11379,g11581,I18813,g29792,g24851,I23709,g14753,g3931,I40967,g5121,I35744,I13478,g21135,g20934,g20392,g8792,g7632,g21487,g30102,g21381,g27797,g25279,g25087,g27720,g14954,g11246,g21988,I23845,I33437,g17503,I26491,g25148,g26585,I34812,g9958,g23984,g19677,g18969,g10324,g28849,g30808,g26978,g8076,g19701,g24802,g13369,g30092,g20417,g26713,g27003,g28474,I27149,I35518,I23766,g30457,g16489,g18826,g20269,I36588,g27371,g14537,g21765,g28374,I21361,g29155,g1960,g20289,g1576,I24340,I31730,g13266,g10044,I36272,g23505,g25405,g13486,g15461,g270,I17681,g12325,I39913,I38330,g1131,g151,g8851,g30097,g1761,g12989,I28038,g27718,g29008,g24469,g23415,g23129,I32686,g23408,g13194,g25647,g24748,g24571,I30116,g29736,g29270,g17189,g21990,g17129,g16392,g1172,g29512,g10300,I17933,g13221,g11389,g11789,g26984,I18205,g15707,g16162,g23100,I34150,g5878,I35437,g8528,g1037,I20791,I38437,g17947,I35715,I40113,g21823,I37296,g17667,g26999,g666,g20647,g8832,g21163,g11588,g13156,g20298,g10709,g28340,I14009,g7337,g27528,g27045,g12064,I33825,g16629,g27950,g29398,I40715,g27197,g25119,g13400,g13127,g23643,I40600,g5999,g1515,I29547,g20182,g2330,g10545,g10081,g14244,g23905,g29344,I17913,g10199,g9747,g26268,I25198,g12142,g5412,g17419,g23291,g28158,I40862,g19194,I35500,I37125,g29857,I36942,g30887,g9752,I33703,g27322,g5753,g18223,I24318,g7848,g3098,g15774,g18842,g22154,g28350,g25180,g29150,g21226,g8239,g4360,I18551,g17145,g23190,g3805,g27149,g28369,g11781,I15466,g5598,g24347,I40170,I38401,g2650,g2981,g26851,I37851,I16939,g11743,g29310,g18170,I38743,I30020,g10679,g29982,g15671,g11917,g28493,g30986,g24098,g19768,I30263,g29077,g25322,I27032,I40021,g26708,g6890,g5972,g2802,g24406,g24916,g2814,g4517,I24916,I37128,I36885,g28163,g24353,I20598,g10571,I26676,g23857,g379,g13963,I18827,I21083,g17183,g7754,g14132,g25209,g18972,g19038,g13218,g28482,g21189,g21800,I33371,g12651,I36915,g18881,I21566,g23478,g1276,g19168,g23458,g17445,g12513,I22626,g21202,g21695,I15651,g12523,g11840,g28321,g9892,g20556,g26900,g12259,g29793,g26979,I17998,I15222,g27939,g182,g8276,g28017,I18280,g26548,I40904,g14233,g12113,g30864,g19480,I38746,g5413,I14957,g1928,g4363,g8013,I20709,g21792,g19852,g1390,g24166,g22157,I38647,g1240,I25089,g24058,g28306,I37311,I40487,g15483,g16551,g28228,I16641,I27107,g25618,g6030,g29641,g21162,g21779,g4721,g4800,I29516,I25189,g19578,I30317,g26960,g18090,g18883,g25189,g30008,g17429,g2857,g18735,I30026,g7964,g10482,g19933,g10086,g17531,g19150,I13742,I24913,I32568,I24538,g22671,I16015,I28767,g19714,g30594,g24834,g22241,I29513,g21039,g21845,g13933,I40558,g26670,g13613,g16764,g10416,g25553,g30644,g25968,g4156,g12159,g15561,I34668,g28113,g7915,g23079,g19104,g403,g22306,g22233,g13336,I33448,g21071,g29615,g8515,g6177,g25352,I31751,g17171,g30227,g26481,g28552,g29572,g29740,g25145,g13853,g15244,g9126,g22936,g27334,g10323,I20444,I26311,g4492,g20587,g1214,g5148,I35673,g7779,g11735,g22038,I40122,g16301,g23938,I35083,g15994,I33358,g14039,g2707,g24237,g27630,g28643,g12654,g4272,I13122,g30894,g6027,g28734,g30731,g20294,g17927,g22195,g14985,I29177,g23543,g30056,g14071,g15268,I38245,g13024,I18013,g29955,g13353,I31769,g30735,g29184,I23103,g13366,g14000,g26840,g28168,I31826,g25588,g16382,g10337,g28048,g27390,g724,g17162,g29519,g13251,g27435,g27562,g5981,I22694,g19847,g30609,I18563,g17752,g24637,g10366,I32391,g5900,I21267,g16047,g5856,I14056,I31165,g22278,g22805,g2864,g12913,g1665,g22122,g12971,g21182,g28267,g29958,g1315,g21076,I23082,I32178,g26489,g29195,I25150,I20685,g28718,g2854,g21243,g25356,g20522,I38668,I34755,g30810,g26014,g12068,g7896,g23982,I38898,g8808,g25401,g29486,g25953,I36981,g30730,I14475,I32286,g28648,g24572,g12118,g17234,g3085,g2208,g5088,g13027,g5642,g22236,g7700,g23900,g21895,I24709,g11771,I17907,I37771,g16829,g16018,g26565,g11358,g24547,g27328,g113,g17159,I37056,g25530,g823,g12204,g20410,g12388,g1645,I27405,g26665,g20057,g23797,g21508,g478,g27308,g28126,g19982,g26398,g17460,g1553,g149,g10883,g6056,I37170,I20376,I41011,g16070,g21773,g16054,I29083,g21027,g17093,g6572,g2246,g13846,g25628,g28711,I34722,g24115,I40140,g7259,g10269,g28624,g10235,g30833,g11,g30865,g25627,g29045,g3963,g6418,g28353,g1399,g16298,g24657,I32617,g26440,g26733,I31589,I29004,g4346,I39764,g21139,g30361,g3937,g8852,g21072,g24833,I23314,I29288,g17193,g13546,g19054,g19664,g451,g152,g26638,g20597,g1868,I15671,g15235,I22842,g23789,g24900,g28703,g18858,g30251,I21952,I40787,g25933,g17969,g29893,I31035,I21149,g21550,g15424,g15845,I34830,g5009,g11014,g21886,I37068,g21066,g16853,g15877,g12790,g23633,g204,g11032,g24285,g12273,g10972,I29669,g10569,g12904,g11468,g9286,g27372,I15909,g5278,I31451,g16057,g23066,g14336,g8510,g4292,g14221,g14214,g14863,I22828,g22173,g14975,I22503,g23198,g28293,g30276,g30510,g28007,g13378,g24952,I13849,I37191,g5996,g10940,I26123,g30437,I37269,g27577,g7730,I13601,g17618,g435,g25387,g22864,I16006,I29981,g28444,g5246,g28443,I40515,g18933,I36099,g19353,g25033,g15596,g10011,g12833,g5888,I36311,g16400,g15857,g9228,g25376,I26320,g24088,g24224,g7573,g19257,g20569,I23760,I34306,I21939,g19241,I25750,g19903,I16372,g24131,I34674,g7845,I37173,g4626,g21995,g10591,I23830,g28414,g24413,I31580,I24454,g5929,g19857,g13364,g10127,g19656,I20625,g21791,I21508,I36224,g15801,g9143,g13242,I35992,I38801,I40475,I26413,g30664,g17674,g844,I36075,g15829,g25295,I25940,g23210,g28053,g24464,g28967,g30339,g23386,g14322,I22515,g29031,g23571,g24560,g11459,g27044,I27062,g11414,I37029,g5990,I18536,g30667,g21092,g29716,I34698,g15652,I29101,g30315,g16239,g23263,g1393,g13941,g22108,I36072,g24303,g25340,g11633,g16626,g18115,g13737,g22596,g8089,g28847,I28813,g4552,I21609,g26393,g22581,g20553,I14532,g11650,g19652,g19884,g10694,g246,g24752,g12324,g22695,g21361,g17333,g18830,g10797,g851,g21398,I32567,I21286,g29627,g26634,I35407,g27336,g8552,g29954,I21638,I34063,g23300,g18854,g9038,I30908,g5610,g26283,I37086,I21404,g16058,g7712,g5814,g19858,I15317,g5800,g14768,g18526,I17771,I39794,g24563,g19705,g22128,I18743,g23467,g11234,g18648,g25105,g27167,I39895,g23483,g9101,g11055,I31286,g5775,g21003,g1958,I26843,g2920,g23544,I31124,g17092,g26447,g12882,g4515,g30899,I30002,I19753,g17301,g5587,g11991,g27063,I16231,I18758,g19382,g23639,g20279,I16270,g10126,g13070,g11249,g18996,g30518,I20622,I20009,g23950,I26972,g20595,g16250,g20386,I31745,g13245,g24758,g30755,g14554,I25138,g4228,g26587,g2267,g30088,I24601,g19333,g21143,I31562,g15655,I14654,I21449,g16430,g24774,g11411,I25132,I18539,g29297,g3207,g4441,g7466,I18560,g18971,I21755,g19689,g22497,g29278,g5813,g28150,g5951,g16163,g1550,g14936,g18478,g20247,g26814,g29445,g30772,g1779,g2997,g15841,g26230,g15196,I22044,g29218,g28339,g4048,g586,I37593,I31805,I36769,g839,g19554,g15265,g8492,I14900,g4865,I31181,I16128,g25337,g12248,g23730,g5401,g731,I20799,g10196,g8253,g16142,g15843,g27329,g28359,g25066,g23802,g10206,g16134,g7615,g26401,g30030,g13224,I40071,I31637,g21410,g2685,g19859,g29164,g25364,g30719,g30807,I24037,g21358,g23204,g27215,g27254,I29351,g30749,g1279,g16515,I34809,g13097,I25294,I40676,I40603,g28285,g9424,g21122,g12688,I30119,g24925,g10728,g20585,g24047,g30673,I37787,I21548,I36420,I23105,I33463,g23531,g4854,g30822,g13241,I32461,I40605,g20356,g11727,g10858,g27464,g1070,I20553,g21091,I31763,I41105,g19093,I18801,g12960,I20264,I35419,g13189,g30203,g12027,g23076,g28494,g8488,g5406,g12151,I40313,g21086,g1066,g13361,g15878,g14467,g26282,g18166,g20926,I24669,I25064,g26594,g19105,g26809,g29400,I25867,g1776,g24439,g28086,I23161,I24194,g16477,I20451,g20043,g20109,g11613,I32409,I36900,g1253,I17872,g20465,g29527,g14301,g18237,g30263,g29273,g8882,g19780,I20673,g5953,g10711,g9102,g8483,I28742,I36476,I32949,g2462,g10272,g25383,g23638,g13991,g17383,g13173,g11499,I23218,g11471,g24345,g16136,I30917,g26637,g5758,I26440,g7522,I37897,g28722,g27951,I16261,g29521,g11327,I20691,I22718,g19308,I40209,g2647,g26931,g21894,g276,g26890,g9633,g23462,g27627,g5773,g14222,g13345,g13176,I14006,g24101,g6221,g6119,g27472,g21137,I18198,g8545,g28755,g15838,g7085,I16465,g5817,g24252,I25495,g13881,g29782,g6887,g1128,g2200,g7265,I35731,g10693,g28484,g29406,g2924,I23908,g25681,I19608,g30080,g21623,I18317,I14865,g16988,g8557,g27900,g19180,g22144,g24215,I16363,I39815,g4456,g18992,g18179,g28700,g8977,I32991,g23193,g22009,g2658,g29213,g2383,g9293,I23056,g24308,g6215,I18411,g13126,g1177,I23430,g26989,g11860,I19750,g16967,g24453,I19526,g1091,I32670,g23330,I39077,I37143,g29725,g14431,g6209,g19752,g444,I35923,I24634,I16289,g22792,I35698,g17842,I22983,g27776,g11638,g12429,g5627,g2113,g11986,I35059,g30563,g20752,g29330,g29484,g18995,g30906,g6212,g9723,g21198,g19022,I34369,g26578,g16110,g2104,I30401,g30778,g22827,g15519,g17181,g16356,g28149,g4052,I26426,g11822,I30754,I38178,g1145,g9212,g29943,g22409,I30260,I39068,I40490,g27409,g4609,g1001,I39136,g11809,g23472,I38752,g5210,g11929,g8576,I18695,I21995,g25272,g18990,I23028,g4870,I29307,g13797,g15782,g9427,I17780,g16602,I29252,g13491,I17140,I17822,I21337,g19159,g11054,g25496,I32647,I32334,g20423,g11709,g30269,g25973,I20743,I35723,g28417,g21359,g19484,I13538,g9501,I27197,g22454,g23097,g28650,g16845,g24174,g12866,g20149,g8424,g13289,g6015,g22203,g19924,I18139,I16283,g15127,g19742,I33246,g1254,I37623,g30700,g26844,g26157,g28379,I25334,I39475,g6193,g20952,g10968,g18245,g29083,g28111,I18389,g29206,I24765,I39945,g28258,I38483,g5190,I16457,I19869,g23847,I14816,g25637,g30026,I27565,I40326,g12080,g13623,g21817,g27065,g30007,g30834,g30732,g18566,g5342,g13518,g1585,g13528,g5636,I18773,g26566,I38924,g10525,I22919,g15852,g2553,g1243,I29881,g11788,g27861,g10255,g12218,g24160,I32490,I32478,g24430,g5703,g22759,I38491,g20193,g10963,I14769,g5864,I27361,g4324,I18734,g10664,g4936,g1211,g12559,g19400,g8473,I32140,g10889,I24236,g2519,I30636,g9623,I33532,g13223,I27917,I15863,g13406,g12451,g23851,g22518,g22991,g7592,g16539,g20554,g4775,g10085,g29808,g24146,g7830,I39121,g10120,g30110,g15324,g29731,I15866,I28273,g978,g27098,g26571,g18900,g30532,g20582,I34535,g25271,I36473,g30512,g21432,g19697,g26876,g28241,g13424,I25971,g26245,g12752,g24506,g26795,I34313,g23870,g4476,g17324,g20739,g24909,I30137,g29109,g20568,g1038,g30379,I40811,g15527,g29640,g16644,g20925,I36483,I24387,g12544,g3179,g216,g12564,g21884,g6781,I29936,I37712,I37065,g11990,g24417,g10805,g17139,g25214,I39892,g25552,I16315,I34080,I29817,g4032,g15760,g22058,g5767,g19531,I32393,I24338,I29203,I40651,g19282,I23019,I34845,g30,g26167,g17269,g29405,g12921,g5971,g16466,g13936,g9755,g19568,g20950,I30601,g3925,g24459,g16445,g23119,g27892,g23246,g25130,I40498,I37080,g3204,g18639,I18253,g17634,g3142,g26672,g22741,g8295,I22581,g30516,g13435,I28521,I18365,g395,I14195,I25386,I37757,g29777,g17850,g23045,I37026,I28181,g6019,I15580,g13550,g18911,g10530,g25880,g17230,g10270,g28706,g2793,I23095,I39539,I33600,I14424,I16134,I23895,g5221,I20382,g5997,g26035,g13131,g19145,g15030,g8230,g23292,g30770,g21124,g25410,g13274,g21292,g894,g11642,I15853,g9401,g13255,I19648,I15484,g25620,g28829,g2239,g27628,g11957,g27307,g8575,g346,g13161,I39853,I35425,g30298,I29566,g2753,I17294,I24992,g29174,g29148,I22759,g3984,I27077,g19694,g10891,g12246,I32098,g19708,g4179,g24795,g28254,g15556,g28018,g21051,g17393,g30672,I16569,g24817,I18614,g28993,g15104,g20690,g22758,g27501,g22253,g838,g25444,g13341,g28177,g22708,g19882,g12943,g2209,g8427,g6067,g12435,I24339,g28096,I33843,g8872,g13755,g11905,g16514,g1839,g30368,g22643,g12186,g29241,I19932,I39348,g23936,g15734,g25221,g21812,g29813,g6117,g15260,g22777,g1372,g12466,I15794,g15813,g17966,g11765,g23592,g8587,I40934,g22428,g15033,I33723,g15171,g27896,g20447,g13011,g19726,g5947,g1695,I37617,g24878,g5777,I36585,I37814,g18441,g16633,g26777,I19898,I30029,I38831,I16785,g14106,g26343,g20555,g10118,g21382,I29591,I40215,I13128,g4575,I21647,I15532,g4038,g13229,I28080,g13511,g18555,g28449,g22865,g24099,I34797,I18256,g13864,I16897,g10165,g10793,g11958,g12478,g24962,g15418,g28676,g21103,g4724,I29462,g30270,I24539,g21615,g8681,g13330,g13983,g18070,g12373,g25011,g21956,g13000,g26873,g23393,g17186,g11972,g23244,g24478,g331,I28825,g28512,g25672,g25166,g17468,g6156,I19924,g30325,I25344,g26214,g10472,g22803,I39840,g30618,g19222,g7157,I23639,g20550,g198,g28022,I33861,g5821,g29382,g19710,g10520,g3101,g15443,g12907,g29704,g16895,g29985,g25259,g21395,g5914,g24051,I32883,g18204,g23118,g21890,g25436,I40766,I15433,g12376,I40886,g28763,g12219,g16458,g16999,I15803,I32468,g19201,g21098,I18473,I26993,I25032,I28994,g8144,g23008,g4962,g30259,g514,I38142,g25020,g25862,g18583,g30072,I18100,I17831,I33460,I24452,g11830,g2066,g30167,g27997,g12481,g29758,I35824,g25213,g15933,g20708,I38936,I40883,g29468,g27008,g7391,g17510,I18590,g19883,g2324,g21196,I30536,I21979,g23671,g16212,g4351,g30781,g15853,g24309,g5704,g10303,g21476,I37494,g611,I25201,g9909,g23280,I14920,I34686,g5397,g13115,g4833,g30357,g21925,g4964,g17058,g27347,I30269,g25907,g23724,g15747,I30326,g5919,g27171,g2984,g12786,g1663,I39423,I15574,g16061,I29317,g29949,g30836,g29197,I15454,g15659,g28167,g11951,g16140,g22296,I37047,g25283,g13401,g22221,g13625,g17523,g29456,g29564,g26439,g148,g13343,I16942,g11690,g17654,g25028,I18611,g22627,g30071,g8820,g10895,g29418,g1636,g20371,g12601,g8983,I29180,g24414,g28005,g9132,I24028,g20380,g20268,g8161,g29978,g17868,I23878,g21407,g8718,I24372,g11740,g30499,g10052,g10161,I30170,I38686,g28460,g9613,g24951,I36093,g13791,g12853,g13164,g12086,g10321,g19756,I27667,g22995,g30311,I18061,I30380,g21809,I22705,g30708,g13485,g16865,I24560,g29964,g28382,g15803,g21694,g29403,g16111,g7972,g7528,g29966,g26993,g30888,g12330,g24338,g25343,g29971,g18986,g27285,g4006,g20315,g4806,g21123,g10842,g17425,g5824,g17624,I40733,g23305,g16676,I26726,g19304,g25183,g12699,I23926,g11160,g5053,g10462,g26896,g18419,g28260,g29821,g11151,g27038,g12275,g30274,g26968,g21390,g11970,g17616,g29264,g27919,g17065,I27549,I18341,g30889,I40197,g8434,I20535,g27689,g26471,I22936,g24447,g30897,g30387,g6200,I30215,g9524,I23943,g26944,g10906,g22387,g885,g10251,g21320,g19227,g1705,g404,g27913,g20999,I36132,g21846,g24239,I16587,g14015,I34990,g19899,g23610,I14605,g19671,g13612,g30744,g11518,g26842,g29364,g25193,g27658,I17715,g26215,I36936,I13119,g24855,g28731,g22107,g28165,I36153,g27228,g11987,g29820,g24293,g28638,I18151,I26868,g19560,g25873,I24093,g29990,g15832,g11157,g9416,g24092,g30968,g28397,I20441,g23887,g6180,g25952,g24495,g28327,g5204,I31592,g20491,g8138,I38764,g7607,g16743,g5071,g25039,g11932,I28189,g11462,I24732,g11208,I24565,I31835,g8704,g19806,I24554,g14286,I29194,I38042,g10184,g29561,g24423,I39240,g9248,g7520,I27577,I18943,I27005,I28443,g26820,g24901,g22589,I35893,I16312,I21825,g29796,g18983,g17682,g25009,g27222,g18502,g15685,I19466,I26028,g20438,I28962,g30788,g518,g26957,g17023,I28494,g26589,g20763,g1594,g20147,g9725,g10454,g30226,I15613,I16608,I16566,g23916,g29932,g26427,g23562,g17275,g5207,I30741,g28768,g22811,g17673,g23769,I32323,I21677,I27122,g27680,g17212,g19078,I34659,g26314,g20718,I35087,I29472,g3069,g17384,g21252,g21362,g26010,g28842,I24481,g3710,g21276,g16276,g24648,g5963,I32874,I22584,g15871,g23546,g177,I15511,g25018,I21796,g29422,g13902,g13293,g30363,g13519,g17556,g4760,I39631,g7335,g1564,g5064,g9730,I22545,g23766,g19303,g12448,g29570,g9808,I39843,I37277,g26278,I18820,g29606,I36744,g11981,g11921,g24527,g23538,g11088,g29284,g7652,g22045,I37158,g23979,g13558,g26545,I39674,g19044,g18224,I15205,g13197,g380,g20697,g19183,g20913,g19146,g18630,g12995,I27253,g1985,g30776,g20722,g24313,g19541,g10328,g30090,g1462,I32895,I24611,g27783,g10653,g30060,I15815,g16682,g8751,g16100,g22403,I33737,g22037,I30104,g26520,g28799,g13774,I27516,g23561,g12533,g19632,g24873,g12538,g27587,g13482,I39349,g9170,I23433,g2156,g19504,g2623,g1956,g25958,g19135,g25354,g23413,I36087,g19620,g20296,g372,g15436,g8722,I17730,I40952,g8899,g12607,g15207,g14016,g28794,g24168,g26636,g24311,g9890,g18217,I34210,g22714,g28910,g23485,g23175,g17924,g16159,g8100,g13513,g16457,g10528,I25001,I22563,g48,g7926,I36705,g28091,g28110,I30191,g23116,I36479,g20383,I31883,I15184,g535,I21933,g26734,g29030,g20381,I24727,I36761,g21254,I30552,g21964,g24302,I18025,g19028,g12191,g12331,g11815,g29980,g25533,I15847,I17483,g25986,g11456,g4829,g10257,g27508,g20601,g16483,I27293,g10387,g26455,g23970,I29345,g26408,I29375,g30841,g25844,I16965,I24717,g17679,I16104,I30810,g1750,g23547,g27107,g29117,g27454,g2760,I28781,I35153,g19454,g20365,I35485,g23908,g28492,g29335,g862,g1419,g20717,g3306,g23401,g17903,g4495,g22182,g29685,I34644,g9013,g2836,g10933,g21756,g29246,g1973,I28959,g28399,g28657,I40291,g26892,g28305,g28919,g2348,g14614,I28330,g15912,g6230,I15271,I27092,g9939,g19950,I32378,I35254,g26801,I35125,g19253,g20354,g20498,g15505,g23894,g28313,g26796,g22077,I33640,g27456,g818,g9902,I18467,g16230,g3201,g19297,g29151,g12535,g21155,g458,g23748,g5898,g27095,I19591,g20991,I15237,g30364,I40700,g10558,g25205,g13114,g18864,I36888,g9232,g17773,I37620,I38018,g12840,g23278,I36533,g27230,I18575,I24171,g20796,g8336,g1782,g10106,g25215,g18258,g30830,g6974,g4026,g21322,g20008,g21219,g2300,g4465,I33535,I26645,g28683,g8531,I30176,I28148,g20775,g3957,g27253,I36647,g10213,g13671,g8382,I26240,I14593,g20107,I30122,g22871,g25164,g20132,g7388,g13455,g17340,g1007,g15382,g12743,g8090,I21259,I17804,g17698,g18942,I14541,g20385,g19571,g21142,g10536,g25053,g5687,g19097,g2327,I25311,g26934,g24509,I28115,g10073,g24448,I36341,g9289,g10176,I26561,g29321,g4260,g11787,g9105,g26612,g19630,g11189,g17853,g2359,I30068,I36496,g27432,I13158,g11934,g27349,g3338,g23146,g5005,g12499,g25334,g15259,g3161,g25661,g26220,g3966,g20145,g267,g27113,g10307,g6901,I31766,I33507,g27235,g7975,g10121,I31784,g26126,g8518,I18106,g24310,g5774,g13082,g16384,I24327,I28206,g9356,g672,g25655,g10747,I14660,g1573,I17843,g21477,I19530,g30900,g12121,I13417,I29445,g22079,I40098,g13205,g16321,g24072,g572,I17042,g21776,g10311,g25257,I38059,g10875,g24403,g26371,g2103,g29424,g30985,g2655,I27318,g26618,I38869,g13257,g28408,g27073,g868,I18722,g16015,g27811,g28421,I18378,g27932,I30486,g9767,g16236,I38480,g24554,g28032,I25571,g21788,g3057,g20249,g15437,I27152,I18166,g23882,g26271,g26793,I28093,g23574,g9419,g23469,g5903,I35470,g28937,I17125,g7578,g24083,g9049,I35667,g30904,g23306,I16723,g22620,g13900,I38477,g5761,I16972,I28876,g3164,g12657,g17758,g23120,g28483,g30373,I27408,g30066,g15902,g3013,g19099,g26114,g30580,I30626,g30898,g22520,g2591,g3246,g28863,g24316,g10365,I39878,g10042,g29234,g24982,g12558,g30552,g2664,g12980,g16154,g19221,I29575,I38169,I32925,I40618,g9523,I23171,g24599,g25994,g23690,g1231,g2013,g19763,g27564,I40266,g26556,g30300,g6146,g13872,I22813,g29276,g2616,g22477,I33485,g25961,I35852,I37939,I18641,g180,g19838,g28344,g9527,g25411,g16841,g18955,I39359,g21599,g10625,I40227,g15411,g26875,I32422,g19618,g4541,g13065,g19782,g8179,g20404,g26595,I20634,I38278,I14688,I21511,g19187,g23892,g4412,g24516,g1757,g12315,g11891,g14352,I26545,g16968,g5918,g13687,g918,g28788,g9128,g18404,g19511,g18841,g28002,g2779,g25431,g19665,g24845,g17914,I39472,g16064,g9094,g23691,g11797,g4564,g30268,g29361,I40808,g13673,g19678,g1896,g30354,g23619,g2361,g2682,g16449,g20902,I36882,g7582,g13059,I14499,g7614,g23983,g7554,I16489,g17632,g9876,g12262,g11017,I29435,g30579,g30284,I30005,I35940,g8757,g13199,g8801,g11404,g10057,g24880,g19317,g9952,g6363,g22434,I28984,I14981,g13104,g26507,g24488,g24923,g7471,g24142,I40628,g19977,g9306,g15459,g11712,g1742,g18919,I16936,g17025,g13089,g29408,I40588,I23125,g13136,I23045,g28948,I29191,g24587,g30346,g308,g4089,g28162,g26574,g26727,g4818,g22699,I16624,I21523,g11521,I33611,I40736,g2733,g14765,g27448,I39532,g30301,I16793,g10009,I35714,g19323,g28194,g20937,g2082,g5693,I31445,g25939,g20291,g3087,g11839,g19911,g19230,g19919,g19901,g18961,g12914,g3972,g5596,g7604,g21082,g14028,g13099,I16930,g24084,g9063,I30868,g5822,I18067,g6017,g9150,g20994,g20628,g23424,g22515,g29546,g26140,g12030,I20959,g11767,g5763,g2222,g21106,g22559,I18282,g30040,I13215,g16591,g5035,g27147,g1136,g4652,g2987,I34156,I13931,g7629,g14966,g5945,g20816,I15873,g23017,g1648,g27201,I17705,g9161,g16198,g21951,g12708,I34316,g13585,g17247,I18799,g13839,g25599,I27038,g23050,g30257,I36111,I33421,g28037,g14165,g18878,I30155,g1395,I16056,g28580,I27209,I37632,g16085,I18548,g16179,g18611,g14691,g4020,g30345,g10494,g13269,g20063,g16252,g30400,g25200,g24728,g13122,I15448,I34916,g27516,g25605,g13160,g11536,I36636,g18331,g3077,g30641,g29110,I37946,I25645,g28491,g13837,g2355,I20050,I29125,g30265,g9641,I16286,g13454,g3941,g22133,g25483,I29046,I18362,g27153,g25291,g12424,g8567,g13895,g17701,g8256,g30256,g28026,g14337,g9041,g1930,g18982,g1222,I39361,g25188,g19522,I14037,g26269,g10221,g17836,g28056,I40294,I28953,I38817,g12408,I22572,I23493,g7736,g13246,g14551,I27002,g11478,g13397,g13399,g5606,I14641,I27537,g30694,I40179,I20514,I39347,g1955,I13098,I39331,I22783,g13098,I23498,g9047,g10010,g27120,g28424,g22744,g20593,g2788,I40534,g18047,g5861,g22213,g25983,g16183,g15441,I40155,g13564,g1029,g12112,g18483,g22506,g162,g23586,g22451,g2510,I25243,g26703,g26652,g10087,g25560,g20342,I14650,g15408,g25573,I33335,g23502,I21780,I31868,I23335,I38833,I34111,g10099,g29928,I35373,g5110,g16650,g30063,g6104,g29106,g18813,I27008,g30976,I33399,I29283,g19217,g1681,I36803,g22692,g23773,g27869,I37793,g16990,g3075,I18127,I36627,I24351,I31781,I26525,g29208,I18620,g142,g29976,g14565,g16583,g26316,g12868,g28749,g835,g10090,I32193,g9484,g29212,I38841,g26466,g20217,g826,g13848,g15787,I36301,g23247,g4532,g30570,g30111,I32539,I32469,g11435,g8769,g173,g23105,g10405,I41096,I19611,g22725,I18320,I32958,g10615,g17447,g18913,g577,g12867,I16357,g27507,g26099,g21781,g28278,g27847,I18494,g18275,g26798,I35079,I35527,g28708,g10937,I34579,I15696,g29805,g30002,g26233,g19475,I33289,I40456,g6289,g21850,g8008,g26043,g22353,g22801,g10962,g21665,g17076,g23184,g19032,g22618,g22295,g23187,g21178,g12212,g18874,g21722,g24928,g23359,g14630,g16558,I37982,g24304,g11209,g30574,g11835,I22640,g19811,g23831,g21610,g1312,g11802,g29236,I33479,I40760,g24595,g28813,I23104,g6281,g28791,g27897,g30085,g18147,g15647,I27215,I33918,I22855,g22194,g2633,g7518,I22667,g24539,I21537,I25692,g21302,g11256,g9953,g10289,g23202,g16092,I22702,I34026,I14984,I26420,g21982,g9776,g18247,g6035,I25772,I35076,g16423,g12546,I28360,g6672,g14176,g30914,g24433,g13445,g1257,g12022,g28207,g22047,g13211,g9199,g13359,g13465,g18587,g18424,g4651,g876,g15887,I32907,g5741,g317,g26426,g29573,g2084,g20326,g19263,g23551,I32175,g16619,g29229,g1161,g24103,I22737,g22338,g19573,g30691,I18716,g24493,g25207,g29096,I23192,g30466,g557,I27593,I29429,I29026,g29768,g22223,g13168,g4956,g25300,g22126,g21424,g2950,I33427,g23238,g305,g29161,g13670,g10231,g13398,g15759,g30568,g10155,I27014,g24949,g10999,g12066,g12886,g29257,g18036,g2778,I17798,g7228,g19214,g28747,g30115,g30134,I25099,g3068,g29781,g29649,g24763,I24306,g13204,g10510,I40697,g9806,g16091,I18350,I38635,g16067,g27446,g19275,g27192,g24097,I31874,g16460,g18886,I16462,g465,I25922,g22298,I32910,g9648,g13467,I36673,g15471,I13907,g16672,g20305,g27524,g28982,I15949,g13913,g26151,I14083,g8631,g22869,I34353,g30138,g15952,g5960,g20048,g2282,g21369,g22090,g21388,g21246,I34716,g12650,I16071,g23873,g22555,g10305,I36679,g27175,g16219,I23599,g19840,g11513,g12004,I15935,g10614,g30790,I24030,I32889,g20138,g771,g12968,g12473,g19254,g10295,g26797,g8711,g22718,g24013,g261,g26802,g626,I15308,g9480,g9534,I18142,I31607,I18305,g29654,I36156,g9894,g30472,g12536,I22679,g515,g21372,g8341,g7990,I27050,g19202,g18430,g16785,g20191,g9366,g10024,I38496,I16325,g21935,I23219,I24292,g733,I38028,g24591,g25289,g26002,I16450,I20132,g13601,I21252,I38193,g27181,I21531,g21557,g26521,g7389,g8665,g6052,I25826,I15523,g960,g13884,g27937,g2554,g23285,g20254,I38510,g18825,g8651,g1030,g30187,g30076,g27497,I18007,I23036,I31697,g18809,I24646,g15623,g5407,g18929,g29232,I25732,g4677,g8791,g30125,g12645,I35449,I34683,g27976,g26575,g25977,g314,I16482,g7766,I28119,g24238,g29520,g19984,g23615,g519,g3240,I14831,I18518,I29797,g23718,g11851,g888,g12339,g900,g27053,I37304,g22842,I38199,I18746,g11510,g27276,g27136,g21564,g28771,I14338,I24234,g24392,g17653,g16081,g17893,g20144,g18025,g26410,g11790,I30329,g16852,g3617,g26016,g5787,I24745,g16855,g16182,g20324,g13348,I24602,g17422,g10061,g17148,I18085,g20606,I14416,g27990,g21199,g29226,I25144,g26750,I21458,g12171,g1116,g18604,I31008,g15658,g11420,g12988,I18370,g19593,g24312,g18837,g29348,g29228,I35521,I23274,g24847,g15399,I18842,g17621,g8250,g25856,g23997,I17645,g2660,g25070,g28669,g11780,g7574,g17408,g19164,g23569,g25174,I19415,g9763,I20021,g29755,g25044,g19269,g23394,g11772,g12269,g4483,g2873,I34974,g13656,I33361,g19291,g15581,g26148,I27170,g19300,I32423,g10887,g24332,g19220,g8516,g22750,I24148,g17190,g16486,g3084,g21448,I14704,g4839,g26620,I38208,I36551,g29609,I24157,I31499,g23171,I30511,g8845,g27814,g9904,g15322,g22225,g18958,g8873,g14316,g8015,g21250,g30804,g9676,g21857,g8311,g7862,g30868,g9883,g17304,g22687,g17715,g30520,I16182,I37626,g23,g488,g28583,g13179,g28795,g8236,g14471,g20323,g13905,I32452,g27915,g19208,I14587,I29903,g789,g26897,g1965,I26898,g14490,g29918,I25921,I16499,g23860,g30479,g11902,g20461,g27963,g8921,g27018,I32424,g19207,g30982,g21172,g26596,g10871,g13226,I32634,g24890,g24517,g8538,g16389,g13870,g19698,I16215,I33304,g531,g1962,g11255,g30501,g29202,I24272,I32597,I19429,g30879,g26768,I35551,g5318,I17753,g22682,g13494,g13488,I37200,I35464,g27754,I18701,I16873,g17226,g23536,g23281,g21052,g10273,g21873,g30496,g530,g8168,g1219,g22693,g10692,I37842,g2776,g20700,g30789,g28954,I21841,g30514,g21711,g23114,g29356,g21816,g26616,g22222,g18906,I37973,I26639,g1934,g26246,g19515,g9584,g10004,g721,g10313,I13990,g22016,g22537,g30448,g26250,g30890,g5765,g28075,g17755,g30322,I15475,g11213,I36459,g25860,g23614,g23829,g27096,g27708,g15566,g15771,g27722,I30398,g24263,I34857,g30341,g29429,I29945,g21309,g27346,I35803,I38770,g30159,g28104,g16578,I35539,I15978,g22290,g27410,g20333,g8339,g15998,I33268,I16101,g9062,g4869,I16156,g18030,I21641,g5789,g19478,I33807,g23418,I21364,I32444,g23234,g21042,g26158,g9488,I23911,g2394,g12961,I36867,g28395,g13033,I23821,g19826,g7815,g4939,I19289,I30651,I32346,I15538,g5778,g39,g7015,I25141,g14298,g27923,g29009,g8329,g27109,g2321,g3235,g20376,g30676,I27900,g8658,g1171,g5759,g19693,g8484,g26085,g30680,g30699,g17967,I25562,I39821,I35099,g20588,I25740,g13047,g23444,g28187,g21167,g17802,I18369,g25064,I35497,g30171,I30221,g30796,g25099,g19384,g27355,g19029,g21544,g23688,g8912,g10641,I25653,g30826,I13140,g5402,g13632,g723,g23265,g27741,g15525,g7347,I31270,g10399,g19181,g15770,g5000,I36502,g27566,g3960,I37176,g29901,g8640,g432,g1525,I34695,I40712,g8381,g29963,g22669,I36237,g28060,g27089,I34444,g2363,g19000,g15410,g14328,I21514,I31742,g9183,I37824,g24161,g25974,g26829,I23981,g20328,g10652,g16141,g16987,I16335,g17390,g24393,g22740,I30654,I36264,I36612,I40173,g27246,g8563,g9438,g30726,g9928,g21748,g16840,g26947,g19411,I14238,g26782,g2428,g2371,g9203,g11890,I29603,g26551,g9774,I24308,I17765,g22191,I17878,g16050,I37356,g26724,g5098,g29360,I25423,g18597,I35146,I38659,I37602,g640,g15353,g30940,g29917,g20458,I21494,g16433,g25249,g8939,g5973,I16918,g17224,I33561,I37330,I25159,g28485,g20064,g24515,g19749,g9093,I15893,g14006,g30686,g24526,g19521,g4107,g9035,g29386,g23440,g29555,g24613,g28841,g12312,g20903,I14017,g18205,g21983,I18491,g23158,g19011,g21397,g12288,g14794,g24870,g19934,I33514,g20228,g7149,g19320,I13916,g29354,g2555,g20531,g16527,g10704,g3241,g26206,g20676,g28033,I23287,g26810,I32535,g1682,g16388,g15823,g18820,g26954,g8706,g12290,g22141,g1784,g7529,g10512,g28302,g21763,g28660,g18893,g30382,g30004,g19231,g30469,g27980,I16131,g24258,I38857,g24958,g28332,g28282,I28966,g19325,g19419,I25216,g26866,I33646,g23070,I29542,g22691,g4656,I32526,I19852,g17767,g21047,g29042,I35701,g9760,I19823,g13935,g15553,I40104,g13579,g12306,I30194,I21900,g17168,g5012,g1654,g21210,g8771,g22980,I23992,g26110,g21391,g21505,I17801,g20583,I25671,g11571,g25268,g28215,g2124,g28487,g1874,g25191,I20583,g16090,g19804,I37614,g24908,g26029,g30411,I29197,g28361,g28914,g10167,g969,g27247,I36358,g13030,g1890,g30901,g27211,g30280,I36454,g891,g13346,g13134,g27986,g19657,g26859,g3948,I31808,I40853,g22310,I18503,I20506,g9004,g8577,g24749,I24758,g27048,g2235,g29340,g13243,g24848,g735,g16943,g18085,g11539,g30537,g5934,g18805,g13906,g26390,g2479,g4275,g19141,g15780,g27025,g25429,g27988,I35515,g17117,g729,g21975,I27395,g24582,g12419,g1051,I28043,g25110,I38626,g30860,g25502,I21241,g17985,g1523,I34002,I14665,g23463,I33990,g12863,I23625,I17311,g14347,g5752,g13052,g30392,g13468,g25688,g28951,g19895,g8632,I32829,g2473,g10441,g14217,g26651,g10322,g8867,g9610,g5989,g23311,g21892,g1402,g17173,g13701,I23142,g4567,g12543,g24226,g8778,I25865,g22247,I38456,g19699,g3093,I26282,I21601,g23764,g26075,I37119,g28050,g22140,g29979,g585,I31250,I24016,g23893,g20904,g24619,I21482,I33717,I22952,g19258,g25514,I38421,g10663,g27493,I40772,g25184,g28996,g29259,I18157,g19904,g11144,g10471,g19252,g20347,g25388,I32150,g17019,g27055,g10804,g28732,g1706,g21093,I15556,I30359,g7715,g25310,I36258,I22823,g27241,I37167,g29948,I21742,g15248,g16222,g1669,g10986,g17482,g26740,g17176,g26718,g1536,g5875,g29509,I38466,I34254,g17398,g19577,g16438,g11522,I32588,g26004,g4912,g30969,I37044,I14675,g8084,g21868,g30470,I32575,I37474,g24861,g21385,I32347,g23152,g549,g24583,g26409,g23998,g5293,g28618,I16041,g22270,g11968,g5410,g21996,g21848,g11237,I33368,I15299,I28975,g26277,g18650,I18500,g21197,g10766,I16110,g4176,g30584,I26874,g13860,g18109,g27883,I28369,g26754,I31505,I31790,I33517,g2794,g12849,g15923,I14378,g19116,g10822,g16859,g21590,g12034,g16622,g18786,I16273,g15046,g23295,g1291,I30392,g24567,I41141,g27558,g28759,g6443,I32898,g13411,g19864,g3649,g28179,g30661,g22367,g19203,g30592,g23138,I29960,g29941,g313,g30698,g9647,g1453,g6085,g24259,I39080,I39625,g15540,I40670,I29969,g24496,I36315,I39324,I16303,g10519,g22841,I15571,g24940,g26319,g11132,I31031,g13611,g17555,g1600,I27739,g21449,g16237,g22062,I38629,g30199,g10646,g11748,g4094,g13414,g27693,g11527,I39788,I34800,g1830,I26182,g24746,g22082,g20901,g9125,g7971,g23103,g22736,g14171,I27173,g20881,g11607,g29248,g23169,g11225,g8562,g30949,g11950,g28840,g13190,g23216,g23681,g12772,g15293,g5396,g29924,g24305,g7623,I20062,g12412,g25467,g15402,I21688,g18645,g25488,g18225,g28319,I15899,g19548,g10527,g21874,g19791,g18938,g20308,g30338,g30721,g11936,g24054,I26508,I22618,g20086,g23909,g19491,g29097,I19321,g15757,g489,g8836,g28652,g15678,g23528,g18788,g30924,g29126,g14752,g27116,I25690,g29299,g15349,I32520,g13538,g5391,I22768,g24603,g24933,g10680,g11783,g18843,g9664,I18115,g26154,g21002,I14246,g12949,I36593,I25120,I31484,I19844,g27585,I37092,g14130,g24798,g11730,g20000,g27802,g15890,I24668,I29963,g24314,g14959,g19452,g16824,g7156,g2568,g25074,g13165,g8785,I16966,I31922,g20462,g27551,g20011,I31889,g20183,g22361,g16697,I30218,g13335,I24522,g22696,g17545,g5769,g797,g27146,g21938,g29811,g20682,g26573,I35452,g22798,g25834,I38064,g1813,g22881,g30593,g30895,I27281,I13959,g26165,g19256,g18466,I27041,g6040,I19618,g24867,g24941,g22866,g24889,I32668,g25022,g29427,g23794,g17878,g29355,g11662,I27131,I16085,g713,g1555,I19833,I23788,g8775,g23710,g29171,g15112,g24865,g11920,g13090,g10116,g30917,g3251,g3024,I15190,g26248,g17202,I23932,g5114,g30139,g28178,g2993,I28913,g26182,g26023,g3897,I34677,g24162,I26661,g29553,I30065,g23275,g4913,g29243,I29001,I34074,g10566,I18271,I41064,g19595,g17051,g22830,g10892,g12909,g29209,g28853,g11831,I39264,g1282,g17607,g12493,I29043,g22621,g28420,g29638,g22979,g13847,g23590,g11841,g29532,g2391,g5072,g17649,g19865,g23676,g4916,g26069,g27283,g20559,g27763,g30096,g13053,I24063,g29839,g30861,g20425,g10596,g26334,g30920,I25541,g13416,g24863,I30242,g27102,g30654,g18578,I25126,I36510,g8440,g9146,I30669,I15859,I34143,g20185,g29956,g4153,g30847,g18569,g27972,g18870,I18103,g19822,g21707,g20306,I39086,I33564,g22536,g30658,g8859,g10363,g10122,g6635,I19756,g26380,g5883,g17315,I27143,I13904,g20921,g10789,g12978,g28707,g2110,g8911,g10408,g15595,I23655,I37752,I14760,I31514,g23609,g23083,I30224,g8537,I35000,g18593,I37305,g23293,g23388,I36060,g19764,g27249,I38405,g18256,I18542,g22833,I21680,I21208,I35503,g1889,g8372,g30842,g5701,g22784,I18731,g26633,I21908,I25078,g13124,g17487,I30881,g27305,g13857,g30350,I30962,g29797,g19070,g7139,I23874,g20393,I39997,g15744,g21482,g22384,g26428,g8391,g479,g11059,g1168,g11079,g9082,g24134,I37800,g28029,g29154,I24576,g29744,I21443,I18302,I17054,g13437,g29319,I14516,I13134,g1763,I14449,g25256,g28152,g24064,g24815,I23608,g7626,g27387,g7936,g7721,g20189,g29935,I17904,I31077,g20113,g23242,g17262,I39017,I22631,I31141,g4573,g27437,g18991,g14442,g16040,g12117,g22229,I24006,g10783,I20909,g29318,g568,g30617,g5507,g30079,g22876,g2270,g25347,g5187,g15003,g2654,g13572,I32285,g2791,g26193,I36527,g28141,I17662,g15493,g6062,g17085,g11066,g24604,g29353,g23974,g18726,g970,g20975,g18803,g9016,g18892,g19110,I17059,I16024,I19808,g29309,g11897,g27462,g26280,g7852,I29174,g21153,g5668,g10218,g23176,g15724,g20786,g8579,g30536,g23409,g2489,I26348,g25725,g20401,g11560,I16578,g17791,g14774,g5736,g11395,g10690,I21354,g2096,g26830,g26351,g11550,I22945,g30885,I14243,g30460,g27563,g13869,g20106,I36499,g7796,g23414,g19608,g8551,g12216,I30857,g19284,g29026,g30447,I19455,g8176,g7655,g24412,g13677,I31496,g8328,g5696,g1810,g2291,I31290,g7345,g11091,g20641,I19452,g10529,I29715,g27367,g4581,g13706,g18949,g21736,g29163,g10943,g1083,g26001,I37978,g9144,I17149,I38698,I31085,g24179,g28945,g30850,g21527,g27910,I30725,g19228,g8947,g2766,g12565,g23778,g8958,g11825,g21102,g12881,g23052,g26808,g29373,I26682,g21069,I21292,I23010,I38214,g15379,g3054,g22063,I32577,g21730,g12169,g26199,I37968,g3036,g10119,I19513,g18880,g13739,g13427,g28077,g29951,I23698,I18405,g6060,g19148,g28916,g25190,g7842,I18145,g11407,g21227,g10331,g12440,g21156,g5041,g8944,g24869,I32345,g24860,g24177,g13539,g30024,g28227,I16581,g14115,I17863,g25685,I24133,I28726,I16870,g16004,g21455,I25633,g13516,I31673,I23839,g25990,g21440,g27766,g29146,g10043,g17461,g19328,g2223,g2151,g26073,g22114,I37113,g29987,I34997,g21973,g23192,g5547,I14574,g858,g25870,g19295,g17619,g28330,g28357,g11210,g23738,g5306,g16415,g533,g10523,g5015,I17658,g29085,I30113,I30911,I19794,g12228,g5252,g22179,g28479,g26136,g28098,g25197,g1924,I38701,g18504,I21923,g10459,g21949,I25811,g19416,g29372,g11763,g210,g23799,g25078,g5889,I30041,g28898,g11669,g22625,g19727,g6284,g27151,I35863,g29778,I25882,g11769,g22049,g27335,I40982,g24245,g10195,g13119,g1152,g22289,g24445,g23002,g13078,g5708,I27399,I30642,I29503,g22975,g8946,g5764,g301,g29800,g11548,g6081,I18626,g25262,g27221,g30033,g10443,I31387,g10481,g25698,g8705,g11836,g20428,g30329,g21379,I36668,I21497,g4079,g28877,I24531,g6227,I28190,g25991,g2211,g22130,g20297,g10294,I33488,g13503,g30334,g25278,g26344,I18359,g11782,g20633,g4598,g19619,g510,g25290,I34647,I31850,g19842,g16469,g2783,g19849,g23106,I21809,I15211,g24514,g17876,g20719,g4369,g26645,g11421,I23806,I28357,I23115,g1426,g21057,g936,g10212,I29525,g28950,g13106,g11520,I23954,I35506,g3110,g10548,I17627,g18023,g15258,g255,g23314,g19896,I33846,I35702,g24441,g30560,g28093,g21159,g11710,g23081,g12698,g28656,g27360,I36105,g10973,I40161,g1903,I23217,g9320,g22098,g2425,I28800,I19160,g9886,g13540,g13549,I19958,g20007,g1957,g2000,I17795,I15879,g9779,I16059,g11584,g25076,I13965,I13190,g18855,I35879,g13622,g29530,g164,g6369,g15343,g28331,g13367,g5676,g4787,g19716,I38728,I36250,g11801,I20631,g20891,I40107,I36848,g5193,g30669,g9644,g26000,I21761,g569,g20211,g25703,g22523,g20995,g22556,g1288,I38931,I17786,g26210,g30814,g23185,g11532,g1897,g28412,I34108,g12482,g11706,g25830,g17892,I30738,g23846,g15872,g17143,g29338,I40940,I29900,I17975,g30765,g30355,g23115,g17919,g18605,g21801,g21720,g1551,g13132,I18683,g11874,g15850,g16940,g14182,g8555,g28835,g15805,g8984,I40254,g18429,I27270,g11778,g12155,g29807,g22219,g22902,I26154,g28525,I30578,g20115,I30722,I23960,g5058,I34207,g16851,I29058,I33614,I38202,g1002,I23403,g2622,I38638,I18082,I14822,g30378,I36653,g15145,g2892,g26011,g29802,g11945,I22745,g17031,g11331,I37891,g19036,g18944,g11882,g12970,g11101,I36738,I20565,g12503,I25147,g8760,g2513,I16876,I24110,g18606,g23518,g15836,I32569,g23022,I20500,g8350,g30542,g22767,g847,I20679,g17661,I40658,I37053,I26796,g11966,g22549,g14910,g23729,g9124,g12534,I34162,g11262,g4332,g29502,g13431,g17100,g17675,g6444,g27265,g29082,g17271,g22101,g14060,g18446,I21998,g30896,I33364,g19783,I30011,I30167,g20875,g234,g26558,g30108,g12972,g25058,g480,g25346,g8823,g10250,I34165,g24874,g2810,g2608,g30610,g19551,g24508,I40629,g23078,g3900,I40667,g296,I13980,g9785,g29929,g12176,g9777,g1270,g27020,I14808,I23510,g3120,g18142,g25349,I41132,g27938,g20586,g6205,g4919,g13250,g18035,g28252,g13498,I35467,g26396,g12234,I30875,g23890,g12389,g22267,g17694,g23937,I25061,g22163,I32697,g15704,g18754,g27188,I19826,g23183,g18810,g29069,I40524,g11529,I22741,g22277,g24036,g11425,g14292,g565,g16495,I14489,g21009,g9588,g19156,g8448,g11871,g352,g27532,I23487,g22516,g19735,g28312,g4000,I18426,g10855,g21541,g19633,g19754,g2830,g26539,g27534,g23235,g12498,I37358,g17746,g8029,I19105,g29413,g9202,g13200,g29683,I31529,g16263,g20441,g26803,I29107,g30775,g20536,g4879,g3460,g21012,I34791,g30059,g2448,g19607,g28796,I29700,g30745,g27124,g20379,I28497,g9893,g17716,g26303,g23452,g25903,g2232,g7782,g28279,g17496,g30849,g11998,I33912,g16187,g12554,g21822,g24057,g5021,I28582,I25358,g605,g30605,g22739,g18074,g29741,g19787,g25124,g27023,g28016,g28324,g19240,I36162,I18392,I30131,g4379,I20652,g23822,g22847,g16019,g25052,g26615,g7658,I17433,g15173,g24778,g6032,g17288,g13526,g24260,g12990,g903,g20248,I18399,g15363,g27309,I37459,g28261,I34321,I37152,g28469,I39148,g21261,g23497,g21378,g16069,g17729,g17327,g24295,g1398,g16835,g26764,I23904,g22444,g19431,I39332,I24258,I31426,g2522,g26753,g20098,g30337,g11582,g23594,I30894,g8558,g30258,g22573,I18692,g29625,g27066,g7549,g29632,g7603,g24218,g12848,g26562,g583,g12441,g5338,g5551,g30883,g1134,g321,g5904,I31547,I14381,I30053,g30006,g8909,g22014,I35809,g2091,g20377,I26999,g7912,g16025,g22268,g25324,I33338,I28500,g2619,g25225,g20220,g22383,g5909,g25452,g21304,g28844,g11692,g20271,g20212,g26538,g17402,g18758,g4315,g10867,g22397,I31694,I23225,g25945,I24436,I29142,I36797,I17734,I29013,g18458,g23923,g26234,I34020,g22667,g21064,g25984,g19943,I18034,g29383,g13138,g22113,g15507,g132,g29961,g4734,I32587,g27373,I15185,g30753,I40919,g27661,g29363,g23849,g14830,g26505,g26425,g29423,g13375,I40754,g18218,I25432,g9075,g25106,g18319,g1090,g5887,g1915,I24555,g2436,g25421,g20227,g26407,I28609,g27019,g16909,g11592,g10423,g27106,I20550,g27032,I20390,I39881,g28729,g13789,g8305,I34851,g20694,g992,g26531,g8458,g23674,I25898,g27076,g21878,g27172,I23067,g30710,I24678,g20793,g7928,g25911,g28758,I40568,g22401,g2273,g11696,g2218,g3059,g836,g4343,g29010,I25426,I14553,g20607,I22901,g9519,g30840,g9569,g19545,g5807,g848,g19213,I13155,I36755,g13212,g1265,g19415,g15788,g29535,g13815,g22232,I30014,g2406,g27366,I25129,g26406,g16814,I40730,g11577,I30476,I33511,g20897,g22746,g22422,g23041,g18617,g29349,I32716,I15896,g27280,g24153,g2234,g20095,g5943,g27125,g25029,g2507,g4185,g30215,g26769,g18523,I28482,g5706,I35491,g28653,g9887,g29088,I24982,I22953,I27246,g17770,g21045,I32679,g19009,g16348,I29093,g29690,g28802,I33589,I17948,g5613,I32854,I24279,g26469,g28244,g725,g29999,g10500,I40164,g17048,g10172,I37131,I37662,I33352,g10659,g24456,I34879,I30062,g15784,I24156,g24178,I16166,I21282,I16850,I18353,I34400,I16244,g805,g22202,g10315,I21249,I16605,g21453,g20137,g2540,g23194,g19298,g24361,g28440,g30459,g20467,I25710,g6115,g11622,I17100,g1258,I15967,g16023,g22654,g2704,g24586,g19132,g14702,I27182,I33411,g30706,g13055,g26766,g9932,g23573,g22480,I26745,g13118,g27130,g4249,g27090,g11834,g26644,g27242,g29661,g18943,I38591,I20425,g23575,I32379,g16506,g18781,g18453,I36042,g27505,g19294,g21787,g852,g10946,I15354,g1082,g20372,g22162,g5243,g6051,g15228,g29132,g9355,g4366,g4752,g18679,g22677,g16411,g15996,I13161,g11541,I25510,g10056,g18852,g24330,I29522,g28415,g2233,g10918,g13209,g27561,I36864,g1435,g5785,g27612,g10296,g15725,g30305,g22886,I37357,I38641,g12057,I41065,I36554,g17560,g15339,g19124,g18522,I21793,g29100,I39573,g21229,g21376,I34114,g8568,g23525,g10826,g11681,g27058,g25972,g27725,I27119,I36468,g1900,g28434,g30321,g11873,I23076,g5427,g29621,g27809,g16293,I33624,g20892,g13840,g22917,g30476,I24544,g18932,g13619,g26482,g11525,g25479,g13510,I17709,g14478,g16093,g16560,g17330,I32922,I36966,g30314,g10559,I21819,I15605,g16105,I38536,g10865,g15880,g24102,g24606,I14731,g24236,g25314,I23442,g4091,g26555,g2252,I27235,g26605,g30967,g23037,g19868,g30919,g15065,g16825,g11705,I16711,g12162,I35003,g3197,g18490,g7973,I36371,I35953,I34327,g29227,I41044,g17259,g15870,I17692,g28641,I32518,g7594,g2093,g13384,I32430,I24437,g9507,g29516,g4753,g22015,g701,g11498,g26723,I20394,g23784,g29541,g30816,g8630,g8324,g22786,g17633,g23283,g28125,g19861,g21454,I35946,g22404,g25126,g17409,g25156,g10582,g21957,g10380,I33573,g8312,g19814,I29036,g24240,g28990,g11504,I25057,g22637,g29263,g29568,g28386,g26103,g18447,I26432,g28255,I28557,g23548,g2883,g29771,g2985,g8321,g776,g15453,I40039,g29279,g10362,g2463,I40531,g13409,g13934,g20534,g24396,I40892,I14615,g29446,g22418,g24556,g21063,I21790,g24771,g5654,g30748,I29280,g20910,g1945,g2809,I31799,I36444,g7739,g21133,I16703,g27298,I24132,I31532,g13116,g17314,g20896,g12939,g28664,g19815,g22873,I14945,g21882,g20157,g14414,g19335,I13433,I24633,I25030,g3188,g26018,I34863,g28625,g15178,g29336,I19432,I25742,g12597,g11912,I23833,g12267,I40634,g21174,I40300,g10103,g24405,g13305,g15210,g11906,I13604,g17862,g13535,g26726,g2938,g17951,I15843,g13389,g11686,I40682,g22080,g16854,g481,I23817,g17499,g28088,g23166,g8375,g13148,g24904,g1011,I17143,I35856,I40685,g21714,g11623,g28008,I40426,g11729,g12040,g5024,g17926,g24523,g20299,g11707,I38223,g8233,I29122,g22028,g26120,g12328,g18863,g20153,g29038,I29954,g20361,I16247,g25949,g28389,g17937,g29159,g2476,g17446,I23084,g5164,g1264,g4438,g16749,I26980,I24453,I23929,g5881,g10047,I24111,g1165,I20697,g18329,I18133,g1218,g21323,g10969,g25026,g16161,g25336,g20192,g22971,g25808,I38515,I39133,g30478,I33472,g2072,g21298,I20049,g7958,g22766,I18962,g27599,g30450,g28176,g25543,I24077,g20406,I39023,g2220,I33136,g11682,I19637,g22608,g12859,g15563,g8816,g25032,I25579,g30533,g27365,g19185,g26183,I22120,I20520,g29308,I26926,I35124,g29525,g24969,g19597,g28300,I24514,g12598,g23111,g22487,I15662,g21537,I32184,g16312,g5272,g16906,g7566,g27258,g4728,g20187,g1272,g25935,g27928,g8378,g29075,g27699,g18124,g24903,I33858,I30496,I35841,g30977,g15491,g17537,g14059,I24943,g11795,g361,g30054,I23436,g14541,g30348,g8507,g5952,I20640,g23331,I26624,g29233,g30881,I33900,g23874,g23372,g19532,I29638,I34752,g27105,g15651,I22881,g26592,I17106,g11988,g23470,g23637,g27767,g17165,g5030,g28635,g3998,I39083,g26915,I23958,g3994,g29455,g8053,g26186,g22180,g26973,g29529,g23006,g26009,g19142,I16984,g19587,g30707,I18114,I24227,g26238,g27304,g7053,g20799,I36873,g13141,g10400,g20634,g29701,g18921,g26646,I23209,g3616,g1913,g13644,g2877,g20513,g26600,g11737,I14547,I38217,g28490,I29294,I40856,I38811,g3239,g12223,g18901,I30404,g8987,g13177,I17689,g30105,I32198,I29484,g1809,g3028,I32645,g2471,g26364,g28105,g7465,g13444,g29180,g21875,I37647,g16484,I31658,g16543,I34803,g25175,g18644,g9391,g4017,g9872,g12415,I40871,I39375,g22272,g11312,g1217,g21795,I34827,g16008,g24038,g2879,I37101,g8147,I30748,g15859,g19084,g21794,I35542,g18486,g30647,I21905,I16814,g23419,I18344,g11745,g26705,g21393,g30360,g22238,g13818,g23049,g29774,I17203,g1777,g861,g26721,g10587,g24862,I37488,g18956,g22659,g29769,g25067,g30728,g29254,g1963,g11566,I16549,I38832,g30253,g13050,g27077,I36290,g10156,g29945,g27357,g14206,I31598,I23348,I16559,g19972,g29454,g29977,g8891,g22115,g27050,g24235,g11511,I21476,g15764,g30061,I15505,g20659,g19599,I25897,g4003,g29136,g16594,g17984,g5895,g29544,I31014,I36870,g8625,g9481,g29221,g16817,I29909,g28693,g20108,I37077,I40955,g24286,g12765,g8103,g29189,g26290,g14027,g14022,g13105,g1140,g8294,g26339,g23207,g8670,I33686,g27786,g3073,g16422,g19239,I28143,g17081,I22972,I13680,I23602,g25139,g1260,g5749,I14976,g22484,I36221,g23922,g13088,g30600,g20783,g12035,g9273,g2375,g8955,g3066,g22402,g29210,g26254,g11803,g19736,g24624,g30065,g28148,g5122,g24333,I27020,I18629,g2975,g9110,g16135,g22868,g710,I38820,g26962,g29022,I16835,g15738,g288,g27701,g17056,g24791,g2807,g22264,g25675,g16907,g26456,g29425,g9241,I16209,I27689,g25557,I23233,g19401,g207,g30335,g2441,g15346,g30534,I20848,g23861,I37514,g5309,g19687,g12119,g21667,g14044,I23374,g2797,I35017,g5034,I40158,g4112,g1300,I28712,g20083,g29554,I23034,I22797,g1870,g4507,g25288,I25681,g3252,I28178,g5872,g14290,g22730,g27702,g25539,g28524,g11656,g9786,g2399,g2524,g11300,I26085,g22312,g23473,g16463,g4064,g16292,g27291,g1306,g20525,g30463,g15170,g21553,g29534,I13977,g24600,I29675,g28320,g1203,I18929,g24694,I36615,g6043,g9127,I31481,g18101,g2366,g2858,I34456,g18183,g7556,g29143,g30023,g30911,g29305,g19839,g11806,g15731,g10271,g21818,g915,g29293,I30792,I27047,I37041,g22224,I30107,g15992,I16779,g23209,g12409,g6116,g10124,g10586,g11561,I15015,g23032,g17137,g20618,g6134,g20625,I38653,g18904,g21872,g11098,I38810,g12552,g23792,g29238,I40817,g17597,g172,g18981,I20688,g10813,g4168,g17896,g24533,I39466,g17182,g30739,I29993,g19061,g20915,I27832,g30973,g26404,g17098,g739,I27225,I28374,I17978,g19315,I22604,g30988,g21651,g26828,g23855,g15105,I13901,I16218,g13290,g15661,g25059,g18554,g27571,g10465,g17268,g7682,g19455,I24179,g10904,g21228,g26845,g2625,g20223,I33700,I24213,g1407,g30057,g22958,g10838,g18873,I20832,g23136,g25817,g28941,g20341,I33711,g1200,g13196,g18895,g27327,g19162,g30465,I18707,g4452,g27198,I20283,g13563,g23255,g20976,I38656,g19357,g19206,I22852,I32646,g12467,g1831,I29389,g21129,g27660,g11620,g4480,g8206,I33286,I20295,g13699,g318,g21611,g7667,g8044,g23745,g6707,g18572,g19628,g15307,g23850,I28896,I24475,g1916,g22843,I29556,I39062,g27054,g25602,g27522,g11824,g26878,I19634,g13079,g13256,I30959,I25938,g4783,I35530,g18346,g30483,g25847,g27311,g23243,g25505,g28679,g24825,I25856,g29528,g9591,g15612,g24907,g15789,g17528,I17960,g1384,I20278,g30575,g8446,I31036,g29080,g26067,g15257,I35106,I29933,g820,g5323,g17144,g2824,g22360,I33801,g1285,I18268,g23589,g30250,I23633,g11268,I18737,I31754,g19108,g28028,I40143,g26778,g26731,g4702,g10008,I30374,I31577,I40748,g16501,g20466,I18659,I33558,g10227,g14,I32548,g27383,g22118,g12217,I32498,g26580,g19131,g20162,g18957,g17282,g16718,g10495,g16467,g30852,g13029,g16290,g29795,g18585,I25857,g13004,g25203,g28309,g1912,g24306,I37638,I40110,g29062,g27480,g28114,g26451,I34132,g9819,I33009,g25724,g19940,g18270,g11852,g17233,I39863,g18060,g18998,g8908,I38740,g29249,g29247,g11347,g13525,g20090,I18455,I14925,g23486,g26953,g13228,I22845,g26054,g2787,g11749,g25569,g18619,g29307,g18261,I36227,I23463,I40868,g23067,I16931,I34980,I18656,g22774,g13036,I25654,g8965,I16472,I28341,g28807,g24534,g5087,I16196,g22269,g26302,I16656,g1155,g4629,g2789,g28094,g18013,g17724,I33232,g22060,g11185,g7906,g26332,g9245,g1921,I30786,I39899,g30010,g22256,g13323,g27734,g801,I31616,I28628,g21598,g10689,g20198,g29447,g17962,I35768,g26685,g8745,g16867,g1346,g8512,I30098,I24586,g12783,g24821,g2254,g15888,g29936,g12333,I34392,g8542,I30023,I35849,g14596,I37725,g20397,g13609,I24625,I20523,I26985,g13893,g29680,g8941,g1511,g3117,g1471,g9770,g26774,g8809,g25402,I26429,g20104,I40976,g11872,g17214,g9727,I24381,g30283,I41010,g23302,g5707,I19718,I17768,g28803,I14343,g16554,g28675,I29585,g24522,g19942,g27751,g18885,g11526,g28466,g21635,g13982,g24281,I36591,g25510,g686,I16954,g19880,g18649,g12265,g9660,g13149,g30031,g5757,g25127,g20485,g23907,g25506,g21157,g10650,g24367,g2398,g15664,g23939,g29452,I18710,g29129,I24278,g25170,g10538,g4329,g11821,g24541,I32356,I17238,g1297,g10886,I25168,I19820,g15808,g14626,g24956,g11126,g8868,g2703,I16147,g21804,g13871,g24082,g18718,I38074,I35762,g24210,I19208,g5908,g2078,g27748,g11994,g25519,g30331,g20133,g24568,g14885,g10049,g20703,g21782,g4659,g20753,g315,I27212,g6631,I28594,g30103,g11993,g13551,g20563,I34806,g1556,g19368,I18338,g16450,g14711,g16861,I37605,g5828,g24876,I40805,g20894,g11804,g7542,I36963,g20616,g3060,g11188,I23172,g27688,g29682,I25338,g18155,g30391,g16046,g4224,g12299,I14934,g28694,g29646,g2648,g5735,g24030,g26485,g10623,g16188,g23552,g30946,I40078,g27031,g351,g13061,g30094,g10825,g18221,g17617,g22099,g30567,g24480,g21001,g16487,g25036,g18370,g5866,g4479,g22074,g27831,g20280,g27110,g13536,I32085,g15396,g26264,g16002,I33621,g30625,g397,g158,g13460,I14778,I26134,g1869,I18787,g18062,g22612,g30293,I35473,g7776,g3521,g15593,I33643,g13451,g8602,g28092,g22935,I38875,g9479,I21377,g11916,g15579,g1909,I28479,g186,g5594,I29987,g5142,g27407,g23139,g29414,g29643,g23094,I30101,g24422,I33873,g30266,I36758,g15245,g19907,I33476,g30591,I36714,I25539,I33316,g10677,g5,g19113,g7224,g12154,g14736,I22730,I36897,g3091,g16712,g27608,I33834,g1746,g12042,g26581,I39828,g22882,g11878,g13674,g19081,g2387,I23667,g15494,g19653,g13303,I39991,g10075,g1137,g28372,g2947,g18131,g24220,g22380,g7868,I34737,g22207,g289,g11928,g24043,g8798,g24731,I30823,g21706,I26654,g11501,g8357,g485,g27970,g22939,g2086,g8578,g13457,g24521,I21479,g8762,g3170,g30908,g20099,g12519,g12756,I30813,g15737,g19774,I37775,g28366,g28191,I32660,g24381,I23763,g11567,g26275,g28702,I37312,g27467,g17735,I38613,g12966,g29517,I34140,g25980,g27985,g5998,g23565,I24226,g15031,I37822,g8910,g7861,g20492,g10585,g13129,g25120,I17300,g26012,g16126,g29483,g16380,I30407,g19935,I37273,g17252,g28495,I19657,g8964,g29691,I25105,g10493,I35297,I36253,g16651,g13073,g15403,g16137,g1703,g19600,g12974,I36781,g26423,I41090,g13851,g24380,g19316,g23429,I16514,g27502,g28308,g7138,g7338,I27338,g24457,g29993,I15568,g23853,g23494,g4898,g7949,g24458,g28328,g26790,g16181,g14894,g5656,g8761,g10388,g5710,g1730,g29658,g1547,g19414,g18450,g16088,g20250,g21594,g27343,I18178,g16391,g8937,g16476,g1979,g12134,g25202,g22563,g2395,g30336,g19747,I40272,g30674,g28063,g5835,I35399,g24035,g22091,g3043,g138,g2610,g13805,I29064,g19760,g24145,I38632,g13700,g28336,g30464,g10745,g20348,I23575,I25846,g20604,g8979,g11035,g16287,I35772,I29478,g30308,g608,g21183,g23618,g28667,g10016,g17610,g2285,g24248,I37089,I39139,I26365,g22797,g19031,I26996,g5230,g27271,g11102,g18297,g2609,g22245,g17658,I15925,g12811,g13130,g16199,g26744,I25018,I31565,g25038,I36951,g17813,g27514,g29435,I38447,g544,g15329,I40167,g8805,I23836,g23595,g19762,g5659,g468,I35172,g20286,I19997,g8968,g19614,g4208,I36957,g3494,g12195,g6638,I39776,g17936,g24107,g14412,g23513,g25629,g22073,I37965,g21696,g12382,I19938,g7557,I20816,g15429,I40946,g24331,g24350,g20336,g23241,g11644,g24630,g12891,g20040,g23891,g11736,g21688,I23075,g2501,g8504,g14577,g26175,g19818,g11829,g15855,I23942,g20346,g21566,I18767,g22104,g5640,g20340,I28447,g29637,g26614,g18189,g22998,g4250,g28045,g5901,g20435,g29669,I26777,I39056,I29942,g5954,I13943,g13915,g11173,I40781,g24151,g24337,g4584,g2369,g28061,g23644,I13239,I36362,g8254,I40230,g19296,g2180,I26407,I37014,g21497,g1997,I29966,I36144,I35994,g11370,g17132,I25406,g25395,g12294,g20378,g16107,I30245,I26237,g414,g26725,g21413,g2559,g16337,g17336,g28095,g12843,I30953,I17200,g11828,g5646,I32297,I16225,g30857,I27194,g27428,g21075,g15247,g27084,I18866,g9057,g22770,g29912,I31676,I27375,g18727,g11481,g21136,I25474,g17736,I13232,g17243,g5852,g2003,g15720,g29458,g25045,g5739,g1953,g12247,I30332,g8027,g1888,g16843,I23567,g21351,I22317,I35890,g23231,I35341,g23313,g4516,g4610,I14799,g30016,g27225,g15284,g708,g24841,I27402,g26461,g529,g23854,g25312,g7579,I25031,g17509,I25102,g19827,g12192,I15784,I29249,g27918,g11876,g24269,g27459,g18989,g24886,I13101,I36598,g30527,g11683,I27328,I33876,g28242,I37746,g28036,g26833,g19563,g30127,g178,g16379,g4868,I40083,g10910,I25666,g26353,I33633,g12890,g22088,g29345,g26756,g6167,g27709,g282,g13280,g21772,g17116,I28191,g26417,I33145,I32335,g8430,g21821,g11955,g11807,I22590,I14513,g12100,g23162,g10383,g26835,g27440,I18124,I25761,g14118,I32156,g6288,I20562,g8304,g9528,g30742,g15129,I19469,g7878,g19651,g20159,g27087,g13425,g29430,g20092,I16766,g13207,I38617,I21787,g16702,g5867,g27001,g28784,g19015,I32985,g24773,g22359,g30320,g17130,I38440,I28949,I24124,g23455,g23464,g14956,g15074,g22997,g26659,g28810,I39418,g8098,g23329,g13215,g30652,g21218,I37260,I37934,g27617,g7869,g4127,g13318,g10104,g10080,g16098,g21008,g29578,I33852,g5070,I14882,g30535,g20334,I33431,g27622,g16065,g19879,I21318,g2089,g12895,g7541,g30211,I24464,g28705,g324,g20019,g22916,g5793,g9794,I18530,g19501,g28486,g29613,g29668,g16570,I23712,g27576,g15321,g9764,g24902,g28085,g30695,g11540,g19075,g22490,I31053,I33390,I15922,g19715,I40002,g28159,g19953,I35509,I13956,g9425,g28690,I40468,g19209,g12935,g19921,g19725,I33831,g27400,g25019,g26174,g8635,I39392,g30319,I23412,g24446,g11953,g29252,I36404,g29495,g21259,g27251,g27166,g19251,g26800,g24479,g13421,g20578,g12006,g19030,I23879,g23492,g19330,I16179,g21245,g13169,g30564,I18058,g16733,I39454,I37008,g8601,g21716,I38843,g18789,g21194,I17070,g15930,I25231,g25319,g5825,I29572,g24754,g30588,g2303,I30938,I31748,g11493,g13568,g21749,g14230,g22578,g27793,I37942,g10258,g30511,g13291,I25303,I26590,g21740,g25233,g29401,g10557,g1661,g27742,g12789,g26701,I16009,g25458,g29190,g2469,g28673,g26382,g5846,g850,g2963,g28623,g26472,I28833,g28834,g17172,g23689,g23092,g573,g10649,I40637,g17042,I33586,g15475,g12003,g20837,I41099,g8626,g28084,g17779,g9100,g19846,g8004,g25121,I25624,I34764,g27338,g24379,I21942,I17813,g12748,I23338,g21674,g19544,g26066,I39411,g29696,I25315,g10260,g21626,g26051,I38196,g19649,g1563,g15176,I33219,I35043,I27011,g281,g4257,g26895,g26295,g21149,I16153,I18043,g13600,g10583,g16572,I13947,g25243,g7888,g24544,g18110,g28498,g24370,I38136,g29664,g24292,g23510,g22335,g8351,g17375,g6425,g21005,g21967,I27068,g9066,g5837,g2560,g25593,g28678,g21301,I27684,g297,g30655,g5772,g1394,g6314,g4171,g19757,I21563,g25735,g16567,g15425,I32725,g2417,I37781,g30653,I29215,g30446,g21195,I37994,I39585,g23482,g24125,g8540,g22184,g14114,g24831,g12062,I24520,g8156,g10015,g5678,g21893,g2374,I38920,g8725,g26794,g13158,g28101,g8853,g23624,g11653,I17653,I27385,I22475,I22836,g12184,g8439,g4447,g16351,I40597,g18918,g24428,g18909,g16611,g25015,g19235,g11827,g4731,g23779,g11303,I30335,g2276,g4620,g24180,g30009,g27780,g19534,g27030,g26497,g5679,I40970,I33864,g2433,g2851,g15043,g28681,g5694,I21726,I34421,g27385,g29302,g15240,g1074,g9815,g27091,g5162,g13262,I16601,g17490,I33810,g28066,I36393,I24166,I25521,I15372,I30575,g15802,g13352,g12220,g5369,g25088,g14273,I36129,g599,I32982,g24681,g23862,g20160,g22150,g7230,g23579,g27801,g10651,g19641,g22186,g5138,I27534,g10182,g25236,g4133,g26049,I37575,g24181,g27714,I36557,g24317,I40317,g24029,g912,g30474,g20134,g10067,g24789,g3942,I15191,g17213,I38471,I23748,g30327,g10539,g11732,g29623,g5235,g11039,g17450,g2116,g28189,I35049,g1914,I21488,g18823,I18800,I29405,g21803,I18064,g20598,I33330,g9954,I36954,g5200,g22275,I34782,I31043,g29869,g26906,g27969,g26543,g19912,g23233,g29923,g28276,g7559,I26401,g10301,g22885,g11808,g13304,g30798,g19576,g1686,g27443,g23669,g9737,I21644,g22178,g25874,I35814,g30933,g2700,g21731,I25240,g9822,I30095,g19731,g22657,g26173,g21517,I17048,g5942,g22655,g16099,I24641,I32586,g10386,g25527,I25135,I40573,g5858,g11799,g30089,g28658,g13433,g9793,g23252,g14601,g9077,g23693,I18190,I24271,g20612,I28693,g19327,g13838,g29191,I33608,g9505,I17677,g12814,g11974,g29583,g17215,I31538,I23530,g12462,I40865,g25231,I38518,g15452,g1048,g12049,I27023,I24502,g18014,g536,g11570,I25280,g2354,I30941,g24978,I28184,I32724,g2642,g20402,g2503,g21876,g12933,g17223,I32583,g19237,I15989,g27539,g26760,g10469,g22239,g28972,g22212,I16444,g10888,g28814,g19792,I35092,g29477,g25895,g10638,g17600,g22175,g16221,g19266,g17114,g19176,g29717,g30648,I32709,g28645,g830,g27326,g21473,I21615,I23144,g10096,g25430,g29072,g10628,g15666,g8455,g27315,g17998,g10070,I29736,I23018,I30525,g13420,g16284,g18328,g13373,I29067,g21356,g25223,g8783,g22201,I17951,g22940,g22315,g22204,I27958,g1675,g9941,g22299,g17476,g19026,g24383,g25267,I40901,I28470,I36609,I37650,g22363,g28775,I16867,g13113,g26662,g28838,g5859,g11535,g14895,g13175,I29625,g26619,g15047,g9091,g24343,g18626,I31478,I32661,g17151,I36766,I31880,g25227,g14135,I21160,g30312,g9521,g2603,g25034,I28123,I37716,g12321,g3398,g20605,g20673,g17463,g23003,g24364,I40640,g27886,g27011,g27000,g23237,g4959,g23864,g2661,g26446,g18352,g29399,g29442,g10422,I16279,g28851,g15320,g28079,g20384,g16177,g28997,g13198,g1071,I13110,I23472,I18566,g1234,I22014,g17246,g30559,I16053,g10725,I21955,I20706,g18102,g484,I21894,g21747,g22790,g7635,g4617,g11794,g21266,g25919,g15819,I39533,g13885,g8411,g30751,g10437,g22069,g593,g21789,g23495,I29168,I25728,g21725,g13922,g23517,g30122,g22747,g13970,g20922,I24738,g559,g10446,g29786,I24487,g22622,g2962,g2574,I27358,g20955,I24362,g15806,g5379,g5770,g9450,I21758,g22249,g27260,g23433,g13446,g19250,g19778,g28911,I32296,g3044,g13174,g4067,g24675,g30569,g20506,I26512,g15825,I38139,I26416,g8918,g11964,g15421,g5647,g11848,g8620,g17449,g26074,g19850,g23299,g5955,g24559,I24363,g13481,g28670,g23423,g7806,g18910,g8840,g3158,I37415,g18602,g21022,g18669,g3134,I24326,g29460,I33903,g19280,g3052,g29804,g25237,g13219,I34993,g29359,g19841,g13879,I14094,I20365,g28289,g26786,g11762,g986,g17949,I30901,g12644,I26923,I27074,g20610,I24973,g7590,g21204,g9033,g14922,g17227,g24938,g4791,g11563,g12173,I21775,g10102,g4973,g13647,g3772,g18207,g15995,g1917,g27289,I20305,I31472,I23448,g25260,g2643,g8177,g15290,g28218,g29973,I18485,I32365,I34746,I31571,I23692,g8432,I40907,I20794,g26194,I37095,g25418,g17180,g27515,g817,g2396,g11938,I31068,g7822,g5605,g30328,g16213,I25554,g20621,g16402,I26931,g1825,g19289,I33265,g2688,I38502,g27590,g30690,I25477,g4558,g11056,g23587,I24361,g20322,I27491,g24165,g9120,g5950,g18556,g29939,I26317,I40913,g22634,g20295,g22810,I14621,I39638,g16849,I26505,g9781,g1457,I16479,g18784,g17115,g17925,g24460,I38232,g21160,g21420,g20594,g13166,g18108,I24290,g2170,g30682,g8541,I20486,g13858,g24297,g14450,g20626,g10934,I35369,g22640,I33396,g28049,I40727,g25852,g19622,g17,I36993,I30594,g9160,g21524,g23839,g17457,g26309,I34848,g24612,I14825,g23126,I39124,g29439,g7855,g13439,g3074,I23383,I30493,g27270,g18897,g2108,g27342,g29068,g24342,g448,I25234,g3167,g13537,g16671,g16413,g6194,g19941,g16803,I32919,g13060,g13458,I38352,g13741,I27838,g1229,g19448,I34710,g9290,g25162,g6184,I23715,g12149,g23020,g30277,g23360,I25618,I15350,I20532,I25165,g13265,g8466,g24760,g13233,g24251,I38148,g5820,I21313,g21414,g24385,g10407,g10726,g8132,g24182,I23008,g426,I41138,g21403,g22836,g22646,g22132,g22341,g29666,g23601,g25143,I21505,g13010,g23230,g1018,g4897,g25585,I36630,g5832,g10570,g17717,I31037,I24071,g28970,I25572,g20468,g882,g13453,I40706,g21770,I27717,g27056,g15509,g8825,I34201,g22543,I25889,I39074,I31088,g5257,g493,g7354,I13971,g4070,I18094,g13074,I26664,I31457,I40432,g7993,g4427,g10560,g24512,g5327,g29699,g28263,g12527,I40044,I34343,g24835,g22102,g29705,g6066,g21963,g14238,I19816,g21251,g7158,I23584,I19929,g13442,g15588,g30021,I24353,g16536,g28051,g4322,g30264,g16452,g30717,g24468,I17783,g14119,g24274,g8508,g13268,g13989,I22282,g29346,I30227,I39035,g1052,I30973,I32677,g26355,g24270,g25055,I33630,g28239,I36302,g8489,g1481,I37808,g25648,g20450,I31553,g26516,g8257,g15528,g19155,g24536,g8074,g21738,g29103,g28704,I15460,g30959,g16109,g26105,g27875,I17989,g3211,g18407,g525,g5957,g8839,g27281,g28271,g30083,I21374,g10018,g26298,g11699,g23558,g28058,g24532,I21881,g26336,g16286,g21396,g26079,g30440,g22656,g10952,g8022,g9592,g10681,g29478,g27292,I26444,I17828,g19151,g5508,g9404,g11537,g27079,g20971,g16571,I37122,g28250,g21565,g12128,g28065,g13032,g11980,g29350,I25377,g26570,g2784,g14186,I38761,g4047,g29631,g42,g7146,g30543,I15398,g7575,g21847,I40310,g26925,g29919,g18290,g30983,g13275,g4451,g1905,I36084,I33469,g21976,g28733,g6304,I29697,g21441,g23885,I16021,g23451,g19623,g27510,g30015,g28433,I32266,g26470,I38450,g1694,g2640,I38453,g15990,I31195,g22680,I31541,g26327,g13856,g30163,I16838,g29203,g13580,g30369,g26205,g12158,g18492,g25330,g21339,g24808,g8513,g3237,g24485,g15971,g21084,I20873,g9780,I19689,g19836,g19885,g30947,g29225,g27521,I20613,g19738,g22613,g2908,I38101,g20914,I34818,I23377,I24206,g17219,g17543,g17341,g4757,g20627,I27176,g11111,g30635,g10414,g21778,g1660,g17942,g26192,g420,I30188,g5745,g14395,I40182,I18277,g22716,g12129,g29577,g30963,g13672,g24562,g21285,g5394,g27685,g11500,g11385,g21989,g21987,g845,g15807,g19013,g1700,g26261,g27917,g26728,I39270,I17928,g29250,I19855,g1501,I28928,g21016,g25328,g22143,g23395,g10391,g23830,g12045,g22628,g30863,g8700,g10392,I32973,g29933,g9351,g12075,I34785,g25073,I21822,g28966,g20665,I15912,g9639,g2297,g29920,g4842,g17397,g10146,g27495,g12421,g25315,g29169,I24695,g11731,g8212,g19748,g14613,I41041,g25885,g10521,g10817,g26576,g28710,I32596,g5419,g26791,g11176,I35689,g11516,I25044,I28789,g20866,I38056,g9338,g30408,g19810,I25412,g25449,g5826,I15810,g30869,g18369,g12147,g21759,g29579,g1486,I33457,g13071,g25196,g17313,g24872,g30220,g11996,g13184,g8062,I14049,g28151,I18435,I23191,g9081,g5801,I39856,g24004,g10130,g20472,g22344,I29999,g21375,g18814,I18192,g24374,I13421,g9225,g15634,g7827,g24027,I23581,g12163,I31727,g22914,g19060,g16662,g28010,g24660,g22317,I21626,I25156,I30779,g15625,g27787,I25192,g23251,g15547,I26025,g30036,g21307,g16473,I40661,g1678,g16102,g21911,I15168,g22970,g5731,g20649,g1664,g1544,g20088,g30844,g29428,g4911,g12596,I20466,I29629,I35883,g27509,g16029,g14033,g28290,g12109,g21732,g29091,I13984,g2364,I15226,g5645,g2357,g20581,I26679,g21686,I30266,g8550,I23113,g5987,I32410,g25964,g16974,g25357,g23640,I35458,g33,g21336,g28080,I22657,I15827,g22852,g26956,g19205,g25386,g23377,g702,g23763,g11231,g13329,g15962,g29947,g28078,g19928,g15185,g19197,g18985,g19700,g28185,I18288,g2249,g30952,g13279,g26063,g17720,I16031,g10166,g28998,g25152,g22636,I31814,I31862,g3461,g22231,g27747,g1867,g26911,g19829,I17184,g28164,g17378,g26707,g18973,g10209,g29665,I32453,g2670,g25150,g27376,g28719,I26472,I23278,I40027,g11992,g13321,g5434,g15143,g26765,g24301,g11704,g20711,g15064,g8901,g19512,g26642,I35301,g27914,g26125,g29280,g29634,g25962,I16027,I30707,g5870,g21483,g857,g29479,g1514,I37917,g28610,g29692,g27775,I33617,g30971,g18622,g12860,I22566,g19555,g28232,g26732,g10533,g27114,g2119,I35404,g8699,g10378,g17838,I21723,g27626,g27154,g18717,g27129,g11135,g13497,g17063,I24465,I22527,g20317,g5067,g25957,g1506,I17837,I31847,g22576,I40572,g19041,I18794,I30212,g2552,g19014,g12749,I38662,g16016,g28378,I14877,g25987,g22547,g28012,I32203,g23348,g29120,I38160,g29791,g13714,I32126,g10381,g2795,g28251,g15714,g23917,g24529,g26557,I14618,g25365,I34464,g7891,g23716,g24561,g7461,I36644,g8194,g20093,I16095,g11947,g22776,g22117,g15374,g20448,I33882,g29970,g25865,g19848,g10475,g4899,I16212,g28629,I24657,g21035,g29086,g17620,g17236,g30692,g5591,I15836,g8707,I29159,g29905,g14213,g24803,g29262,g12819,g12252,g11595,g6513,I17840,g24152,I14163,g17200,g6777,g10074,I18287,g7460,g22170,g20535,g5979,g7558,g9453,g16471,g16844,I25021,g22476,g28121,I36246,g27450,g20996,g28238,g7769,g19182,g11382,g10109,g20738,g28133,g11587,g19876,g25321,g30475,g17265,g25582,g16073,I15278,I20529,I14802,I19736,I17721,g10368,g30068,g30934,g16011,I23190,g2362,g21334,g3048,g15722,I23454,g26678,I17854,g18190,I32109,g25241,g8847,g30649,g15161,g17544,g12446,I31130,I36687,I32678,g20345,I31463,g20277,g11431,I35136,I36524,g29089,g1925,g9006,g16074,I29663,g5925,I39936,g6166,g30725,g22639,g18007,g29023,g27724,g19821,g10995,g28115,g22987,I25816,g28315,g21502,g4644,I32137,g24081,g14201,g19939,g5361,g2210,g21373,g17839,g11573,g27205,g8522,g5911,g22875,g17155,g27695,g2442,g30843,I15559,g30687,g24318,g29897,g1237,g19223,I22982,I21739,I28047,g29462,g20430,g10537,g28497,g4925,I20858,g29713,g30412,g30750,I17599,g24622,g14958,g20735,g452,g365,g3678,g4295,I39873,g15496,I33995,g10290,g15415,g25192,g4641,I23605,g19777,g10924,g18164,I25597,g17191,g16842,I37912,I37999,I19711,I34964,g16066,I22988,I40949,g5092,I33402,g20442,I25258,g30112,g28478,I18476,g12052,g12343,g23727,g4512,g20985,g16302,g29490,g863,g29216,g5923,I40627,I36789,g2845,g12445,g16705,I25595,g19441,g23399,g22061,I37137,g27185,g11585,g18120,g1543,g30118,I16827,I31907,g23080,I23406,I32511,g29511,I18761,g30487,g14099,g13417,g9131,g22248,g4205,g5848,g8527,g16417,g10851,g4201,g21842,g5420,g15521,g19388,g5663,I24325,g11297,g26055,g5241,g17913,g22598,g22851,g26041,g11674,I24537,g3337,g21271,g2516,g15761,g19906,g23866,g25923,I37410,g19647,g10746,I14848,g15739,g21742,I21569,g21290,I32308,g23660,g1175,I31832,g19471,g25929,g7910,g25944,g19016,g26013,g28081,I31943,g22220,g29944,g23260,g1412,g21888,I37584,g27165,I16203,g19386,g28298,g867,g23720,g17121,g1267,I34680,I40224,g19481,I28068,I29116,I32928,g19636,g228,g16989,g27810,I25253,g5424,I16321,g26818,g29751,I14182,g28317,I30200,g15826,I29918,g25471,I32719,g283,g13143,g25770,g13152,g5984,g26229,g29461,I33968,I36927,g13270,I41019,g8973,g11879,g2458,g2606,g15726,g18922,g19172,g21761,g10133,g22234,g1235,g24349,g4970,g23826,g29700,I40462,g19023,g12898,g18977,g1922,I40991,g25060,g8556,g18568,g10063,g11918,g16938,g16266,I32506,g21188,g4508,g27588,g20591,I13910,g19604,g11025,I25791,g447,g29139,I39398,g5932,I21865,g18514,I33434,g14718,g19200,g19767,g22706,g22768,I30563,I40604,I24374,g10642,g19812,g20571,g24519,g24159,g25741,g11805,g20446,g394,I40251,g4862,g20443,g14048,g9622,g23179,g27138,g21269,g29926,g21815,g22035,g18379,g27746,g8797,g28555,I23504,g20006,I37038,g9604,g15218,g279,g10197,g25222,g1976,I17992,I30614,g23664,I23207,I17910,g12994,g24820,g20596,g20602,I21037,g11937,I40679,g28024,I20682,I37238,g18004,g30530,I24595,g19565,I28527,g8870,I23661,g15959,g15040,g11190,g27021,I35044,I35872,I20351,I36601,g15317,I22974,g9103,g25404,g29472,I36283,g12038,g20085,g20445,g18011,g25217,g13327,g21917,g5056,g30128,g29630,g24708,g18832,g2803,g25041,g5728,g20050,I39367,I40320,g19091,g14131,I13366,I25561,I37104,g22953,g23584,I34266,g29616,g26272,g10153,g6309,g28924,g20002,g22787,g27394,g25172,I35829,g1712,g24598,g181,g8614,I35058,I21351,I30586,g23493,g2336,I31027,g29314,g26187,I19401,g30371,g5242,g15236,g14525,g18406,g23622,g21346,g8580,g16426,g290,g21609,g25182,g10507,g11847,g12059,g7078,g10373,g5218,g17047,g13560,I20032,I19485,g5473,I32635,g5863,g13094,I32952,g28619,g25450,g10772,I37894,g25177,g7694,g23741,g19058,g27732,g24183,g9303,g23182,g15488,I31469,g24538,I20407,g5326,g9497,I29827,g7358,g17630,g29510,I35461,g1671,g10513,g4797,g12857,g3151,g14234,I24444,g26025,g19624,I40961,g1754,g29119,I18214,g26606,g1491,I25207,g28097,g16639,g21419,g17807,g23099,I36906,I34788,I20048,g8560,g16788,g20119,g26019,g29542,g25012,g12940,g29547,g5948,I29539,g10225,g1303,g29312,g12705,g19970,g8826,g29806,g8447,g12253,I17834,g21640,g9936,g27150,I38486,g19592,g10630,g30477,g10850,I27185,g19869,g13642,I19507,I39164,I37005,g13298,I41108,g15237,g14618,g27178,I18136,g29760,I22687,g29676,g17303,g5754,g17511,I35545,g12438,g11863,g30404,g29942,I17789,g8676,I36230,I32462,I21658,g2492,g28398,g27559,g13026,I28009,g18994,I18206,g18634,g7639,g26546,g2953,I19542,g19233,g21363,g21881,g8637,g26717,g26714,g13894,g20989,g28837,g9115,g15476,g19817,g19930,g1898,g24772,g26850,g10082,g9374,g14438,g28400,g2530,g8662,g11784,g18414,I21711,g24067,g5855,g27451,I24677,g10168,g15470,I30161,g24046,g26082,g7576,g19035,I33198,g21774,g13621,g22050,g21017,I39577,I16306,I19865,I33504,g29815,g18902,g19957,g27085,I33182,g23825,g23852,g24761,g22624,I24299,g5854,g5937,g10327,g28456,I14306,g21312,g26040,g20429,I38665,I29418,g30729,g29244,g27589,g27935,g8088,g2727,g12984,g8536,g12439,g22844,g10448,g25157,I29055,g6064,g1215,I21137,I14091,I33324,g8810,g16049,I22954,g25360,g17050,g9078,I13913,g23262,g29953,I24493,g18894,g26480,g3113,g4095,g12379,I24743,g10835,I30308,g23344,g11779,g7760,g24287,g30461,I16541,I35455,g19740,g20178,g20567,g9226,g12198,g1397,g16343,I19307,I31892,g20916,I37578,g22670,g27998,I23490,g4705,g26087,g26044,I33689,g8813,g19167,g1273,g1411,g17835,g27991,g30375,I23066,g26836,g13557,g28161,g27779,I18386,I39032,g6430,I24923,g5423,g18474,g7880,g21402,g11774,g20419,I13125,g11741,g4282,g1255,g6980,g7841,I38707,g1702,g20415,g15849,I29972,g23782,g18987,g28358,g2602,g21627,g30642,g27229,g15034,I19449,g22003,g30941,g24564,g21802,g28701,g19334,g9640,g17022,g20188,g967,g20517,g5390,g8924,g1417,g8613,g9898,I34707,g23214,g3071,g16453,g27864,g11758,g23284,g26745,g30091,g25369,g27794,g105,g1749,I18704,I23857,I32067,I28130,I32937,g30191,g13107,I18262,g23879,g23613,g22151,g16387,I32092,g7531,I19836,g10329,g20139,I23143,g2565,g26986,I34118,g1224,g25000,g5543,g6427,g14297,g7540,I38348,g8724,I25050,I17670,g22065,g12256,g16383,g10801,g10604,g9629,g19017,g19087,g11811,g23736,g21324,g10631,I18824,g2190,g24105,g11114,g28616,g30347,g19981,g19931,I32265,I22316,g5319,I34077,g26789,g27140,I23179,g29140,g20600,g8553,g21341,I39848,I30236,g24028,g19719,I34180,I23317,I38885,I19886,I37875,g10637,I14668,g14402,g14991,g8678,g19324,I40435,I15958,g28462,I16092,I14446,I17370,g25890,g9441,I32251,g20648,I33003,I38812,g23835,g29374,I36243,g25063,g1078,g27657,g30891,g20614,g2638,g715,g23180,g4143,g10316,g10908,I16002,g4549,g15409,g22297,g18141,g18363,g19971,g30662,I27927,g27010,I32538,g16233,g2294,I19560,g23217,g8904,I23725,g17209,g4203,g12181,I32860,g28761,g24826,g29237,I18686,g24429,g2912,g28741,I35905,g19674,g13249,g1271,g23143,g11926,I32851,I14478,g23767,g20613,g2160,g26834,g28883,I19374,g9098,g24839,g860,I20643,I24307,g5714,g11810,g20016,g16877,g1142,g6711,g10224,g25379,g30950,g21306,g2636,I24196,g23048,g25664,g18963,g28377,g28222,g29673,g12821,g10729,g5153,g13201,g170,g1513,I39835,g28039,I14602,g14378,g1391,I32388,g5873,g26622,g15866,g29317,I40194,g13035,g12263,g23605,I21926,g28118,g27631,g28962,g28236,g11003,g18840,g5296,g29301,g30289,I40016,g29735,g30486,I26630,g523,I18557,I21392,g11579,g11663,g23227,I36307,g30249,I18554,I33249,I15359,g26529,g29269,I17901,g27594,g25928,g30769,g28112,g1268,g16185,I18593,g22366,g27578,g28188,g933,g29927,g29453,g15830,I27191,g29765,I29915,g13962,g29316,g14153,g24163,g15094,I39168,g9184,g19160,g13039,I27332,g24079,g29762,g5548,I22539,I29119,g27255,I16694,g2390,g12920,g26263,g22254,g29885,I40203,g20020,g24552,g9873,g29644,g17718,I35035,g19219,g10765,g2528,g29698,I33188,g23269,g29104,g391,g17542,I14766,g5185,g12852,g1532,I25888,g29651,I21190,g18744,g6100,g17824,g2740,I40269,g9119,I20359,I18644,g28889,g22772,g26260,g27243,g25930,g11552,g18165,g21249,I31535,g11933,I18521,I39916,g24420,g22100,g29624,I35007,I15313,g26729,g6189,g5615,g10468,g13422,g26860,g5411,I28506,g25246,g20103,g30981,g18308,g16371,g30471,I32615,I20886,g26137,g4115,g22649,g16775,g24597,g30505,g24939,g19161,I14104,g21080,I19377,g11907,g15340,g28745,g5797,g17216,g16474,g25056,g19690,g10077,I16309,g23553,I33408,g6942,g13139,I39939,g18960,g29440,I17206,I22671,g21427,g16863,g17799,g28773,g19034,g23597,g30954,g26584,g23353,g1662,g1949,g11324,g29526,I16062,g4073,I33655,g10675,g17696,g21946,g24924,g16189,g23271,g27312,g17055,g16289,I37885,I14472,g28470,g16218,g23904,g13816,I22884,I30632,g20574,I39463,g22753,g7718,I30607,g27026,I25532,I26476,g24997,g3198,g11768,g18543,I32695,g18899,g22633,I24186,g1221,g21090,g23434,g312,g12996,g28031,I23173,g27396,I17225,I31266,g10435,g13548,g21849,g11643,I17972,g24827,g20631,I15584,g18355,g8708,g7533,g24404,g13862,I38821,g5893,g23607,I18674,g19875,g19543,g240,g10354,I24566,g20560,I31841,g27062,g11941,g26653,I27779,g27726,g3210,g17652,I32943,g24809,g16781,g12329,g17598,g10463,g2237,g5665,g3100,g26588,g19786,I13149,g13475,g11720,I18308,g28651,g30774,g2917,I29852,g1418,g12938,g18240,g25797,g28713,g4955,g25206,I35957,g8878,I25985,g865,I31544,g30955,g30407,I22284,g30820,g2998,I21119,I21580,I40116,g27926,I17673,g15763,I23264,I25839,g23239,g15464,g11866,g13360,g16491,g28607,I29975,g4520,g20772,g15603,g21659,g23659,g13077,g29084,I37179,I19645,g16174,g30048,g30179,g1404,g5182,g11410,g20579,g16265,I36690,I34671,g27005,g27074,g20562,g17086,g27240,g21060,I32189,g6157,g20537,g20993,g29448,g4076,g19585,I29077,g16820,I34692,g2241,g4150,g18780,g27009,g20810,I33466,g27266,g12136,g18521,g18965,g27134,g9630,g1115,g4058,I23323,I22999,g24717,g4529,g27316,g23630,I40450,g26178,I38003,g5776,g897,g15115,I31628,g8717,g20769,g14291,g1929,g3147,I36117,g28102,I39818,I18052,I20595,g25071,g19290,g27279,g8221,g26772,g4933,g30224,g8673,g3806,g5556,g28272,I14027,g28464,g12692,g25853,g6623,g30296,g27282,g12091,g16954,g30825,g9632,g29992,g9669,g8824,g29618,g29173,I35961,I23345,g8843,g1666,g28297,g4307,g12017,g18866,I22530,I17942,g23088,g23132,g18951,g6637,I36438,I24639,g27955,I27365,I16034,g30768,I24632,I20417,g12689,g26289,g9027,I28229,g22246,g28042,g30377,g19870,g19244,g21981,g19520,g20325,g13676,g25245,g30403,g24377,I40757,g18354,I22893,g26730,g5831,I29339,g24009,g7703,g165,g26168,g26437,I31778,g15495,I20658,g25264,g28441,I25623,g13450,g18848,g373,I19412,g29315,I40739,g8024,g22362,I36271,g2333,g7900,g1672,I15493,g19886,g22097,g9187,I37950,g28692,g401,g30923,g20883,g1413,I23521,g5853,I20448,g27582,g2790,I35431,g22340,g19265,g23127,g19179,g29799,g1534,g15139,g16857,I23035,g18153,g29214,g5795,g28147,g19021,I27614,g29508,g24537,I40146,I24500,g27122,g24641,g26702,g25490,g30027,g21879,g28403,g29357,g30223,g29968,I16123,g21887,g13066,I14917,g15179,g5985,g6162,g14746,g16403,g13796,I32704,g22165,g12043,g6441,g11472,g27131,g30681,I14624,g4029,I25721,g10907,I32355,I36066,I23478,g16133,g26843,I38958,g10744,g4691,g7353,g15271,g26741,g21284,I35036,g2306,g28342,g23742,g22139,I40307,g28688,g14725,g21746,I39926,I40584,g21353,g10624,g717,g29610,I23967,I35416,g21310,g28709,g537,I30928,g5711,I30467,g26498,I17849,g20963,g16238,g19680,g23616,g11862,g10376,g23364,g24034,g10792,g24491,g20150,g28296,g13419,g17582,I29310,g9913,g24530,g28365,g23889,g24262,g14454,g4828,g29272,g29371,I25533,g17599,g4779,I40611,g11817,g17150,g18188,g27684,g23911,g15754,g28230,g711,g22294,g12759,I27382,g25992,g9056,g13517,I34961,I37059,I31021,g853,g27715,g10818,g12798,g28229,g18405,g26345,I18438,g17197,g2631,g25242,g29064,g16427,g30660,g3111,g1554,g17387,g23145,g21308,g26221,g19890,g22209,g12776,I39325,g15095,g10280,I24608,g23021,g26955,g27275,g5788,g28684,g24610,g23516,g27046,g23273,g8102,I29235,g21970,I35915,g3097,g23279,g27057,g15144,I26455,g28932,g11008,g2673,I31574,I34740,g705,g28269,g22265,g13850,g5936,g26680,I25580,g27762,I29490,g15254,g24921,g28288,g15486,I26437,g23563,g27525,g19305,g29983,I24596,g8215,g8827,g26667,g23167,I22771,I35141,g16655,I31475,g9108,g27931,g2632,I30891,I21560,I31454,g23636,g29657,I29395,I27275,g25394,g13178,I15481,g15723,g19502,g18497,g5819,g17410,g23036,g12002,g26276,I32961,I32153,g25596,I34761,g12691,g5084,g24444,I28076,g22966,g17798,I37641,I39002,g16866,g6016,I32491,g5341,I38827,g11559,g26294,g23229,I35964,g29787,g8565,g532,g24757,g3250,I13745,g20118,I31121,g27145,g10037,I38187,I16185,g25144,g29500,g15604,g5213,g4204,g8564,g11392,g15537,g17567,g21010,g27535,I39930,g866,g27196,g24378,I30017,g10369,g23435,I30158,g6098,g24208,I22506,g11922,g29147,I30128,I36711,g11575,I39368,g21121,g19188,g10266,g27572,g30922,I29948,g21377,g23258,g9326,g13261,g5876,g22334,g2109,g28137,g4489,I33567,g15262,g21421,g22526,g11845,g28116,g29940,g25040,I27749,g28687,g18432,g23629,g29881,g8018,g6977,g18692,g30247,g17300,I18464,g28715,g11915,g19505,g14252,g26547,g7709,I18581,g20977,g23549,g25160,g14520,g26415,g30506,g25399,g2590,g10298,g19144,g24250,g570,g12279,g20900,g23533,I27379,g27905,g30288,g27550,g19770,I36321,g6832,g28463,g12436,g8763,g438,I37659,g20920,I25573,g19542,g11895,g10996,I36621,g23739,g9384,g4688,I35876,g25086,I18402,I26532,g15177,I40236,g25252,g26533,g18665,g13145,g8120,I29246,g26163,g13443,g24824,g16485,g5224,I35334,g20858,g21961,I35014,g29311,g8433,I30071,I40091,g9636,g10062,I40275,g16390,g19772,g20273,g25069,g15357,I35681,g11031,g5622,I15915,g28175,g26106,I17857,g27447,g23476,I26558,I30368,g22577,g24418,g26677,g21871,g11900,g18806,I37266,g15639,g5885,I31005,g16540,g19314,g30787,g20364,I18587,g20967,g20312,g22907,g26017,g22153,I31511,g7545,g15699,g20948,I14034,g24465,I31625,I20571,I21612,g18937,g8548,g189,g8869,g5400,I14874,g18862,g5906,g21423,g11048,g15717,I38680,g10256,g2624,g13271,g11361,g25466,g5827,g27303,g25779,g9117,I22551,g5609,g12450,g12485,g23898,g30572,g15323,g18024,I37394,g541,g10730,g8554,I25325,I32133,g12908,I24015,I20490,g12352,g10145,g29450,g18195,g28393,g24212,g29145,g150,g21125,I40200,g2219,g19042,g23623,g24558,g17046,g13834,g15577,g27771,g20388,g10219,g23599,g8696,g1512,g28435,g29211,I40263,g10319,I32964,I30991,g8821,g8396,g13135,g16042,I37569,g17464,g2342,g4780,g16123,g22357,g30827,g18531,I20577,I29209,g1697,I16200,I37149,g23298,g8499,g9387,g24887,I17881,I36724,g20507,g22068,I25781,I34665,I16117,g29432,g30439,g30937,I14191,g22584,I39803,g21208,g23084,I33327,g22307,g8068,g15560,g16346,g24663,I30353,I36150,g19092,g29207,I40521,I32281,g6897,I28755,g3833,g29718,g7352,I38758,g26977,g25165,I22964,g18980,g15834,g11641,g17281,g16051,I36354,g13463,g23672,g24877,g22039,g29671,g13788,g26081,g25969,g27466,g29790,I25778,g24132,g24363,g18400,g25546,g117,g8766,g16686,g1053,g13112,g10705,g25185,g9061,g30394,I16486,g26983,g26825,g11813,g19313,g29709,g27002,I29687,g28642,I25054,I19628,g24525,g22764,g23173,g28737,g27839,g19590,I35975,g12289,g21724,g22001,g27143,I29369,g28209,g921,g11179,I31162,g18891,g21330,g28307,g23307,g25051,g21067,g16031,I35716,g5836,I25809,I31718,I24317,g21241,g29060,I24078,I32210,I30864,g23188,g24415,g23213,g16128,g4985,g24346,g14359,g19096,I33539,g28153,g21496,g30926,g26887,g19248,I21666,g2842,I16159,I21813,g25368,g24141,I23527,g17475,g22458,I36507,I34767,I34689,g5834,I15620,g8828,I18482,g26070,g11896,g25023,g12060,g20349,g15903,g12251,g11773,g21004,g17797,g20281,I33816,g15721,I33804,g26995,g7664,g23226,I25195,g22493,g20440,g18038,g24402,g16493,g3064,g11515,g23201,g1938,g19779,I23539,g9911,g8180,g19279,g846,I21096,g22308,I32560,g25640,I39948,I19426,I38713,g21415,I36513,I36776,I30293,I28217,g22284,I29087,g2817,g29491,g16625,g16014,g8459,g30444,g26967,g25135,g13654,g12923,I24466,g13267,I21321,I15946,g26391,g20992,g13412,g24849,g6053,g21316,g30297,I41053,g2244,I34836,g5075,g27324,I23163,g19584,I23920,I38157,I26051,g27103,g3103,g19873,I23409,g28867,g6626,I39044,g5730,g2561,g26118,I22690,g23867,g26032,I20131,g5618,g25461,g22835,g734,I30254,g25738,g24307,g27707,I39785,g4301,g23221,I20379,g29411,g12522,I15869,I18671,I38275,g29231,g1206,g26996,g633,I37023,g23225,I31622,g26972,I30976,g23358,I18049,g29166,g11512,g25138,g29092,I32576,g28172,g3099,g25270,I40829,g320,I32892,g22920,g4386,g29766,I36808,g26552,g17948,g1639,g4544,g30507,g5865,g4857,g11899,g21181,g22552,g30727,g21065,g26902,g7476,I37871,g21861,g14158,g17203,g23223,I13207,g9383,g30821,g27850,g2581,g1871,g23896,g30832,I38842,g22583,I37155,I14885,g26367,g1612,g24407,I17750,I26621,g160,I34121,I14775,g2426,g22733,I20619,g28936,g1261,g12340,g22742,g28023,g19453,g23128,g21020,g14212,g29853,I27288,g28349,g9121,g716,g19503,I24055,g12430,g18851,g1227,g17741,I35319,g28370,g30696,g28674,g27889,g5426,g20484,g28839,g175,g18725,g5249,g26776,g20565,g18584,g10014,I20610,g23863,g25125,I24253,g9149,g21061,I14634,g11698,I21949,g26313,g20620,g22867,I36894,g21315,g24000,I16300,g23317,I24744,g29763,g16456,g22328,I23114,g22675,g13045,I33984,g23684,g30095,g2801,g1209,I20823,g28082,I25821,g12892,I16915,g29101,I33282,I19472,g23786,g28385,g22046,g5018,g16062,g20161,I18241,g25065,g29093,g22945,g11422,g25194,g13434,g12449,g18353,I16590,g4509,g11819,g23441,g27419,g6222,g13157,g12847,g15446,g15109,g20449,g26710,g15019,g4415,g23304,I16881,g5719,g13043,g29582,g18872,g23170,g842,g26656,g18763,g25255,g24888,g11551,g18653,I36126,g23685,g9173,g966,g30064,g12447,I16141,I38734,g30282,g21597,g12122,I34957,g10413,g22650,g21046,g17353,g26050,g29215,I35524,I22869,g21031,g29835,I39951,g9933,g12999,g24467,I18458,g620,I34967,I38104,g23845,g12201,g27769,g5916,g24818,g6061,g9649,I16252,g11963,g17874,g29550,g17000,g1107,g20749,I15392,g11078,I32499,g19482,g27711,g15941,g323,g30126,g26679,g26244,I31760,g26884,I36090,g19670,I23739,I28515,g9816,g19616,g25226,g924,g27959,g26247,g22025,I33257,g29370,g27112,g19312,g24466,g22081,g5896,g29489,g29138,I19777,g11965,I39761,g10723,g19855,g29420,g8224,I38940,I25810,g9080,g20001,g12476,g18491,g10332,g10988,I13173,I38620,g26792,I38119,g5677,g2786,I25711,I29402,g28351,I16782,g8794,g16158,I20430,g11542,g9906,g15018,g28475,I37134,g24207,g26384,g23663,I13922,g9106,I13940,g18388,g17297,I36046,I15277,I25383,g3975,g23955,I25415,g11744,g14684,g29388,g19887,I29727,g2523,g13469,g10767,g22196,g19147,g11785,I18250,g11956,I19961,I18223,I26934,g4778,I36407,g26027,g22210,g19157,g23189,g19745,g8000,g22464,g27817,g25579,I35711,g27259,I17939,g20490,I25977,I16114,I21534,g10627,g20539,g930,g28171,I36081,g16323,g21780,g5675,g9426,I13116,g4269,g22600,g23014,g9924,I40820,I13152,g5978,g6057,g26928,g23603,I40847,g25353,g5949,I35759,g24231,g28311,g13095,g23734,g5078,g17486,g28661,I40790,g13121,g8594,I37901,g15638,g21903,g942,g29551,g29466,I24694,g13042,g3253,g17208,g13489,g22356,I31904,g12965,I25607,I30299,g6149,I23733,I18755,g12547,g27323,g11837,g26815,g8164,g5614,g11826,g15932,g28352,g1677,I39385,g11946,I32380,I38035,I18835,I18172,g30818,g14960,g10526,g19799,g2607,g2536,g27686,g133,g27203,g18845,I31152,g25851,g1862,I17963,I21730,I31928,g30252,g24275,g7892,g870,g25646,g27158,g21775,I25004,I29016,g26905,g24294,g12185,g28243,g4711,g25043,g17084,g24836,g26542,g2165,g30555,g18772,g19807,g16528,g23250,I23065,g21068,g22262,g13344,g25075,g27027,I32167,I19211,g20965,g18783,g16924,I33828,I30519,g26668,g16599,g26512,g24356,g11903,g147,g26698,g7877,I31796,I25820,g14023,g10286,I30841,g13144,g15592,I30257,I25829,g21877,g28582,g17670,g10708,g21912,I31071,g29523,I19803,I38190,g15682,g30953,g30370,g11973,g27199,g10438,I19503,g18590,g23680,g18879,I40578,I40673,g30216,I30790,g5715,g5667,g12055,g22197,g27830,I21747,g27216,g13181,I20526,g21650,g26030,g21880,g26747,g26755,I30077,g19888,g11997,g10639,I21064,g8714,g29261,g5038,g24233,g17563,g3990,I17103,I21381,g26474,g10079,g10144,g29557,g1008,g24387,g15449,I38602,g22717,g9968,g954,g285,g24623,g6367,g26281,I39922,g2418,g23774,g27455,g304,I29996,I17297,I36078,g10763,g22762,g16000,I33680,g26129,g30381,g30011,g4908,g27773,I15183,g17648,g9440,g28047,I36571,g24793,g8569,g30877,g24355,g30503,g22376,I13320,g20146,g17900,g26752,g427,g6103,I32042,g30123,g28472,g28410,I36300,I30047,I30860,g12695,I40101,g27846,g24419,g21867,g11438,g13263,g29387,g7809,g12146,g20493,g534,g8001,I15623,I17737,g12292,g23212,g5750,g22845,g24267,I22860,I31257,g543,I14637,g1176,I13820,g17526,g14090,g26883,g758,g29552,I30598,g23542,g21041,g24499,g15650,I33894,g12944,g30912,g23199,g5135,g21762,g9319,g29732,I20504,I22521,I34946,g16075,g25771,I30816,g9888,g19100,g4891,g10542,g26650,g15197,I24485,g13999,g1829,g21786,g17749,g23728,g16370,g27903,I25210,g19796,g18484,g25667,g22343,g23074,I37804,I33551,I33849,g11870,I37790,g21928,I22707,g3995,g27858,g18968,g22720,I18599,I19759,g20399,g23007,I38710,g30703,g16310,g21177,g9137,I38342,g26716,I33695,g3182,I23046,I23751,g19059,g2039,g7142,g2903,g2645,g12912,g19566,g27256,I25560,g9903,g16462,g25745,g16442,g1526,I31065,g27936,g21808,g9895,g1089,g26416,g26373,g6055,g23511,g27012,g27119,g28416,g1256,g21425,g28356,g28212,g24401,g21258,g13021,g6713,g26091,g30780,g24543,g22250,I23553,g28581,g26649,I34168,g20067,g9809,g1416,g2978,I29098,g28157,I36667,g2651,g18964,g11984,g10220,I23009,g24475,g11373,g12952,g18812,g1597,g14175,g29652,g21666,g17248,g8200,g28099,g28899,g10395,g27244,I40654,I40594,g23259,I33000,I40643,g14228,I30230,I27727,I36663,g26342,g23301,g15766,g22309,g11163,g15867,g24280,g2694,g14371,g25384,g12876,g29952,g24373,I39014,g14001,g20572,I23999,g27723,g26341,g11092,g1745,g5786,g4424,g27204,g18853,g4098,g21677,g21107,g26352,g23793,I30092,g19277,g24278,g1024,I16163,g27108,I32129,g27361,I38505,g30752,g29426,g18152,g30677,I13934,g18656,g3061,g5335,g16341,I31523,g22566,I17666,g20757,g28920,g26826,I20431,I16627,g27973,I39806,g13635,g16472,I25429,I35900,g1088,I40880,g16012,g1378,g24766,g29219,g20197,g30389,g30522,I31715,I39154,I39237,I40688,g15531,I36972,I25802,g24271,g8863,I30689,g6517,g16529,g25229,g30044,g9442,I40742,g19744,I35756,g10866,g19871,g17796,I20328,g15844,I30320,g26997,g25811,g17294,I32625,g20589,g30492,I33593,g5104,g18603,g12107,I28096,g25261,g13466,g27297,g29304,g9003,g20841,I16735,I30531,g11141,g29368,g27186,g23914,g12235,g14256,g18765,I27531,g21180,g20827,g21112,g30632,g19329,g2206,g20669,I18028,g30797,g30353,I26377,g24106,g23593,I40537,g22651,g29803,g16939,g19918,g20545,g20878,g26301,I37050,g30875,I36948,g3919,g2612,g26743,g25342,g14194,I20547,g23208,g4997,g24400,g16659,g21883,g23620,g27731,g22701,I24263,I37182,g14011,g24504,g3194,g9635,g15314,g9868,g20094,g8400,g2256,g12161,g15835,I25717,g5145,I31733,g23308,g12494,g20136,g15680,g23376,g18573,I25673,g349,g23746,g24221,g12477,g19271,g8915,g10261,g30771,g7963,g23309,g30493,I30925,g21690,I41102,g18296,g19052,g12120,I35886,g22227,g28432,I15806,g30870,g2582,g7548,g25684,I18470,g22632,g4662,g4401,g12608,g1151,I33819,g6135,g25717,g25523,g29784,g23042,g24078,g21044,g27565,g24492,g5959,g21021,g25623,g10320,I22651,I14712,g7482,g30025,g29160,g15389,g26048,g26816,g10401,g11892,g24126,g27049,g22174,g1244,g1205,g22281,g8369,g29002,I34395,g15243,g30876,g16802,I38462,g1056,I31102,g27805,g21343,g15901,g20058,g2360,I35389,I18163,g23686,g19820,g19672,g22314,g21969,g5395,I26481,g1114,I36530,I19859,g23726,g26325,g19184,g27358,g25366,g26613,g28567,I30888,g22192,g21025,g26501,g6099,g12926,g12998,g26872,I24647,g27296,g11364,I19739,I29459,g16178,g17965,g25263,g28556,g27632,g19932,g3997,g25240,I28323,g30799,g22048,I20324,g25333,g29053,g18368,g20898,g28612,g13022,g587,I23392,g19080,g11734,g27193,g5650,g23030,I15577,I28346,g28257,g1164,g1946,g13868,g5815,g30397,g21452,g4685,I34405,g23877,I22820,g25773,I37502,g30960,I27733,g19112,g428,g2081,I29243,g3135,g5421,I22524,g21586,g18246,g26005,I33670,g15118,g11530,g17474,g1466,g25976,I23466,g16360,g20366,g24069,g1951,g8460,g4836,g17737,I39919,I29223,g9889,g11971,g2228,g24442,g17021,g17691,g3095,g9025,I24319,g11904,g19346,g23836,g22431,g22041,g30497,I29132,g26597,g22313,g10293,g19856,g19389,g11290,g10419,g13072,g21470,g24592,g13328,g30931,I27125,g1054,I17486,g20314,g25590,g15037,g10671,g29300,I19595,I20676,g16139,g23406,g27395,I38804,g28119,g12822,I40465,g21233,I29588,g25932,g8028,g8363,I33683,g30873,g24545,g1537,g1723,g17399,g30410,g10617,I35904,g28057,g29608,g22106,g20927,g22155,I21551,g30147,I28003,I28727,g12993,g30936,g5004,I32295,g21253,I27278,g17024,g14068,g20570,g11844,g30498,g28411,I33168,g30872,g29635,g10117,g5697,I34909,g7619,g30916,I24215,g252,g26308,g5683,g21040,g24241,g30754,g15017,g18079,g11979,g9726,g11332,g999,I15800,g28859,I21012,g24989,g9603,g13351,I18605,g25499,g25198,g25049,g17149,g13297,I36536,g24776,g5751,g23319,g679,I29641,g5729,g5662,g27743,I14857,g8529,g25103,g10810,g29054,g5167,I36650,g14280,g26770,g14737,g22558,I38163,g19412,I14609,I18810,g24819,I16332,g12470,g25329,I40958,g11854,g1541,I33961,I24486,I16138,I19174,g19051,g13602,g9468,g13001,g2874,g27694,g20874,g29464,g12452,g20632,g27332,g2393,I14739,g23013,g989,I32248,g1562,g13092,g29260,g30087,g5089,g2133,g20487,g2792,I34433,g24589,g23218,g10262,g15251,g2250,g16108,g27583,g29313,I31112,I36347,g9733,g13308,I40931,I39540,I39340,g1409,g22257,g21806,I32480,g12005,g18539,g21355,g23576,g25403,I18488,g19138,g10929,g22244,I26458,g29694,g14669,g20288,g9112,g26759,g9626,g29889,g16492,g10911,I37334,I24415,g28499,g9581,I39047,g22551,I28518,g24454,g8861,g17131,g18105,g19552,g10394,I38434,g23303,g27034,g24854,I33542,g25784,g24683,g11820,g14642,g19523,g11823,g4246,I30713,I39145,I18326,I25644,I13801,g26941,g26318,g8025,I16524,I16826,g18795,g21062,g28015,I29135,g4221,g7751,I38671,g24217,g16039,g26909,g27968,g1527,g12804,g19863,I35791,g10876,g18003,g15487,I29336,g10629,g30489,g14472,g29402,I24626,g29358,g29473,g17354,g11051,I39985,I39773,g19498,g25802,I34244,g5946,g13865,g25859,I21407,g25116,g27075,g26823,I25723,g14097,g17601,g28375,g30221,g20190,I19915,g28013,I17156,g20813,g27735,g10228,g27217,g21646,g16797,g7858,I31133,I16234,g21203,I40826,g23621,g6676,I24950,I26396,g5346,g4214,I29978,g29684,g19605,I24112,g13260,g10714,g21184,g1918,g1676,g5879,I19905,I30844,g1886,g22761,I36563,g29812,I13655,g4832,g28649,I18232,I30695,g29840,I16681,g21011,g25413,g18395,g21263,g4647,g28640,g10105,I33482,g5057,g22804,g5902,g30133,g29395,I26369,g28423,I27065,g28003,I23893,I16880,g12079,g6084,g22806,I27155,g11263,g27135,g12504,g9010,g10310,g21671,I38282,I34096,g9159,g5149,g22337,g15797,I39029,I40784,g26448,g30957,g30175,g30077,I15830,I40527,I30948,g2095,I22989,g7610,g11002,I34728,g5702,g10205,g19854,g24549,g17428,g13317,g24777,g5802,g18930,g25940,g8521,g19837,I40152,g23151,g18212,I28766,g28979,I16341,I22800,g5626,g27924,I18668,g19570,g29688,g25370,g24505,g23098,g30395,g2821,g24253,g11630,g10724,I34086,I36618,g24110,I40059,g26608,g9099,g26709,g12808,g22027,g19089,g19718,g24219,g13395,g12490,g22834,g16220,g4182,g13193,I21045,g4220,g28744,I25655,g5992,I25308,I16644,g27290,g15337,g4905,g28127,g29239,g11887,g6438,g2772,g13187,g11497,g13750,g30812,g26746,g22273,g21207,g26379,g23149,g19381,g7706,I29536,g14829,g30733,g7424,g27703,g7911,g22731,I16832,I13804,g12893,g19476,g7527,g24431,I22022,g23537,g27834,I18187,g2611,g22614,g28609,I36257,g24261,g83,g109,g6130,g20502,I29550,g4111,I19598,g12268,g23140,g12020,g24804,g27549,I34029,g23973,I17051,g12291,g19272,g13918,I19797,g28893,g17201,g27194,g4526,g10094,g13117,g12486,g23082,I25683,g16935,I40877,g22230,I39902,g25204,g15390,g23557,g27239,g4888,g11492,I36975,g1195,g15904,I36990,g11842,g302,g9957,I32439,g10589,I36432,g19107,g5771,g30944,I34650,g17045,g15758,I32445,I18432,g8093,g12880,g12604,g30806,g20451,I17889,g20127,g16001,g18333,g25946,g25286,g14637,g8083,g19572,g12457,g982,I24388,I36417,g19226,I21297,g25176,g27152,I27221,g8574,g21634,g19702,I29229,I34009,g26749,g26767,g26867,g5760,g3079,g2261,g30254,g27060,g10831,g2811,g1772,I37297,I21862,g25707,g20746,g11816,g2138,g11129,I18295,g13003,g5234,g29482,g27478,I19605,g22161,g30116,I16354,g26598,I24587,g11145,g22336,g15326,g24482,g1816,g29536,g26869,I25847,I24603,g7134,I31871,g21945,g8255,g26026,I28435,g9605,I32081,I15262,I29921,g28322,g1923,I24036,g30551,g17395,g19663,I23968,g11786,g859,g10749,I25773,I28792,g26383,I32528,g22647,g1406,I17012,g21950,g11306,I14442,g22304,g4202,g17875,I13968,g22509,g25400,g21752,I30803,I29672,I26195,g2933,g11930,g16127,g5343,g23040,g2312,g19345,g29063,g18401,g26553,g28677,I24103,g10660,g1067,g19615,g5922,g1609,g5986,g29098,I27488,g13031,I14891,g9761,I34128,g22127,g28266,g13634,I32844,g10309,g18967,g16285,g28680,g30445,g20382,g5061,g18542,g303,g19103,g26629,I40709,g28035,g24830,g24322,g26076,g26969,I28210,g15130,g4254,g16586,I34704,g13206,g2392,g22678,g16813,g538,g30762,I35360,I31417,g29567,g22145,g8449,g1887,g18222,g7583,g2477,g9044,g13461,g2992,g23865,I25792,g11020,g28089,g23679,g2309,g1186,g9912,g30683,g499,I23341,g17594,g20499,g17118,g26819,g25305,I21452,I34385,g23795,I16193,I30305,g20464,g20742,I35042,g20500,I29313,g20962,g4708,g7742,g18728,g23261,I35945,g11961,I39127,g17761,g29467,g13764,g26189,g22198,g27391,I18199,I36008,g8605,g24762,g3006,g16459,g18623,g12180,I31685,g26265,g22026,g9461,g12051,g4283,I21830,g4016,I23651,I32901,g19264,g9287,I36390,g28986,g23665,g24837,g4082,I25800,g709,g13390,g23642,g18037,g22146,I35944,I25516,I13677,g4538,I26500,I19573,g28347,I35410,I27335,g27855,g8689,g20241,g11494,g30438,g19843,g27463,g24866,g10497,g17812,g13234,g28419,I24716,g27163,g28214,g24216,I29656,g21605,g24816,g26758,g26715,g15096,g15762,g14342,g13565,g22002,g25981,g18831,g12747,g19111,I25041,g20973,g13368,g22570,g10784,g7923,g5917,g22586,g22266,g973,g11877,I25320,g3078,g11880,g20974,I29073,g9923,g5713,g7785,g15842,g30393,I26538,g17514,g25142,I29475,g10238,g15048,g18884,g23712,g19666,g26628,g20158,g23168,g12156,g10150,g7083,g4603,g121,g26090,I31667,I39809,g22218,g2991,g20945,g19008,I27972,g24001,g1542,I27672,I34986,g513,g21577,g20964,g9019,g18719,I34656,g21140,g21974,g29656,g24576,g21737,g9955,g21329,g21962,g30984,I36996,g8802,g16253,g25010,g11716,I18004,g27712,g8543,I32325,I18653,g27425,g15827,g16761,g7974,I20839,I15204,g2676,g2009,g15308,g4769,g29288,g30546,g5375,g5126,g28468,g8667,I30954,g25133,I18420,g18890,I30365,g18435,g28452,I30074,I14113,g26882,g24127,g17576,g11700,g26457,g19634,I24546,I23424,g28740,g7733,g24243,g30586,g29127,g29611,g27231,I35834,g29816,g27036,g17887,g12816,g27483,I17701,g10778,g22208,I23863,g25493,g21429,g20427,g15812,g9118,g18244,g28268,g28226,I38716,I25567,g30399,g27132,g12981,g7646,g27379,I35020,I37203,g12039,g4860,I17860,g6751,g1982,g23715,g8045,g11533,I29600,g10613,I22925,g26664,g30622,g17369,g21445,g30001,I16562,I21992,I36289,g27224,g28697,g11506,g21255,I18217,g26641,g29470,I24298,g23069,g27340,g30656,g2780,g30693,g18088,g22880,g29107,I34758,g24875,g15355,I34453,g16009,g11671,g17439,g12791,I30125,g17451,g18824,I28159,g24753,g28663,g15225,g25487,g30583,I19784,g16884,g1530,g15219,g30292,g16300,g6912,g8931,I24005,g24357,g1415,g12642,g29292,g24750,g5163,I27303,I17698,I29559,g5349,g16964,g24455,I28201,g13914,g2549,g5101,g19236,g18947,g15950,g29848,g28055,g5746,g20623,I17641,I16879,I34233,g30571,g15142,g8502,g23211,g27728,g1420,g25327,g22737,g19695,g25540,g30756,g18586,g18836,g28083,g24566,g12087,I15469,g28551,g28686,g24920,g10154,g24782,g11546,g4623,I14413,I17866,g27613,g21760,I23894,g15499,g13002,g23153,g22379,g30862,I29372,I27992,I35859,g11627,I23244,I40565,g23596,g12973,I18375,g10901,g6632,g30838,g20476,g24299,I18184,g24175,g1199,I22946,I23824,g15999,g10312,g11967,g5422,g28190,g25787,g496,g29639,g13487,g26540,g16393,g3951,I36147,g12510,g21758,g13120,g20456,g26549,I24512,g28655,I36577,g19533,g13331,I39647,I24426,I34051,I24394,g10432,I14631,g27094,g24376,g13370,g24770,g16546,I30508,g18635,g8755,g1845,I40571,g10360,I14571,I27766,g22066,g27553,g22713,g29515,g30326,g19106,g25091,g29178,g11596,I30716,g13326,g19949,g27264,I39401,g18787,g1961,I30344,I38088,g26572,g1950,I20802,g7532,g7999,g26579,I33382,I26112,g2605,g408,g28422,g28388,g28685,g25936,g12366,g11453,g12690,g9449,I32970,g16005,g16498,g19238,I14599,g2564,I39234,g11901,I17895,g29463,g11287,g1642,I23842,I30776,g14408,g10532,I15616,g10445,I36779,I17792,g26374,I31940,I18515,g27542,g13479,g28246,g11386,g22125,g20826,g19356,I24102,I36879,g977,g30383,I19972,g388,g29194,g24937,g29499,I27188,g23318,g19177,g26349,g10966,g28413,g23919,I25635,g14502,g2229,g8494,g2480,g28155,I24408,g21870,g27299,g5366,g15854,g14650,g16770,g12545,g28584,g4405,g12054,g27427,g27156,g22879,g7745,g22872,g20732,I14295,I30347,g10340,I20497,I33649,g2900,g21960,g25274,g12103,g10486,g5882,I40555,I40979,I20476,I23371,I15918,g28034,g12021,g24584,g13873,g14464,I38767,g27667,g28406,g6898,I34172,g24965,g5938,I40841,g26232,g29094,g25117,g20542,g15978,g26346,g14032,g25151,g6426,g14559,I36069,g29612,g9921,g20186,g13313,g23205,g12555,g1624,g740,I24619,g6065,g9926,I25848,g291,g16241,g19163,g24973,g16048,g27070,g23203,I31910,I30847,g7079,g22874,g22235,g24123,I24612,g19952,g27310,I18016,g11598,I17557,g25988,g5961,g7676,I38097,g24093,g2444,g23095,g25565,g2466,g11318,I25371,g6038,I35434,g1880,I29456,I31144,g29681,g20373,g13069,g23858,I31700,I23559,g28314,I21586,g578,g24070,g991,g10994,I18662,g27321,g13142,g26222,g1792,g25299,g22382,g24368,g28329,I23808,g16030,I35123,g8684,I34662,g29291,g10905,g7856,I16169,g2827,g13020,g15022,I37863,g20013,g2986,I18055,g2175,I29660,g19784,g21262,g3866,I18037,g25484,g17339,I39333,g16395,g780,g23296,I33440,I38360,g27250,g12561,g2833,g17255,g25892,g30907,I36984,g23165,g213,g23856,g27101,g1059,g25515,g23945,g30964,I25855,g13852,g26532,g11294,g19775,g30783,g15188,g21404,I29448,g7799,I37635,I15212,g22644,g24607,g21018,g19648,I29151,g23743,g8465,g23402,g5830,I36912,g23591,g26683,g1560,g13849,g10444,I29265,g10936,g14703,g22385,I35022,I14143,I29007,g21777,g26304,I29930,g19354,g26389,g4922,I40441,g1352,I39071,g4348,I20589,I29632,g22595,g2090,g12076,g26748,g1098,g4339,g7802,g26279,g23064,I25682,g17865,I32112,g11444,I27206,I26615,g19660,g11969,g5988,g7833,g12794,g19326,I28111,g1748,g28451,g1476,g28428,I36135,g2470,g28682,g17222,g23107,g6087,g4421,g4486,g18311,I23235,I24513,g14775,I25612,g5504,g18689,g15282,g11182,g29754,g17506,I36574,g4101,I23132,I25700,I16098,g26700,g4430,g24473,g23489,g10186,g4873,g2118,g27121,g18835,I30056,g21931,g16041,g11982,I36447,g17122,g28617,g30613,g22259,g22279,g16089,g30018,g26400,g23339,g13675,g350,g749,g12082,g28338,g1685,g20321,g26226,I27228,g29112,g22724,I20462,I33006,g5431,g2454,I15599,g29099,g3063,g23177,I34277,g24704,g24489,g732,g14052,g24147,g1690,g23606,I25904,g18756,g27033,g24653,g20015,g20822,I24553,g26347,g300,g17635,g30380,g24813,g15606,g30951,g16513,g1651,g13867,I21655,I36256,I13868,g23509,g4437,I14519,g8532,g8209,g20387,g21739,g8703,g29416,I23518,g23972,g542,g18934,g29834,g22527,g10580,I37484,I32880,g24871,I36633,g4197,I29481,g24408,g30621,g25997,g24723,I30663,I32669,g15080,g25634,g20672,g24518,g22129,g10821,I31601,g9670,g29672,g21958,I13211,g720,g30738,g1808,g10676,g9097,g20135,g14053,g2105,g18917,g11169,I36382,g11503,g29728,g30970,g24436,I21691,g24411,g28394,g13102,I28541,g322,I31679,I36516,g24593,g24372,g10078,g15508,g26424,g7826,g13637,g21113,g5334,g5438,g18916,g28779,g24059,g12231,g27168,g28337,g9111,g4967,g13295,g24720,g19889,g134,g22138,g29540,g19171,g92,g834,I37961,g5378,g23155,I38704,g9498,g4130,g22635,g15454,g11538,g8417,I19488,I20805,g23124,g27223,I27257,g24784,I19587,g27527,I38408,g6033,g26062,I31595,g19270,g8296,I37765,g19712,g28004,I17969,g27180,g8153,g5944,I35072,g23174,g11962,I13504,g7950,g6028,g15824,g16350,g2571,g28871,I24149,g30553,g2483,g101,g6204,g14091,I29984,I16517,I23923,I30032,g17161,g9880,I21806,g8181,g26804,g30566,I37386,I35906,g2580,g19788,g3086,g7927,g9096,g19010,g16446,I17825,g11760,g20087,g988,g19318,g14385,g21120,g29703,g18121,I15169,I31865,g21514,I25228,I16318,g26788,g13155,g8443,g29095,g27912,g21230,g12941,g16758,I16661,g16643,g24100,g20980,I23020,g25887,I24228,g841,g7925,I31934,g15847,g26559,I32916,I14020,g21971,g1192,I29378,g4124,g13626,g5803,g18821,g20609,I20649,I22900,I41123,I25291,I30501,g21869,g22124,I32333,g13075,g11330,g13339,g18371,g14067,I35011,g29193,g30028,g17220,g18931,g2594,g7901,g9471,g13438,I30979,g21321,g5292,g5969,g28046,I13275,g26599,g176,g24056,g11583,g7757,I39065,g28146,g28030,g28647,g11219,g24443,g2247,g7823,g29167,g8905,I24704,g8940,I29863,g23969,g20422,g23604,g25149,g19717,g10100,I38916,I19774,g29959,g28221,g24805,g21533,g5977,I34824,g17030,g28955,g28316,g29533,g17097,g20370,g27218,I20655,g7834,g26654,g20580,g27569,g16535,I23162,g30614,g25081,I16747,g27872,g18838,g29076,g13946,g27404,g1220,g25179,g11909,g9092,I32310,g24850,g833,g2679,g15868,g25385,g22260,g20012,I23198,I38623,g13493,g9133,g10859,g22546,I25071,I29033,g5716,g30704,g10516,I25037,g19175,g1795,I38866,g28108,g28418,g29073,g16336,g14904,g16878,g906,I14069,I14628,g21073,g30839,I21694,I29562,g25118,g125,g12272,g18785,g10066,I25890,g26113,I31919,I34135,g26577,g21352,g26046,g10185,I32057,g19196,I29104,I34017,g15711,g27503,g17855,g29118,g30892,I20386,g528,g19045,g8135,g28944,g5844,I23181,I26910,g3104,g12871,I29010,g23539,g19724,g19881,I17916,g27838,g26554,g17529,I39641,I23807,g26166,g13495,g28445,g5635,g12407,I29415,g1668,I21432,g2142,I35897,g26340,g20505,g14268,I29129,g18976,g24282,g30098,g1174,g28043,g3050,g20436,g14546,g15392,g28220,g9364,g30502,g24779,g623,g26891,g30362,I16074,I25183,g813,g30684,I18635,I31436,I18509,g27697,g15970,I31856,g15510,g27278,I17373,g10107,I21844,g30760,g704,g20970,g21104,g19954,g319,g10467,g25348,g21864,g21400,g13064,g19062,g9022,g26350,g15897,g12085,I35440,g13347,g14955,g28054,g20318,I17756,g16722,g1387,g8835,g9026,I25701,g21968,I28455,I31091,I16176,g29168,g30295,g21458,g30965,I18506,g12065,I35034,g13529,g28174,g19102,g13292,g17394,g29513,g24672,g29465,g3677,g26422,g3105,g21211,g29988,g26582,g2697,g12179,g13459,I29951,g10173,g30055,g14007,g10515,I36582,g18876,g29134,g22131,I23556,g2556,g26056,g9123,g17352,I29090,g2527,g20283,g2,I29301,g24812,g2848,I17066,g4471,g8347,g25068,I39261,g2969,g26121,I29927,g11309,I17981,g21741,g13283,g29549,g13294,g10217,I27056,g30803,g23061,g17166,g20455,I18969,g25016,g20779,g12274,I18229,I21329,g20292,g22494,g30248,g5688,g26541,g29647,I19533,g2799,g28264,g28459,g24223,g26495,g23236,g29662,g8846,g24462,g22906,g146,g11666,g2720,g22626,g12130,g12431,g28915,g24080,g11589,g23843,g29697,I31691,g4717,g25363,g18061,g11021,I18079,g24636,g16461,g13028,g18999,g1000,g18782,g28156,g1005,I40288,g19199,g28429,g20407,g30678,g4436,g16026,I14384,g12033,g10431,g18953,g27540,g1216,I15636,I38107,g23942,g15198,g4263,g25998,I32400,g8340,g29303,g26464,g30388,g13100,g29727,g1101,g30867,I28013,I28034,g23895,g14773,g12242,g2227,g29441,g23016,I24726,g18827,g4982,I24389,g762,g4671,g25266,g15426,g29142,g30639,g7838,I23055,g11777,g28087,g13068,I37185,I30832,g8844,g26762,g19468,I16720,I27059,g88,I20310,I36891,g4693,g11818,g16211,I39252,I18497,g28323,g26211,I15876,g11355,g4861,g8065,g7638,g30519,g10849,g23315,I34363,g24957,g21399,g9365,g25744,g24574,g24853,g27575,g8097,I38241,I33954,I14786,g26921,I25914,g15753,I23682,g4061,g5592,g16020,g28120,g29451,g11846,I34068,g27422,I38014,g19975,g23692,I33867,g27331,I26913,g29670,g10748,g11746,g29995,g20421,g12521,g14249,g16401,g23254,g17785,I27321,g13080,g7670,g8894,g12815,g9174,g29678,I15445,g14366,g29780,g1424,g24644,g23770,g5816,g5179,g14592,g22280,g27141,g17585,I24494,I41050,I28488,g30014,g19569,g23906,I33906,g20683,g6161,g951,g20408,I29939,I27416,g13299,g28874,g28540,g30823,g3002,I38725,I20455,g30815,g25061,g27232,g24300,g3094,I34770,I13501,I28981,I13999,g27017,g25129,g1358,g12600,g19064,I34866,g6183,g19948,g15545,g17713,I39038,g18537,I38459,g8948,g714,g19809,g2592,I19654,g28553,g11894,g23731,g22365,I15230,g21927,g8467,I39404,I21554,g19299,g450,g429,I18461,g24230,I30185,I41126,g21019,g14229,g1339,I39089,g13657,g3132,g24883,g30608,g30668,I37590,g29217,g28294,g24768,g28778,I17922,I14525,I23253,g28488,g24745,I34479,I22414,g4601,g19215,g27320,I29530,I25899,I32509,g20156,g16103,g25520,I20580,g20592,g10983,g20437,g23918,g17825,I25872,g24066,g14881,g22870,g5935,g27295,I37110,I26708,g26761,g25790,I17892,I30050,g21495,g16640,g23157,g1113,g20357,I28512,g2098,I16504,I38428,g24964,I18638,g21344,I16511,g11069,g22672,g22727,g26719,g17240,I37188,g19828,I30383,g14041,g28224,g13646,g29524,I17727,g16311,I40221,g27333,g25518,I39323,I35799,g15585,g25254,g7227,g27704,I17807,g25658,g4418,g5804,g19556,g719,I39800,g8547,g30629,I14709,g10436,I40191,g4668,g5352,g12013,g29287,g22172,I32877,I40242,I40444,I21491,g29565,I31232,g24739,I21708,I27017,g19101,g25948,I13197,g13133,g11893,g4928,g9962,g20684,g26392,I31949,I20667,g19758,g1422,g582,I36604,I22918,I16258,g1385,g12125,I30314,I16854,g26661,g8643,g24780,g23682,g27999,g13063,g27595,g24767,g56,g4736,g11685,g2812,g28132,g20285,g22300,g8452,I40054,I24291,I15657,g23723,I23588,g13172,g23147,g27678,g17001,g19348,g23031,g7553,g22339,g14102,g2046,g9583,g30779,g7697,g9048,I21520,g1252,g19037,g28390,g24510,g28109,g29326,g21902,g2818,g16180,I21108,g17342,g28122,g10612,g24394,g12215,g12425,g25723,g22342,I13224,I28305,I14948,g10442,g25296,g21810,g24397,I16993,I30931,I34183,g20693,g3136,g20575,g19575,g12444,I32994,g12266,g18869,g26853,g29141,g14092,g26366,g30740,g2944,g9067,g26544,g27792,g5623,g21825,I31853,g21050,I30086,g1069,g28371,g12178,g30332,g25891,I37813,g26806,g21179,g20924,I30751,g15989,g16217,g25826,g11284,I19800,g24090,g15594,g10214,g10980,g22901,g20790,g1693,g26262,g21480,g22587,g5924,g23585,I16684,g17968,g3108,I31688,I16726,g11691,g19242,I14942,g28427,g909,g12850,g30303,g27770,g15263,g24906,g3305,g24832,g13214,g29027,g26699,I39407,g2587,I39369,g1778,g11594,g28476,I27621,g25024,g23943,I16593,g30396,g27314,I16611,g13643,g5664,g1819,g15755,g5823,g18860,I36718,I17995,g23272,g12979,I31213,g10367,g3934,g4340,I23152,g4948,g15580,g16425,g29183,g21083,g8784,g13499,g17882,g8285,g2667,g29505,I31062,g1783,g24461,g15136,g15578,g30736,I17159,g8533,g15407,g1531,g16448,I16360,I28473,g18690,I18784,I15971,g10754,g23521,g21015,g10101,g24585,g1630,g25714,g29266,g8811,I33840,g21926,g22271,g29436,g24434,I30203,g22503,I37280,g26007,g30746,g16454,g21965,g30053,g13240,g26235,g20947,I41129,I35422,g21175,g7587,g29389,g11855,g179,g17645,I23398,g4335,g506,I18725,g6905,I23421,I25074,g27543,g30330,g8395,g1516,g13058,g27671,g7772,g16804,g23268,g10113,I16664,g28067,g1765,g6643,I23074,g10045,g22609,g9621,g20725,g8677,g20218,g27823,g23071,g14098,g20418,g26682,g18923,I28061,I24594,g9407,g30306,g26738,I26006,I24655,g4347,g23801,g30104,g5385,g16860,g20923,g25123,g12537,g29327,g6776,g1861,g3996,g27082,g13101,g27384,g15785,g10038,I38151,g24256,I16900,g20331,I31082,g5684,g23566,g22686,g22319,g27580,g12249,I25246,g22440,g28154,g22674,g10534,g18833,g26473,g453,I36708,g1657,I39635,g29559,I34749,g19027,g15615,I31649,g23156,g2240,g27117,g10226,g15516,I30272,g13648,g16201,g1618,I39276,g12782,g6519,g17059,g23164,g26307,g29074,I27083,g30939,g6170,g6675,g1954,I24399,g21843,g17527,I18191,g23461,g30494,g24844,I17919,g11315,g27268,g30989,g11651,g28064,g12781,g8360,g18552,g20617,I23791,g27200,g10352,g14668,g26525,I13896,g1894,g24687,g29347,g30317,g21225,g11562,g21920,g29663,g3133,g1944,g13576,I15472,g23089,g15151,g30851,g9034,g16692,g24273,g27042,I37629,I26266,I31520,g12106,g2318,g28277,g23670,g11985,g26433,I36291,g23709,I22676,I18479,g25776,I38229,I38878,g22473,g10403,I24158,g27207,g30539,g21580,g4979,g16970,g13943,g28892,g4121,I32626,g19224,I38692,g21661,I13962,g13645,g8693,g29410,I40495,g3978,g2389,g22276,g26237,g30508,I29323,g2800,g20780,g20479,I16012,I22752,g27655,I34238,g24122,g2429,g29444,I28564,g13817,g27142,g24014,g30482,I28027,g28334,I39151,g4882,g26697,g11919,I38321,g30905,g21522,g23410,g8748,g28726,g8026,g19603,g30962,g18846,g16229,g25375,I28314,g15846,I15192,g15506,g4725,g12160,I15499,I26892,I26651,g28909,g2339,g13669,g19095,I23941,g25796,g2115,g30734,g1546,g4475,g15618,I14134,I40075,g8974,g14062,g6188,g25877,g12442,I38863,g18286,g1294,g545,g20561,I18226,I34473,g16120,g28975,g26326,I22136,g26172,g14259,I21127,g2088,g24148,g753,g19229,g8524,g15848,g26450,I23982,g580,g629,I14402,g25378,I40504,g20177,g21094,g27408,g6054,g8892,g1319,g3083,g7897,g14573,I33676,g30854,g11761,g16119,I27755,g23439,g6145,g13649,g1125,g28855,g12434,g25109,g29177,g20374,g4951,g18867,g4035,g20424,g7538,I24966,g20526,g12453,I28051,g23453,g16451,g22185,g29930,g30022,g9756,g19902,I23123,I26612,I36234,I39770,g9787,g26188,g6945,g28751,g4632,I29019,I36063,g6305,g27489,I38172,g26751,I39550,g17348,g13581,I24689,g26690,I37116,I28450,g26312,I22990,g15474,g28527,g4376,I37796,I25691,g25341,g28286,g19925,g30554,g25793,I34241,I36411,I19563,g21528,I40176,g17988,g15274,g8123,g30130,g16616,g16575,g20184,I25399,g18966,I18347,g8431,g10556,I14052,g16036,I21632,g2106,g10808,g730,I32402,g9925,I18838,I32871,g2878,g20629,g22825,g8059,g12875,I25114,g21277,g17554,I21888,g8666,g14849,g23634,g25758,g3410,g10433,g1245,g25372,g8898,g13978,g22954,g26901,g12432,g29331,g22763,g30628,g10351,g17974,g19281,I21178,I18211,g19862,g1866,g24899,I31946,I27146,g12951,g22826,I18332,I40131,g13009,g12844,g28262,g9109,g21820,g4976,g24799,g8245,g21490,g17278,I20744,g25253,g15828,g4885,g10325,g16359,g1084,I26354,g1877,g23172,I38166,g20123,g27157,g19761,g6037,g14205,g12437,I23368,g17062,I17228,I18088,I24214,g29282,g21000,g16291,g30724,I31631,g10862,g1202,I32267,I22973,I38175,g29369,g22400,g7303,I38695,g21096,g13589,g20687,g27431,g10013,g17366,g24528,g10353,g17707,I31712,I22587,g145,g29179,g10288,g28396,g17989,g23009,g27730,I32710,I21897,g23248,I27158,I37815,g2010,g15572,g21128,g27238,g18415,I30146,g22756,g22123,I25549,g5176,g30805,g2584,g21643,g21033,g2972,g30802,I41012,g6978,I37481,I23501,g26568,I38032,I36945,g28764,g7580,g27977,g4266,g20452,g30069,g16200,g21618,g8287,g26493,I37906,g25158,g12041,g30581,g6036,g26663,I13974,g5905,g27263,I35930,g2397,g15701,g22934,I41114,I32116,g16251,g1535,I21246,I27250,g16197,I27167,I28031,I30302,g25419,g26987,I34977,g6163,g29111,g30374,g15106,g11898,g26021,g29306,g10974,g27492,g13123,g1859,g20728,g2120,g20624,g30845,g27692,g1533,g29298,g19905,g21217,g8972,g4696,g19637,g10890,g28882,g23039,I36108,g5552,g21049,g10496,g13125,g25507,I31703,g14374,g30458,g10848,I34971,g30310,g19691,g17082,I38674,I29582,g5201,g1701,g2214,I27785,g17175,g22054,I30377,I30686,g21283,g22705,g1396,g1266,I16556,g16879,I37656,g30443,g5546,I14860,g1860,g7426,g29176,I36752,g9076,g22005,g30831,I27098,g15204,I33415,I15629,g23722,g30467,g10299,g23257,g5081,I18323,g25031,g22166,g22915,I25751,g11629,g27183,g19722,g26354,g24369,g26569,g30853,g29365,I40447,I38258,g22557,g23578,g28405,g3999,g18811,I37508,g16910,g5512,I33312,g25453,I23329,I13179,g29377,g26590,I22063,g14766,g6294,I19345,g30585,I37323,g509,g18753,I35512,g11624,g22252,g16416,g2659,g617,I33708,I40769,g1194,g12024,g12560,g21757,g29756,g30372,I28126,g15679,g22560,g8468,g12148,g21655,g30866,g29039,I26078,I40459,g28380,g28906,g19001,g25691,g27301,g29049,g23282,I32940,g20956,g8770,g22282,g29938,g11166,g15681,g15574,g30101,I27104,g30651,I13095,g19287,g30540,g11586,g18861,g14144,g25451,g26107,g27981,g7819,I29606,I40889,g10691,I25047,I15463,I30838,g1832,g23096,g23800,g1753,I37928,g29394,g22287,g30670,g8172,g2147,g4044,g4592,g8525,g20389,g20416,g22030,g1545,g2644,g9931,g21007,I38046,g18877,g27236,I24530,g5304,I38722,g22665,I21855,g4824,I18281,g10843,g21959,g8907,g14024,g8159,g20369,g3049,g2775,g8933,g27261,g21681,g19430,I33885,g19189,g18647,g25720,g8523,g1911,g4963,g29748,g15351,g8498,g2714,g28256,g27302,g27213,g4606,g18984,g18997,g30942,g26348,g27518,g11702,g19309,g28069,g20131,g10961,g25077,g21006,g29016,I14973,g15942,g24323,g25814,g29759,g28284,g25273,I24427,I20541,g27176,g1735,g30758,g23668,g26068,I26340,I29154,I16741,g23400,g27964,I20604,I33570,I18235,g24114,g25230,g30219,g5970,I20410,I14502,g3304,g24929,g10931,g19914,I15239,g12332,g12392,I25492,g25037,g17028,g12456,I29183,g8385,g13588,I40478,g30716,g19602,g10599,g24375,g13272,g24339,I14559,I23658,g24823,I29712,g23824,I36960,g19773,I31757,g14724,g25234,I40185,g23266,I27218,g24596,I27110,I15457,g30401,g25668,g10125,g11931,g17138,g22242,I24725,g21222,g22785,I30611,I36123,g28833,I26567,I18584,g27865,I24091,I40664,g21270,g28836,g29915,g21360,I16276,I36486,g8303,g30500,g24810,g22615,g26821,g13128,I20517,g27683,g19753,g27987,g7996,g15922,I23754,I21852,g4217,g28166,I32624,g22648,g487,I23742,g13702,g15350,g23818,g4930,g11557,I32931,g23025,g10370,g14811,g15338,g26626,I37920,I24235,I29304,g3114,I19569,I14839,g25013,I37596,g23719,g4380,g9229,I37164,g24575,I26231,I19226,g5362,g26632,g29916,g12295,g10839,g21606,g581,I25111,g26249,g4110,g17142,g4743,g15913,g17363,g28438,g20044,I23513,I20414,g19805,g27698,g1846,I25880,g28978,I22886,g28716,g13562,g21947,I18665,g5851,I13182,g26084,g2384,g27513,I32181,g15336,g25311,g10581,g23056,g29113,g2424,g28949,I25913,I23208,g27086,g12768,g30275,I27705,g12232,g29921,g464,g26722,g28384,g163,g23556,I26571,I29741,g2345,g10593,I39360,g16559,g23197,g25882,g27727,g9465,g18970,g16028,g25309,g21518,g19927,I24710,g18295,g15791,g2533,g29294,g25798,g5141,g1075,I22775,g8160,I39160,g10021,g9811,g24736,I18070,g28248,g29342,g11556,g24410,g10541,g20538,g23112,g27470,g19319,g1193,g10847,g27486,g27272,I18698,g16053,g5927,g11148,I29320,I30763,g17695,g1326,g5330,g12077,I30870,g26258,g4357,I16677,g23484,g6018,g157,I36786,I18719,I28765,g12955,g16432,g23144,g2456,g8191,I32857,g28217,g19449,I19667,g22757,g23195,I31302,g11085,I29442,I17740,g10440,g8293,g23028,I30648,g19347,I18368,g22694,I27772,g30143,g11867,I31709,g10276,g6630,I30080,g27177,g2774,g16033,g25050,g10384,I30735,g7899,g579,g17871,g9965,g26604,g5983,g10302,g1908,I18073,g13054,I14647,g23772,g11495,I31898,g19210,g29019,g15900,g13561,g8497,I36493,g5320,g17094,g26365,g22788,g5216,I21165,g24073,g4147,g29996,g21054,g11935,g23524,I34153,g29514,I34854,g3247,g13901,g5720,g26694,g25168,I28019,g28727,I26357,I22019,g16832,g30561,I29912,g11832,g18629,I23701,I15932,g11120,g299,I15822,I17957,I15369,I21936,I30389,g10703,g384,I13925,g2224,g12063,g7591,g29149,g12959,g16447,g12460,g29721,g27529,g8284,I22509,g30713,I31838,g28579,g25700,I36327,g21715,g25941,g13787,g25993,g26096,g25136,g17360,I23358,g4453,g25224,I23564,I27920,g15869,I25456,I27711,g25619,g19519,g13859,g27552,I38396,g24324,g5113,g13171,g1204,g13573,I40850,g29772,g30882,g821,g2495,I34102,g30490,g18875,g20842,g15740,I25712,I39246,I38272,g9423,I23673,g28245,g30299,g26130,g1931,I36684,g28199,g19355,g21032,g3065,g25027,I27391,g10377,I34071,I35554,g11441,I27086,g13324,g24497,g13504,g19781,g2593,g3248,g602,I27388,g21158,g24945,I24346,g24167,I36999,g6197,I32687,g24857,g8879,I24125,I23570,g1196,g22824,g24633,g7837,g15049,g20089,g19893,I15964,g11976,g22738,g7872,g24864,I25733,g29497,I27116,g1421,g11766,g10710,g2805,g20051,g15480,g13248,g16694,g10357,g28578,g21954,g21900,g20679,g25046,g30943,g20558,g7688,I31526,I35031,g10727,g28654,g26036,I23785,g26885,g10498,g26171,g13620,g11496,g945,g15520,I40257,g12502,g29849,g24897,g27080,g23403,g26315,g26886,I37140,g566,g27413,g29343,g24852,g16027,g26038,g27530,g27827,g7336,g13945,g16186,g27765,g1948,I33974,I35494,g20519,I19829,I25731,I30356,g22585,g4162,g28240,g23901,g486,I14584,g1760,I19342,g13413,g10330,g24149,g21687,g20766,g27682,g15438,I30869,g25155,g15889,g8472,g29946,g1937,I36939,g358,g29873,g29341,g24257,g14309,g19301,g24548,g24801,I40260,g12992,I14535,g29437,I19516,g700,g5279,g28363,g5649,g20053,I29622,I38524,g22013,g15631,g13819,I33813,g26530,g9487,I25300,g20969,I31274,I25782,g11022,g15052,g13140,I16714,g27691,g12801,I26846,g11770,g16455,g15573,g26807,g3010,I29262,I23309,g13524,g25825,g19383,g23564,g29198,g19306,g8397,g30267,g3922,g343,g12009,I18019,I23234,g11612,g19688,g2221,g18567,g4674,g4314,g11684,g28880,g10048,g12098,g17372,g22187,I25831,g22645,g21481,g1410,g24581,g21866,g22149,g699,I31670,g19547,g25057,I36924,g25335,g17156,g19063,I18356,I23364,g20400,g10485,g15246,I29872,g8535,g8559,I25123,g10095,g30958,I25540,g2114,g12102,g17351,I20568,g16414,g26910,g1158,g10457,g28695,g13040,g490,g4611,I39258,g30000,I16958,I39767,g9104,I13143,g11590,g12349,g14086,g29485,g20021,I37324,g3124,g3493,g22105,g27690,g2432,g21371,g25199,g30309,g27234,I33154,g11277,g16063,I38080,g25169,g30035,g11776,g30718,g19667,g369,g30927,g29385,g20877,g2539,g16998,g25706,g10555,g17814,g29434,g13507,I37846,g27719,g21024,g8971,g5159,g8997,g15332,g27022,I34469,g2351,I40303,g1316,g28404,I13104,g29622,g20944,I25081,g20327,g8414,g10055,g5845,I18452,g9884,g13410,I16338,g10439,g7763,I20863,g12224,I34099,g22089,I38975,g19559,I16107,I40587,I36978,g22771,I21629,g1529,I21736,g4225,g27713,g2546,g19983,g19978,g10396,g21921,g6046,g8566,I22536,g27104,g14390,I36138,g22903,I29506,g23459,I31235,g27994,I37032,g6293,g13278,I15680,g1680,I33321,g4684,I30290,g974,I32164,g27123,g4444,I29924,I38609,g26681,g30017,g13462,I16047,I39050,I21595,g5768,g24487,g27942,g5857,g5150,I15839,g30260,g24012,I18113,g19067,g24113,g29695,g1775,g831,I29145,g26164,g15811,g16386,g30697,I34124,g25244,g11534,g23245,g11344,g13952,g29581,g11617,I35678,g10382,I24656,I36659,g9341,g24352,I17762,g11348,g16006,g10868,g287,I15626,g12175,g26506,I40928,g15879,g29538,g22715,g19549,g16264,g25351,g8622,I17966,g1731,g222,I30994,g26216,g19598,g25211,g26293,g16322,g27449,g1768,I27029,g29569,I17527,g722,g9242,g28014,g18652,I13937,g28767,g10263,g18277,g1092,I30311,g17570,g30859,g12108,I25096,I19921,I34734,I38731,I25838,g29156,I30617,g22358,g13048,g17307,g21899,I40988,g22274,g21077,I19733,g30587,g24124,I38125,g25708,g15741,I21989,g21721,I20100,I38378,g11095,g24209,I30386,g972,g25938,g29337,I34505,g28281,I37295,I18740,g29001,g5283,g10379,g20457,g2100,g12883,g29157,I24092,g12174,g26386,g3102,g8493,g29788,g12270,g11450,g22142,g7162,g30666,g24272,g30132,g28987,g11216,g27755,I14529,g2451,I17363,I31817,g26914,g20644,g1807,I34833,g4165,g21244,g5862,I14842,I20670,g18927,g21349,g7420,g25470,g4772,I15975,g19546,g5740,g26131,I39008,g22217,I33300,I21918,I13236,I27311,I39255,g28458,I24696,g30573,g17540,g18667,g26441,g16985,I23676,g30800,g5156,I14357,I30679,I29162,g1582,I18777,g13436,g30365,g28402,I27095,g22305,g30932,g25699,g22603,g1679,g5689,g25764,g28391,g6086,g19245,g19125,g24664,g20611,g23612,g23583,g417,g30261,g23554,g29507,g10670,I23854,g13285,g26414,I32696,g29636,g984,I15267,g28409,g13432,g16470,g28473,g26003,g30961,g14008,g29362,g12378,g6232,g8403,g23559,I24053,I29277,I33580,I28978,g12454,I14219,g28259,g24751,g29046,I17712,g23297,g5874,g7879,g21851,g4535,I37880,g11611,g16905,g2097,g13034,I18175,g16034,g17573,g24893,g23871,g24577,g27337,g24842,I23542,g17990,g22984,I25923,g10991,g20640,g20893,g24386,I15995,g1804,g10060,g24326,g28387,g17111,g8437,g24424,g29438,g4092,I18623,g13855,g23325,g28526,g12114,g554,g22292,g24242,g15756,g28169,g13418,g19055,g20619,I36280,g30935,g29563,g21380,g4338,g23427,g8526,g30237,g258,g2380,I25213,g28554,g24143,I40125,I24409,I36120,g12942,g5920,g21885,g26593,I21838,g23999,I20601,g7263,g5975,g19033,g17020,g19675,g20352,g2929,g25536,g10573,g2248,g23277,I31115,g20830,I33891,g2615,I32479,g15644,I15526,g11889,I20574,I21878,g19094,g27729,g16996,g21447,I38071,I18854,g17774,g17764,I30035,g7953,g19679,I15535,g18857,g11943,g21340,g26657,g25331,I33501,g10292,I15429,g11274,g19746,I13218,g30218,g25943,g19307,g16497,g15220,g20405,g8333,I21271,g19212,I35446,I25283,g5818,I26464,g11123,I19025,g10192,I33307,g30151,g22709,I33405,g10479,g7595,g12153,I28503,I38499,g13447,I28743,I35064,g18324,g18850,I20483,g23827,g6783,g5980,g29240,g27574,g5737,g17685,g24682,I27822,g26052,g16739,g29187,g26855,g9050,g22789,I24567,g28748,g25615,g19267,g28881,g1724,g10788,g1045,I18780,g13836,I32309,g5389,g548,g25566,g27174,g15222,g28699,I19549,I29906,I18857,g20655,I31664,g24211,g10834,g19109,g20052,g27541,g27164,g18231,I23983,I30791,g29925,g30880,I34195,I35837,g10735,g7642,g26083,g11243,I33013,g12157,g7606,g16494,I16438,g4015,g19154,g23550,I35376,g10402,g10415,g19090,g26950,g22169,g16282,g29449,g5469,g5933,g28100,g29267,g2504,g20662,g16385,g21422,g17508,I23794,I28000,I34358,g26849,g27570,I19621,g24095,g19596,g12211,I38474,g30602,g2253,I38947,I24474,g8906,I37291,I24613,g26033,g17541,g10371,I16241,g22592,g19553,g28671,g26432,I15304,g30711,g27984,g27785,I38128,g8938,g3046,g24797,g22530,g9140,g29391,I24753,g20652,I27419,I15238,g10076,g13103,g5700,g25021,g29981,g7685,g19557,g28721,g1423,g21813,g11543,g11572,g21593,g29334,g596,g13394,g6153,I37020,g12829,g28437,I29841,g477,g16003,I16700,g1615,I35067,g30093,g28025,g8949,I19303,I40763,g29975,g23953,g3056,I23545,g30793,g19681,g21764,g26299,g22591,I29569,I31604,g19739,g29188,g14177,g17057,I31205,g24486,I15833,g29922,g5416,I20334,I34296,g27927,g30468,I38220,g2934,g237,g17135,g20112,g10007,g24249,g26971,g24290,g14497,g27604,g10171,g15817,g29537,g23200,g8617,g22263,g20054,g4142,g2225,g25749,I28090,g24425,g25821,g19564,g4545,g7622,g21819,I32443,g21411,g13396,g26145,g30701,g17015,g12139,g9919,g14507,g30531,g28453,g25350,g25937,I37497,g18688,I36731,I33343,g4398,I37146,g14963,g28219,g5312,I23782,I19479,g20940,I23415,g30217,g29775,g3072,I28247,g10661,g29562,g576,g411,g22839,g28746,g11857,g18236,g13958,g26039,g25362,g23222,I31775,I15983,g22183,g23468,I38854,I24894,g5639,g19249,g19211,I21277,g12377,g20310,I37736,g4136,g27245,g7009,g2583,g29829,g29162,g20809,g10284,I32934,g25886,g4211,g23113,g3055,g26208,g12007,g26648,g27339,g8486,g507,g28273,I39541,g20953,g12115,g22237,g16969,g24435,g24398,g17192,g26092,g10967,g3191,g19046,I27827,I32988,g17318,g5275,g3070,I27089,g26150,g8779,I23611,g15172,g2526,g26213,g20819,g22540,g19790,g13559,g19417,I32561,g1122,g11004,g5811,g7342,g15809,g28383,g18844,g1439,g22286,g17588,g21602,I14066,g24060,g6435,g8354,I36465,g8330,I29040,g26209,I37608,g16082,I14014,g26207,g7875,g30675,g29281,I40775,g24811,g28270,I27080,g19020,g18431,g24340,g8980,g20337,I37729,g22899,g30785,g7488,I22560,I25862,g25248,g24898,I26871,g29390,I23029,g5976,g10478,g19720,g4159,g16995,g11603,g9463,I23976,g22425,g5333,g8197,I29052,g28848,g29548,I25162,g30766,I29070,g5894,I28318,g405,g26020,g22799,g29268,g17479,g11952,g5107,g23065,g9757,g10158,I19877,g12099,I40691,g8774,g26358,g13087,g1836,I40559,g22838,g4692,I25605,g18469,I16653,g12293,g11616,g19456,g1952,g24266,I39797,g28760,g15492,g23324,g27359,g27465,g22749,I31931,g18935,g26687,g25161,g5790,g18975,g4994,g11717,I26171,g30062,g15820,g13150,g21569,g13154,g20805,I15955,g29152,g18174,g29650,I35926,I21974,g21350,g5717,I30997,I18001,g1939,g5123,I19631,g3650,g13997,g22112,I21720,g10492,g30945,g12967,g4118,g5315,g20114,I15565,g3773,I19862,g20343,g27949,g29659,g6678,g10012,g27538,g11036,I13221,g11502,I38181,g13111,g17859,g16007,g26257,g23842,g27061,g25332,g3139,g29607,I25783,g29679,g25131,g12900,I37599,I15543,I28335,I33909,g30582,I15890,g22599,g20608,g12116,g27313,g4735,g20120,g16596,g11949,I23689,g26561,g11376,g7539,I22512,g23848,I32284,I41038,g19797,g1738,g22228,I38369,I38038,g10470,g11875,g11910,g11652,g30558,g23687,g18358,I25672,g22726,g26270,g4763,g28477,g23454,I30483,g30915,g14606,g12530,I31056,g5199,g11678,g19260,g16953,g18808,g26160,I39157,g25824,g24144,I33205,g25163,g7484,I15986,I23524,I33385,g29102,g28785,g27784,g8856,I22663,g10283,g20412,I29500,g423,I27585,I25557,g17566,g27237,I33798,I21982,g11564,I34159,g20335,g11508,g17901,g3969,I20429,g16850,g25371,g1704,g18974,g13239,g25216,g27586,g15810,g16068,g1855,I32604,g30342,I30623,g19165,I28432,g8252,g29271,g29153,I29519,g24320,g21326,I32470,I18010,I29465,I36800,g16421,I29619,g2966,g12053,g20833,I27949,g2245,g22381,I32419,g249,I36693,g21192,g25140,g26292,g23335,g23673,g23015,g1036,I23445,I36792,g20990,g22318,g19352,g30938,g2255,I30660,I31655,g9782,I35750,g30722,g24846,g8888,g24792,g19540,g19056,I27134,g16424,g19874,g24279,g15467,g28738,g11574,g29032,I31706,g3554,I36560,g21700,g1667,g30117,g28903,I15882,g18330,g12239,g20351,g18898,I35021,g3981,g14321,g2365,g21619,I35313,g22364,g26362,g12023,g26631,g22398,g7455,I32979,g19650,g23047,g17194,g20928,g25979,g15675,g29459,g9323,g19283,g23276,I22548,g8862,g20413,g19025,g17091,g9790,g26686,g20469,g22412,g21078,g29909,g11205,g29642,g471,g13547,g28123,I14734,g13512,g819,g22729,g13162,g22989,g16324,g15851,g22700,g11491,g27736,g1392,g23832,I33790,g21498,I40703,g4498,I28467,g16017,I15553,g28040,I31820,I14868,g25389,g15899,g6136,I16961,g20478,g13316,g16313,I32159,g28804,g4395,I18578,g19500,I20465,g9216,I15167,g1670,g11519,I30149,g18096,g18130,g22181,g12187,g24858,g29914,g24255,I24401,g18654,g19655,g29911,I35283,g30828,I25489,I35741,g2656,g26864,I18169,g6048,g24555,g13356,g28672,I37768,g286,I22683,g6838,I37319,g1180,g30550,g16055,g21467,g17877,g27401,g30262,g26673,g2502,g7349,g10949,g10524,g12152,I15992,g21081,g27118,g19451,I31490,g2796,g12245,g19276,g30491,I29366,g10434,g16223,g24133,g17991,g2604,I20820,g29488,g19118,g20577,g18637,I22630,g25181,g17979,I30470,I30323,g27191,g26813,g29687,I18265,I30547,I34388,I28380,g23570,g30207,g1141,g6943,I37098,g28326,g13736,g29989,I28137,g28348,g30302,g27882,g19729,I22569,g12026,I35482,I40694,I40751,g21446,g22610,g25772,g22057,g29726,g29128,g14677,g29376,g24950,g10036,g16342,g8478,g24055,g4754,I37991,g201,I34839,g19121,g16024,g28354,g26212,g26324,g29290,g22103,I25534,g30324,g28247,g25861,I18677,g767,g23290,g11659,g3244,I39243,g12088,I14763,g9354,g17272,g15786,g12233,g27072,g12916,g7192,I30878,g3018,g15783,g29404,g11398,g23316,I38951,I16328,g1603,I36741,g5868,g27227,I16811,I25219,I28972,g2092,g18678,g8,g18618,I21420,g27717,g14884,I13194,g13108,I22062,I38386,g26627,g21576,g74,g26787,g25355,g26047,g30052,g1538,g17551,g20760,g4501,g24711,g13408,g26335,g5297,g8469,I33627,g23545,g15804,g28301,g25841,I39053,g9773,g10314,I31844,g19589,g2447,g18856,g10764,g27187,I30589,I39026,g24476,g13374,g9582,I13316,g2478,g13137,I25643,g1828,g17950,g19853,g22704,g19676,I37083,g27603,g11608,g27300,g19255,g29653,g25643,g19741,I22926,g13599,I15645,I24582,g23512,g27144,g28442,g659,g30871,g26675,g27267,g29379,I22937,g25210,g23711,g23059,g8482,I34198,g5727,g24882,g12097,I33495,g30930,g1966,g11591,I24459,g22900,I26497,g25301,g20936,g25697,I24703,g13608,g5912,g22075,g18201,g21939,g4298,g13456,g5403,g20246,g141,g26609,g18265,g10506,g29910,g13478,g14776,g18058,g23560,I22810,g28170,g10398,g23910,g25048,g20879,g28044,g10829,g10123,g325,g630,g2080,g3062,g9400,I30341,I18429,I14888,I17816,g16647,g8934,g29629,g26874,g24550,g30777,I19318,g30646,I31487,g27906,g20979,g30878,g1167,g1567,I18408,I31787,I22611,g11883,I34921,g1904,g26623,g23572,g30120,g26643,g13192,g5709,g21622,g1910,g12934,g15698,g9260,I30480,g26805,g28211,I17945,g21863,g25954,g29960,g20222,I27179,g18849,g24234,I19813,g1683,g2598,g28450,g30272,g26363,g24077,I23775,g20025,g11011,g402,g10297,g29130,g2861,I19624,g564,g24395,g15182,g11942,g12071,g2251,I35727,I20836,I32913,g45,I26276,g16566,g10987,g13186,I38548,I34220,g5372,I34743,g23776,g983,g2238,g4188,g4848,g28073,I39386,g20304,g9891,I37986,g27179,g14767,g28826,g2734,g8544,g24579,I32688,g21138,g1852,g25443,g20972,g13091,g21913,I15549,g20355,g12207,g21631,g21319,g28931,g29503,g29242,I26541,g5408,g23954,g13025,I31159,I36102,g30544,g29539,g17228,g15833,I24265,g29322,I39267,g23093,I36545,I16344,I16018,g28071,g2867,g5939,g10424,g22206,g7329,g22723,g11170,g9506,I33673,g18547,I13775,g18337,g7812,I22763,I38851,I36052,I14002,g22216,I21769,I33278,I37107,I39866,I20538,g19713,g10932,g16112,I19767,g18314,g16420,I26966,g8719,g26434,g856,g23878,I27264,g1762,g156,g12094,g14183,g25995,g26647,g26735,I19615,g17099,g7581,I40248,g21300,I14538,g29710,g13208,g19048,I31517,g26625,g24244,g2264,g25005,g13426,g30343,g20363,I22998,g1964,g18063,g21303,g22448,g27555,g4409,g4375,I37074,g8726,g26028,g4404,g15412,g26534,g22332,I36639,g13974,g22116,g131,g5638,g1430,g5358,g27621,g30081,g22711,I20355,I35708,g1606,g28287,g16984,I16763,g23141,g3076,g28724,g16335,g23125,g11028,g29984,I40721,g4595,g2079,I22518,g24065,I18527,I35053,g22796,I16744,g26858,g19259,g17637,g20061,g20918,g27481,I23917,g11728,I24178,g29135,g11911,g15442,g18988,g21193,g19490,g26333,g29626,g25947,g30979,g8654,I40589,g12472,g11703,g27386,I21340,g3365,I35413,g30323,g1230,g4278,I28248,g25999,g22942,I16987,g21811,I16476,g11490,g15729,g11814,g20287,g5880,g1139,g1988,g29798,g3522,g1801,g8877,g11869,g23568,g18907,g23046,g25008,g16347,g21944,g17912,g30874,g61,g20630,g21074,g9058,g22754,I13950,g8780,g30106,g19872,g18598,g25561,I29226,g15876,g366,g22437,I23622,g8487,g10093,I25459,g19178,I26535,g14079,g9439,g30545,I17151,g23087,g28523,g1633,I26819,I25084,g16309,g20403,I32708,g27526,g8511,g30978,g3123,g20776,I27695,g1110,g2959,g26938,g30485,g28117,g21043,I30350,g26583,g25963,g7673,g23240,g6310,I35993,g29617,g13023,g22679,g15502,I32633,g20463,g13404,g4433,g18939,I26334,g22215,g8388,g25454,g785,g8500,g30367,g18334,I32609,g22031,I30152,g9095,g29558,g29412,g12250,g20880,g4023,I27352,g16991,g22512,g15822,g3928,g21678,I29421,I38068,g13883,I16990,g25147,g13863,g23385,g21148,g1012,g11597,g25827,g13861,I28100,g8421,g29457,g28461,g19322,I40802,g18865,g21087,g9116,g21972,g30245,I20586,I29579,g4231,I33596,g2870,I36490,I19404,I17819,g29392,I34815,g24474,g28355,g976,g13273,g22795,I39832,g16894,I28219,g13610,I30766,g23368,I22789,I14612,g28611,g18561,g26865,I23395,I33498,g5967,g22255,I40874,I18274,g9662,I32411,g879,g8169,g10203,g12318,g10204,g12081,g551,g26601,g15264,I33726,g10430,g12837,g19755,I24300,g19216,I18689,g24399,g16052,g10112,g18169,g25318,g2746,g29660,g27028,I19557,g7919,g20124,g26824,g27426,g11959,g12962,g6142,I13089,I40581,I32074,g4372,g13044,g28027,g15534,g8056,I17984,g12305,I31559,I28272,g24409,I32120,g18281,g8928,g13882,g16823,I23729,g18839,g11725,I22786,g4139,g22200,g22055,g22258,I23093,I31613,g16778,g8075,g4354,I27203,I36676,g12443,g1798,I26667,g2808,g19047,g10574,I40832,g13527,I29408,g30013,g28471,g5593,g26144,g24421,g7143,g17080,g24111,I29333,g24384,g13062,g21108,g27716,g1524,g19734,g10514,I22866,g19900,g5382,g9758,I40438,g15283,g18390,g27139,g1345,I20646,g14609,g29384,g19723,I23460,g508,g16358,g6512,g24071,I14811,I18220,I30179,g18948,I20479,I15677,g13210,I38122,g30082,g20658,g6039,g29133,g14413,g25669,I16347,g12471,I39622,g13880,I37011,g25755,g20477,g27756,g9749,g29005,g17591,g21119,g2107,g26385,g25630,g16608,g27318,I28491,g2207,I38077,g9905,g20459,g11576,g27341,I25660,g19170,g12369,g15794,g4665,g15435,g16242,I38689,g21161,g26711,g19285,g26059,g17697,g6298,g10333,g22211,g24096,g27,g21327,g11240,g1579,g3053,g20707,I27343,g13636,g21766,g27212,I27026,I27372,g30078,I41093,g5974,g7691,g24540,g10522,g30925,g28186,g17157,g20806,I23851,I30639,g5217,g24975,g28431,I27868,g20590,g28447,g27353,g3127,I18329,g12991,g23791,g558,g16419,g30636,g26737,I32320,g10157,I38339,I24280,I26337,g18847,I24382,g21647,g19730,I25866,g30723,g9585,g24416,g15385,g13703,g27733,I33888,g12899,g13878,g3040,I20299,g19588,I15998,I20493,g12426,I17875,I22599,g2990,I30044,g11447,g19640,I40973,I36918,g21311,g27330,g10706,g11693,g11222,g25212,g4175,I18990,g22732,g16369,g737,g18882,g9196,I31556,g3566,I13107,g10977,g17079,g21860,g2379,I35937,g30495,g25445,g10508,g2094,I39130,g13381,g12036,g5756,I21962,g6836,g30058,I27164,g29220,I25442,g29818,g7924,g5601,g10773,I24718,g24742,g5263,g28223,g25047,I15490,g17128,g28074,g5808,g15325,g29325,g8659,g24382,g23349,g11726,g28006,g28634,g17225,g26357,I36367,I36930,g25426,g18915,g25218,g22415,g8572,g7475,g5685,g24129,g27768,g16381,g2781,I40086,g16881,g1408,I36521,g27992,g25062,g27904,g23477,g18868,g25338,g12455,g6486,g387,g25732,g3722,g12326,g1248,g15221,g12775,g21654,I38848,I15245,g16043,g7727,g15126,g24427,I39059,g11138,I36337,g17413,g9145,g10921,g1517,g5718,I22726,I30059,I30800,I18204,g19247,g17229,g26479,g16152,g15858,g23820,g20917,I23279,g22152,g1496,g30279,I23256,g27097,I22025,g24788,g17017,I37644,g27173,I18791,g17627,I38999,g1041,g454,g13892,g5809,g7792,g23675,g19789,g21085,I23769,g25137,I33855,g25457,g16488,g27189,g12874,g28750,I22981,g30893,g11708,g29633,I23094,g13147,g728,I37760,g12518,g14329,g30356,g8099,I29165,g26381,g24695,I25606,g26438,g13490,g12825,I27137,g28362,g873,g30659,g9367,g29256,g29333,g5941,g29192,g698,g14580,I23451,g21056,g9083,g23133,g20394,g29861,g25154,g30918,g18503,g2117,g4104,g21338,g1104,g13501,g5877,g24735,g14883,g22311,g28009,I27300,I40218,g30715,I23243,g19668,g15710,g18959,I24144,g19190,g25219,g9084,g19696,g17631,g19261,g28595,I35428,g15376,I38184,g13220,g13227,g13969,g4740,g20433,g11505,I38755,g9922,g9711,g11545,g26217,g28762,g18691,I35355,I20421,I26528,g27989,g14061,g28200,g10480,g12124,g28940,g21034,g22850,g30884,g10404,g24276,I31724,I17209,g26780,g11565,I25463,I27308,g28923,g17217,g29172,g7521,g3047,g23117,g10662,g19635,g5286,g10152,g15423,I27658,I36450,I16267,g19192,g16913,g12915,g22470,I31937,I35686,g16010,g25412,I14644,g28659,I24545,I19482,g27037,g21529,g10114,g30349,g30313,g22710,g29498,I23457,I25939,g13332,g5363,g15821,g13631,g1835,g30702,g19186,g11428,g25729,g27092,g21699,g574,g29230,g14797,g1148,g23567,g3112,g29783,g1967,g25085,g5655,I23866,g25361,g16665,g26586,g7724,I30089,g8506,I28464,g29108,I35868,g23340,g12089,g11865,g29481,g8952,g11063,g17136,I34230,g21147,g6139,g21682,g24511,g17321,g6024,g11636,g12418,g26881,g26736,g11569,I16150,g23940,I30287,g15602,g21313,g19530,g5233,I35351,g16171,I38807,g14327,g9518,g357,g29277,g10198,g16614,I15244,g11939,g22684,g17530,I31859,I14249,g11697,g11742,I26593,g20311,g28448,g25339,g18940,g12744,g12830,g2839,I34083,I25994,g29131,I27243,g22638,g2388,g25195,I33260,g2085,g7613,g5748,I21705,g17090,g10201,g24329,g4591,g13232,g21026,I33545,g19286,g2440,g171,g840,g25153,g1842,g2782,I39011,g16480,g7333,g22793,g28717,g15375,g19798,I26627,g26445,g20998,g27662,g27051,g5132,I36240,g5806,g28208,g22177,g13051,g21859,g20486,g27356,g5913,I30504,I30757,g9673,g20278,g16106,g9371,g13926,g3126,g17310,g27081,g1405,g5033,I39469,g843,g11661,g11621,g17291,I40910,g19173,g17430,I20694,I38111,g17302,g23496,g17345,I22963,I15256,I25177,g16240,g16468,g309,I13919,g4614,g3109,g28935,g8407,g18804,I28162,g30737,g8561,g5269,g13484,g19945,g28318,g9531,g10456,g20367,I13953,g10174,I25762,I23057,g2195,I24764,I20616,g21345,g30528,g15920,g17754,g13159,I40724,g15750,g8690,g21367,I21256,I40745,I32659,I28152,I39690,g19769,g10549,g19915,I14149,g30689,g19152,g28292,g19733,I24763,g7423,g29487,g27764,g3238,g19910,g28850,g7876,g18128,g16632,I25174,g9215,g15133,I15019,I35383,g15352,I15850,g27277,g23150,g23713,g21392,g8509,g23178,g29997,g8501,g12461,I21426,g25247,g12209,g18871,I31721,g27956,g19926,I30914,I16453,I36721,g30987,g13605,g2443,I31736,g8612,g5003,g21751,g4683,I37194,g20454,g2589,g30795,g27111,g24822,g17218,g18950,g29295,g12353,I36702,g9927,g15354,g23232,g1699,g4851,g23159,g30304,g27656,I25840,g27922,I40471,g16132,g10372,g5680,g28823,I13430,I32324,g16357,g14486,I28969,g12922,I19771,I41120,g1135,I36426,g19743,g28291,I34189,g24432,I24577,g36,g22226,g13038,g18548,g16993,g10531,g23058,I40233,g15599,g16431,g30903,g23944,g144,g21169,g23033,I38238,g18307,g13180,g2646,g4587,g5095,g25975,g25589,g153,g364,g2804,g24277,I39142,g22251,g22083,I20458,g24108,g23526,g11554,I37471,g24437,g16475,g21793,I35844,g25228,g19234,g9107,g10222,g27208,I25108,g21573,g28439,g129,g28234,g9443,I33128,g1698,I30143,g8317,I24054,I18148,g27584,g12531,g19193,g20504,g26775,g8327,g10814,g20307,g15641,I19360,g24296,g17016,I24195,I16776,g22641,g14148,g29366,g17442,I40453,g19218,I38235,g16131,g30556,g29476,I35968,g23186,g27547,g19149,g3106,I40149,g8129,g5926,I34461,g21865,g15765,I16044,g26243,g27115,g22461,g15393,g18807,I36441,g4174,g22188,g25475,g17520,g8505,I23670,g30525,g23582,g18519,g17854,g3940,g18707,g5399,g22164,g25549,g30541,I34653,g7462,g8932,I20544,g5958,g9139,g12214,g155,g10389,g12177,I29271,g17270,I29023,I40994,I24648,g25950,I36728,I13146,g15458,I23227,g793,g5991,I18650,I18040,g10869,g18924,I41047,g19944,g20216,I31000,g17049,g5590,g2472,g24769,g10017,g12058,g30441,g13093,g29407,g4561,g10600,I39534,I33355,g23055,g6059,g20102,g15304,g3618,g25320,g24351,I30829,g23790,I30239,g12363,g18796,g16153,g24691,g23142,I20505,g6068,g5238,g30452,g5425,g26320,g26674,I40925,g22291,I21884,g23289,g16045,g19499,g9335,g12308,g22148,g24254,g829,g706,g18140,g24289,g1166,g24627,g23735,g27962,I36141,g13046,g23678,g8246,g15856,g28426,g26102,g14320,I40835,I30544,g28283,g17012,g24588,g19819,g29419,g29828,g963,I27942,I28476,g14558,g29677,g18257,g5404,g7857,I28649,g26693,I14596,g21030,g27820,g18129,g9916,I30516,I22593,g25678,I18449,g29757,g2372,g990,g11800,g22676,I20398,g3107,g11859,g12858,I16144,g22303,g10249,g22606,I31652,g5755,g6058,g23823,g28725,g7748,g28275,g22168,g837,I27035,g4942,g16130,g16254,I29509,I30209,I20810,I18046,g17676,I27969,g9464,g10643,g19243,g23381,g20431,I18097,g939,g27774,g23627,g27206,g29433,I18076,g21907,g27382,g18508,I24662,I31466,g24053,g10707,g26080,g9871,g24366,g20743,I36969,I38205,g20242,g24359,I18817,I36462,g24438,g22021,g21260,g25122,g28253,g11764,I30281,g26959,I38677,g26181,I33529,g26490,I24443,g8539,I14990,I25528,g30782,g18302,g29785,I18022,g9138,g11721,g26688,I27267,g21889,g27161,g16679,g17837,g20882,g19012,g382,g4234,g13325,I37823,I23199,I14951,I28754,I40481,g25746,g11914,g16044,I33636,g10035,g14459,g27047,g11940,g28730,g24885,g26086,g29531,I30769,g19802,g20350,g22629,g27506,g25978,g455,I30905,g4821,g11775,g26998,g7898,I30164,I37858,g26852,g8655,g19024,g26564,g4049,g11599,g24472,g29480,I17150,g22331,g20391,g28107,g13541,I16068,I29030,I13892,I31253,I33662,g703,g27666,I24264,g25258,g5415,g26985,g8517,g4286,g24800,I24123,I17846,g30454,g30032,g26195,g3185,g30436,I16538,I40560,g15670,g13386,g30255,g25178,g29655,g15287,g30246,g8546,g17207,g13614,g20603,g23941,g5658,g7193,g21036,g23768,g5611,g2059,g8474,g19951,g27148,I32527,g16013,g30794,g9302,I39812,g30980,g18520,g30318,g18926,I23888,g30316,g27269,g23051,g29972,g26773,g11509,g19369,g23611,g1588,g20501,g29251,I36213,g11733,g19158,I41035,g3878,g9666,I36217,g5008,I23507,I39376,g2373,g25187,I25915,g10193,g25576,I30692,g28303,g20941,g20221,g26042,I26494,g20302,I19937,g27294,I36032,g1540,g21670,g19225,g12711,g3080,I15938,g2101,g5915,g30183,g13449,g14419,g15921,g26980,I25204,g15055,g19246,g10223,g9722,g25838,g11547,g22985,g28637,g13183,g11723,g5651,g19703,g29381,g17416,g17204,I24640,g4699,g21439,I31925,I17936,g12012,g18341,g11722,g23828,g28430,g10455,g18941,g29035,I19702,g22189,I32401,I21435,g10809,g1520,g30817,I23418,g20884,g21805,g24747,I31901,g14040,g25102,g30131,g14529,g21099,g21658,g29258,g79,g22800,I15213,I37581,I28524,g11568,g22243,g13927,g2806,g16636,g2111,I18647,g22316,g948,g19550,I27346,g14493,g30019,I27101,g13081,g13167,g26202,g10285,g27798,g21953,g13355,I34032,g17507,g30902,I37467,g6141,g30824,g20163,g16520,I19576,g22582,g23662,g12123,g27908,g24213,g29998,g18925,g24358,I27113,g24388,g23714,g8344,g25438,g16923,g1942,I29326,I34411,g8463,g18636,I14544,g23392,I35777,g22832,g4794,I30701,I30854,I34274,I13928,I32726,g15997,g28886,g12836,g12101,g24471,g8183,g12542,g25208,I20117,g8978,g11694,g29415,I34901,g22597,g2217,g10282,g11861,g5812,I18608,I19380,g20164,g5705,g19444,g30643,g2376,I15961,g6025,I22533,I18752,g20414,g24783,g15296,g15021,g17992,g30462,g12145,g25437,I16120,g21028,g8519,g14524,g17258,g1269,g8141,g24228,g30966,g3088,g1262,I15942,g11884,I24428,g28090,g21342,g16418,g29986,I37854,g27738,g10003,g8286,I27984,g12420,g11923,g2288,I35695,g30287,I19271,g15234,I14590,g9342,I22444,g25167,g17604,g25833,I36780,g10453,g18643,g24500,g15360,g18828,g516,g17753,I17043,g8178,g20966,g9114,g27262,I32510,g9665,g8925,I16796,I23000,g13076,g1732,I39377,g25951,g2315,g26300,I15442,g28790,g21790,g29393,I40484,I14459,g12894,g5115,I19787,g20943,g30538,I34449,g21906,g15550,g27348,g24787,I32607,g28501,g29522,g22623,g27133,I21803,g19759,g24246,g15665,g23060,I15329,g13502,g30948,g5799,g8874,g10877,g9422,I18441,I22917,I40420,I18770,g19278,g18952,g22293,g27209,I25578,I24679,g19617,I38881,I28174,g18794,g20954,g5266,I17278,g28367,I41017,g22396,I25665,g23310,g10830,g18200,I30395,I25506,g15356,I18289,I30284,I25664,g1,g13340,I17649,g15949,I25355,g24164,g168,g22922,I20844,g25281,g21723,g294,g23725,I38094,g5428,g20850,I31502,g5227,g1528,g7679,I18749,g23215,I21262,g27504,g29474,g18912,g13185,I26383,I19901,g21536,g25186,g29283,I25819,g3125,g25781,g19562,I32451,g18699,g23161,g29518,g23249,g29801,g26045,I35780,g25996,I36539,g13492,I37426,g6000,g12050,g280,g7605,g12931,g26602,g25201,g19088,g30359,g25417,g28971,g22567,g24104,g29833,g5899,g27907,g19824,I31310,g2185,I23591,g30601,g17710,g18905,g17485,g1786,g24222,g22092,g8101,g8406,I13092,I16469,I25222,g23683,g21234,g23661,g30886,g16595,g19851,g10854,g29560,I38822,g25294,I23772,g4504,g22193,g29144,g21796,g21048,g26691,g27482,g3058,I29110,g26974,g29789,I23695,g25606,g28489,g28216,g8203,g10304,g28021,g30557,g474,I24038,g9309,g24712,g23075,g27293,I37232,I17774,g1865,g27160,g2618,I29990,g27137,I23124,g16429,I17724,g28500,g27381,g29504,I39339,g13264,g13440,g23264,g9634,g13182,I14073,I24532,g28376,g28233,I13578,g17448,g18206,g19204,g12084,I36749,g11672,g4085,g27496,g10872,g28304,g9870,g16481,g584,g27004,g13320,I24273,g27252,g23777,g27345,I20700,I39249,g9778,g27791,I20637,g24319,g24616,g28630,g21176,I15517,g23600,I39909,g10898,g21708,I18108,g16965,g22992,g29245,I29897,g25763,g27159,g2400,g26981,g20439,g22033,g660,g21401,g21855,I20664,I25596,g24283,I21959,g8150,g23077,g2498,g26822,g7967,g19830,g10590,g24520,g4523,I37740,g25934,g4389,I36732,g19302,g2356,g18448,g13225,g28059,g6041,g19057,g26513,g12193,g1006,g16184,I29802,g27533,g22483,g21807,g26640,g26982,g22988,I39942,g28457,g19477,I23996,I30362,g20496,g19808,g5418,g1004,I30673,I24150,g3045,g29994,g12327,g29201,g19673,I25092,I23266,I26895,I36568,g5849,g15873,g19936,g9766,g19654,g12135,g28854,g27471,g809,g20330,g16971,g231,g15020,g5732,g30665,g12820,g30409,g6131,I28087,g10451,g15718,g26877,g20836,g16880,g22642,I32146,g29320,I24352,g24507,g28213,g1003,g22533,g20368,I31136,g13322,g24859,g16523,g26692,g29200,g29574,g17500,g18048,g16368,I19642,g24494,g30241,g28728,g24265,g10535,I34041,I24380,g19929,g26361,g20409,I29439,I39391,g11228,g16791,g28959,g19765,g28310,I25389,g30451,I24187,g25025,g5798,I31682,g1570,g26832,g29181,g15305,g29693,g9520,I37611,g2457,g1718,g28845,g25238,I33915,g4737,g25132,g9580,g4055,I36542,g10046,g10870,g26022,g16129,I25264,I27128,g22660,I26220,g9765,I36159,g29965,I14550,g11948,g21685,g27484,g12463,g16283,g9810,I33554,g11341,g7895,g20480,g30529,g1389,g26550,g29332,g25609,I32547,g29543,g1119,g8418,g17396,g23717,g20426,g21771,g30975,g27248,g21856,g11853,g17493,g7152,g10567,g11600,g29937,g13500,g12901,g23844,g8475,g16934,I32492,g27436,g12008,g5641,g17719,g27286,g12515,g13057,g4578,I15546,I25617,g23626,g25280,g28041,g19766,I18569,g27210,I40718,I19602,g23428,g1060,g11975,g24963,g13833,g6896,g13170,I37924,g19007,g29545,g21111,I39341,g12797,I30826,I24188,g2020,I38345,g21144,I18524,g20332,I18130,I24207,g15175,g24268,I41018,g20473,g6220,g5907,g130,g15831,g14657,g18536,I36733,g2597,g12553,g22685,g10594,g13824,I17746,g18436,I25702,g28076,g832,g19050,g25752,g9288,g17018,g5869,g28817,I21301,g1068,g11995,g24391,g21948,g7970,g20420,g4749,I25445,g17993,g27029,I16050,g19591,g23872,g24214,g22004,g16862,g692,g6173,g13953,g16097,I27232,g11724,g22809,I31823,I16650,g19662,g8218,I37702,I38091,I29148,g29285,g28225,g30020,g11885,g23899,g28038,I19986,g12505,g13552,I25525,g12551,g30484,I18121,I17925,g9009,g26811,g26429,g28528,g7989,I18533,g23057,I15779,g10164,g26635,g8242,g16345,I14937,g13655,g398,g28639,g27916,g21242,g20453,g20503,g23913,I29049,g24068,I23200,g17776,g19098,g7560,I21398,g16404,I34204,g29817,g14332,g4243,I22554,g24868,g24594,g8485,I35057,I29432,g29175,g23448,g13252,g7534,g20938,I30206,g7328,g2226,g20014,g2486,I13228,g29708,g23181,g19813,g26817,I16221,g22134,g30562,I18181,g19418,g13866,I16082,I36423,g26607,g29877,I18680,g19785,g29396,I29383,g28052,g28455,I22715,g16262,I29206,I39041,g22721,g15793,I25117,g22999,g13971,I34719,g13835,g24569,g20666,I29426,g28436,g1789,g6290,g5928,g23631,I16172,g29770,g9746,g8302,g29469,g30456,g2562,I21429,g26494,g30435,g28928,g23320,g9920,g20284,I33418,g15261,g16590,g27737,g9227,g2777,g27344,I31127,g25562,g28666,g30129,g8793,g25265,g7916,g17237,g15591,g9595,g21053,g21117,g1739,I26461,g19379,I31793,I35983,g14123,I32431,I28249,I35028,g21461,g7478,g17357,g2377,g27162,I27314,g13049,g24580,g14423,I16633,I26115,g29667,g10912,I40823,g2785,g27233,g24638,g23137,g22076,g23721,g28335,I34776,g15839,g24501,g19574,I32519,g16728,g27088,g17902,g30913,g22707,g24759,g14570,g367,g21134,g15032,g8636,g7530,I13242,g5860,g28173,I30952,g5173,I23645,g10361,g5260,g28496,g20729,g21164,I27200,g24176,I24104,g22288,g29205,g20557,I35364,g7962,g30405,I18602,g27672,I27285,I26596,g10279,g21209,g968,g6063,g15366,g5956,I28461,g23160,g10385,g10605,g26846,g23196,g30523,g18920,g24856,I19545,g10477,g10678,g28106,I31568,g21966,g30333,g4809,g25030,I34059,I39414,g22661,I24438,g185,I28271,I28065,g27195,g2773,I22912,I25067,I23133,g13441,g21862,g17578,g23460,g3774,g30813,g22887,I25771,I25153,I23226,g4788,g27214,g13284,I21075,g19524,g5027,g25054,g29614,g13992,g29289,g13705,g174,g26449,g4894,g24974,g22171,I20033,g28193,I15451,g29471,g16444,g3945,I17060,g26696,g25915,g10194,I21871,g12282,I33583,g12611,g28333,I15887,g13415,I21415,g21457,g19350,g6083,g5305,g16836,g1039,I13169,g18666,g987,I16857,g10572,g8014,I28072,I33692,I13137,g9446,I35933,g2421,I33652,g738,g11514,g24656,g3128,I16736,I35796,I17030,g70,g8009,g15790,I27161,g26191,g1095,I29957,g12221,g16966,I21395,g24150,g22059,g12044,g3245,g25094,g27257,g927,I38606,g29747,g24993,I28988,g10291,I40297,g10909,g10626,g21238,g27706,I16292,g20754,g25112,I40844,g9277,g22611,I17027,g29375,I22962,I14280,g24128,I19971,g29443,I19500,g1223,I26285,g30222,I31226,g25985,g8752,g11524,g9005,g18936,I15288,g13515,I21289,g24570,g22911,I27426,g19467,I17632,g15544,I37653,g17973,g8649,g19018,I36903,g13342,g28897,I19722,g13530,g16325,g25942,g30307,I37778,g17124,g30743,g6216,I27369,g12354,g12105,g20911,g15477,g24452,I31895,I14568,g21267,g24668,g10406,g26676,g29556,I28084,I28997,g1085,g14483,g27517,g135,g5196,g13213,I28218,I30140,I26816,g1332,g4041,I33659,I25768,g22020,g22666,g26356,g8278,g27760,g27202,g22261,g11117,g19191,g9745,g17734,g29844,g21501,g10779,g10645,I34713,g29170,g24794,g20411,I37197,g12539,g5921,g23819,g18553,g25850,I23619,I16065,I39384,g29496,g12742,I30278,g1895,g17249,g4289,g25931,g15440,g10170,I15487,g13309,I34105,g5962,g24477,I38683,g9734,I23959,I34438,g13483,g27925,g10935,I17869,I33667,I29392,g6045,g30290,g8627,I14897,g4655,I30728,g653,g20432,I38860,g9910,g10915,g17433,g15640,g10326,g27629,g18226,g2941,g26311,I37956,g11798,I38650,g11558,g16794,g11199,g2083,g4474,g575,g12520,I40134,I14783,g8481,g16412,g354,I18154,g29397,I29354,g17064,g10211,g21389,I26469,g25989,g12078,g25835,g29275,I26695,g6082,g11528,g29934,I25763,I26574,g19494,g15605,g30029,g10588,g9065,g27696,g25104,g28529,g1621,I27240,g28368,g7013,g3155,g29186,g15898,g11660,g30442,g28691,I32540,g9807,g17382,g30757,g27679,I28741,g24321,I36330,I40429,I29399,g13954,g28481,g15439,I40943,g4827,g26119,g21357,g25393,g1858,g3051,g29761,g11264,g22588,g28401,g25462,I40793,g25631,g30759,g18389,g996,g29286,I30922,g26015,I25374,g12025,g13907,I25225,g16113,g10169,I14819,g7141,g9663,g22658,g22728,g15730,g5886,g28480,g30565,g28696,I17122,g28465,I40066,I38007,g21314,g30228,g20460,g4602,g6301,g17959,g13704,I14496,I31886,g1991,g17688,g1063,g562,g19079,g18638,I33520,g11417,g20622,g22044,I13186,I38905,g30233,g2279,g26563,g22794,g16170,g30705,g30856,g7957,g2588,g6020,I27071,I26690,g19704,g23577,g20982,g20599,I15478,I20022,g27946,I21389,g11843,g13429,g11401,g16864,g25304,g8860,g28662,I38085,I34192,g30084,g3254,g5129,g14360,g30801,g13505,I36876,g28723,g20840,g30070,g20045,g28280,g10796,I21598,I31011,I17759,I29493,g24440,g27083,g20935,g19321,g24130,g5597,g8490,I34860,g8387,g26504,g12194,I28365,I38380,g18505,g23432,g11868,g18059,g21428,g29628,g19561,g11202,g18509,g29576,g28846,I26947,g21152,I40985,g20444,g25146,g12930,g15931,g26961,g10683,g24371,g13624,g30747,g25377,g16708,I35116,g11954,I22318,g16654,g6021,g24490,g19413,I31298,I32500,I36909,g30124,g2258,g27674,g9762,g30974,g21130,g13153,I33714,g22702,g28068,g21932,I31877,g27909,I21326,I40137,I14755,g23783,g20949,g22773,I20559,g21491,g18465,g590,g30829,g21328,g28145,g27673,g18053,I25015,g30273,I16967,g20471,I28351,g30119,g20968,g1138,I15562,g1733,g30517,g9812,g18903,I24205,I30110,g1970,g15524,g29950,g30663,g30390,g13582,g20282,g30402,I38379,I27422,g26477,g15460,g30509,g25042,I31074,g20316,g30366,g4845,g21438,g15993,I34794,g11989,g6031,g4144,I38154,g5255,g18755,I25486,g12302,g30549,g6431,I24476,g12210,I40032,g10568,g12548,g8031,I18238,g10616,g8570,I18197,I24445,g13109,g9462,g1400,g23029,g23287,g26970,g28346,g20290,g21636,g1833,I13176,g520,g30515,g13998,g2956,g23796,g24551,g16656,I35488,g23555,I16552,I18423,g22812,g29223,g4325,g30281,g24206,g26918,g5355,g29814,g23135,I30371,g24502,I31244,g8961,g26251,g24879,g24229,g29506,g26779,g15128,g11045,g22769,I15206,g20396,I32642,g18313,g30767,I20320,I41117,g1403,I35783,I25616,I19894,g11864,I28235,g15691,g26190,g5910,g19771,g14113,g822,I39906,g2599,I38145,g19987,g28606,g28070,g273,g995,g16848,g21105,g29819,g6044,g26785,g6641,g13496,g25072,g29367,I16544,I32357,g25524,g20111,g23270,I24368,g17235,g12213,g22093,I25395,I17081,g20329,g12307,g22846,g1444,I31583,g29421,I35443,g10058,g25805,g20912,g97,g353,g7570,g12346,I17097,I41111,g19195,g29776,g7562,g13598,g6448,g29222,g29686,g21735,I34779,g21173,g11711,I27897,g26837,g11154,g23785,g25282,g30597,g12506,I36296,I28133,g1899,g27319,g19390,g11944,g12264,I34476,g19349,I23154,I29533,g6080,g26660,I25237,g21914,g9310,I41066,g18822,g27182,I26642,g21116,g4570,I25752,g25313,g1183,g13286,I15590,g22167,g13903,g30344,g11687,g26291,g27059,g13110,g10458,g26958,I36933,I13113,I34701,I17009,g6118,I30944,g20270,g16478,g11713,g27806,g1044,g461,I25830,I18414,I35821,I32886,g10374,g24781,I36987,g18383,g25232,g26671,I23679,g15562,g29575,g18012,I35548,I40898,g20038,g29571,g22590,g13633,g22683,g22619,g23501,g869,g25014,I40964,g27364,g16094,I39791,g27284,I40501,g24531,g22775,g13790,g24912,g8893,g18834,g26239,g21364,g21370,I15276,I37303,g11531,g17788,g20714,g23888,I39825,g23677,g15513,I39457,g4304,I37002,g22455,g5118,g8571,g7348,g23023,g25017,I15602,g9000,I40507,g12769,I23860,g12070,g27879,g1734,I32546,I25351,g7865,g12370,g22760,I19539,g10259,g18670,g9390,I20703,g18646,g27710,I18512,I32868,g28739,g16856,g30578,g20081,I34725,g21023,I40838,g10644,g1009,g25173,I29238,g12197,I40510,g28011,I40895,g3834,g19043,g30449,g27721,I40922,I38539,I31913,g26771,g3243,I31050,I18728,I39691,g19913,I18160,g27184,g23667,g27071,g28231,g29475,g9090,g2099,g3092,g5256,I36267,g5871,g24790,g23771,I34773,g25927,I20556,g4237,g21354,g27126,g22029,g20,g11675,g19380,I26990,I30985,g27568,g15769,g18993,g29967,g26669,g16615,I24417,g19631,g7661,I39005,g5810,g12532,g11913,g6014,I29451,g19457,I31772,g27052,g26658,g11701,g10682,g25881,g2427,g14747,g1785,g25409,g21639,I32559,g8817,g4468,g26442,g12056,g24838,g1947,g26399,g11367,g29204,I22885,g20005,g19040,g23886,I33377,g4720,g24605,g30107,I20813,g28360,I40239,g23191,g22147,g27219,g20942,g19128,g30351,g21268,g29619,g23666,I14993,g16243,I31282,g27554,g12487,g9908,I38363,g3067,g5744,g22735,g28644,g27799,g16479,g11719,g4929,g24052,I30083,g26739,I23131,g26783,g26763,g16278,g8788,I29690,g19737,g4191,g8534,g4954,g27700,g192,g20105,g18896,I37379,g20997,g1250,g21029,g16736,I24029,g24755,g19483,g10595,g25513,g5762,g22034,g17436,g22445,I38599,g23740,g5050,g12780,I24702,g8990,I24684,g3176,g23420,I40937,g21991,g16725,g16032,g24884,I40814,g225,g25159,I25588,g12828,g29724,g9064,g18351,I39020,g10509,g7849,I33732,g14745,I25272,g2798,I32143,g18743,I32847,g26617,g21589,g23224,g6034,g15667,g9857,I18444,g1055,g19586,g23148,g22550,I38024,g23508,g25035,g7922,g29767,g5621,g20919,g30928,g18464,g17285,g5966,I18764,g16767,I34641,I30275,g21055,I26599,g25269,g1834,I22947,g28958,g24003,g23219,g19629,I24667,g17815,I24624,I27349,g26621,g10674,g10232,g24315,g16056,I31508,g8822,g52,g24578,g23038,g2649,g20344,I33157,g17714,I18617,g8885,I39889,g30712,g26684,g28072,g11796,I17954,I31640,g29974,I24247,g19198,I34091,g13191,I25402,I30296,g1386,g28843,g11553,g23897,g22986,g5712,g28299,I29613,g26560,g368,g13244,g26639,I23027,I31460,g29296,g24796,g2628,I38838,I33424,g12196,g16138,g27681,I26564,g28206,g26567,g18276,g28192,g19860,g15635,I21868,g30005,I20031,g20615,I30338,g1414,g20573,I22578,g21278,I23257,g27772,I28550,I39689,g19621,g6226,g8842,g15624,g17158,I27053,g1727,g7459,I34842,g12807,g19709,I24407,I37161,g17856,g13296,g12643,g16035,g1259,g15777,g27581,g14355,g24288,g13203,g22712,g29380,g20899,g5604,I13203,g11108,g26935,g13506,g7479,I33491,I16238,g9869,g5890,g10499,g16443,g24756,g29810,g10473,g30791,g21305,I22755,g11637,g6022,g18091,g13163,g25626,I27044,I16521,g13202,g16439,g3366,g12854,g13096,I22557,I23351,g17640,g11908,I19872,g25250,g29827,g18829,g7643,g2525,g27043,g8650,g1201,g10175,g11695,g6079,I38412,g2691,g9257,g10409,g316,I16206,I36921,g29057,I33837,g7483,g10460,g4009,g3236,g4680,I28956,g25612,g10517,g8573,I30782,g567,I35533,g16072,I23745,g22064,I22632,I38211,g18962,g7616,g14795,g25111,g13041,g26236,g15781,g2657,g24037,g21844,g23617,I18632,g13428,g7140,g24335,I24062,I24180,I16532,I24285,g27523,g449,g28446,g24775,g28712,g30406,g13740,g20939,g14957,g7555,g20470,g26259,g23608,g17548,g23110,g23267,I40796,g11670,I40188,g23294,g24291,g24450,I15856,g2563,I14030,I21310,g17221,g30709,I14298,g30109,g15201,I41135,g23598,I15818,I22803,g19166,I15771,I18572,I23047,g24089,g10375,g17782,g12172,g30286,g20576,g26397,g25251,g29090,I30248,g17664,g29501,I26916,g20022,g718,g2378,g30809,g28720,I13165,g4650,g5417,I32976,I35737,g28900,g21521,g23737,g30671,g7577,I16697,g27220,g22663,g25476,I21274,g25323,I34056,I39886,I39933,g10450,I28991,g29739,g24922,g21235,g30229,g13237,I39870,g26061,g30340,g24498,I38594,g12061,g21141,g1689,g29339,g8313,g29931,g25235,g736,g28852,I22028,I35974,I27355,I14562,g20885,g169,g21726,g10308,g2026,g22996,I29212,g13571,g15148,I32608,g22283,I23292,g20049,g11007,g30398,g24365,g9607,g26812,g23154,g9901,g9759,g30645,g2617,g8829,I31829,g26060,g26655,g11718,g5634,g28345,g12166,g30524,g28772,g22333,g29185,g14514,g28714,g30195,I20592,I16630,g13151,I14577,g29764,g8491,g25472,g23438,g9276,g20637,g381,g5398,I23966,g20148,I18545,I29348,g15700,g29648,g19639,g10397,g5897,g19638,I15012,g19268,g10210,g13845,g26781,I37587,g1425,g12000,g25134,g4902,g21689,g20983,I36096,g18720,g21070,I18107,I38909,I24588,g24362,g9879,g30811,g26868,g11647,g9795,g29329,g2129,g25767,g21293,g15719,g20080,g30480,g11838,I25171,I27646,g23765,g25128,I20339,I15326,g17704,g10065,I24752,g20946,g5289,g14124,g13786,I39859,g11593,g26508,g20272,g14764,g11555,I31916,g26223,g18538,g28103,g30714,g28636,g16719,g30657,g17557,g10151,g13756,g25277,g10189,g30547,g25762,g27705,g6026,g19626,I28753,g30784,g27024,g13904,g614,I22902,g13430,g25982,g30521,g23968,g26611,g6140,g15688,g30481,g27475,g29013,I30251,I17898,g24327,g27759,g28646,g18485,g19728,I24017,I36114,I17637,I27260,g3173,g4876,g22829,g2006,g27099,g18154,g5414,I33526,g27687,g4093,g13423,g1561,g23068,g27579,g29061,g19117,g16992,g23274,g8438,g20039,g27485,I23636,g27007,g2230,g27761,g17454,g6574,g18463,g1010,g4766,g26603,g27274,g30285,I20745,I32432,g22722,I26714,I15902,g9940,g24344,g19825,g27971,g9122,g13319,g13942,g17534,g28325,g19627,g28789,g26317,g17123,g2236,I29080,I21661,I37284,g550,I21461,g17029,g16277,g7795,g27498,I32967,g21444,g26159,g15800,g154,g30453,g1210,g20584,g21814,g30548,g25554,g14107,g2641,g14976,g5405,g10606,I29724,I33374,g30099,g24354,g24676,g1769,g24140,g11858,g19351,g23798,g23256,g23971,I27140,g10252,g19776,g11465,I18396,g9073,I27761,g264,I18298,I19030,I15610,g28754,g21299,g25482,g23288,I23180,g19019,g1764,g1627,g26008,g2653,g295,g985,g27273,I14565,I15246,I33879,g27548,g30376,g21523,g16858,g17847,g15093,g5833,g22949,g26712,g10598,g11578,I18713,I20661,I32835,I24575,I35976,I30008,g8996,g22408,g7976,g1696,I24251,g22681,g22042,g16428,I31643,g16830,I16296,g21079,g21325,g29620,g1994,g12945,g27325,g20518,g26695,I37572,g8841,g21426,g25287,I16598,g28237,g8688,g10179,g143,g20353,I37665,g15388,g25780,g20117,g19795,g13514,g5940,g22036,g21554,g18651,g26037,I25741,g12285,g11432,g298,g10059,g5692,g26231,I36860,g10511,g29378,g9301,g1263,I22163,g29050,g9885,g22386,g28249,g30741,g9134,g12296,g21572,g20062,g159,g25463,I18845,g21435,g19262,g9631,I40212,I14834,g15840,g1040,g19358,g23206,g18084,g30155,g5884,I23277,g21118,g22703,g13825,g22190,g30504,g21858,g23694,g9263,g27035,g16831,I14556,g22840,g3032,I32370,g13476,g1558,g5766,g24449,g5409,g11082,g17795,g19661,g15569,g8900,g23915,I22064,I28169,I23475,g10787,g26854,g10393,g28274,g26630,I24521,g9961,g16490,g23532,g8897,g11351,g22043,g20984,g18908,I33603,g26757,g14263,g18616,g18928,g29182,I15642,g10147,I15787,g13407,g13056,g25220,g30455,g13195,I30489,I33822,g27414,g16986,g219,g22214,g2087,I30797,g10183,g22443,g23024,g441,g20825,g22837,g21337,I36592,g29105,g17471,g18312,g12271,g11291,g16482,g30114,g27190,g23407,g3249,I29635,g13300,g22831,g15660,g16160,I19996,g19692,g29779,g18278,g29087,g20390,g24091,I38355,I25966,I13652,g20802,g8687,I24076,g22285,I19891,g30638,g26,g25967,g27824,I17884,g29645,g517,I38719,g24264,I22542,g22517,g16299,g24328,g16349,g29324,g18764,I35703,g28124,I21304,g864,g19803,g1388,g4012,I40916,g29137,g12067,g23527,g20082,g15526,g13067,I35347,g28983,I34146,g27016,g30909,g30473,g13738,g20293,g30225,g13944,I33999,g12433,I19274,g4786,g9956,I39628,g27531,g30910,I17743,g9775,g25239,g24109,I21772,g27567,g28963,g9504,g10800,I30560,g17577,g20481,g4548,I22875,g25899,g28062,I40206,g7788,I18311,I36379,g10287,g17655,g13310,g11888,g19143,g24481,I22924,g5995,g5280,I17061,I24416,g5170,I37400,g20434,I24252,g24225,g13391,g10306,I38226,I33577,I22699,I31802,g13354,I34428,g15557,g30294,I13246,g22990,g27155,g24284,g26689,g24513,g11628,I36772,g2935,I25365,I34731,g1552,g21955,g12001,g26288,g24905,g18089,I16493,g4803,g15092,g27494,g9079,I40614,g16288,I14742,g10880,g11927,g27868,I28509,g5666,I24049,g4240,I19510,g22690,g27842,g18655,g28665,g29158,I33297,g24336,g10447,g3129,I23265,I18381,g15818,g23632,g22205,g11278,g29224,g24881,g21418,g26034,g29969,g17405,g26742,I16432,I31493,I38250,g19288,g30637,I31024,I29496,g23001,I35536,g24553,g22743,g11281,g9522,g30067,I21577,g1539,g4310,g29962,g30835,g10466,I25180,g27397,g19420,g16846,g21703,g25711,g12969,g24033,g29199,g195,g13222,g15231,g19450,g24463,g1236,g19711,g16997,g24341,g28783,g13854,g971,g21095,I37784,I18247,g23641,g22941,g23775,g2543,g29265,I16037,g14139,g19567,g10928,I19315,g24565,g18945,I20828,g1557,g29809,g28689,g26706,g17083,g4251,g20895,g19976,I16228,g20091,g28832,g5850,g12646,I20628,I29468,g16071,g26405,I28728,g17160,g4714,I14928,g23312,I26960,I40799,g24524,g23837,g2529,g27911,g1401,g15622,g26861,g26964,g13146,g15306,g10474,I40647,I30038,g29580,I17685,g28608,I38049,g27006,g10846,I18335,g30688,I31739,g28235,g20140,g20704,g20564,I34983,I24373,g23253,g10064,g12385,g13477,g26196,g16101,I34044,g23838,g25422,I40051,I16089,g29566,g15991,g571,I37071,I32997,I33016,g29794,g27546,g23912,g2102,g27226,I30965,g12507,g16507,I35095,I32556,g14837,I32102,g15391,g2257,g15404,g25694,I13131,g7346,g25004,g22755,g19732,g1849,g27288,I30988,I16507,g2040,g17954,g11812,g2439,g11507,g8079,I38737,g12932,g22802,g25115,g10584,I18091,g26006,g25096,g17830,g6201,g27952,g1684,g23481,g14420,g12762,g21494,g12170,g30086,g24611,g17775,g22673,I40423,g6102,g29823,g27945,I29357,g8866,g23588,g29165,g2033,g30956,g10601,g27287,g12647,I38011,I36397,g9074,g21660,g20303,g2052,g19169,g20116,I25634,g12090,g12150,g1081,I16190,g24121,g10108,I25625,g21799,I31586,g21612,I28671,g24573,g22719,I30182,g12514,g10597,I16759,I39279,g9724,g9661,g6023,g11271,g24700,g7477,g10334,g9907,g19721,g11856,I23648,g10208,I40008,g6101,g21901,g5044,g8394,g27560,g11999,g26827,g21891,I22706,g15951,g20497,g11321,g19894,g21561,g22962,g29253,g29081,g10476,I22382,g7600,g337,g19558,g20986,g22548,g27573,g3096,g30121,I28458,g16505,g20313,g5968,I27324,g21214,g8503,I23386,g10518,g6894,g20516,g20398,g30679,g8227,g15792,g12069,g7561,I14715,g10592,g23580,g16809,g20951,g13957,g30855,I16079,g21943,g2930,g12851,g27965,g5047,g20255,g15335,g8871,g19053,g25095,I36270,g15837,g5794,g30837,g8514,I27976,I32369,g2455,g25306,g25141,g22240,I23880,g27993,I34425,g10673,g28407,g12208,I29360,g22056,g24247,g22828,g30358,g25869,g21154,g22748,g22921,I30173,I18596,g28925,g17465,g24232,g744,I29220,I30233,I18259,g2231,g16367,I17235,g28894,g27078,g15981,g29274,g29431,I25500,I19747,g29328,g12048,I15593,g20084,g23747,g1448,g18668,g849,g6190,I20852,I16255,g4945,I24501,g20978,g12495,I41024,g25818,g11747,g17462,g20110,g28373,g21952,I27411,g22067,g23602,g22607,I13987,g24470,g10927,g11544,g24590,I25801,g20219,I30568,g24227,I20347,I31109,g14584,g15609,g28265,g10281,g11252,g24535,g28698,g27354,I22283,g26799,g23220,I33548,g30278,I37252,g20375,g8366,g18757,g10412,g24002,g26966,g1173,g10207,g6047,g22399,I24400,g17579,g23500,I34872,g707,g376,g20566,I33870,g3242,I24751,g26922,I31646,I30676,g23357,I29259,g1959,g20309,g25868,I32955,g11354,g24390,g6042,g24298,g15628,I23578,g1309,g29689,I32946,g25171,g11042,g29196,I21674,I24131,g26310,g7649,g1228,g21456,g26994,g15174,I31610,g29417,g10672,g2370,g4574,g17174,g8277,g23821,g1822,g15311,g12755,g30291,g8621,g26831,g30113,I40997,g27064,g29235,I40119,g3954,g21489,g11523,I35479,g12524,g8850,g18332,g24389,g10041,I29653,I19552,g27843,g18708,g6568,g10202,g11881,I26940,I22575,g4318,g21486,I38872,g13480,g13037,g8182,g13247,g19669,I28057,g22087,g14381,g26610,g26031,g5628,I19883,g21530,I40518,g28128,g28735,g161,I32904,g21750,g5982,g22199,I21446,g5630,I18244,g29255,I24495,g727,g2358,I38053,g1251,g26496,g28820,I38391,g8945,g21374,g8723,g29822,g19625,g19594,g21558,g24325,g29702,g21412,g29957,I37322,g27100,g26963,g5847,g11759,g15160,g27790,g24652,I37313,I36666,g4555,g30513,I18314,g9368,g2112,g24094,g19232,g11259,I18417,g26053,g23859,g8107,g30792,g13990,g5829,g30764,g12104,g11791,g28392,g10640,g22948,g11960,I32170,g26988,I19523,g23123,g24814,g22791,g30650,I24507,g24546,g17517,g22500,g22765,g28668,g19387,I34821,I30134,g24557,g10452,I25722,I36314,g29773,g30352,g22032,I27297,g4194,g25392,I20467,g23628,g5186,I31811,I23153,I29386,g22156,g28467,g11673,g12037,I36316,I13993,g20362,I39393,I19240,I23242,g11475,g2888,g18374,I18031,g15546,g21488,g16673,g21628,I23380,g15694,g2205,I21583,g23228,I29274,g20789,g9606,g21540,g19385,I19847,g1893,g14207,I36656,I14580,g23471,g26478,g19049,g30720,I24711,g524,I22938,g8993,g26666,I25881,g30763,g4281,g18815,g12362,g30271,g21394,g24840,I25186,g28341,g27854,g30848,g2813,I23326,I13200,I32595,g18946,g21824,g21980,g12336,g284,g19153,I25249,g30640,g25082,g23012,I40542,g24503,g22467,I19195,I16264,g65,g4406,I37228,g957,g30100,g28782,g18107,g15582,g21368,g17177,g24426,I23361,g27479,g26240,I19119,I38749,I32487,g342,g23635,g9382,g30034,g7195,g20395,g20360,g30786,g6636,g23286,g11606,g23581,g17381,g23803,g646,g8756,g26704,I40778,g10540,I28155,g27317,g1747,g1559,g23625,g13405,I32460,g21331,g26024,g27370,I15654,I20607,g4326,g10364,I33293,g14882,g30488,g25761,I35109,g13385,I37566,g16607,g11265,g11105,g29323,g29991,g30929,g23387,g24451,g24360,g975,g15422,g11886,I15345,g6908,g25652,g16994,g2639,I31661,g10229,g26720,I35919,g30685,g27093,g27659,g24986,I29610,g8549,g21335,g11549,g17613,g28454,g15814,g30819,I14040,I33347,g28364,I26198,g10230,g20876,I17303,g14831,g23163,g1365,I28485,g17636,g20981,g2412,g25367,g18914,I31634,g19039,I25790,I33445,g13188,g4383,I31550,g30012,g22664,g24542,g20512,I34012,g17794,g21097,g19816,I19582,g16104,g14796,I36696,g8071,g13238,I32392,g10930,g18106,I33897,g16908,g14719,g8520,g1591,g22405,g26624,I29812,g981,g13724,I17429,g26143,g28381,g6421,I26388,g243,I31188,g26841,g10115,g18954,g14685,g726,g12225,g30846,g16344,g23000,g12702,g14690,I40859,I13575,I31619,g10464,g2459,g5298,g29065,g29913,g3987,g24334,g12997,g26488,g13452,g30526,g19606,I23083,g13448,g28160,g22662,I38644,g11517,g28736,I19952,g6029,g28425,g19823,g26372,g19920,I37017,g8530,g396,g30761,g12083,I28107,g18449,g24348,g13365,g21291,g12599,g27800,I19791,g5805,g29409,I35394,I35817,I40128,g8126,g16847,I28103,g27415,g5301,g23744,g12222,g28774,g15672,g16693,g30858,g9748,g23104,g21168,g17738,g9264,g22734,g26965,I37868,g28210,g19601,g14641,g30972,I24007,g22040,g13464,I39982,g1033,g8646,g11983,g22668,g26387,g22745,g5631,g13886,g11833,g11580,g18859,g23134,g8386,g22000;
//# 28 inputs
//# 106 outputs
//# 1636 D-type flipflops
//# 13470 inverters
//# 8709 gates (4154 ANDs + 2050 NANDs + 226 ORs + 2279 NORs)
//
//
//
  MSFF DFF_0(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2814),.DATA(g16475));
  MSFF DFF_1(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2817),.DATA(g20571));
  MSFF DFF_2(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2933),.DATA(g20588));
  MSFF DFF_3(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2950),.DATA(g21951));
  MSFF DFF_4(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2883),.DATA(g23315));
  MSFF DFF_5(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2888),.DATA(g24423));
  MSFF DFF_6(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2896),.DATA(g25175));
  MSFF DFF_7(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2892),.DATA(g26019));
  MSFF DFF_8(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2903),.DATA(g26747));
  MSFF DFF_9(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2900),.DATA(g27237));
  MSFF DFF_10(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2908),.DATA(g27715));
  MSFF DFF_11(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2912),.DATA(g24424));
  MSFF DFF_12(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2917),.DATA(g25174));
  MSFF DFF_13(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2924),.DATA(g26020));
  MSFF DFF_14(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2920),.DATA(g26746));
  MSFF DFF_15(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2984),.DATA(g19061));
  MSFF DFF_16(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2985),.DATA(g19060));
  MSFF DFF_17(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2930),.DATA(g19062));
  MSFF DFF_18(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2929),.DATA(g2930));
  MSFF DFF_19(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2879),.DATA(g16494));
  MSFF DFF_20(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2934),.DATA(g16476));
  MSFF DFF_21(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2935),.DATA(g16477));
  MSFF DFF_22(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2938),.DATA(g16478));
  MSFF DFF_23(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2941),.DATA(g16479));
  MSFF DFF_24(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2944),.DATA(g16480));
  MSFF DFF_25(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2947),.DATA(g16481));
  MSFF DFF_26(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2953),.DATA(g16482));
  MSFF DFF_27(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2956),.DATA(g16483));
  MSFF DFF_28(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2959),.DATA(g16484));
  MSFF DFF_29(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2962),.DATA(g16485));
  MSFF DFF_30(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2963),.DATA(g16486));
  MSFF DFF_31(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2966),.DATA(g16487));
  MSFF DFF_32(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2969),.DATA(g16488));
  MSFF DFF_33(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2972),.DATA(g16489));
  MSFF DFF_34(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2975),.DATA(g16490));
  MSFF DFF_35(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2978),.DATA(g16491));
  MSFF DFF_36(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2981),.DATA(g16492));
  MSFF DFF_37(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2874),.DATA(g16493));
  MSFF DFF_38(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1506),.DATA(g20572));
  MSFF DFF_39(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1501),.DATA(g20573));
  MSFF DFF_40(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1496),.DATA(g20574));
  MSFF DFF_41(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1491),.DATA(g20575));
  MSFF DFF_42(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1486),.DATA(g20576));
  MSFF DFF_43(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1481),.DATA(g20577));
  MSFF DFF_44(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1476),.DATA(g20578));
  MSFF DFF_45(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1471),.DATA(g20579));
  MSFF DFF_46(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2877),.DATA(g23313));
  MSFF DFF_47(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2861),.DATA(g21960));
  MSFF DFF_48(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g813),.DATA(g2861));
  MSFF DFF_49(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2864),.DATA(g21961));
  MSFF DFF_50(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g809),.DATA(g2864));
  MSFF DFF_51(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2867),.DATA(g21962));
  MSFF DFF_52(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g805),.DATA(g2867));
  MSFF DFF_53(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2870),.DATA(g21963));
  MSFF DFF_54(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g801),.DATA(g2870));
  MSFF DFF_55(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2818),.DATA(g21947));
  MSFF DFF_56(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g797),.DATA(g2818));
  MSFF DFF_57(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2821),.DATA(g21948));
  MSFF DFF_58(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g793),.DATA(g2821));
  MSFF DFF_59(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2824),.DATA(g21949));
  MSFF DFF_60(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g789),.DATA(g2824));
  MSFF DFF_61(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2827),.DATA(g21950));
  MSFF DFF_62(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g785),.DATA(g2827));
  MSFF DFF_63(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2830),.DATA(g23312));
  MSFF DFF_64(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2873),.DATA(g2830));
  MSFF DFF_65(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2833),.DATA(g21952));
  MSFF DFF_66(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g125),.DATA(g2833));
  MSFF DFF_67(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2836),.DATA(g21953));
  MSFF DFF_68(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g121),.DATA(g2836));
  MSFF DFF_69(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2839),.DATA(g21954));
  MSFF DFF_70(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g117),.DATA(g2839));
  MSFF DFF_71(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2842),.DATA(g21955));
  MSFF DFF_72(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g113),.DATA(g2842));
  MSFF DFF_73(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2845),.DATA(g21956));
  MSFF DFF_74(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g109),.DATA(g2845));
  MSFF DFF_75(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2848),.DATA(g21957));
  MSFF DFF_76(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g105),.DATA(g2848));
  MSFF DFF_77(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2851),.DATA(g21958));
  MSFF DFF_78(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g101),.DATA(g2851));
  MSFF DFF_79(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2854),.DATA(g21959));
  MSFF DFF_80(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g97),.DATA(g2854));
  MSFF DFF_81(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2858),.DATA(g23316));
  MSFF DFF_82(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2857),.DATA(g2858));
  MSFF DFF_83(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2200),.DATA(g20587));
  MSFF DFF_84(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2195),.DATA(g20585));
  MSFF DFF_85(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2190),.DATA(g20586));
  MSFF DFF_86(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2185),.DATA(g20584));
  MSFF DFF_87(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2180),.DATA(g20583));
  MSFF DFF_88(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2175),.DATA(g20582));
  MSFF DFF_89(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2170),.DATA(g20581));
  MSFF DFF_90(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2165),.DATA(g20580));
  MSFF DFF_91(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2878),.DATA(g23314));
  MSFF DFF_92(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3129),.DATA(g13475));
  MSFF DFF_93(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3117),.DATA(g3129));
  MSFF DFF_94(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3109),.DATA(g3117));
  MSFF DFF_95(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3210),.DATA(g20630));
  MSFF DFF_96(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3211),.DATA(g20631));
  MSFF DFF_97(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3084),.DATA(g20632));
  MSFF DFF_98(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3085),.DATA(g20609));
  MSFF DFF_99(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3086),.DATA(g20610));
  MSFF DFF_100(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3087),.DATA(g20611));
  MSFF DFF_101(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3091),.DATA(g20612));
  MSFF DFF_102(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3092),.DATA(g20613));
  MSFF DFF_103(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3093),.DATA(g20614));
  MSFF DFF_104(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3094),.DATA(g20615));
  MSFF DFF_105(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3095),.DATA(g20616));
  MSFF DFF_106(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3096),.DATA(g20617));
  MSFF DFF_107(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3097),.DATA(g26751));
  MSFF DFF_108(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3098),.DATA(g26752));
  MSFF DFF_109(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3099),.DATA(g26753));
  MSFF DFF_110(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3100),.DATA(g29163));
  MSFF DFF_111(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3101),.DATA(g29164));
  MSFF DFF_112(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3102),.DATA(g29165));
  MSFF DFF_113(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3103),.DATA(g30120));
  MSFF DFF_114(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3104),.DATA(g30121));
  MSFF DFF_115(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3105),.DATA(g30122));
  MSFF DFF_116(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3106),.DATA(g30941));
  MSFF DFF_117(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3107),.DATA(g30942));
  MSFF DFF_118(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3108),.DATA(g30943));
  MSFF DFF_119(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3155),.DATA(g20618));
  MSFF DFF_120(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3158),.DATA(g20619));
  MSFF DFF_121(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3161),.DATA(g20620));
  MSFF DFF_122(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3164),.DATA(g20621));
  MSFF DFF_123(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3167),.DATA(g20622));
  MSFF DFF_124(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3170),.DATA(g20623));
  MSFF DFF_125(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3173),.DATA(g20624));
  MSFF DFF_126(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3176),.DATA(g20625));
  MSFF DFF_127(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3179),.DATA(g20626));
  MSFF DFF_128(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3182),.DATA(g20627));
  MSFF DFF_129(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3185),.DATA(g20628));
  MSFF DFF_130(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3088),.DATA(g20629));
  MSFF DFF_131(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3191),.DATA(g27717));
  MSFF DFF_132(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3194),.DATA(g28316));
  MSFF DFF_133(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3197),.DATA(g28317));
  MSFF DFF_134(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3198),.DATA(g28318));
  MSFF DFF_135(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3201),.DATA(g28704));
  MSFF DFF_136(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3204),.DATA(g28705));
  MSFF DFF_137(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3207),.DATA(g28706));
  MSFF DFF_138(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3188),.DATA(g29463));
  MSFF DFF_139(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3133),.DATA(g29656));
  MSFF DFF_140(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3132),.DATA(g28698));
  MSFF DFF_141(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3128),.DATA(g29166));
  MSFF DFF_142(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3127),.DATA(g28697));
  MSFF DFF_143(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3126),.DATA(g28315));
  MSFF DFF_144(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3125),.DATA(g28696));
  MSFF DFF_145(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3124),.DATA(g28314));
  MSFF DFF_146(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3123),.DATA(g28313));
  MSFF DFF_147(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3120),.DATA(g28695));
  MSFF DFF_148(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3114),.DATA(g28694));
  MSFF DFF_149(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3113),.DATA(g28693));
  MSFF DFF_150(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3112),.DATA(g28312));
  MSFF DFF_151(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3110),.DATA(g28311));
  MSFF DFF_152(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3111),.DATA(g28310));
  MSFF DFF_153(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3139),.DATA(g29461));
  MSFF DFF_154(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3136),.DATA(g28701));
  MSFF DFF_155(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3134),.DATA(g28700));
  MSFF DFF_156(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3135),.DATA(g28699));
  MSFF DFF_157(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3151),.DATA(g29462));
  MSFF DFF_158(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3142),.DATA(g28703));
  MSFF DFF_159(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3147),.DATA(g28702));
  MSFF DFF_160(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g185),.DATA(g29657));
  MSFF DFF_161(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g138),.DATA(g13405));
  MSFF DFF_162(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g135),.DATA(g138));
  MSFF DFF_163(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g165),.DATA(g135));
  MSFF DFF_164(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g130),.DATA(g24259));
  MSFF DFF_165(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g131),.DATA(g24260));
  MSFF DFF_166(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g129),.DATA(g24261));
  MSFF DFF_167(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g133),.DATA(g24262));
  MSFF DFF_168(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g134),.DATA(g24263));
  MSFF DFF_169(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g132),.DATA(g24264));
  MSFF DFF_170(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g142),.DATA(g24265));
  MSFF DFF_171(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g143),.DATA(g24266));
  MSFF DFF_172(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g141),.DATA(g24267));
  MSFF DFF_173(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g145),.DATA(g24268));
  MSFF DFF_174(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g146),.DATA(g24269));
  MSFF DFF_175(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g144),.DATA(g24270));
  MSFF DFF_176(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g148),.DATA(g24271));
  MSFF DFF_177(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g149),.DATA(g24272));
  MSFF DFF_178(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g147),.DATA(g24273));
  MSFF DFF_179(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g151),.DATA(g24274));
  MSFF DFF_180(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g152),.DATA(g24275));
  MSFF DFF_181(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g150),.DATA(g24276));
  MSFF DFF_182(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g154),.DATA(g24277));
  MSFF DFF_183(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g155),.DATA(g24278));
  MSFF DFF_184(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g153),.DATA(g24279));
  MSFF DFF_185(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g157),.DATA(g24280));
  MSFF DFF_186(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g158),.DATA(g24281));
  MSFF DFF_187(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g156),.DATA(g24282));
  MSFF DFF_188(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g160),.DATA(g24283));
  MSFF DFF_189(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g161),.DATA(g24284));
  MSFF DFF_190(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g159),.DATA(g24285));
  MSFF DFF_191(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g163),.DATA(g24286));
  MSFF DFF_192(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g164),.DATA(g24287));
  MSFF DFF_193(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g162),.DATA(g24288));
  MSFF DFF_194(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g169),.DATA(g26679));
  MSFF DFF_195(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g170),.DATA(g26680));
  MSFF DFF_196(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g168),.DATA(g26681));
  MSFF DFF_197(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g172),.DATA(g26682));
  MSFF DFF_198(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g173),.DATA(g26683));
  MSFF DFF_199(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g171),.DATA(g26684));
  MSFF DFF_200(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g175),.DATA(g26685));
  MSFF DFF_201(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g176),.DATA(g26686));
  MSFF DFF_202(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g174),.DATA(g26687));
  MSFF DFF_203(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g178),.DATA(g26688));
  MSFF DFF_204(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g179),.DATA(g26689));
  MSFF DFF_205(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g177),.DATA(g26690));
  MSFF DFF_206(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g186),.DATA(g30506));
  MSFF DFF_207(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g189),.DATA(g30507));
  MSFF DFF_208(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g192),.DATA(g30508));
  MSFF DFF_209(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g231),.DATA(g30842));
  MSFF DFF_210(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g234),.DATA(g30843));
  MSFF DFF_211(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g237),.DATA(g30844));
  MSFF DFF_212(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g195),.DATA(g30836));
  MSFF DFF_213(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g198),.DATA(g30837));
  MSFF DFF_214(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g201),.DATA(g30838));
  MSFF DFF_215(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g240),.DATA(g30845));
  MSFF DFF_216(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g243),.DATA(g30846));
  MSFF DFF_217(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g246),.DATA(g30847));
  MSFF DFF_218(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g204),.DATA(g30509));
  MSFF DFF_219(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g207),.DATA(g30510));
  MSFF DFF_220(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g210),.DATA(g30511));
  MSFF DFF_221(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g249),.DATA(g30515));
  MSFF DFF_222(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g252),.DATA(g30516));
  MSFF DFF_223(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g255),.DATA(g30517));
  MSFF DFF_224(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g213),.DATA(g30512));
  MSFF DFF_225(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g216),.DATA(g30513));
  MSFF DFF_226(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g219),.DATA(g30514));
  MSFF DFF_227(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g258),.DATA(g30518));
  MSFF DFF_228(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g261),.DATA(g30519));
  MSFF DFF_229(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g264),.DATA(g30520));
  MSFF DFF_230(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g222),.DATA(g30839));
  MSFF DFF_231(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g225),.DATA(g30840));
  MSFF DFF_232(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g228),.DATA(g30841));
  MSFF DFF_233(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g267),.DATA(g30848));
  MSFF DFF_234(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g270),.DATA(g30849));
  MSFF DFF_235(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g273),.DATA(g30850));
  MSFF DFF_236(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g92),.DATA(g25983));
  MSFF DFF_237(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g88),.DATA(g26678));
  MSFF DFF_238(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g83),.DATA(g27189));
  MSFF DFF_239(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g79),.DATA(g27683));
  MSFF DFF_240(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g74),.DATA(g28206));
  MSFF DFF_241(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g70),.DATA(g28673));
  MSFF DFF_242(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g65),.DATA(g29131));
  MSFF DFF_243(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g61),.DATA(g29413));
  MSFF DFF_244(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g56),.DATA(g29627));
  MSFF DFF_245(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g52),.DATA(g29794));
  MSFF DFF_246(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g180),.DATA(g20555));
  MSFF DFF_247(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g182),.DATA(g180));
  MSFF DFF_248(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g181),.DATA(g182));
  MSFF DFF_249(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g276),.DATA(g13406));
  MSFF DFF_250(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g405),.DATA(g276));
  MSFF DFF_251(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g401),.DATA(g405));
  MSFF DFF_252(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g309),.DATA(g11496));
  MSFF DFF_253(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g354),.DATA(g28207));
  MSFF DFF_254(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g343),.DATA(g28208));
  MSFF DFF_255(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g346),.DATA(g28209));
  MSFF DFF_256(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g369),.DATA(g28210));
  MSFF DFF_257(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g358),.DATA(g28211));
  MSFF DFF_258(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g361),.DATA(g28212));
  MSFF DFF_259(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g384),.DATA(g28213));
  MSFF DFF_260(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g373),.DATA(g28214));
  MSFF DFF_261(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g376),.DATA(g28215));
  MSFF DFF_262(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g398),.DATA(g28216));
  MSFF DFF_263(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g388),.DATA(g28217));
  MSFF DFF_264(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g391),.DATA(g28218));
  MSFF DFF_265(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g408),.DATA(g29414));
  MSFF DFF_266(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g411),.DATA(g29415));
  MSFF DFF_267(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g414),.DATA(g29416));
  MSFF DFF_268(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g417),.DATA(g29631));
  MSFF DFF_269(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g420),.DATA(g29632));
  MSFF DFF_270(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g423),.DATA(g29633));
  MSFF DFF_271(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g427),.DATA(g29417));
  MSFF DFF_272(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g428),.DATA(g29418));
  MSFF DFF_273(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g426),.DATA(g29419));
  MSFF DFF_274(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g429),.DATA(g27684));
  MSFF DFF_275(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g432),.DATA(g27685));
  MSFF DFF_276(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g435),.DATA(g27686));
  MSFF DFF_277(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g438),.DATA(g27687));
  MSFF DFF_278(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g441),.DATA(g27688));
  MSFF DFF_279(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g444),.DATA(g27689));
  MSFF DFF_280(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g448),.DATA(g28674));
  MSFF DFF_281(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g449),.DATA(g28675));
  MSFF DFF_282(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g447),.DATA(g28676));
  MSFF DFF_283(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g312),.DATA(g29795));
  MSFF DFF_284(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g313),.DATA(g29796));
  MSFF DFF_285(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g314),.DATA(g29797));
  MSFF DFF_286(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g315),.DATA(g30851));
  MSFF DFF_287(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g316),.DATA(g30852));
  MSFF DFF_288(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g317),.DATA(g30853));
  MSFF DFF_289(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g318),.DATA(g30710));
  MSFF DFF_290(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g319),.DATA(g30711));
  MSFF DFF_291(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g320),.DATA(g30712));
  MSFF DFF_292(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g322),.DATA(g29628));
  MSFF DFF_293(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g323),.DATA(g29629));
  MSFF DFF_294(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g321),.DATA(g29630));
  MSFF DFF_295(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g403),.DATA(g27191));
  MSFF DFF_296(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g404),.DATA(g27192));
  MSFF DFF_297(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g402),.DATA(g27193));
  MSFF DFF_298(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g450),.DATA(g11509));
  MSFF DFF_299(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g451),.DATA(g450));
  MSFF DFF_300(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g452),.DATA(g11510));
  MSFF DFF_301(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g453),.DATA(g452));
  MSFF DFF_302(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g454),.DATA(g11511));
  MSFF DFF_303(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g279),.DATA(g454));
  MSFF DFF_304(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g280),.DATA(g11491));
  MSFF DFF_305(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g281),.DATA(g280));
  MSFF DFF_306(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g282),.DATA(g11492));
  MSFF DFF_307(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g283),.DATA(g282));
  MSFF DFF_308(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g284),.DATA(g11493));
  MSFF DFF_309(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g285),.DATA(g284));
  MSFF DFF_310(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g286),.DATA(g11494));
  MSFF DFF_311(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g287),.DATA(g286));
  MSFF DFF_312(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g288),.DATA(g11495));
  MSFF DFF_313(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g289),.DATA(g288));
  MSFF DFF_314(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g290),.DATA(g13407));
  MSFF DFF_315(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g291),.DATA(g290));
  MSFF DFF_316(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g299),.DATA(g19012));
  MSFF DFF_317(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g305),.DATA(g23148));
  MSFF DFF_318(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g308),.DATA(g23149));
  MSFF DFF_319(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g297),.DATA(g23150));
  MSFF DFF_320(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g296),.DATA(g23151));
  MSFF DFF_321(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g295),.DATA(g23152));
  MSFF DFF_322(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g294),.DATA(g23153));
  MSFF DFF_323(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g304),.DATA(g19016));
  MSFF DFF_324(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g303),.DATA(g19015));
  MSFF DFF_325(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g302),.DATA(g19014));
  MSFF DFF_326(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g301),.DATA(g19013));
  MSFF DFF_327(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g300),.DATA(g25130));
  MSFF DFF_328(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g298),.DATA(g27190));
  MSFF DFF_329(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g342),.DATA(g11497));
  MSFF DFF_330(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g349),.DATA(g342));
  MSFF DFF_331(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g350),.DATA(g11498));
  MSFF DFF_332(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g351),.DATA(g350));
  MSFF DFF_333(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g352),.DATA(g11499));
  MSFF DFF_334(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g353),.DATA(g352));
  MSFF DFF_335(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g357),.DATA(g11500));
  MSFF DFF_336(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g364),.DATA(g357));
  MSFF DFF_337(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g365),.DATA(g11501));
  MSFF DFF_338(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g366),.DATA(g365));
  MSFF DFF_339(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g367),.DATA(g11502));
  MSFF DFF_340(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g368),.DATA(g367));
  MSFF DFF_341(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g372),.DATA(g11503));
  MSFF DFF_342(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g379),.DATA(g372));
  MSFF DFF_343(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g380),.DATA(g11504));
  MSFF DFF_344(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g381),.DATA(g380));
  MSFF DFF_345(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g382),.DATA(g11505));
  MSFF DFF_346(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g383),.DATA(g382));
  MSFF DFF_347(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g387),.DATA(g11506));
  MSFF DFF_348(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g394),.DATA(g387));
  MSFF DFF_349(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g395),.DATA(g11507));
  MSFF DFF_350(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g396),.DATA(g395));
  MSFF DFF_351(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g397),.DATA(g11508));
  MSFF DFF_352(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g324),.DATA(g397));
  MSFF DFF_353(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g325),.DATA(g13408));
  MSFF DFF_354(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g331),.DATA(g325));
  MSFF DFF_355(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g337),.DATA(g331));
  MSFF DFF_356(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g545),.DATA(g13419));
  MSFF DFF_357(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g551),.DATA(g545));
  MSFF DFF_358(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g550),.DATA(g551));
  MSFF DFF_359(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g554),.DATA(g23160));
  MSFF DFF_360(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g557),.DATA(g20556));
  MSFF DFF_361(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g510),.DATA(g20557));
  MSFF DFF_362(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g513),.DATA(g16467));
  MSFF DFF_363(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g523),.DATA(g513));
  MSFF DFF_364(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g524),.DATA(g523));
  MSFF DFF_365(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g564),.DATA(g11512));
  MSFF DFF_366(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g569),.DATA(g564));
  MSFF DFF_367(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g570),.DATA(g11515));
  MSFF DFF_368(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g571),.DATA(g570));
  MSFF DFF_369(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g572),.DATA(g11516));
  MSFF DFF_370(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g573),.DATA(g572));
  MSFF DFF_371(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g574),.DATA(g11517));
  MSFF DFF_372(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g565),.DATA(g574));
  MSFF DFF_373(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g566),.DATA(g11513));
  MSFF DFF_374(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g567),.DATA(g566));
  MSFF DFF_375(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g568),.DATA(g11514));
  MSFF DFF_376(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g489),.DATA(g568));
  MSFF DFF_377(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g474),.DATA(g13409));
  MSFF DFF_378(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g481),.DATA(g474));
  MSFF DFF_379(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g485),.DATA(g481));
  MSFF DFF_380(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g486),.DATA(g24292));
  MSFF DFF_381(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g487),.DATA(g24293));
  MSFF DFF_382(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g488),.DATA(g24294));
  MSFF DFF_383(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g455),.DATA(g25139));
  MSFF DFF_384(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g458),.DATA(g25131));
  MSFF DFF_385(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g461),.DATA(g25132));
  MSFF DFF_386(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g477),.DATA(g25136));
  MSFF DFF_387(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g478),.DATA(g25137));
  MSFF DFF_388(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g479),.DATA(g25138));
  MSFF DFF_389(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g480),.DATA(g24289));
  MSFF DFF_390(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g484),.DATA(g24290));
  MSFF DFF_391(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g464),.DATA(g24291));
  MSFF DFF_392(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g465),.DATA(g25133));
  MSFF DFF_393(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g468),.DATA(g25134));
  MSFF DFF_394(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g471),.DATA(g25135));
  MSFF DFF_395(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g528),.DATA(g16468));
  MSFF DFF_396(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g535),.DATA(g528));
  MSFF DFF_397(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g542),.DATA(g535));
  MSFF DFF_398(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g543),.DATA(g19021));
  MSFF DFF_399(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g544),.DATA(g543));
  MSFF DFF_400(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g548),.DATA(g23159));
  MSFF DFF_401(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g549),.DATA(g19022));
  MSFF DFF_402(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g499),.DATA(g549));
  MSFF DFF_403(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g558),.DATA(g19023));
  MSFF DFF_404(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g559),.DATA(g558));
  MSFF DFF_405(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g576),.DATA(g28219));
  MSFF DFF_406(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g577),.DATA(g28220));
  MSFF DFF_407(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g575),.DATA(g28221));
  MSFF DFF_408(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g579),.DATA(g28222));
  MSFF DFF_409(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g580),.DATA(g28223));
  MSFF DFF_410(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g578),.DATA(g28224));
  MSFF DFF_411(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g582),.DATA(g28225));
  MSFF DFF_412(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g583),.DATA(g28226));
  MSFF DFF_413(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g581),.DATA(g28227));
  MSFF DFF_414(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g585),.DATA(g28228));
  MSFF DFF_415(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g586),.DATA(g28229));
  MSFF DFF_416(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g584),.DATA(g28230));
  MSFF DFF_417(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g587),.DATA(g25985));
  MSFF DFF_418(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g590),.DATA(g25986));
  MSFF DFF_419(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g593),.DATA(g25987));
  MSFF DFF_420(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g596),.DATA(g25988));
  MSFF DFF_421(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g599),.DATA(g25989));
  MSFF DFF_422(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g602),.DATA(g25990));
  MSFF DFF_423(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g614),.DATA(g29135));
  MSFF DFF_424(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g617),.DATA(g29136));
  MSFF DFF_425(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g620),.DATA(g29137));
  MSFF DFF_426(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g605),.DATA(g29132));
  MSFF DFF_427(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g608),.DATA(g29133));
  MSFF DFF_428(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g611),.DATA(g29134));
  MSFF DFF_429(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g490),.DATA(g27194));
  MSFF DFF_430(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g493),.DATA(g27195));
  MSFF DFF_431(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g496),.DATA(g27196));
  MSFF DFF_432(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g506),.DATA(g8284));
  MSFF DFF_433(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g507),.DATA(g24295));
  MSFF DFF_434(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g508),.DATA(g19017));
  MSFF DFF_435(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g509),.DATA(g19018));
  MSFF DFF_436(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g514),.DATA(g19019));
  MSFF DFF_437(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g515),.DATA(g19020));
  MSFF DFF_438(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g516),.DATA(g23158));
  MSFF DFF_439(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g517),.DATA(g23157));
  MSFF DFF_440(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g518),.DATA(g23156));
  MSFF DFF_441(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g519),.DATA(g23155));
  MSFF DFF_442(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g520),.DATA(g23154));
  MSFF DFF_443(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g525),.DATA(g520));
  MSFF DFF_444(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g529),.DATA(g13410));
  MSFF DFF_445(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g530),.DATA(g13411));
  MSFF DFF_446(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g531),.DATA(g13412));
  MSFF DFF_447(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g532),.DATA(g13413));
  MSFF DFF_448(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g533),.DATA(g13414));
  MSFF DFF_449(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g534),.DATA(g13415));
  MSFF DFF_450(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g536),.DATA(g13416));
  MSFF DFF_451(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g537),.DATA(g13417));
  MSFF DFF_452(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g538),.DATA(g25984));
  MSFF DFF_453(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g541),.DATA(g13418));
  MSFF DFF_454(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g623),.DATA(g13420));
  MSFF DFF_455(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g626),.DATA(g623));
  MSFF DFF_456(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g629),.DATA(g626));
  MSFF DFF_457(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g630),.DATA(g20558));
  MSFF DFF_458(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g659),.DATA(g21943));
  MSFF DFF_459(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g640),.DATA(g23161));
  MSFF DFF_460(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g633),.DATA(g24296));
  MSFF DFF_461(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g653),.DATA(g25140));
  MSFF DFF_462(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g646),.DATA(g25991));
  MSFF DFF_463(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g660),.DATA(g26691));
  MSFF DFF_464(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g672),.DATA(g27197));
  MSFF DFF_465(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g666),.DATA(g27690));
  MSFF DFF_466(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g679),.DATA(g28231));
  MSFF DFF_467(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g686),.DATA(g28677));
  MSFF DFF_468(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g692),.DATA(g29138));
  MSFF DFF_469(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g699),.DATA(g23162));
  MSFF DFF_470(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g700),.DATA(g23163));
  MSFF DFF_471(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g698),.DATA(g23164));
  MSFF DFF_472(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g702),.DATA(g23165));
  MSFF DFF_473(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g703),.DATA(g23166));
  MSFF DFF_474(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g701),.DATA(g23167));
  MSFF DFF_475(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g705),.DATA(g23168));
  MSFF DFF_476(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g706),.DATA(g23169));
  MSFF DFF_477(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g704),.DATA(g23170));
  MSFF DFF_478(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g708),.DATA(g23171));
  MSFF DFF_479(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g709),.DATA(g23172));
  MSFF DFF_480(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g707),.DATA(g23173));
  MSFF DFF_481(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g711),.DATA(g23174));
  MSFF DFF_482(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g712),.DATA(g23175));
  MSFF DFF_483(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g710),.DATA(g23176));
  MSFF DFF_484(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g714),.DATA(g23177));
  MSFF DFF_485(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g715),.DATA(g23178));
  MSFF DFF_486(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g713),.DATA(g23179));
  MSFF DFF_487(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g717),.DATA(g23180));
  MSFF DFF_488(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g718),.DATA(g23181));
  MSFF DFF_489(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g716),.DATA(g23182));
  MSFF DFF_490(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g720),.DATA(g23183));
  MSFF DFF_491(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g721),.DATA(g23184));
  MSFF DFF_492(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g719),.DATA(g23185));
  MSFF DFF_493(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g723),.DATA(g23186));
  MSFF DFF_494(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g724),.DATA(g23187));
  MSFF DFF_495(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g722),.DATA(g23188));
  MSFF DFF_496(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g726),.DATA(g23189));
  MSFF DFF_497(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g727),.DATA(g23190));
  MSFF DFF_498(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g725),.DATA(g23191));
  MSFF DFF_499(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g729),.DATA(g23192));
  MSFF DFF_500(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g730),.DATA(g23193));
  MSFF DFF_501(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g728),.DATA(g23194));
  MSFF DFF_502(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g732),.DATA(g23195));
  MSFF DFF_503(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g733),.DATA(g23196));
  MSFF DFF_504(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g731),.DATA(g23197));
  MSFF DFF_505(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g735),.DATA(g26692));
  MSFF DFF_506(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g736),.DATA(g26693));
  MSFF DFF_507(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g734),.DATA(g26694));
  MSFF DFF_508(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g738),.DATA(g24297));
  MSFF DFF_509(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g739),.DATA(g24298));
  MSFF DFF_510(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g737),.DATA(g24299));
  MSFF DFF_511(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g826),.DATA(g13421));
  MSFF DFF_512(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g823),.DATA(g826));
  MSFF DFF_513(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g853),.DATA(g823));
  MSFF DFF_514(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g818),.DATA(g24300));
  MSFF DFF_515(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g819),.DATA(g24301));
  MSFF DFF_516(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g817),.DATA(g24302));
  MSFF DFF_517(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g821),.DATA(g24303));
  MSFF DFF_518(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g822),.DATA(g24304));
  MSFF DFF_519(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g820),.DATA(g24305));
  MSFF DFF_520(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g830),.DATA(g24306));
  MSFF DFF_521(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g831),.DATA(g24307));
  MSFF DFF_522(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g829),.DATA(g24308));
  MSFF DFF_523(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g833),.DATA(g24309));
  MSFF DFF_524(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g834),.DATA(g24310));
  MSFF DFF_525(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g832),.DATA(g24311));
  MSFF DFF_526(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g836),.DATA(g24312));
  MSFF DFF_527(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g837),.DATA(g24313));
  MSFF DFF_528(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g835),.DATA(g24314));
  MSFF DFF_529(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g839),.DATA(g24315));
  MSFF DFF_530(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g840),.DATA(g24316));
  MSFF DFF_531(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g838),.DATA(g24317));
  MSFF DFF_532(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g842),.DATA(g24318));
  MSFF DFF_533(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g843),.DATA(g24319));
  MSFF DFF_534(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g841),.DATA(g24320));
  MSFF DFF_535(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g845),.DATA(g24321));
  MSFF DFF_536(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g846),.DATA(g24322));
  MSFF DFF_537(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g844),.DATA(g24323));
  MSFF DFF_538(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g848),.DATA(g24324));
  MSFF DFF_539(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g849),.DATA(g24325));
  MSFF DFF_540(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g847),.DATA(g24326));
  MSFF DFF_541(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g851),.DATA(g24327));
  MSFF DFF_542(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g852),.DATA(g24328));
  MSFF DFF_543(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g850),.DATA(g24329));
  MSFF DFF_544(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g857),.DATA(g26696));
  MSFF DFF_545(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g858),.DATA(g26697));
  MSFF DFF_546(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g856),.DATA(g26698));
  MSFF DFF_547(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g860),.DATA(g26699));
  MSFF DFF_548(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g861),.DATA(g26700));
  MSFF DFF_549(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g859),.DATA(g26701));
  MSFF DFF_550(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g863),.DATA(g26702));
  MSFF DFF_551(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g864),.DATA(g26703));
  MSFF DFF_552(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g862),.DATA(g26704));
  MSFF DFF_553(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g866),.DATA(g26705));
  MSFF DFF_554(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g867),.DATA(g26706));
  MSFF DFF_555(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g865),.DATA(g26707));
  MSFF DFF_556(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g873),.DATA(g30521));
  MSFF DFF_557(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g876),.DATA(g30522));
  MSFF DFF_558(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g879),.DATA(g30523));
  MSFF DFF_559(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g918),.DATA(g30860));
  MSFF DFF_560(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g921),.DATA(g30861));
  MSFF DFF_561(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g924),.DATA(g30862));
  MSFF DFF_562(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g882),.DATA(g30854));
  MSFF DFF_563(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g885),.DATA(g30855));
  MSFF DFF_564(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g888),.DATA(g30856));
  MSFF DFF_565(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g927),.DATA(g30863));
  MSFF DFF_566(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g930),.DATA(g30864));
  MSFF DFF_567(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g933),.DATA(g30865));
  MSFF DFF_568(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g891),.DATA(g30524));
  MSFF DFF_569(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g894),.DATA(g30525));
  MSFF DFF_570(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g897),.DATA(g30526));
  MSFF DFF_571(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g936),.DATA(g30530));
  MSFF DFF_572(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g939),.DATA(g30531));
  MSFF DFF_573(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g942),.DATA(g30532));
  MSFF DFF_574(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g900),.DATA(g30527));
  MSFF DFF_575(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g903),.DATA(g30528));
  MSFF DFF_576(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g906),.DATA(g30529));
  MSFF DFF_577(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g945),.DATA(g30533));
  MSFF DFF_578(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g948),.DATA(g30534));
  MSFF DFF_579(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g951),.DATA(g30535));
  MSFF DFF_580(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g909),.DATA(g30857));
  MSFF DFF_581(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g912),.DATA(g30858));
  MSFF DFF_582(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g915),.DATA(g30859));
  MSFF DFF_583(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g954),.DATA(g30866));
  MSFF DFF_584(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g957),.DATA(g30867));
  MSFF DFF_585(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g960),.DATA(g30868));
  MSFF DFF_586(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g780),.DATA(g25992));
  MSFF DFF_587(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g776),.DATA(g26695));
  MSFF DFF_588(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g771),.DATA(g27198));
  MSFF DFF_589(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g767),.DATA(g27691));
  MSFF DFF_590(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g762),.DATA(g28232));
  MSFF DFF_591(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g758),.DATA(g28678));
  MSFF DFF_592(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g753),.DATA(g29139));
  MSFF DFF_593(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g749),.DATA(g29420));
  MSFF DFF_594(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g744),.DATA(g29634));
  MSFF DFF_595(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g740),.DATA(g29798));
  MSFF DFF_596(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g868),.DATA(g20559));
  MSFF DFF_597(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g870),.DATA(g868));
  MSFF DFF_598(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g869),.DATA(g870));
  MSFF DFF_599(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g963),.DATA(g13422));
  MSFF DFF_600(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1092),.DATA(g963));
  MSFF DFF_601(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1088),.DATA(g1092));
  MSFF DFF_602(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g996),.DATA(g11523));
  MSFF DFF_603(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1041),.DATA(g28233));
  MSFF DFF_604(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1030),.DATA(g28234));
  MSFF DFF_605(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1033),.DATA(g28235));
  MSFF DFF_606(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1056),.DATA(g28236));
  MSFF DFF_607(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1045),.DATA(g28237));
  MSFF DFF_608(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1048),.DATA(g28238));
  MSFF DFF_609(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1071),.DATA(g28239));
  MSFF DFF_610(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1060),.DATA(g28240));
  MSFF DFF_611(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1063),.DATA(g28241));
  MSFF DFF_612(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1085),.DATA(g28242));
  MSFF DFF_613(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1075),.DATA(g28243));
  MSFF DFF_614(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1078),.DATA(g28244));
  MSFF DFF_615(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1095),.DATA(g29421));
  MSFF DFF_616(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1098),.DATA(g29422));
  MSFF DFF_617(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1101),.DATA(g29423));
  MSFF DFF_618(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1104),.DATA(g29638));
  MSFF DFF_619(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1107),.DATA(g29639));
  MSFF DFF_620(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1110),.DATA(g29640));
  MSFF DFF_621(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1114),.DATA(g29424));
  MSFF DFF_622(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1115),.DATA(g29425));
  MSFF DFF_623(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1113),.DATA(g29426));
  MSFF DFF_624(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1116),.DATA(g27692));
  MSFF DFF_625(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1119),.DATA(g27693));
  MSFF DFF_626(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1122),.DATA(g27694));
  MSFF DFF_627(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1125),.DATA(g27695));
  MSFF DFF_628(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1128),.DATA(g27696));
  MSFF DFF_629(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1131),.DATA(g27697));
  MSFF DFF_630(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1135),.DATA(g28679));
  MSFF DFF_631(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1136),.DATA(g28680));
  MSFF DFF_632(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1134),.DATA(g28681));
  MSFF DFF_633(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g999),.DATA(g29799));
  MSFF DFF_634(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1000),.DATA(g29800));
  MSFF DFF_635(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1001),.DATA(g29801));
  MSFF DFF_636(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1002),.DATA(g30869));
  MSFF DFF_637(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1003),.DATA(g30870));
  MSFF DFF_638(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1004),.DATA(g30871));
  MSFF DFF_639(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1005),.DATA(g30713));
  MSFF DFF_640(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1006),.DATA(g30714));
  MSFF DFF_641(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1007),.DATA(g30715));
  MSFF DFF_642(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1009),.DATA(g29635));
  MSFF DFF_643(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1010),.DATA(g29636));
  MSFF DFF_644(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1008),.DATA(g29637));
  MSFF DFF_645(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1090),.DATA(g27206));
  MSFF DFF_646(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1091),.DATA(g27207));
  MSFF DFF_647(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1089),.DATA(g27208));
  MSFF DFF_648(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1137),.DATA(g11536));
  MSFF DFF_649(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1138),.DATA(g1137));
  MSFF DFF_650(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1139),.DATA(g11537));
  MSFF DFF_651(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1140),.DATA(g1139));
  MSFF DFF_652(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1141),.DATA(g11538));
  MSFF DFF_653(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g966),.DATA(g1141));
  MSFF DFF_654(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g967),.DATA(g11518));
  MSFF DFF_655(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g968),.DATA(g967));
  MSFF DFF_656(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g969),.DATA(g11519));
  MSFF DFF_657(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g970),.DATA(g969));
  MSFF DFF_658(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g971),.DATA(g11520));
  MSFF DFF_659(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g972),.DATA(g971));
  MSFF DFF_660(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g973),.DATA(g11521));
  MSFF DFF_661(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g974),.DATA(g973));
  MSFF DFF_662(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g975),.DATA(g11522));
  MSFF DFF_663(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g976),.DATA(g975));
  MSFF DFF_664(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g977),.DATA(g13423));
  MSFF DFF_665(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g978),.DATA(g977));
  MSFF DFF_666(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g986),.DATA(g19024));
  MSFF DFF_667(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g992),.DATA(g27200));
  MSFF DFF_668(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g995),.DATA(g27201));
  MSFF DFF_669(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g984),.DATA(g27202));
  MSFF DFF_670(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g983),.DATA(g27203));
  MSFF DFF_671(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g982),.DATA(g27204));
  MSFF DFF_672(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g981),.DATA(g27205));
  MSFF DFF_673(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g991),.DATA(g19028));
  MSFF DFF_674(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g990),.DATA(g19027));
  MSFF DFF_675(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g989),.DATA(g19026));
  MSFF DFF_676(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g988),.DATA(g19025));
  MSFF DFF_677(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g987),.DATA(g25141));
  MSFF DFF_678(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g985),.DATA(g27199));
  MSFF DFF_679(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1029),.DATA(g11524));
  MSFF DFF_680(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1036),.DATA(g1029));
  MSFF DFF_681(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1037),.DATA(g11525));
  MSFF DFF_682(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1038),.DATA(g1037));
  MSFF DFF_683(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1039),.DATA(g11526));
  MSFF DFF_684(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1040),.DATA(g1039));
  MSFF DFF_685(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1044),.DATA(g11527));
  MSFF DFF_686(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1051),.DATA(g1044));
  MSFF DFF_687(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1052),.DATA(g11528));
  MSFF DFF_688(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1053),.DATA(g1052));
  MSFF DFF_689(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1054),.DATA(g11529));
  MSFF DFF_690(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1055),.DATA(g1054));
  MSFF DFF_691(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1059),.DATA(g11530));
  MSFF DFF_692(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1066),.DATA(g1059));
  MSFF DFF_693(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1067),.DATA(g11531));
  MSFF DFF_694(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1068),.DATA(g1067));
  MSFF DFF_695(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1069),.DATA(g11532));
  MSFF DFF_696(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1070),.DATA(g1069));
  MSFF DFF_697(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1074),.DATA(g11533));
  MSFF DFF_698(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1081),.DATA(g1074));
  MSFF DFF_699(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1082),.DATA(g11534));
  MSFF DFF_700(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1083),.DATA(g1082));
  MSFF DFF_701(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1084),.DATA(g11535));
  MSFF DFF_702(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1011),.DATA(g1084));
  MSFF DFF_703(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1012),.DATA(g13424));
  MSFF DFF_704(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1018),.DATA(g1012));
  MSFF DFF_705(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1024),.DATA(g1018));
  MSFF DFF_706(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1231),.DATA(g13435));
  MSFF DFF_707(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1237),.DATA(g1231));
  MSFF DFF_708(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1236),.DATA(g1237));
  MSFF DFF_709(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1240),.DATA(g23198));
  MSFF DFF_710(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1243),.DATA(g20560));
  MSFF DFF_711(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1196),.DATA(g20561));
  MSFF DFF_712(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1199),.DATA(g16469));
  MSFF DFF_713(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1209),.DATA(g1199));
  MSFF DFF_714(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1210),.DATA(g1209));
  MSFF DFF_715(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1250),.DATA(g11539));
  MSFF DFF_716(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1255),.DATA(g1250));
  MSFF DFF_717(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1256),.DATA(g11542));
  MSFF DFF_718(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1257),.DATA(g1256));
  MSFF DFF_719(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1258),.DATA(g11543));
  MSFF DFF_720(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1259),.DATA(g1258));
  MSFF DFF_721(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1260),.DATA(g11544));
  MSFF DFF_722(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1251),.DATA(g1260));
  MSFF DFF_723(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1252),.DATA(g11540));
  MSFF DFF_724(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1253),.DATA(g1252));
  MSFF DFF_725(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1254),.DATA(g11541));
  MSFF DFF_726(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1176),.DATA(g1254));
  MSFF DFF_727(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1161),.DATA(g13425));
  MSFF DFF_728(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1168),.DATA(g1161));
  MSFF DFF_729(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1172),.DATA(g1168));
  MSFF DFF_730(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1173),.DATA(g24333));
  MSFF DFF_731(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1174),.DATA(g24334));
  MSFF DFF_732(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1175),.DATA(g24335));
  MSFF DFF_733(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1142),.DATA(g25150));
  MSFF DFF_734(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1145),.DATA(g25142));
  MSFF DFF_735(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1148),.DATA(g25143));
  MSFF DFF_736(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1164),.DATA(g25147));
  MSFF DFF_737(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1165),.DATA(g25148));
  MSFF DFF_738(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1166),.DATA(g25149));
  MSFF DFF_739(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1167),.DATA(g24330));
  MSFF DFF_740(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1171),.DATA(g24331));
  MSFF DFF_741(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1151),.DATA(g24332));
  MSFF DFF_742(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1152),.DATA(g25144));
  MSFF DFF_743(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1155),.DATA(g25145));
  MSFF DFF_744(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1158),.DATA(g25146));
  MSFF DFF_745(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1214),.DATA(g16470));
  MSFF DFF_746(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1221),.DATA(g1214));
  MSFF DFF_747(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1228),.DATA(g1221));
  MSFF DFF_748(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1229),.DATA(g19033));
  MSFF DFF_749(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1230),.DATA(g1229));
  MSFF DFF_750(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1234),.DATA(g27217));
  MSFF DFF_751(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1235),.DATA(g19034));
  MSFF DFF_752(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1186),.DATA(g1235));
  MSFF DFF_753(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1244),.DATA(g19035));
  MSFF DFF_754(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1245),.DATA(g1244));
  MSFF DFF_755(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1262),.DATA(g28245));
  MSFF DFF_756(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1263),.DATA(g28246));
  MSFF DFF_757(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1261),.DATA(g28247));
  MSFF DFF_758(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1265),.DATA(g28248));
  MSFF DFF_759(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1266),.DATA(g28249));
  MSFF DFF_760(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1264),.DATA(g28250));
  MSFF DFF_761(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1268),.DATA(g28251));
  MSFF DFF_762(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1269),.DATA(g28252));
  MSFF DFF_763(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1267),.DATA(g28253));
  MSFF DFF_764(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1271),.DATA(g28254));
  MSFF DFF_765(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1272),.DATA(g28255));
  MSFF DFF_766(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1270),.DATA(g28256));
  MSFF DFF_767(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1273),.DATA(g25994));
  MSFF DFF_768(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1276),.DATA(g25995));
  MSFF DFF_769(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1279),.DATA(g25996));
  MSFF DFF_770(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1282),.DATA(g25997));
  MSFF DFF_771(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1285),.DATA(g25998));
  MSFF DFF_772(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1288),.DATA(g25999));
  MSFF DFF_773(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1300),.DATA(g29143));
  MSFF DFF_774(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1303),.DATA(g29144));
  MSFF DFF_775(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1306),.DATA(g29145));
  MSFF DFF_776(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1291),.DATA(g29140));
  MSFF DFF_777(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1294),.DATA(g29141));
  MSFF DFF_778(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1297),.DATA(g29142));
  MSFF DFF_779(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1177),.DATA(g27209));
  MSFF DFF_780(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1180),.DATA(g27210));
  MSFF DFF_781(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1183),.DATA(g27211));
  MSFF DFF_782(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1192),.DATA(g8293));
  MSFF DFF_783(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1193),.DATA(g24336));
  MSFF DFF_784(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1194),.DATA(g19029));
  MSFF DFF_785(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1195),.DATA(g19030));
  MSFF DFF_786(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1200),.DATA(g19031));
  MSFF DFF_787(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1201),.DATA(g19032));
  MSFF DFF_788(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1202),.DATA(g27216));
  MSFF DFF_789(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1203),.DATA(g27215));
  MSFF DFF_790(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1204),.DATA(g27214));
  MSFF DFF_791(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1205),.DATA(g27213));
  MSFF DFF_792(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1206),.DATA(g27212));
  MSFF DFF_793(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1211),.DATA(g1206));
  MSFF DFF_794(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1215),.DATA(g13426));
  MSFF DFF_795(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1216),.DATA(g13427));
  MSFF DFF_796(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1217),.DATA(g13428));
  MSFF DFF_797(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1218),.DATA(g13429));
  MSFF DFF_798(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1219),.DATA(g13430));
  MSFF DFF_799(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1220),.DATA(g13431));
  MSFF DFF_800(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1222),.DATA(g13432));
  MSFF DFF_801(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1223),.DATA(g13433));
  MSFF DFF_802(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1224),.DATA(g25993));
  MSFF DFF_803(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1227),.DATA(g13434));
  MSFF DFF_804(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1309),.DATA(g13436));
  MSFF DFF_805(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1312),.DATA(g1309));
  MSFF DFF_806(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1315),.DATA(g1312));
  MSFF DFF_807(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1316),.DATA(g20562));
  MSFF DFF_808(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1345),.DATA(g21944));
  MSFF DFF_809(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1326),.DATA(g23199));
  MSFF DFF_810(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1319),.DATA(g24337));
  MSFF DFF_811(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1339),.DATA(g25151));
  MSFF DFF_812(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1332),.DATA(g26000));
  MSFF DFF_813(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1346),.DATA(g26708));
  MSFF DFF_814(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1358),.DATA(g27218));
  MSFF DFF_815(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1352),.DATA(g27698));
  MSFF DFF_816(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1365),.DATA(g28257));
  MSFF DFF_817(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1372),.DATA(g28682));
  MSFF DFF_818(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1378),.DATA(g29146));
  MSFF DFF_819(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1385),.DATA(g23200));
  MSFF DFF_820(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1386),.DATA(g23201));
  MSFF DFF_821(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1384),.DATA(g23202));
  MSFF DFF_822(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1388),.DATA(g23203));
  MSFF DFF_823(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1389),.DATA(g23204));
  MSFF DFF_824(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1387),.DATA(g23205));
  MSFF DFF_825(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1391),.DATA(g23206));
  MSFF DFF_826(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1392),.DATA(g23207));
  MSFF DFF_827(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1390),.DATA(g23208));
  MSFF DFF_828(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1394),.DATA(g23209));
  MSFF DFF_829(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1395),.DATA(g23210));
  MSFF DFF_830(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1393),.DATA(g23211));
  MSFF DFF_831(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1397),.DATA(g23212));
  MSFF DFF_832(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1398),.DATA(g23213));
  MSFF DFF_833(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1396),.DATA(g23214));
  MSFF DFF_834(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1400),.DATA(g23215));
  MSFF DFF_835(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1401),.DATA(g23216));
  MSFF DFF_836(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1399),.DATA(g23217));
  MSFF DFF_837(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1403),.DATA(g23218));
  MSFF DFF_838(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1404),.DATA(g23219));
  MSFF DFF_839(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1402),.DATA(g23220));
  MSFF DFF_840(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1406),.DATA(g23221));
  MSFF DFF_841(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1407),.DATA(g23222));
  MSFF DFF_842(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1405),.DATA(g23223));
  MSFF DFF_843(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1409),.DATA(g23224));
  MSFF DFF_844(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1410),.DATA(g23225));
  MSFF DFF_845(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1408),.DATA(g23226));
  MSFF DFF_846(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1412),.DATA(g23227));
  MSFF DFF_847(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1413),.DATA(g23228));
  MSFF DFF_848(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1411),.DATA(g23229));
  MSFF DFF_849(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1415),.DATA(g23230));
  MSFF DFF_850(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1416),.DATA(g23231));
  MSFF DFF_851(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1414),.DATA(g23232));
  MSFF DFF_852(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1418),.DATA(g23233));
  MSFF DFF_853(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1419),.DATA(g23234));
  MSFF DFF_854(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1417),.DATA(g23235));
  MSFF DFF_855(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1421),.DATA(g26709));
  MSFF DFF_856(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1422),.DATA(g26710));
  MSFF DFF_857(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1420),.DATA(g26711));
  MSFF DFF_858(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1424),.DATA(g24338));
  MSFF DFF_859(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1425),.DATA(g24339));
  MSFF DFF_860(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1423),.DATA(g24340));
  MSFF DFF_861(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1520),.DATA(g13437));
  MSFF DFF_862(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1517),.DATA(g1520));
  MSFF DFF_863(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1547),.DATA(g1517));
  MSFF DFF_864(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1512),.DATA(g24341));
  MSFF DFF_865(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1513),.DATA(g24342));
  MSFF DFF_866(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1511),.DATA(g24343));
  MSFF DFF_867(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1515),.DATA(g24344));
  MSFF DFF_868(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1516),.DATA(g24345));
  MSFF DFF_869(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1514),.DATA(g24346));
  MSFF DFF_870(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1524),.DATA(g24347));
  MSFF DFF_871(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1525),.DATA(g24348));
  MSFF DFF_872(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1523),.DATA(g24349));
  MSFF DFF_873(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1527),.DATA(g24350));
  MSFF DFF_874(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1528),.DATA(g24351));
  MSFF DFF_875(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1526),.DATA(g24352));
  MSFF DFF_876(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1530),.DATA(g24353));
  MSFF DFF_877(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1531),.DATA(g24354));
  MSFF DFF_878(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1529),.DATA(g24355));
  MSFF DFF_879(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1533),.DATA(g24356));
  MSFF DFF_880(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1534),.DATA(g24357));
  MSFF DFF_881(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1532),.DATA(g24358));
  MSFF DFF_882(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1536),.DATA(g24359));
  MSFF DFF_883(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1537),.DATA(g24360));
  MSFF DFF_884(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1535),.DATA(g24361));
  MSFF DFF_885(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1539),.DATA(g24362));
  MSFF DFF_886(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1540),.DATA(g24363));
  MSFF DFF_887(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1538),.DATA(g24364));
  MSFF DFF_888(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1542),.DATA(g24365));
  MSFF DFF_889(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1543),.DATA(g24366));
  MSFF DFF_890(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1541),.DATA(g24367));
  MSFF DFF_891(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1545),.DATA(g24368));
  MSFF DFF_892(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1546),.DATA(g24369));
  MSFF DFF_893(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1544),.DATA(g24370));
  MSFF DFF_894(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1551),.DATA(g26713));
  MSFF DFF_895(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1552),.DATA(g26714));
  MSFF DFF_896(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1550),.DATA(g26715));
  MSFF DFF_897(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1554),.DATA(g26716));
  MSFF DFF_898(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1555),.DATA(g26717));
  MSFF DFF_899(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1553),.DATA(g26718));
  MSFF DFF_900(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1557),.DATA(g26719));
  MSFF DFF_901(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1558),.DATA(g26720));
  MSFF DFF_902(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1556),.DATA(g26721));
  MSFF DFF_903(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1560),.DATA(g26722));
  MSFF DFF_904(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1561),.DATA(g26723));
  MSFF DFF_905(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1559),.DATA(g26724));
  MSFF DFF_906(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1567),.DATA(g30536));
  MSFF DFF_907(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1570),.DATA(g30537));
  MSFF DFF_908(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1573),.DATA(g30538));
  MSFF DFF_909(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1612),.DATA(g30878));
  MSFF DFF_910(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1615),.DATA(g30879));
  MSFF DFF_911(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1618),.DATA(g30880));
  MSFF DFF_912(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1576),.DATA(g30872));
  MSFF DFF_913(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1579),.DATA(g30873));
  MSFF DFF_914(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1582),.DATA(g30874));
  MSFF DFF_915(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1621),.DATA(g30881));
  MSFF DFF_916(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1624),.DATA(g30882));
  MSFF DFF_917(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1627),.DATA(g30883));
  MSFF DFF_918(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1585),.DATA(g30539));
  MSFF DFF_919(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1588),.DATA(g30540));
  MSFF DFF_920(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1591),.DATA(g30541));
  MSFF DFF_921(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1630),.DATA(g30545));
  MSFF DFF_922(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1633),.DATA(g30546));
  MSFF DFF_923(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1636),.DATA(g30547));
  MSFF DFF_924(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1594),.DATA(g30542));
  MSFF DFF_925(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1597),.DATA(g30543));
  MSFF DFF_926(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1600),.DATA(g30544));
  MSFF DFF_927(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1639),.DATA(g30548));
  MSFF DFF_928(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1642),.DATA(g30549));
  MSFF DFF_929(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1645),.DATA(g30550));
  MSFF DFF_930(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1603),.DATA(g30875));
  MSFF DFF_931(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1606),.DATA(g30876));
  MSFF DFF_932(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1609),.DATA(g30877));
  MSFF DFF_933(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1648),.DATA(g30884));
  MSFF DFF_934(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1651),.DATA(g30885));
  MSFF DFF_935(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1654),.DATA(g30886));
  MSFF DFF_936(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1466),.DATA(g26001));
  MSFF DFF_937(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1462),.DATA(g26712));
  MSFF DFF_938(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1457),.DATA(g27219));
  MSFF DFF_939(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1453),.DATA(g27699));
  MSFF DFF_940(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1448),.DATA(g28258));
  MSFF DFF_941(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1444),.DATA(g28683));
  MSFF DFF_942(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1439),.DATA(g29147));
  MSFF DFF_943(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1435),.DATA(g29427));
  MSFF DFF_944(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1430),.DATA(g29641));
  MSFF DFF_945(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1426),.DATA(g29802));
  MSFF DFF_946(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1562),.DATA(g20563));
  MSFF DFF_947(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1564),.DATA(g1562));
  MSFF DFF_948(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1563),.DATA(g1564));
  MSFF DFF_949(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1657),.DATA(g13438));
  MSFF DFF_950(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1786),.DATA(g1657));
  MSFF DFF_951(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1782),.DATA(g1786));
  MSFF DFF_952(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1690),.DATA(g11550));
  MSFF DFF_953(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1735),.DATA(g28259));
  MSFF DFF_954(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1724),.DATA(g28260));
  MSFF DFF_955(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1727),.DATA(g28261));
  MSFF DFF_956(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1750),.DATA(g28262));
  MSFF DFF_957(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1739),.DATA(g28263));
  MSFF DFF_958(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1742),.DATA(g28264));
  MSFF DFF_959(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1765),.DATA(g28265));
  MSFF DFF_960(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1754),.DATA(g28266));
  MSFF DFF_961(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1757),.DATA(g28267));
  MSFF DFF_962(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1779),.DATA(g28268));
  MSFF DFF_963(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1769),.DATA(g28269));
  MSFF DFF_964(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1772),.DATA(g28270));
  MSFF DFF_965(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1789),.DATA(g29434));
  MSFF DFF_966(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1792),.DATA(g29435));
  MSFF DFF_967(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1795),.DATA(g29436));
  MSFF DFF_968(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1798),.DATA(g29645));
  MSFF DFF_969(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1801),.DATA(g29646));
  MSFF DFF_970(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1804),.DATA(g29647));
  MSFF DFF_971(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1808),.DATA(g29437));
  MSFF DFF_972(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1809),.DATA(g29438));
  MSFF DFF_973(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1807),.DATA(g29439));
  MSFF DFF_974(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1810),.DATA(g27700));
  MSFF DFF_975(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1813),.DATA(g27701));
  MSFF DFF_976(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1816),.DATA(g27702));
  MSFF DFF_977(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1819),.DATA(g27703));
  MSFF DFF_978(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1822),.DATA(g27704));
  MSFF DFF_979(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1825),.DATA(g27705));
  MSFF DFF_980(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1829),.DATA(g28684));
  MSFF DFF_981(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1830),.DATA(g28685));
  MSFF DFF_982(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1828),.DATA(g28686));
  MSFF DFF_983(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1693),.DATA(g29803));
  MSFF DFF_984(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1694),.DATA(g29804));
  MSFF DFF_985(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1695),.DATA(g29805));
  MSFF DFF_986(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1696),.DATA(g30887));
  MSFF DFF_987(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1697),.DATA(g30888));
  MSFF DFF_988(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1698),.DATA(g30889));
  MSFF DFF_989(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1699),.DATA(g30716));
  MSFF DFF_990(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1700),.DATA(g30717));
  MSFF DFF_991(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1701),.DATA(g30718));
  MSFF DFF_992(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1703),.DATA(g29642));
  MSFF DFF_993(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1704),.DATA(g29643));
  MSFF DFF_994(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1702),.DATA(g29644));
  MSFF DFF_995(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1784),.DATA(g27221));
  MSFF DFF_996(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1785),.DATA(g27222));
  MSFF DFF_997(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1783),.DATA(g27223));
  MSFF DFF_998(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1831),.DATA(g11563));
  MSFF DFF_999(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1832),.DATA(g1831));
  MSFF DFF_1000(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1833),.DATA(g11564));
  MSFF DFF_1001(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1834),.DATA(g1833));
  MSFF DFF_1002(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1835),.DATA(g11565));
  MSFF DFF_1003(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1660),.DATA(g1835));
  MSFF DFF_1004(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1661),.DATA(g11545));
  MSFF DFF_1005(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1662),.DATA(g1661));
  MSFF DFF_1006(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1663),.DATA(g11546));
  MSFF DFF_1007(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1664),.DATA(g1663));
  MSFF DFF_1008(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1665),.DATA(g11547));
  MSFF DFF_1009(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1666),.DATA(g1665));
  MSFF DFF_1010(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1667),.DATA(g11548));
  MSFF DFF_1011(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1668),.DATA(g1667));
  MSFF DFF_1012(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1669),.DATA(g11549));
  MSFF DFF_1013(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1670),.DATA(g1669));
  MSFF DFF_1014(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1671),.DATA(g13439));
  MSFF DFF_1015(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1672),.DATA(g1671));
  MSFF DFF_1016(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1680),.DATA(g19036));
  MSFF DFF_1017(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1686),.DATA(g29428));
  MSFF DFF_1018(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1689),.DATA(g29429));
  MSFF DFF_1019(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1678),.DATA(g29430));
  MSFF DFF_1020(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1677),.DATA(g29431));
  MSFF DFF_1021(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1676),.DATA(g29432));
  MSFF DFF_1022(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1675),.DATA(g29433));
  MSFF DFF_1023(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1685),.DATA(g19040));
  MSFF DFF_1024(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1684),.DATA(g19039));
  MSFF DFF_1025(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1683),.DATA(g19038));
  MSFF DFF_1026(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1682),.DATA(g19037));
  MSFF DFF_1027(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1681),.DATA(g25152));
  MSFF DFF_1028(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1679),.DATA(g27220));
  MSFF DFF_1029(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1723),.DATA(g11551));
  MSFF DFF_1030(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1730),.DATA(g1723));
  MSFF DFF_1031(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1731),.DATA(g11552));
  MSFF DFF_1032(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1732),.DATA(g1731));
  MSFF DFF_1033(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1733),.DATA(g11553));
  MSFF DFF_1034(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1734),.DATA(g1733));
  MSFF DFF_1035(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1738),.DATA(g11554));
  MSFF DFF_1036(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1745),.DATA(g1738));
  MSFF DFF_1037(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1746),.DATA(g11555));
  MSFF DFF_1038(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1747),.DATA(g1746));
  MSFF DFF_1039(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1748),.DATA(g11556));
  MSFF DFF_1040(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1749),.DATA(g1748));
  MSFF DFF_1041(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1753),.DATA(g11557));
  MSFF DFF_1042(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1760),.DATA(g1753));
  MSFF DFF_1043(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1761),.DATA(g11558));
  MSFF DFF_1044(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1762),.DATA(g1761));
  MSFF DFF_1045(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1763),.DATA(g11559));
  MSFF DFF_1046(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1764),.DATA(g1763));
  MSFF DFF_1047(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1768),.DATA(g11560));
  MSFF DFF_1048(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1775),.DATA(g1768));
  MSFF DFF_1049(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1776),.DATA(g11561));
  MSFF DFF_1050(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1777),.DATA(g1776));
  MSFF DFF_1051(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1778),.DATA(g11562));
  MSFF DFF_1052(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1705),.DATA(g1778));
  MSFF DFF_1053(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1706),.DATA(g13440));
  MSFF DFF_1054(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1712),.DATA(g1706));
  MSFF DFF_1055(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1718),.DATA(g1712));
  MSFF DFF_1056(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1925),.DATA(g13451));
  MSFF DFF_1057(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1931),.DATA(g1925));
  MSFF DFF_1058(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1930),.DATA(g1931));
  MSFF DFF_1059(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1934),.DATA(g23236));
  MSFF DFF_1060(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1937),.DATA(g20564));
  MSFF DFF_1061(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1890),.DATA(g20565));
  MSFF DFF_1062(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1893),.DATA(g16471));
  MSFF DFF_1063(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1903),.DATA(g1893));
  MSFF DFF_1064(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1904),.DATA(g1903));
  MSFF DFF_1065(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1944),.DATA(g11566));
  MSFF DFF_1066(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1949),.DATA(g1944));
  MSFF DFF_1067(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1950),.DATA(g11569));
  MSFF DFF_1068(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1951),.DATA(g1950));
  MSFF DFF_1069(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1952),.DATA(g11570));
  MSFF DFF_1070(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1953),.DATA(g1952));
  MSFF DFF_1071(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1954),.DATA(g11571));
  MSFF DFF_1072(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1945),.DATA(g1954));
  MSFF DFF_1073(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1946),.DATA(g11567));
  MSFF DFF_1074(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1947),.DATA(g1946));
  MSFF DFF_1075(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1948),.DATA(g11568));
  MSFF DFF_1076(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1870),.DATA(g1948));
  MSFF DFF_1077(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1855),.DATA(g13441));
  MSFF DFF_1078(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1862),.DATA(g1855));
  MSFF DFF_1079(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1866),.DATA(g1862));
  MSFF DFF_1080(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1867),.DATA(g24374));
  MSFF DFF_1081(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1868),.DATA(g24375));
  MSFF DFF_1082(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1869),.DATA(g24376));
  MSFF DFF_1083(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1836),.DATA(g25161));
  MSFF DFF_1084(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1839),.DATA(g25153));
  MSFF DFF_1085(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1842),.DATA(g25154));
  MSFF DFF_1086(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1858),.DATA(g25158));
  MSFF DFF_1087(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1859),.DATA(g25159));
  MSFF DFF_1088(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1860),.DATA(g25160));
  MSFF DFF_1089(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1861),.DATA(g24371));
  MSFF DFF_1090(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1865),.DATA(g24372));
  MSFF DFF_1091(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1845),.DATA(g24373));
  MSFF DFF_1092(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1846),.DATA(g25155));
  MSFF DFF_1093(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1849),.DATA(g25156));
  MSFF DFF_1094(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1852),.DATA(g25157));
  MSFF DFF_1095(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1908),.DATA(g16472));
  MSFF DFF_1096(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1915),.DATA(g1908));
  MSFF DFF_1097(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1922),.DATA(g1915));
  MSFF DFF_1098(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1923),.DATA(g19045));
  MSFF DFF_1099(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1924),.DATA(g1923));
  MSFF DFF_1100(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1928),.DATA(g29445));
  MSFF DFF_1101(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1929),.DATA(g19046));
  MSFF DFF_1102(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1880),.DATA(g1929));
  MSFF DFF_1103(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1938),.DATA(g19047));
  MSFF DFF_1104(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1939),.DATA(g1938));
  MSFF DFF_1105(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1956),.DATA(g28271));
  MSFF DFF_1106(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1957),.DATA(g28272));
  MSFF DFF_1107(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1955),.DATA(g28273));
  MSFF DFF_1108(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1959),.DATA(g28274));
  MSFF DFF_1109(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1960),.DATA(g28275));
  MSFF DFF_1110(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1958),.DATA(g28276));
  MSFF DFF_1111(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1962),.DATA(g28277));
  MSFF DFF_1112(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1963),.DATA(g28278));
  MSFF DFF_1113(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1961),.DATA(g28279));
  MSFF DFF_1114(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1965),.DATA(g28280));
  MSFF DFF_1115(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1966),.DATA(g28281));
  MSFF DFF_1116(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1964),.DATA(g28282));
  MSFF DFF_1117(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1967),.DATA(g26003));
  MSFF DFF_1118(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1970),.DATA(g26004));
  MSFF DFF_1119(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1973),.DATA(g26005));
  MSFF DFF_1120(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1976),.DATA(g26006));
  MSFF DFF_1121(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1979),.DATA(g26007));
  MSFF DFF_1122(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1982),.DATA(g26008));
  MSFF DFF_1123(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1994),.DATA(g29151));
  MSFF DFF_1124(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1997),.DATA(g29152));
  MSFF DFF_1125(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2000),.DATA(g29153));
  MSFF DFF_1126(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1985),.DATA(g29148));
  MSFF DFF_1127(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1988),.DATA(g29149));
  MSFF DFF_1128(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1991),.DATA(g29150));
  MSFF DFF_1129(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1871),.DATA(g27224));
  MSFF DFF_1130(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1874),.DATA(g27225));
  MSFF DFF_1131(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1877),.DATA(g27226));
  MSFF DFF_1132(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1886),.DATA(g8302));
  MSFF DFF_1133(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1887),.DATA(g24377));
  MSFF DFF_1134(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1888),.DATA(g19041));
  MSFF DFF_1135(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1889),.DATA(g19042));
  MSFF DFF_1136(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1894),.DATA(g19043));
  MSFF DFF_1137(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1895),.DATA(g19044));
  MSFF DFF_1138(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1896),.DATA(g29444));
  MSFF DFF_1139(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1897),.DATA(g29443));
  MSFF DFF_1140(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1898),.DATA(g29442));
  MSFF DFF_1141(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1899),.DATA(g29441));
  MSFF DFF_1142(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1900),.DATA(g29440));
  MSFF DFF_1143(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1905),.DATA(g1900));
  MSFF DFF_1144(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1909),.DATA(g13442));
  MSFF DFF_1145(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1910),.DATA(g13443));
  MSFF DFF_1146(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1911),.DATA(g13444));
  MSFF DFF_1147(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1912),.DATA(g13445));
  MSFF DFF_1148(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1913),.DATA(g13446));
  MSFF DFF_1149(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1914),.DATA(g13447));
  MSFF DFF_1150(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1916),.DATA(g13448));
  MSFF DFF_1151(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1917),.DATA(g13449));
  MSFF DFF_1152(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1918),.DATA(g26002));
  MSFF DFF_1153(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1921),.DATA(g13450));
  MSFF DFF_1154(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2003),.DATA(g13452));
  MSFF DFF_1155(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2006),.DATA(g2003));
  MSFF DFF_1156(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2009),.DATA(g2006));
  MSFF DFF_1157(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2010),.DATA(g20566));
  MSFF DFF_1158(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2039),.DATA(g21945));
  MSFF DFF_1159(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2020),.DATA(g23237));
  MSFF DFF_1160(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2013),.DATA(g24378));
  MSFF DFF_1161(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2033),.DATA(g25162));
  MSFF DFF_1162(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2026),.DATA(g26009));
  MSFF DFF_1163(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2040),.DATA(g26725));
  MSFF DFF_1164(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2052),.DATA(g27227));
  MSFF DFF_1165(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2046),.DATA(g27706));
  MSFF DFF_1166(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2059),.DATA(g28283));
  MSFF DFF_1167(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2066),.DATA(g28687));
  MSFF DFF_1168(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2072),.DATA(g29154));
  MSFF DFF_1169(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2079),.DATA(g23238));
  MSFF DFF_1170(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2080),.DATA(g23239));
  MSFF DFF_1171(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2078),.DATA(g23240));
  MSFF DFF_1172(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2082),.DATA(g23241));
  MSFF DFF_1173(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2083),.DATA(g23242));
  MSFF DFF_1174(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2081),.DATA(g23243));
  MSFF DFF_1175(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2085),.DATA(g23244));
  MSFF DFF_1176(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2086),.DATA(g23245));
  MSFF DFF_1177(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2084),.DATA(g23246));
  MSFF DFF_1178(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2088),.DATA(g23247));
  MSFF DFF_1179(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2089),.DATA(g23248));
  MSFF DFF_1180(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2087),.DATA(g23249));
  MSFF DFF_1181(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2091),.DATA(g23250));
  MSFF DFF_1182(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2092),.DATA(g23251));
  MSFF DFF_1183(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2090),.DATA(g23252));
  MSFF DFF_1184(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2094),.DATA(g23253));
  MSFF DFF_1185(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2095),.DATA(g23254));
  MSFF DFF_1186(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2093),.DATA(g23255));
  MSFF DFF_1187(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2097),.DATA(g23256));
  MSFF DFF_1188(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2098),.DATA(g23257));
  MSFF DFF_1189(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2096),.DATA(g23258));
  MSFF DFF_1190(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2100),.DATA(g23259));
  MSFF DFF_1191(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2101),.DATA(g23260));
  MSFF DFF_1192(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2099),.DATA(g23261));
  MSFF DFF_1193(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2103),.DATA(g23262));
  MSFF DFF_1194(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2104),.DATA(g23263));
  MSFF DFF_1195(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2102),.DATA(g23264));
  MSFF DFF_1196(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2106),.DATA(g23265));
  MSFF DFF_1197(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2107),.DATA(g23266));
  MSFF DFF_1198(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2105),.DATA(g23267));
  MSFF DFF_1199(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2109),.DATA(g23268));
  MSFF DFF_1200(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2110),.DATA(g23269));
  MSFF DFF_1201(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2108),.DATA(g23270));
  MSFF DFF_1202(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2112),.DATA(g23271));
  MSFF DFF_1203(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2113),.DATA(g23272));
  MSFF DFF_1204(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2111),.DATA(g23273));
  MSFF DFF_1205(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2115),.DATA(g26726));
  MSFF DFF_1206(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2116),.DATA(g26727));
  MSFF DFF_1207(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2114),.DATA(g26728));
  MSFF DFF_1208(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2118),.DATA(g24379));
  MSFF DFF_1209(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2119),.DATA(g24380));
  MSFF DFF_1210(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2117),.DATA(g24381));
  MSFF DFF_1211(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2214),.DATA(g13453));
  MSFF DFF_1212(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2211),.DATA(g2214));
  MSFF DFF_1213(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2241),.DATA(g2211));
  MSFF DFF_1214(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2206),.DATA(g24382));
  MSFF DFF_1215(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2207),.DATA(g24383));
  MSFF DFF_1216(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2205),.DATA(g24384));
  MSFF DFF_1217(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2209),.DATA(g24385));
  MSFF DFF_1218(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2210),.DATA(g24386));
  MSFF DFF_1219(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2208),.DATA(g24387));
  MSFF DFF_1220(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2218),.DATA(g24388));
  MSFF DFF_1221(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2219),.DATA(g24389));
  MSFF DFF_1222(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2217),.DATA(g24390));
  MSFF DFF_1223(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2221),.DATA(g24391));
  MSFF DFF_1224(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2222),.DATA(g24392));
  MSFF DFF_1225(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2220),.DATA(g24393));
  MSFF DFF_1226(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2224),.DATA(g24394));
  MSFF DFF_1227(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2225),.DATA(g24395));
  MSFF DFF_1228(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2223),.DATA(g24396));
  MSFF DFF_1229(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2227),.DATA(g24397));
  MSFF DFF_1230(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2228),.DATA(g24398));
  MSFF DFF_1231(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2226),.DATA(g24399));
  MSFF DFF_1232(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2230),.DATA(g24400));
  MSFF DFF_1233(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2231),.DATA(g24401));
  MSFF DFF_1234(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2229),.DATA(g24402));
  MSFF DFF_1235(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2233),.DATA(g24403));
  MSFF DFF_1236(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2234),.DATA(g24404));
  MSFF DFF_1237(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2232),.DATA(g24405));
  MSFF DFF_1238(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2236),.DATA(g24406));
  MSFF DFF_1239(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2237),.DATA(g24407));
  MSFF DFF_1240(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2235),.DATA(g24408));
  MSFF DFF_1241(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2239),.DATA(g24409));
  MSFF DFF_1242(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2240),.DATA(g24410));
  MSFF DFF_1243(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2238),.DATA(g24411));
  MSFF DFF_1244(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2245),.DATA(g26730));
  MSFF DFF_1245(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2246),.DATA(g26731));
  MSFF DFF_1246(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2244),.DATA(g26732));
  MSFF DFF_1247(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2248),.DATA(g26733));
  MSFF DFF_1248(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2249),.DATA(g26734));
  MSFF DFF_1249(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2247),.DATA(g26735));
  MSFF DFF_1250(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2251),.DATA(g26736));
  MSFF DFF_1251(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2252),.DATA(g26737));
  MSFF DFF_1252(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2250),.DATA(g26738));
  MSFF DFF_1253(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2254),.DATA(g26739));
  MSFF DFF_1254(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2255),.DATA(g26740));
  MSFF DFF_1255(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2253),.DATA(g26741));
  MSFF DFF_1256(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2261),.DATA(g30551));
  MSFF DFF_1257(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2264),.DATA(g30552));
  MSFF DFF_1258(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2267),.DATA(g30553));
  MSFF DFF_1259(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2306),.DATA(g30896));
  MSFF DFF_1260(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2309),.DATA(g30897));
  MSFF DFF_1261(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2312),.DATA(g30898));
  MSFF DFF_1262(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2270),.DATA(g30890));
  MSFF DFF_1263(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2273),.DATA(g30891));
  MSFF DFF_1264(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2276),.DATA(g30892));
  MSFF DFF_1265(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2315),.DATA(g30899));
  MSFF DFF_1266(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2318),.DATA(g30900));
  MSFF DFF_1267(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2321),.DATA(g30901));
  MSFF DFF_1268(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2279),.DATA(g30554));
  MSFF DFF_1269(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2282),.DATA(g30555));
  MSFF DFF_1270(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2285),.DATA(g30556));
  MSFF DFF_1271(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2324),.DATA(g30560));
  MSFF DFF_1272(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2327),.DATA(g30561));
  MSFF DFF_1273(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2330),.DATA(g30562));
  MSFF DFF_1274(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2288),.DATA(g30557));
  MSFF DFF_1275(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2291),.DATA(g30558));
  MSFF DFF_1276(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2294),.DATA(g30559));
  MSFF DFF_1277(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2333),.DATA(g30563));
  MSFF DFF_1278(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2336),.DATA(g30564));
  MSFF DFF_1279(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2339),.DATA(g30565));
  MSFF DFF_1280(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2297),.DATA(g30893));
  MSFF DFF_1281(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2300),.DATA(g30894));
  MSFF DFF_1282(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2303),.DATA(g30895));
  MSFF DFF_1283(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2342),.DATA(g30902));
  MSFF DFF_1284(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2345),.DATA(g30903));
  MSFF DFF_1285(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2348),.DATA(g30904));
  MSFF DFF_1286(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2160),.DATA(g26010));
  MSFF DFF_1287(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2156),.DATA(g26729));
  MSFF DFF_1288(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2151),.DATA(g27228));
  MSFF DFF_1289(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2147),.DATA(g27707));
  MSFF DFF_1290(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2142),.DATA(g28284));
  MSFF DFF_1291(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2138),.DATA(g28688));
  MSFF DFF_1292(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2133),.DATA(g29155));
  MSFF DFF_1293(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2129),.DATA(g29446));
  MSFF DFF_1294(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2124),.DATA(g29648));
  MSFF DFF_1295(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2120),.DATA(g29806));
  MSFF DFF_1296(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2256),.DATA(g20567));
  MSFF DFF_1297(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2258),.DATA(g2256));
  MSFF DFF_1298(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2257),.DATA(g2258));
  MSFF DFF_1299(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2351),.DATA(g13454));
  MSFF DFF_1300(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2480),.DATA(g2351));
  MSFF DFF_1301(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2476),.DATA(g2480));
  MSFF DFF_1302(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2384),.DATA(g11577));
  MSFF DFF_1303(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2429),.DATA(g28285));
  MSFF DFF_1304(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2418),.DATA(g28286));
  MSFF DFF_1305(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2421),.DATA(g28287));
  MSFF DFF_1306(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2444),.DATA(g28288));
  MSFF DFF_1307(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2433),.DATA(g28289));
  MSFF DFF_1308(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2436),.DATA(g28290));
  MSFF DFF_1309(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2459),.DATA(g28291));
  MSFF DFF_1310(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2448),.DATA(g28292));
  MSFF DFF_1311(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2451),.DATA(g28293));
  MSFF DFF_1312(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2473),.DATA(g28294));
  MSFF DFF_1313(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2463),.DATA(g28295));
  MSFF DFF_1314(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2466),.DATA(g28296));
  MSFF DFF_1315(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2483),.DATA(g29447));
  MSFF DFF_1316(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2486),.DATA(g29448));
  MSFF DFF_1317(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2489),.DATA(g29449));
  MSFF DFF_1318(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2492),.DATA(g29652));
  MSFF DFF_1319(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2495),.DATA(g29653));
  MSFF DFF_1320(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2498),.DATA(g29654));
  MSFF DFF_1321(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2502),.DATA(g29450));
  MSFF DFF_1322(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2503),.DATA(g29451));
  MSFF DFF_1323(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2501),.DATA(g29452));
  MSFF DFF_1324(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2504),.DATA(g27708));
  MSFF DFF_1325(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2507),.DATA(g27709));
  MSFF DFF_1326(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2510),.DATA(g27710));
  MSFF DFF_1327(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2513),.DATA(g27711));
  MSFF DFF_1328(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2516),.DATA(g27712));
  MSFF DFF_1329(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2519),.DATA(g27713));
  MSFF DFF_1330(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2523),.DATA(g28689));
  MSFF DFF_1331(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2524),.DATA(g28690));
  MSFF DFF_1332(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2522),.DATA(g28691));
  MSFF DFF_1333(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2387),.DATA(g29807));
  MSFF DFF_1334(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2388),.DATA(g29808));
  MSFF DFF_1335(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2389),.DATA(g29809));
  MSFF DFF_1336(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2390),.DATA(g30905));
  MSFF DFF_1337(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2391),.DATA(g30906));
  MSFF DFF_1338(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2392),.DATA(g30907));
  MSFF DFF_1339(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2393),.DATA(g30719));
  MSFF DFF_1340(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2394),.DATA(g30720));
  MSFF DFF_1341(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2395),.DATA(g30721));
  MSFF DFF_1342(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2397),.DATA(g29649));
  MSFF DFF_1343(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2398),.DATA(g29650));
  MSFF DFF_1344(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2396),.DATA(g29651));
  MSFF DFF_1345(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2478),.DATA(g27230));
  MSFF DFF_1346(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2479),.DATA(g27231));
  MSFF DFF_1347(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2477),.DATA(g27232));
  MSFF DFF_1348(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2525),.DATA(g11590));
  MSFF DFF_1349(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2526),.DATA(g2525));
  MSFF DFF_1350(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2527),.DATA(g11591));
  MSFF DFF_1351(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2528),.DATA(g2527));
  MSFF DFF_1352(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2529),.DATA(g11592));
  MSFF DFF_1353(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2354),.DATA(g2529));
  MSFF DFF_1354(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2355),.DATA(g11572));
  MSFF DFF_1355(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2356),.DATA(g2355));
  MSFF DFF_1356(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2357),.DATA(g11573));
  MSFF DFF_1357(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2358),.DATA(g2357));
  MSFF DFF_1358(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2359),.DATA(g11574));
  MSFF DFF_1359(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2360),.DATA(g2359));
  MSFF DFF_1360(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2361),.DATA(g11575));
  MSFF DFF_1361(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2362),.DATA(g2361));
  MSFF DFF_1362(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2363),.DATA(g11576));
  MSFF DFF_1363(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2364),.DATA(g2363));
  MSFF DFF_1364(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2365),.DATA(g13455));
  MSFF DFF_1365(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2366),.DATA(g2365));
  MSFF DFF_1366(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2374),.DATA(g19048));
  MSFF DFF_1367(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2380),.DATA(g30314));
  MSFF DFF_1368(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2383),.DATA(g30315));
  MSFF DFF_1369(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2372),.DATA(g30316));
  MSFF DFF_1370(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2371),.DATA(g30317));
  MSFF DFF_1371(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2370),.DATA(g30318));
  MSFF DFF_1372(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2369),.DATA(g30319));
  MSFF DFF_1373(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2379),.DATA(g19052));
  MSFF DFF_1374(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2378),.DATA(g19051));
  MSFF DFF_1375(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2377),.DATA(g19050));
  MSFF DFF_1376(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2376),.DATA(g19049));
  MSFF DFF_1377(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2375),.DATA(g25163));
  MSFF DFF_1378(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2373),.DATA(g27229));
  MSFF DFF_1379(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2417),.DATA(g11578));
  MSFF DFF_1380(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2424),.DATA(g2417));
  MSFF DFF_1381(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2425),.DATA(g11579));
  MSFF DFF_1382(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2426),.DATA(g2425));
  MSFF DFF_1383(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2427),.DATA(g11580));
  MSFF DFF_1384(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2428),.DATA(g2427));
  MSFF DFF_1385(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2432),.DATA(g11581));
  MSFF DFF_1386(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2439),.DATA(g2432));
  MSFF DFF_1387(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2440),.DATA(g11582));
  MSFF DFF_1388(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2441),.DATA(g2440));
  MSFF DFF_1389(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2442),.DATA(g11583));
  MSFF DFF_1390(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2443),.DATA(g2442));
  MSFF DFF_1391(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2447),.DATA(g11584));
  MSFF DFF_1392(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2454),.DATA(g2447));
  MSFF DFF_1393(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2455),.DATA(g11585));
  MSFF DFF_1394(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2456),.DATA(g2455));
  MSFF DFF_1395(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2457),.DATA(g11586));
  MSFF DFF_1396(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2458),.DATA(g2457));
  MSFF DFF_1397(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2462),.DATA(g11587));
  MSFF DFF_1398(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2469),.DATA(g2462));
  MSFF DFF_1399(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2470),.DATA(g11588));
  MSFF DFF_1400(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2471),.DATA(g2470));
  MSFF DFF_1401(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2472),.DATA(g11589));
  MSFF DFF_1402(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2399),.DATA(g2472));
  MSFF DFF_1403(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2400),.DATA(g13456));
  MSFF DFF_1404(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2406),.DATA(g2400));
  MSFF DFF_1405(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2412),.DATA(g2406));
  MSFF DFF_1406(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2619),.DATA(g13467));
  MSFF DFF_1407(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2625),.DATA(g2619));
  MSFF DFF_1408(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2624),.DATA(g2625));
  MSFF DFF_1409(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2628),.DATA(g23274));
  MSFF DFF_1410(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2631),.DATA(g20568));
  MSFF DFF_1411(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2584),.DATA(g20569));
  MSFF DFF_1412(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2587),.DATA(g16473));
  MSFF DFF_1413(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2597),.DATA(g2587));
  MSFF DFF_1414(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2598),.DATA(g2597));
  MSFF DFF_1415(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2638),.DATA(g11593));
  MSFF DFF_1416(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2643),.DATA(g2638));
  MSFF DFF_1417(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2644),.DATA(g11596));
  MSFF DFF_1418(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2645),.DATA(g2644));
  MSFF DFF_1419(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2646),.DATA(g11597));
  MSFF DFF_1420(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2647),.DATA(g2646));
  MSFF DFF_1421(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2648),.DATA(g11598));
  MSFF DFF_1422(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2639),.DATA(g2648));
  MSFF DFF_1423(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2640),.DATA(g11594));
  MSFF DFF_1424(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2641),.DATA(g2640));
  MSFF DFF_1425(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2642),.DATA(g11595));
  MSFF DFF_1426(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2564),.DATA(g2642));
  MSFF DFF_1427(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2549),.DATA(g13457));
  MSFF DFF_1428(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2556),.DATA(g2549));
  MSFF DFF_1429(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2560),.DATA(g2556));
  MSFF DFF_1430(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2561),.DATA(g24415));
  MSFF DFF_1431(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2562),.DATA(g24416));
  MSFF DFF_1432(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2563),.DATA(g24417));
  MSFF DFF_1433(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2530),.DATA(g25172));
  MSFF DFF_1434(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2533),.DATA(g25164));
  MSFF DFF_1435(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2536),.DATA(g25165));
  MSFF DFF_1436(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2552),.DATA(g25169));
  MSFF DFF_1437(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2553),.DATA(g25170));
  MSFF DFF_1438(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2554),.DATA(g25171));
  MSFF DFF_1439(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2555),.DATA(g24412));
  MSFF DFF_1440(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2559),.DATA(g24413));
  MSFF DFF_1441(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2539),.DATA(g24414));
  MSFF DFF_1442(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2540),.DATA(g25166));
  MSFF DFF_1443(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2543),.DATA(g25167));
  MSFF DFF_1444(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2546),.DATA(g25168));
  MSFF DFF_1445(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2602),.DATA(g16474));
  MSFF DFF_1446(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2609),.DATA(g2602));
  MSFF DFF_1447(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2616),.DATA(g2609));
  MSFF DFF_1448(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2617),.DATA(g19057));
  MSFF DFF_1449(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2618),.DATA(g2617));
  MSFF DFF_1450(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2622),.DATA(g30325));
  MSFF DFF_1451(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2623),.DATA(g19058));
  MSFF DFF_1452(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2574),.DATA(g2623));
  MSFF DFF_1453(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2632),.DATA(g19059));
  MSFF DFF_1454(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2633),.DATA(g2632));
  MSFF DFF_1455(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2650),.DATA(g28297));
  MSFF DFF_1456(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2651),.DATA(g28298));
  MSFF DFF_1457(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2649),.DATA(g28299));
  MSFF DFF_1458(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2653),.DATA(g28300));
  MSFF DFF_1459(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2654),.DATA(g28301));
  MSFF DFF_1460(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2652),.DATA(g28302));
  MSFF DFF_1461(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2656),.DATA(g28303));
  MSFF DFF_1462(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2657),.DATA(g28304));
  MSFF DFF_1463(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2655),.DATA(g28305));
  MSFF DFF_1464(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2659),.DATA(g28306));
  MSFF DFF_1465(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2660),.DATA(g28307));
  MSFF DFF_1466(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2658),.DATA(g28308));
  MSFF DFF_1467(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2661),.DATA(g26012));
  MSFF DFF_1468(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2664),.DATA(g26013));
  MSFF DFF_1469(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2667),.DATA(g26014));
  MSFF DFF_1470(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2670),.DATA(g26015));
  MSFF DFF_1471(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2673),.DATA(g26016));
  MSFF DFF_1472(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2676),.DATA(g26017));
  MSFF DFF_1473(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2688),.DATA(g29159));
  MSFF DFF_1474(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2691),.DATA(g29160));
  MSFF DFF_1475(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2694),.DATA(g29161));
  MSFF DFF_1476(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2679),.DATA(g29156));
  MSFF DFF_1477(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2682),.DATA(g29157));
  MSFF DFF_1478(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2685),.DATA(g29158));
  MSFF DFF_1479(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2565),.DATA(g27233));
  MSFF DFF_1480(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2568),.DATA(g27234));
  MSFF DFF_1481(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2571),.DATA(g27235));
  MSFF DFF_1482(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2580),.DATA(g8311));
  MSFF DFF_1483(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2581),.DATA(g24418));
  MSFF DFF_1484(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2582),.DATA(g19053));
  MSFF DFF_1485(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2583),.DATA(g19054));
  MSFF DFF_1486(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2588),.DATA(g19055));
  MSFF DFF_1487(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2589),.DATA(g19056));
  MSFF DFF_1488(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2590),.DATA(g30324));
  MSFF DFF_1489(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2591),.DATA(g30323));
  MSFF DFF_1490(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2592),.DATA(g30322));
  MSFF DFF_1491(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2593),.DATA(g30321));
  MSFF DFF_1492(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2594),.DATA(g30320));
  MSFF DFF_1493(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2599),.DATA(g2594));
  MSFF DFF_1494(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2603),.DATA(g13458));
  MSFF DFF_1495(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2604),.DATA(g13459));
  MSFF DFF_1496(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2605),.DATA(g13460));
  MSFF DFF_1497(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2606),.DATA(g13461));
  MSFF DFF_1498(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2607),.DATA(g13462));
  MSFF DFF_1499(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2608),.DATA(g13463));
  MSFF DFF_1500(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2610),.DATA(g13464));
  MSFF DFF_1501(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2611),.DATA(g13465));
  MSFF DFF_1502(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2612),.DATA(g26011));
  MSFF DFF_1503(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2615),.DATA(g13466));
  MSFF DFF_1504(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2697),.DATA(g13468));
  MSFF DFF_1505(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2700),.DATA(g2697));
  MSFF DFF_1506(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2703),.DATA(g2700));
  MSFF DFF_1507(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2704),.DATA(g20570));
  MSFF DFF_1508(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2733),.DATA(g21946));
  MSFF DFF_1509(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2714),.DATA(g23275));
  MSFF DFF_1510(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2707),.DATA(g24419));
  MSFF DFF_1511(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2727),.DATA(g25173));
  MSFF DFF_1512(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2720),.DATA(g26018));
  MSFF DFF_1513(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2734),.DATA(g26742));
  MSFF DFF_1514(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2746),.DATA(g27236));
  MSFF DFF_1515(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2740),.DATA(g27714));
  MSFF DFF_1516(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2753),.DATA(g28309));
  MSFF DFF_1517(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2760),.DATA(g28692));
  MSFF DFF_1518(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2766),.DATA(g29162));
  MSFF DFF_1519(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2773),.DATA(g23276));
  MSFF DFF_1520(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2774),.DATA(g23277));
  MSFF DFF_1521(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2772),.DATA(g23278));
  MSFF DFF_1522(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2776),.DATA(g23279));
  MSFF DFF_1523(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2777),.DATA(g23280));
  MSFF DFF_1524(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2775),.DATA(g23281));
  MSFF DFF_1525(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2779),.DATA(g23282));
  MSFF DFF_1526(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2780),.DATA(g23283));
  MSFF DFF_1527(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2778),.DATA(g23284));
  MSFF DFF_1528(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2782),.DATA(g23285));
  MSFF DFF_1529(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2783),.DATA(g23286));
  MSFF DFF_1530(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2781),.DATA(g23287));
  MSFF DFF_1531(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2785),.DATA(g23288));
  MSFF DFF_1532(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2786),.DATA(g23289));
  MSFF DFF_1533(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2784),.DATA(g23290));
  MSFF DFF_1534(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2788),.DATA(g23291));
  MSFF DFF_1535(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2789),.DATA(g23292));
  MSFF DFF_1536(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2787),.DATA(g23293));
  MSFF DFF_1537(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2791),.DATA(g23294));
  MSFF DFF_1538(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2792),.DATA(g23295));
  MSFF DFF_1539(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2790),.DATA(g23296));
  MSFF DFF_1540(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2794),.DATA(g23297));
  MSFF DFF_1541(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2795),.DATA(g23298));
  MSFF DFF_1542(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2793),.DATA(g23299));
  MSFF DFF_1543(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2797),.DATA(g23300));
  MSFF DFF_1544(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2798),.DATA(g23301));
  MSFF DFF_1545(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2796),.DATA(g23302));
  MSFF DFF_1546(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2800),.DATA(g23303));
  MSFF DFF_1547(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2801),.DATA(g23304));
  MSFF DFF_1548(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2799),.DATA(g23305));
  MSFF DFF_1549(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2803),.DATA(g23306));
  MSFF DFF_1550(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2804),.DATA(g23307));
  MSFF DFF_1551(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2802),.DATA(g23308));
  MSFF DFF_1552(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2806),.DATA(g23309));
  MSFF DFF_1553(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2807),.DATA(g23310));
  MSFF DFF_1554(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2805),.DATA(g23311));
  MSFF DFF_1555(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2809),.DATA(g26743));
  MSFF DFF_1556(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2810),.DATA(g26744));
  MSFF DFF_1557(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2808),.DATA(g26745));
  MSFF DFF_1558(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2812),.DATA(g24420));
  MSFF DFF_1559(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2813),.DATA(g24421));
  MSFF DFF_1560(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2811),.DATA(g24422));
  MSFF DFF_1561(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3054),.DATA(g23317));
  MSFF DFF_1562(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3079),.DATA(g23318));
  MSFF DFF_1563(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3080),.DATA(g21965));
  MSFF DFF_1564(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3043),.DATA(g29453));
  MSFF DFF_1565(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3044),.DATA(g29454));
  MSFF DFF_1566(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3045),.DATA(g29455));
  MSFF DFF_1567(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3046),.DATA(g29456));
  MSFF DFF_1568(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3047),.DATA(g29457));
  MSFF DFF_1569(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3048),.DATA(g29458));
  MSFF DFF_1570(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3049),.DATA(g29459));
  MSFF DFF_1571(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3050),.DATA(g29460));
  MSFF DFF_1572(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3051),.DATA(g29655));
  MSFF DFF_1573(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3052),.DATA(g29972));
  MSFF DFF_1574(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3053),.DATA(g29973));
  MSFF DFF_1575(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3055),.DATA(g29974));
  MSFF DFF_1576(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3056),.DATA(g29975));
  MSFF DFF_1577(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3057),.DATA(g29976));
  MSFF DFF_1578(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3058),.DATA(g29977));
  MSFF DFF_1579(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3059),.DATA(g29978));
  MSFF DFF_1580(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3060),.DATA(g29979));
  MSFF DFF_1581(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3061),.DATA(g30119));
  MSFF DFF_1582(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3062),.DATA(g30908));
  MSFF DFF_1583(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3063),.DATA(g30909));
  MSFF DFF_1584(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3064),.DATA(g30910));
  MSFF DFF_1585(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3065),.DATA(g30911));
  MSFF DFF_1586(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3066),.DATA(g30912));
  MSFF DFF_1587(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3067),.DATA(g30913));
  MSFF DFF_1588(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3068),.DATA(g30914));
  MSFF DFF_1589(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3069),.DATA(g30915));
  MSFF DFF_1590(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3070),.DATA(g30940));
  MSFF DFF_1591(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3071),.DATA(g30980));
  MSFF DFF_1592(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3072),.DATA(g30981));
  MSFF DFF_1593(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3073),.DATA(g30982));
  MSFF DFF_1594(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3074),.DATA(g30983));
  MSFF DFF_1595(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3075),.DATA(g30984));
  MSFF DFF_1596(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3076),.DATA(g30985));
  MSFF DFF_1597(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3077),.DATA(g30986));
  MSFF DFF_1598(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3078),.DATA(g30987));
  MSFF DFF_1599(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2997),.DATA(g30989));
  MSFF DFF_1600(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2993),.DATA(g26748));
  MSFF DFF_1601(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2998),.DATA(g27238));
  MSFF DFF_1602(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3006),.DATA(g25177));
  MSFF DFF_1603(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3002),.DATA(g26021));
  MSFF DFF_1604(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3013),.DATA(g26750));
  MSFF DFF_1605(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3010),.DATA(g27239));
  MSFF DFF_1606(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3024),.DATA(g27716));
  MSFF DFF_1607(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3018),.DATA(g24425));
  MSFF DFF_1608(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3028),.DATA(g25176));
  MSFF DFF_1609(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3036),.DATA(g26022));
  MSFF DFF_1610(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3032),.DATA(g26749));
  MSFF DFF_1611(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3040),.DATA(g16497));
  MSFF DFF_1612(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2986),.DATA(g3040));
  MSFF DFF_1613(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2987),.DATA(g16495));
  MSFF DFF_1614(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g48),.DATA(g20595));
  MSFF DFF_1615(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g45),.DATA(g20596));
  MSFF DFF_1616(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g42),.DATA(g20597));
  MSFF DFF_1617(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g39),.DATA(g20598));
  MSFF DFF_1618(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g27),.DATA(g20599));
  MSFF DFF_1619(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g30),.DATA(g20600));
  MSFF DFF_1620(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g33),.DATA(g20601));
  MSFF DFF_1621(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g36),.DATA(g20602));
  MSFF DFF_1622(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g3083),.DATA(g20603));
  MSFF DFF_1623(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g26),.DATA(g20604));
  MSFF DFF_1624(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2992),.DATA(g21966));
  MSFF DFF_1625(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g23),.DATA(g20605));
  MSFF DFF_1626(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g20),.DATA(g20606));
  MSFF DFF_1627(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g17),.DATA(g20607));
  MSFF DFF_1628(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g11),.DATA(g20608));
  MSFF DFF_1629(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g14),.DATA(g20589));
  MSFF DFF_1630(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g5),.DATA(g20590));
  MSFF DFF_1631(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g8),.DATA(g20591));
  MSFF DFF_1632(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2),.DATA(g20592));
  MSFF DFF_1633(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2990),.DATA(g20593));
  MSFF DFF_1634(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g2991),.DATA(g21964));
  MSFF DFF_1635(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1),.DATA(g20594));
//
  NOT NOT1_0(.VSS(VSS),.VDD(VDD),.Y(I13089),.A(g563));
  NOT NOT1_1(.VSS(VSS),.VDD(VDD),.Y(g562),.A(I13089));
  NOT NOT1_2(.VSS(VSS),.VDD(VDD),.Y(I13092),.A(g1249));
  NOT NOT1_3(.VSS(VSS),.VDD(VDD),.Y(g1248),.A(I13092));
  NOT NOT1_4(.VSS(VSS),.VDD(VDD),.Y(I13095),.A(g1943));
  NOT NOT1_5(.VSS(VSS),.VDD(VDD),.Y(g1942),.A(I13095));
  NOT NOT1_6(.VSS(VSS),.VDD(VDD),.Y(I13098),.A(g2637));
  NOT NOT1_7(.VSS(VSS),.VDD(VDD),.Y(g2636),.A(I13098));
  NOT NOT1_8(.VSS(VSS),.VDD(VDD),.Y(I13101),.A(g1));
  NOT NOT1_9(.VSS(VSS),.VDD(VDD),.Y(g3235),.A(I13101));
  NOT NOT1_10(.VSS(VSS),.VDD(VDD),.Y(I13104),.A(g2));
  NOT NOT1_11(.VSS(VSS),.VDD(VDD),.Y(g3236),.A(I13104));
  NOT NOT1_12(.VSS(VSS),.VDD(VDD),.Y(I13107),.A(g5));
  NOT NOT1_13(.VSS(VSS),.VDD(VDD),.Y(g3237),.A(I13107));
  NOT NOT1_14(.VSS(VSS),.VDD(VDD),.Y(I13110),.A(g8));
  NOT NOT1_15(.VSS(VSS),.VDD(VDD),.Y(g3238),.A(I13110));
  NOT NOT1_16(.VSS(VSS),.VDD(VDD),.Y(I13113),.A(g11));
  NOT NOT1_17(.VSS(VSS),.VDD(VDD),.Y(g3239),.A(I13113));
  NOT NOT1_18(.VSS(VSS),.VDD(VDD),.Y(I13116),.A(g14));
  NOT NOT1_19(.VSS(VSS),.VDD(VDD),.Y(g3240),.A(I13116));
  NOT NOT1_20(.VSS(VSS),.VDD(VDD),.Y(I13119),.A(g17));
  NOT NOT1_21(.VSS(VSS),.VDD(VDD),.Y(g3241),.A(I13119));
  NOT NOT1_22(.VSS(VSS),.VDD(VDD),.Y(I13122),.A(g20));
  NOT NOT1_23(.VSS(VSS),.VDD(VDD),.Y(g3242),.A(I13122));
  NOT NOT1_24(.VSS(VSS),.VDD(VDD),.Y(I13125),.A(g23));
  NOT NOT1_25(.VSS(VSS),.VDD(VDD),.Y(g3243),.A(I13125));
  NOT NOT1_26(.VSS(VSS),.VDD(VDD),.Y(I13128),.A(g26));
  NOT NOT1_27(.VSS(VSS),.VDD(VDD),.Y(g3244),.A(I13128));
  NOT NOT1_28(.VSS(VSS),.VDD(VDD),.Y(I13131),.A(g27));
  NOT NOT1_29(.VSS(VSS),.VDD(VDD),.Y(g3245),.A(I13131));
  NOT NOT1_30(.VSS(VSS),.VDD(VDD),.Y(I13134),.A(g30));
  NOT NOT1_31(.VSS(VSS),.VDD(VDD),.Y(g3246),.A(I13134));
  NOT NOT1_32(.VSS(VSS),.VDD(VDD),.Y(I13137),.A(g33));
  NOT NOT1_33(.VSS(VSS),.VDD(VDD),.Y(g3247),.A(I13137));
  NOT NOT1_34(.VSS(VSS),.VDD(VDD),.Y(I13140),.A(g36));
  NOT NOT1_35(.VSS(VSS),.VDD(VDD),.Y(g3248),.A(I13140));
  NOT NOT1_36(.VSS(VSS),.VDD(VDD),.Y(I13143),.A(g39));
  NOT NOT1_37(.VSS(VSS),.VDD(VDD),.Y(g3249),.A(I13143));
  NOT NOT1_38(.VSS(VSS),.VDD(VDD),.Y(I13146),.A(g42));
  NOT NOT1_39(.VSS(VSS),.VDD(VDD),.Y(g3250),.A(I13146));
  NOT NOT1_40(.VSS(VSS),.VDD(VDD),.Y(I13149),.A(g45));
  NOT NOT1_41(.VSS(VSS),.VDD(VDD),.Y(g3251),.A(I13149));
  NOT NOT1_42(.VSS(VSS),.VDD(VDD),.Y(I13152),.A(g48));
  NOT NOT1_43(.VSS(VSS),.VDD(VDD),.Y(g3252),.A(I13152));
  NOT NOT1_44(.VSS(VSS),.VDD(VDD),.Y(I13155),.A(g51));
  NOT NOT1_45(.VSS(VSS),.VDD(VDD),.Y(g3253),.A(I13155));
  NOT NOT1_46(.VSS(VSS),.VDD(VDD),.Y(I13158),.A(g165));
  NOT NOT1_47(.VSS(VSS),.VDD(VDD),.Y(g3254),.A(I13158));
  NOT NOT1_48(.VSS(VSS),.VDD(VDD),.Y(I13161),.A(g308));
  NOT NOT1_49(.VSS(VSS),.VDD(VDD),.Y(g3304),.A(I13161));
  NOT NOT1_50(.VSS(VSS),.VDD(VDD),.Y(g3305),.A(g305));
  NOT NOT1_51(.VSS(VSS),.VDD(VDD),.Y(I13165),.A(g401));
  NOT NOT1_52(.VSS(VSS),.VDD(VDD),.Y(g3306),.A(I13165));
  NOT NOT1_53(.VSS(VSS),.VDD(VDD),.Y(g3337),.A(g309));
  NOT NOT1_54(.VSS(VSS),.VDD(VDD),.Y(I13169),.A(g550));
  NOT NOT1_55(.VSS(VSS),.VDD(VDD),.Y(g3338),.A(I13169));
  NOT NOT1_56(.VSS(VSS),.VDD(VDD),.Y(g3365),.A(g499));
  NOT NOT1_57(.VSS(VSS),.VDD(VDD),.Y(I13173),.A(g629));
  NOT NOT1_58(.VSS(VSS),.VDD(VDD),.Y(g3366),.A(I13173));
  NOT NOT1_59(.VSS(VSS),.VDD(VDD),.Y(I13176),.A(g630));
  NOT NOT1_60(.VSS(VSS),.VDD(VDD),.Y(g3398),.A(I13176));
  NOT NOT1_61(.VSS(VSS),.VDD(VDD),.Y(I13179),.A(g853));
  NOT NOT1_62(.VSS(VSS),.VDD(VDD),.Y(g3410),.A(I13179));
  NOT NOT1_63(.VSS(VSS),.VDD(VDD),.Y(I13182),.A(g995));
  NOT NOT1_64(.VSS(VSS),.VDD(VDD),.Y(g3460),.A(I13182));
  NOT NOT1_65(.VSS(VSS),.VDD(VDD),.Y(g3461),.A(g992));
  NOT NOT1_66(.VSS(VSS),.VDD(VDD),.Y(I13186),.A(g1088));
  NOT NOT1_67(.VSS(VSS),.VDD(VDD),.Y(g3462),.A(I13186));
  NOT NOT1_68(.VSS(VSS),.VDD(VDD),.Y(g3493),.A(g996));
  NOT NOT1_69(.VSS(VSS),.VDD(VDD),.Y(I13190),.A(g1236));
  NOT NOT1_70(.VSS(VSS),.VDD(VDD),.Y(g3494),.A(I13190));
  NOT NOT1_71(.VSS(VSS),.VDD(VDD),.Y(g3521),.A(g1186));
  NOT NOT1_72(.VSS(VSS),.VDD(VDD),.Y(I13194),.A(g1315));
  NOT NOT1_73(.VSS(VSS),.VDD(VDD),.Y(g3522),.A(I13194));
  NOT NOT1_74(.VSS(VSS),.VDD(VDD),.Y(I13197),.A(g1316));
  NOT NOT1_75(.VSS(VSS),.VDD(VDD),.Y(g3554),.A(I13197));
  NOT NOT1_76(.VSS(VSS),.VDD(VDD),.Y(I13200),.A(g1547));
  NOT NOT1_77(.VSS(VSS),.VDD(VDD),.Y(g3566),.A(I13200));
  NOT NOT1_78(.VSS(VSS),.VDD(VDD),.Y(I13203),.A(g1689));
  NOT NOT1_79(.VSS(VSS),.VDD(VDD),.Y(g3616),.A(I13203));
  NOT NOT1_80(.VSS(VSS),.VDD(VDD),.Y(g3617),.A(g1686));
  NOT NOT1_81(.VSS(VSS),.VDD(VDD),.Y(I13207),.A(g1782));
  NOT NOT1_82(.VSS(VSS),.VDD(VDD),.Y(g3618),.A(I13207));
  NOT NOT1_83(.VSS(VSS),.VDD(VDD),.Y(g3649),.A(g1690));
  NOT NOT1_84(.VSS(VSS),.VDD(VDD),.Y(I13211),.A(g1930));
  NOT NOT1_85(.VSS(VSS),.VDD(VDD),.Y(g3650),.A(I13211));
  NOT NOT1_86(.VSS(VSS),.VDD(VDD),.Y(g3677),.A(g1880));
  NOT NOT1_87(.VSS(VSS),.VDD(VDD),.Y(I13215),.A(g2009));
  NOT NOT1_88(.VSS(VSS),.VDD(VDD),.Y(g3678),.A(I13215));
  NOT NOT1_89(.VSS(VSS),.VDD(VDD),.Y(I13218),.A(g2010));
  NOT NOT1_90(.VSS(VSS),.VDD(VDD),.Y(g3710),.A(I13218));
  NOT NOT1_91(.VSS(VSS),.VDD(VDD),.Y(I13221),.A(g2241));
  NOT NOT1_92(.VSS(VSS),.VDD(VDD),.Y(g3722),.A(I13221));
  NOT NOT1_93(.VSS(VSS),.VDD(VDD),.Y(I13224),.A(g2383));
  NOT NOT1_94(.VSS(VSS),.VDD(VDD),.Y(g3772),.A(I13224));
  NOT NOT1_95(.VSS(VSS),.VDD(VDD),.Y(g3773),.A(g2380));
  NOT NOT1_96(.VSS(VSS),.VDD(VDD),.Y(I13228),.A(g2476));
  NOT NOT1_97(.VSS(VSS),.VDD(VDD),.Y(g3774),.A(I13228));
  NOT NOT1_98(.VSS(VSS),.VDD(VDD),.Y(g3805),.A(g2384));
  NOT NOT1_99(.VSS(VSS),.VDD(VDD),.Y(I13232),.A(g2624));
  NOT NOT1_100(.VSS(VSS),.VDD(VDD),.Y(g3806),.A(I13232));
  NOT NOT1_101(.VSS(VSS),.VDD(VDD),.Y(g3833),.A(g2574));
  NOT NOT1_102(.VSS(VSS),.VDD(VDD),.Y(I13236),.A(g2703));
  NOT NOT1_103(.VSS(VSS),.VDD(VDD),.Y(g3834),.A(I13236));
  NOT NOT1_104(.VSS(VSS),.VDD(VDD),.Y(I13239),.A(g2704));
  NOT NOT1_105(.VSS(VSS),.VDD(VDD),.Y(g3866),.A(I13239));
  NOT NOT1_106(.VSS(VSS),.VDD(VDD),.Y(I13242),.A(g2879));
  NOT NOT1_107(.VSS(VSS),.VDD(VDD),.Y(g3878),.A(I13242));
  NOT NOT1_108(.VSS(VSS),.VDD(VDD),.Y(g3897),.A(g2950));
  NOT NOT1_109(.VSS(VSS),.VDD(VDD),.Y(I13246),.A(g2987));
  NOT NOT1_110(.VSS(VSS),.VDD(VDD),.Y(g3900),.A(I13246));
  NOT NOT1_111(.VSS(VSS),.VDD(VDD),.Y(g3919),.A(g3080));
  NOT NOT1_112(.VSS(VSS),.VDD(VDD),.Y(g3922),.A(g150));
  NOT NOT1_113(.VSS(VSS),.VDD(VDD),.Y(g3925),.A(g155));
  NOT NOT1_114(.VSS(VSS),.VDD(VDD),.Y(g3928),.A(g157));
  NOT NOT1_115(.VSS(VSS),.VDD(VDD),.Y(g3931),.A(g171));
  NOT NOT1_116(.VSS(VSS),.VDD(VDD),.Y(g3934),.A(g176));
  NOT NOT1_117(.VSS(VSS),.VDD(VDD),.Y(g3937),.A(g178));
  NOT NOT1_118(.VSS(VSS),.VDD(VDD),.Y(g3940),.A(g408));
  NOT NOT1_119(.VSS(VSS),.VDD(VDD),.Y(g3941),.A(g455));
  NOT NOT1_120(.VSS(VSS),.VDD(VDD),.Y(g3942),.A(g699));
  NOT NOT1_121(.VSS(VSS),.VDD(VDD),.Y(g3945),.A(g726));
  NOT NOT1_122(.VSS(VSS),.VDD(VDD),.Y(g3948),.A(g835));
  NOT NOT1_123(.VSS(VSS),.VDD(VDD),.Y(g3951),.A(g840));
  NOT NOT1_124(.VSS(VSS),.VDD(VDD),.Y(g3954),.A(g842));
  NOT NOT1_125(.VSS(VSS),.VDD(VDD),.Y(g3957),.A(g856));
  NOT NOT1_126(.VSS(VSS),.VDD(VDD),.Y(g3960),.A(g861));
  NOT NOT1_127(.VSS(VSS),.VDD(VDD),.Y(g3963),.A(g863));
  NOT NOT1_128(.VSS(VSS),.VDD(VDD),.Y(g3966),.A(g1526));
  NOT NOT1_129(.VSS(VSS),.VDD(VDD),.Y(g3969),.A(g1531));
  NOT NOT1_130(.VSS(VSS),.VDD(VDD),.Y(g3972),.A(g1533));
  NOT NOT1_131(.VSS(VSS),.VDD(VDD),.Y(g3975),.A(g1552));
  NOT NOT1_132(.VSS(VSS),.VDD(VDD),.Y(g3978),.A(g1554));
  NOT NOT1_133(.VSS(VSS),.VDD(VDD),.Y(g3981),.A(g2217));
  NOT NOT1_134(.VSS(VSS),.VDD(VDD),.Y(g3984),.A(g2222));
  NOT NOT1_135(.VSS(VSS),.VDD(VDD),.Y(g3987),.A(g2224));
  NOT NOT1_136(.VSS(VSS),.VDD(VDD),.Y(g3990),.A(g2245));
  NOT NOT1_137(.VSS(VSS),.VDD(VDD),.Y(I13275),.A(g2848));
  NOT NOT1_138(.VSS(VSS),.VDD(VDD),.Y(g3993),.A(I13275));
  NOT NOT1_139(.VSS(VSS),.VDD(VDD),.Y(g3994),.A(g2848));
  NOT NOT1_140(.VSS(VSS),.VDD(VDD),.Y(g3995),.A(g3064));
  NOT NOT1_141(.VSS(VSS),.VDD(VDD),.Y(g3996),.A(g3073));
  NOT NOT1_142(.VSS(VSS),.VDD(VDD),.Y(g3997),.A(g45));
  NOT NOT1_143(.VSS(VSS),.VDD(VDD),.Y(g3998),.A(g23));
  NOT NOT1_144(.VSS(VSS),.VDD(VDD),.Y(g3999),.A(g3204));
  NOT NOT1_145(.VSS(VSS),.VDD(VDD),.Y(g4000),.A(g153));
  NOT NOT1_146(.VSS(VSS),.VDD(VDD),.Y(g4003),.A(g158));
  NOT NOT1_147(.VSS(VSS),.VDD(VDD),.Y(g4006),.A(g160));
  NOT NOT1_148(.VSS(VSS),.VDD(VDD),.Y(g4009),.A(g174));
  NOT NOT1_149(.VSS(VSS),.VDD(VDD),.Y(g4012),.A(g179));
  NOT NOT1_150(.VSS(VSS),.VDD(VDD),.Y(g4015),.A(g411));
  NOT NOT1_151(.VSS(VSS),.VDD(VDD),.Y(g4016),.A(g417));
  NOT NOT1_152(.VSS(VSS),.VDD(VDD),.Y(g4017),.A(g427));
  NOT NOT1_153(.VSS(VSS),.VDD(VDD),.Y(g4020),.A(g700));
  NOT NOT1_154(.VSS(VSS),.VDD(VDD),.Y(g4023),.A(g702));
  NOT NOT1_155(.VSS(VSS),.VDD(VDD),.Y(g4026),.A(g727));
  NOT NOT1_156(.VSS(VSS),.VDD(VDD),.Y(g4029),.A(g838));
  NOT NOT1_157(.VSS(VSS),.VDD(VDD),.Y(g4032),.A(g843));
  NOT NOT1_158(.VSS(VSS),.VDD(VDD),.Y(g4035),.A(g845));
  NOT NOT1_159(.VSS(VSS),.VDD(VDD),.Y(g4038),.A(g859));
  NOT NOT1_160(.VSS(VSS),.VDD(VDD),.Y(g4041),.A(g864));
  NOT NOT1_161(.VSS(VSS),.VDD(VDD),.Y(g4044),.A(g866));
  NOT NOT1_162(.VSS(VSS),.VDD(VDD),.Y(g4047),.A(g1095));
  NOT NOT1_163(.VSS(VSS),.VDD(VDD),.Y(g4048),.A(g1142));
  NOT NOT1_164(.VSS(VSS),.VDD(VDD),.Y(g4049),.A(g1385));
  NOT NOT1_165(.VSS(VSS),.VDD(VDD),.Y(g4052),.A(g1412));
  NOT NOT1_166(.VSS(VSS),.VDD(VDD),.Y(g4055),.A(g1529));
  NOT NOT1_167(.VSS(VSS),.VDD(VDD),.Y(g4058),.A(g1534));
  NOT NOT1_168(.VSS(VSS),.VDD(VDD),.Y(g4061),.A(g1536));
  NOT NOT1_169(.VSS(VSS),.VDD(VDD),.Y(g4064),.A(g1550));
  NOT NOT1_170(.VSS(VSS),.VDD(VDD),.Y(g4067),.A(g1555));
  NOT NOT1_171(.VSS(VSS),.VDD(VDD),.Y(g4070),.A(g1557));
  NOT NOT1_172(.VSS(VSS),.VDD(VDD),.Y(g4073),.A(g2220));
  NOT NOT1_173(.VSS(VSS),.VDD(VDD),.Y(g4076),.A(g2225));
  NOT NOT1_174(.VSS(VSS),.VDD(VDD),.Y(g4079),.A(g2227));
  NOT NOT1_175(.VSS(VSS),.VDD(VDD),.Y(g4082),.A(g2246));
  NOT NOT1_176(.VSS(VSS),.VDD(VDD),.Y(g4085),.A(g2248));
  NOT NOT1_177(.VSS(VSS),.VDD(VDD),.Y(I13316),.A(g2836));
  NOT NOT1_178(.VSS(VSS),.VDD(VDD),.Y(g4088),.A(I13316));
  NOT NOT1_179(.VSS(VSS),.VDD(VDD),.Y(g4089),.A(g2836));
  NOT NOT1_180(.VSS(VSS),.VDD(VDD),.Y(I13320),.A(g2864));
  NOT NOT1_181(.VSS(VSS),.VDD(VDD),.Y(g4090),.A(I13320));
  NOT NOT1_182(.VSS(VSS),.VDD(VDD),.Y(g4091),.A(g2864));
  NOT NOT1_183(.VSS(VSS),.VDD(VDD),.Y(g4092),.A(g3074));
  NOT NOT1_184(.VSS(VSS),.VDD(VDD),.Y(g4093),.A(g33));
  NOT NOT1_185(.VSS(VSS),.VDD(VDD),.Y(g4094),.A(g3207));
  NOT NOT1_186(.VSS(VSS),.VDD(VDD),.Y(g4095),.A(g130));
  NOT NOT1_187(.VSS(VSS),.VDD(VDD),.Y(g4098),.A(g156));
  NOT NOT1_188(.VSS(VSS),.VDD(VDD),.Y(g4101),.A(g161));
  NOT NOT1_189(.VSS(VSS),.VDD(VDD),.Y(g4104),.A(g163));
  NOT NOT1_190(.VSS(VSS),.VDD(VDD),.Y(g4107),.A(g177));
  NOT NOT1_191(.VSS(VSS),.VDD(VDD),.Y(g4110),.A(g414));
  NOT NOT1_192(.VSS(VSS),.VDD(VDD),.Y(g4111),.A(g420));
  NOT NOT1_193(.VSS(VSS),.VDD(VDD),.Y(g4112),.A(g428));
  NOT NOT1_194(.VSS(VSS),.VDD(VDD),.Y(g4115),.A(g698));
  NOT NOT1_195(.VSS(VSS),.VDD(VDD),.Y(g4118),.A(g703));
  NOT NOT1_196(.VSS(VSS),.VDD(VDD),.Y(g4121),.A(g705));
  NOT NOT1_197(.VSS(VSS),.VDD(VDD),.Y(g4124),.A(g725));
  NOT NOT1_198(.VSS(VSS),.VDD(VDD),.Y(g4127),.A(g841));
  NOT NOT1_199(.VSS(VSS),.VDD(VDD),.Y(g4130),.A(g846));
  NOT NOT1_200(.VSS(VSS),.VDD(VDD),.Y(g4133),.A(g848));
  NOT NOT1_201(.VSS(VSS),.VDD(VDD),.Y(g4136),.A(g862));
  NOT NOT1_202(.VSS(VSS),.VDD(VDD),.Y(g4139),.A(g867));
  NOT NOT1_203(.VSS(VSS),.VDD(VDD),.Y(g4142),.A(g1098));
  NOT NOT1_204(.VSS(VSS),.VDD(VDD),.Y(g4143),.A(g1104));
  NOT NOT1_205(.VSS(VSS),.VDD(VDD),.Y(g4144),.A(g1114));
  NOT NOT1_206(.VSS(VSS),.VDD(VDD),.Y(g4147),.A(g1386));
  NOT NOT1_207(.VSS(VSS),.VDD(VDD),.Y(g4150),.A(g1388));
  NOT NOT1_208(.VSS(VSS),.VDD(VDD),.Y(g4153),.A(g1413));
  NOT NOT1_209(.VSS(VSS),.VDD(VDD),.Y(g4156),.A(g1532));
  NOT NOT1_210(.VSS(VSS),.VDD(VDD),.Y(g4159),.A(g1537));
  NOT NOT1_211(.VSS(VSS),.VDD(VDD),.Y(g4162),.A(g1539));
  NOT NOT1_212(.VSS(VSS),.VDD(VDD),.Y(g4165),.A(g1553));
  NOT NOT1_213(.VSS(VSS),.VDD(VDD),.Y(g4168),.A(g1558));
  NOT NOT1_214(.VSS(VSS),.VDD(VDD),.Y(g4171),.A(g1560));
  NOT NOT1_215(.VSS(VSS),.VDD(VDD),.Y(g4174),.A(g1789));
  NOT NOT1_216(.VSS(VSS),.VDD(VDD),.Y(g4175),.A(g1836));
  NOT NOT1_217(.VSS(VSS),.VDD(VDD),.Y(g4176),.A(g2079));
  NOT NOT1_218(.VSS(VSS),.VDD(VDD),.Y(g4179),.A(g2106));
  NOT NOT1_219(.VSS(VSS),.VDD(VDD),.Y(g4182),.A(g2223));
  NOT NOT1_220(.VSS(VSS),.VDD(VDD),.Y(g4185),.A(g2228));
  NOT NOT1_221(.VSS(VSS),.VDD(VDD),.Y(g4188),.A(g2230));
  NOT NOT1_222(.VSS(VSS),.VDD(VDD),.Y(g4191),.A(g2244));
  NOT NOT1_223(.VSS(VSS),.VDD(VDD),.Y(g4194),.A(g2249));
  NOT NOT1_224(.VSS(VSS),.VDD(VDD),.Y(g4197),.A(g2251));
  NOT NOT1_225(.VSS(VSS),.VDD(VDD),.Y(I13366),.A(g2851));
  NOT NOT1_226(.VSS(VSS),.VDD(VDD),.Y(g4200),.A(I13366));
  NOT NOT1_227(.VSS(VSS),.VDD(VDD),.Y(g4201),.A(g2851));
  NOT NOT1_228(.VSS(VSS),.VDD(VDD),.Y(g4202),.A(g42));
  NOT NOT1_229(.VSS(VSS),.VDD(VDD),.Y(g4203),.A(g20));
  NOT NOT1_230(.VSS(VSS),.VDD(VDD),.Y(g4204),.A(g3188));
  NOT NOT1_231(.VSS(VSS),.VDD(VDD),.Y(g4205),.A(g131));
  NOT NOT1_232(.VSS(VSS),.VDD(VDD),.Y(g4208),.A(g133));
  NOT NOT1_233(.VSS(VSS),.VDD(VDD),.Y(g4211),.A(g159));
  NOT NOT1_234(.VSS(VSS),.VDD(VDD),.Y(g4214),.A(g164));
  NOT NOT1_235(.VSS(VSS),.VDD(VDD),.Y(g4217),.A(g354));
  NOT NOT1_236(.VSS(VSS),.VDD(VDD),.Y(g4220),.A(g423));
  NOT NOT1_237(.VSS(VSS),.VDD(VDD),.Y(g4221),.A(g426));
  NOT NOT1_238(.VSS(VSS),.VDD(VDD),.Y(g4224),.A(g429));
  NOT NOT1_239(.VSS(VSS),.VDD(VDD),.Y(g4225),.A(g701));
  NOT NOT1_240(.VSS(VSS),.VDD(VDD),.Y(g4228),.A(g706));
  NOT NOT1_241(.VSS(VSS),.VDD(VDD),.Y(g4231),.A(g708));
  NOT NOT1_242(.VSS(VSS),.VDD(VDD),.Y(g4234),.A(g818));
  NOT NOT1_243(.VSS(VSS),.VDD(VDD),.Y(g4237),.A(g844));
  NOT NOT1_244(.VSS(VSS),.VDD(VDD),.Y(g4240),.A(g849));
  NOT NOT1_245(.VSS(VSS),.VDD(VDD),.Y(g4243),.A(g851));
  NOT NOT1_246(.VSS(VSS),.VDD(VDD),.Y(g4246),.A(g865));
  NOT NOT1_247(.VSS(VSS),.VDD(VDD),.Y(g4249),.A(g1101));
  NOT NOT1_248(.VSS(VSS),.VDD(VDD),.Y(g4250),.A(g1107));
  NOT NOT1_249(.VSS(VSS),.VDD(VDD),.Y(g4251),.A(g1115));
  NOT NOT1_250(.VSS(VSS),.VDD(VDD),.Y(g4254),.A(g1384));
  NOT NOT1_251(.VSS(VSS),.VDD(VDD),.Y(g4257),.A(g1389));
  NOT NOT1_252(.VSS(VSS),.VDD(VDD),.Y(g4260),.A(g1391));
  NOT NOT1_253(.VSS(VSS),.VDD(VDD),.Y(g4263),.A(g1411));
  NOT NOT1_254(.VSS(VSS),.VDD(VDD),.Y(g4266),.A(g1535));
  NOT NOT1_255(.VSS(VSS),.VDD(VDD),.Y(g4269),.A(g1540));
  NOT NOT1_256(.VSS(VSS),.VDD(VDD),.Y(g4272),.A(g1542));
  NOT NOT1_257(.VSS(VSS),.VDD(VDD),.Y(g4275),.A(g1556));
  NOT NOT1_258(.VSS(VSS),.VDD(VDD),.Y(g4278),.A(g1561));
  NOT NOT1_259(.VSS(VSS),.VDD(VDD),.Y(g4281),.A(g1792));
  NOT NOT1_260(.VSS(VSS),.VDD(VDD),.Y(g4282),.A(g1798));
  NOT NOT1_261(.VSS(VSS),.VDD(VDD),.Y(g4283),.A(g1808));
  NOT NOT1_262(.VSS(VSS),.VDD(VDD),.Y(g4286),.A(g2080));
  NOT NOT1_263(.VSS(VSS),.VDD(VDD),.Y(g4289),.A(g2082));
  NOT NOT1_264(.VSS(VSS),.VDD(VDD),.Y(g4292),.A(g2107));
  NOT NOT1_265(.VSS(VSS),.VDD(VDD),.Y(g4295),.A(g2226));
  NOT NOT1_266(.VSS(VSS),.VDD(VDD),.Y(g4298),.A(g2231));
  NOT NOT1_267(.VSS(VSS),.VDD(VDD),.Y(g4301),.A(g2233));
  NOT NOT1_268(.VSS(VSS),.VDD(VDD),.Y(g4304),.A(g2247));
  NOT NOT1_269(.VSS(VSS),.VDD(VDD),.Y(g4307),.A(g2252));
  NOT NOT1_270(.VSS(VSS),.VDD(VDD),.Y(g4310),.A(g2254));
  NOT NOT1_271(.VSS(VSS),.VDD(VDD),.Y(g4313),.A(g2483));
  NOT NOT1_272(.VSS(VSS),.VDD(VDD),.Y(g4314),.A(g2530));
  NOT NOT1_273(.VSS(VSS),.VDD(VDD),.Y(g4315),.A(g2773));
  NOT NOT1_274(.VSS(VSS),.VDD(VDD),.Y(g4318),.A(g2800));
  NOT NOT1_275(.VSS(VSS),.VDD(VDD),.Y(I13417),.A(g2839));
  NOT NOT1_276(.VSS(VSS),.VDD(VDD),.Y(g4321),.A(I13417));
  NOT NOT1_277(.VSS(VSS),.VDD(VDD),.Y(g4322),.A(g2839));
  NOT NOT1_278(.VSS(VSS),.VDD(VDD),.Y(I13421),.A(g2867));
  NOT NOT1_279(.VSS(VSS),.VDD(VDD),.Y(g4323),.A(I13421));
  NOT NOT1_280(.VSS(VSS),.VDD(VDD),.Y(g4324),.A(g2867));
  NOT NOT1_281(.VSS(VSS),.VDD(VDD),.Y(g4325),.A(g36));
  NOT NOT1_282(.VSS(VSS),.VDD(VDD),.Y(g4326),.A(g181));
  NOT NOT1_283(.VSS(VSS),.VDD(VDD),.Y(g4329),.A(g129));
  NOT NOT1_284(.VSS(VSS),.VDD(VDD),.Y(g4332),.A(g134));
  NOT NOT1_285(.VSS(VSS),.VDD(VDD),.Y(g4335),.A(g162));
  NOT NOT1_286(.VSS(VSS),.VDD(VDD),.Y(I13430),.A(g101));
  NOT NOT1_287(.VSS(VSS),.VDD(VDD),.Y(g4338),.A(I13430));
  NOT NOT1_288(.VSS(VSS),.VDD(VDD),.Y(I13433),.A(g105));
  NOT NOT1_289(.VSS(VSS),.VDD(VDD),.Y(g4339),.A(I13433));
  NOT NOT1_290(.VSS(VSS),.VDD(VDD),.Y(g4340),.A(g343));
  NOT NOT1_291(.VSS(VSS),.VDD(VDD),.Y(g4343),.A(g369));
  NOT NOT1_292(.VSS(VSS),.VDD(VDD),.Y(g4346),.A(g432));
  NOT NOT1_293(.VSS(VSS),.VDD(VDD),.Y(g4347),.A(g438));
  NOT NOT1_294(.VSS(VSS),.VDD(VDD),.Y(g4348),.A(g704));
  NOT NOT1_295(.VSS(VSS),.VDD(VDD),.Y(g4351),.A(g709));
  NOT NOT1_296(.VSS(VSS),.VDD(VDD),.Y(g4354),.A(g711));
  NOT NOT1_297(.VSS(VSS),.VDD(VDD),.Y(g4357),.A(g729));
  NOT NOT1_298(.VSS(VSS),.VDD(VDD),.Y(g4360),.A(g819));
  NOT NOT1_299(.VSS(VSS),.VDD(VDD),.Y(g4363),.A(g821));
  NOT NOT1_300(.VSS(VSS),.VDD(VDD),.Y(g4366),.A(g847));
  NOT NOT1_301(.VSS(VSS),.VDD(VDD),.Y(g4369),.A(g852));
  NOT NOT1_302(.VSS(VSS),.VDD(VDD),.Y(g4372),.A(g1041));
  NOT NOT1_303(.VSS(VSS),.VDD(VDD),.Y(g4375),.A(g1110));
  NOT NOT1_304(.VSS(VSS),.VDD(VDD),.Y(g4376),.A(g1113));
  NOT NOT1_305(.VSS(VSS),.VDD(VDD),.Y(g4379),.A(g1116));
  NOT NOT1_306(.VSS(VSS),.VDD(VDD),.Y(g4380),.A(g1387));
  NOT NOT1_307(.VSS(VSS),.VDD(VDD),.Y(g4383),.A(g1392));
  NOT NOT1_308(.VSS(VSS),.VDD(VDD),.Y(g4386),.A(g1394));
  NOT NOT1_309(.VSS(VSS),.VDD(VDD),.Y(g4389),.A(g1512));
  NOT NOT1_310(.VSS(VSS),.VDD(VDD),.Y(g4392),.A(g1538));
  NOT NOT1_311(.VSS(VSS),.VDD(VDD),.Y(g4395),.A(g1543));
  NOT NOT1_312(.VSS(VSS),.VDD(VDD),.Y(g4398),.A(g1545));
  NOT NOT1_313(.VSS(VSS),.VDD(VDD),.Y(g4401),.A(g1559));
  NOT NOT1_314(.VSS(VSS),.VDD(VDD),.Y(g4404),.A(g1795));
  NOT NOT1_315(.VSS(VSS),.VDD(VDD),.Y(g4405),.A(g1801));
  NOT NOT1_316(.VSS(VSS),.VDD(VDD),.Y(g4406),.A(g1809));
  NOT NOT1_317(.VSS(VSS),.VDD(VDD),.Y(g4409),.A(g2078));
  NOT NOT1_318(.VSS(VSS),.VDD(VDD),.Y(g4412),.A(g2083));
  NOT NOT1_319(.VSS(VSS),.VDD(VDD),.Y(g4415),.A(g2085));
  NOT NOT1_320(.VSS(VSS),.VDD(VDD),.Y(g4418),.A(g2105));
  NOT NOT1_321(.VSS(VSS),.VDD(VDD),.Y(g4421),.A(g2229));
  NOT NOT1_322(.VSS(VSS),.VDD(VDD),.Y(g4424),.A(g2234));
  NOT NOT1_323(.VSS(VSS),.VDD(VDD),.Y(g4427),.A(g2236));
  NOT NOT1_324(.VSS(VSS),.VDD(VDD),.Y(g4430),.A(g2250));
  NOT NOT1_325(.VSS(VSS),.VDD(VDD),.Y(g4433),.A(g2255));
  NOT NOT1_326(.VSS(VSS),.VDD(VDD),.Y(g4436),.A(g2486));
  NOT NOT1_327(.VSS(VSS),.VDD(VDD),.Y(g4437),.A(g2492));
  NOT NOT1_328(.VSS(VSS),.VDD(VDD),.Y(g4438),.A(g2502));
  NOT NOT1_329(.VSS(VSS),.VDD(VDD),.Y(g4441),.A(g2774));
  NOT NOT1_330(.VSS(VSS),.VDD(VDD),.Y(g4444),.A(g2776));
  NOT NOT1_331(.VSS(VSS),.VDD(VDD),.Y(g4447),.A(g2801));
  NOT NOT1_332(.VSS(VSS),.VDD(VDD),.Y(I13478),.A(g2854));
  NOT NOT1_333(.VSS(VSS),.VDD(VDD),.Y(g4450),.A(I13478));
  NOT NOT1_334(.VSS(VSS),.VDD(VDD),.Y(g4451),.A(g2854));
  NOT NOT1_335(.VSS(VSS),.VDD(VDD),.Y(g4452),.A(g17));
  NOT NOT1_336(.VSS(VSS),.VDD(VDD),.Y(g4453),.A(g132));
  NOT NOT1_337(.VSS(VSS),.VDD(VDD),.Y(g4456),.A(g309));
  NOT NOT1_338(.VSS(VSS),.VDD(VDD),.Y(g4465),.A(g346));
  NOT NOT1_339(.VSS(VSS),.VDD(VDD),.Y(g4468),.A(g358));
  NOT NOT1_340(.VSS(VSS),.VDD(VDD),.Y(g4471),.A(g384));
  NOT NOT1_341(.VSS(VSS),.VDD(VDD),.Y(g4474),.A(g435));
  NOT NOT1_342(.VSS(VSS),.VDD(VDD),.Y(g4475),.A(g441));
  NOT NOT1_343(.VSS(VSS),.VDD(VDD),.Y(g4476),.A(g576));
  NOT NOT1_344(.VSS(VSS),.VDD(VDD),.Y(g4479),.A(g587));
  NOT NOT1_345(.VSS(VSS),.VDD(VDD),.Y(g4480),.A(g707));
  NOT NOT1_346(.VSS(VSS),.VDD(VDD),.Y(g4483),.A(g712));
  NOT NOT1_347(.VSS(VSS),.VDD(VDD),.Y(g4486),.A(g714));
  NOT NOT1_348(.VSS(VSS),.VDD(VDD),.Y(g4489),.A(g730));
  NOT NOT1_349(.VSS(VSS),.VDD(VDD),.Y(g4492),.A(g732));
  NOT NOT1_350(.VSS(VSS),.VDD(VDD),.Y(g4495),.A(g869));
  NOT NOT1_351(.VSS(VSS),.VDD(VDD),.Y(g4498),.A(g817));
  NOT NOT1_352(.VSS(VSS),.VDD(VDD),.Y(g4501),.A(g822));
  NOT NOT1_353(.VSS(VSS),.VDD(VDD),.Y(g4504),.A(g850));
  NOT NOT1_354(.VSS(VSS),.VDD(VDD),.Y(I13501),.A(g789));
  NOT NOT1_355(.VSS(VSS),.VDD(VDD),.Y(g4507),.A(I13501));
  NOT NOT1_356(.VSS(VSS),.VDD(VDD),.Y(I13504),.A(g793));
  NOT NOT1_357(.VSS(VSS),.VDD(VDD),.Y(g4508),.A(I13504));
  NOT NOT1_358(.VSS(VSS),.VDD(VDD),.Y(g4509),.A(g1030));
  NOT NOT1_359(.VSS(VSS),.VDD(VDD),.Y(g4512),.A(g1056));
  NOT NOT1_360(.VSS(VSS),.VDD(VDD),.Y(g4515),.A(g1119));
  NOT NOT1_361(.VSS(VSS),.VDD(VDD),.Y(g4516),.A(g1125));
  NOT NOT1_362(.VSS(VSS),.VDD(VDD),.Y(g4517),.A(g1390));
  NOT NOT1_363(.VSS(VSS),.VDD(VDD),.Y(g4520),.A(g1395));
  NOT NOT1_364(.VSS(VSS),.VDD(VDD),.Y(g4523),.A(g1397));
  NOT NOT1_365(.VSS(VSS),.VDD(VDD),.Y(g4526),.A(g1415));
  NOT NOT1_366(.VSS(VSS),.VDD(VDD),.Y(g4529),.A(g1513));
  NOT NOT1_367(.VSS(VSS),.VDD(VDD),.Y(g4532),.A(g1515));
  NOT NOT1_368(.VSS(VSS),.VDD(VDD),.Y(g4535),.A(g1541));
  NOT NOT1_369(.VSS(VSS),.VDD(VDD),.Y(g4538),.A(g1546));
  NOT NOT1_370(.VSS(VSS),.VDD(VDD),.Y(g4541),.A(g1735));
  NOT NOT1_371(.VSS(VSS),.VDD(VDD),.Y(g4544),.A(g1804));
  NOT NOT1_372(.VSS(VSS),.VDD(VDD),.Y(g4545),.A(g1807));
  NOT NOT1_373(.VSS(VSS),.VDD(VDD),.Y(g4548),.A(g1810));
  NOT NOT1_374(.VSS(VSS),.VDD(VDD),.Y(g4549),.A(g2081));
  NOT NOT1_375(.VSS(VSS),.VDD(VDD),.Y(g4552),.A(g2086));
  NOT NOT1_376(.VSS(VSS),.VDD(VDD),.Y(g4555),.A(g2088));
  NOT NOT1_377(.VSS(VSS),.VDD(VDD),.Y(g4558),.A(g2206));
  NOT NOT1_378(.VSS(VSS),.VDD(VDD),.Y(g4561),.A(g2232));
  NOT NOT1_379(.VSS(VSS),.VDD(VDD),.Y(g4564),.A(g2237));
  NOT NOT1_380(.VSS(VSS),.VDD(VDD),.Y(g4567),.A(g2239));
  NOT NOT1_381(.VSS(VSS),.VDD(VDD),.Y(g4570),.A(g2253));
  NOT NOT1_382(.VSS(VSS),.VDD(VDD),.Y(g4573),.A(g2489));
  NOT NOT1_383(.VSS(VSS),.VDD(VDD),.Y(g4574),.A(g2495));
  NOT NOT1_384(.VSS(VSS),.VDD(VDD),.Y(g4575),.A(g2503));
  NOT NOT1_385(.VSS(VSS),.VDD(VDD),.Y(g4578),.A(g2772));
  NOT NOT1_386(.VSS(VSS),.VDD(VDD),.Y(g4581),.A(g2777));
  NOT NOT1_387(.VSS(VSS),.VDD(VDD),.Y(g4584),.A(g2779));
  NOT NOT1_388(.VSS(VSS),.VDD(VDD),.Y(g4587),.A(g2799));
  NOT NOT1_389(.VSS(VSS),.VDD(VDD),.Y(I13538),.A(g2870));
  NOT NOT1_390(.VSS(VSS),.VDD(VDD),.Y(g4590),.A(I13538));
  NOT NOT1_391(.VSS(VSS),.VDD(VDD),.Y(g4591),.A(g2870));
  NOT NOT1_392(.VSS(VSS),.VDD(VDD),.Y(g4592),.A(g361));
  NOT NOT1_393(.VSS(VSS),.VDD(VDD),.Y(g4595),.A(g373));
  NOT NOT1_394(.VSS(VSS),.VDD(VDD),.Y(g4598),.A(g398));
  NOT NOT1_395(.VSS(VSS),.VDD(VDD),.Y(g4601),.A(g444));
  NOT NOT1_396(.VSS(VSS),.VDD(VDD),.Y(g4602),.A(g525));
  NOT NOT1_397(.VSS(VSS),.VDD(VDD),.Y(g4603),.A(g577));
  NOT NOT1_398(.VSS(VSS),.VDD(VDD),.Y(g4606),.A(g579));
  NOT NOT1_399(.VSS(VSS),.VDD(VDD),.Y(g4609),.A(g590));
  NOT NOT1_400(.VSS(VSS),.VDD(VDD),.Y(g4610),.A(g596));
  NOT NOT1_401(.VSS(VSS),.VDD(VDD),.Y(g4611),.A(g710));
  NOT NOT1_402(.VSS(VSS),.VDD(VDD),.Y(g4614),.A(g715));
  NOT NOT1_403(.VSS(VSS),.VDD(VDD),.Y(g4617),.A(g717));
  NOT NOT1_404(.VSS(VSS),.VDD(VDD),.Y(g4620),.A(g728));
  NOT NOT1_405(.VSS(VSS),.VDD(VDD),.Y(g4623),.A(g733));
  NOT NOT1_406(.VSS(VSS),.VDD(VDD),.Y(g4626),.A(g735));
  NOT NOT1_407(.VSS(VSS),.VDD(VDD),.Y(g4629),.A(g820));
  NOT NOT1_408(.VSS(VSS),.VDD(VDD),.Y(g4632),.A(g996));
  NOT NOT1_409(.VSS(VSS),.VDD(VDD),.Y(g4641),.A(g1033));
  NOT NOT1_410(.VSS(VSS),.VDD(VDD),.Y(g4644),.A(g1045));
  NOT NOT1_411(.VSS(VSS),.VDD(VDD),.Y(g4647),.A(g1071));
  NOT NOT1_412(.VSS(VSS),.VDD(VDD),.Y(g4650),.A(g1122));
  NOT NOT1_413(.VSS(VSS),.VDD(VDD),.Y(g4651),.A(g1128));
  NOT NOT1_414(.VSS(VSS),.VDD(VDD),.Y(g4652),.A(g1262));
  NOT NOT1_415(.VSS(VSS),.VDD(VDD),.Y(g4655),.A(g1273));
  NOT NOT1_416(.VSS(VSS),.VDD(VDD),.Y(g4656),.A(g1393));
  NOT NOT1_417(.VSS(VSS),.VDD(VDD),.Y(g4659),.A(g1398));
  NOT NOT1_418(.VSS(VSS),.VDD(VDD),.Y(g4662),.A(g1400));
  NOT NOT1_419(.VSS(VSS),.VDD(VDD),.Y(g4665),.A(g1416));
  NOT NOT1_420(.VSS(VSS),.VDD(VDD),.Y(g4668),.A(g1418));
  NOT NOT1_421(.VSS(VSS),.VDD(VDD),.Y(g4671),.A(g1563));
  NOT NOT1_422(.VSS(VSS),.VDD(VDD),.Y(g4674),.A(g1511));
  NOT NOT1_423(.VSS(VSS),.VDD(VDD),.Y(g4677),.A(g1516));
  NOT NOT1_424(.VSS(VSS),.VDD(VDD),.Y(g4680),.A(g1544));
  NOT NOT1_425(.VSS(VSS),.VDD(VDD),.Y(I13575),.A(g1476));
  NOT NOT1_426(.VSS(VSS),.VDD(VDD),.Y(g4683),.A(I13575));
  NOT NOT1_427(.VSS(VSS),.VDD(VDD),.Y(I13578),.A(g1481));
  NOT NOT1_428(.VSS(VSS),.VDD(VDD),.Y(g4684),.A(I13578));
  NOT NOT1_429(.VSS(VSS),.VDD(VDD),.Y(g4685),.A(g1724));
  NOT NOT1_430(.VSS(VSS),.VDD(VDD),.Y(g4688),.A(g1750));
  NOT NOT1_431(.VSS(VSS),.VDD(VDD),.Y(g4691),.A(g1813));
  NOT NOT1_432(.VSS(VSS),.VDD(VDD),.Y(g4692),.A(g1819));
  NOT NOT1_433(.VSS(VSS),.VDD(VDD),.Y(g4693),.A(g2084));
  NOT NOT1_434(.VSS(VSS),.VDD(VDD),.Y(g4696),.A(g2089));
  NOT NOT1_435(.VSS(VSS),.VDD(VDD),.Y(g4699),.A(g2091));
  NOT NOT1_436(.VSS(VSS),.VDD(VDD),.Y(g4702),.A(g2109));
  NOT NOT1_437(.VSS(VSS),.VDD(VDD),.Y(g4705),.A(g2207));
  NOT NOT1_438(.VSS(VSS),.VDD(VDD),.Y(g4708),.A(g2209));
  NOT NOT1_439(.VSS(VSS),.VDD(VDD),.Y(g4711),.A(g2235));
  NOT NOT1_440(.VSS(VSS),.VDD(VDD),.Y(g4714),.A(g2240));
  NOT NOT1_441(.VSS(VSS),.VDD(VDD),.Y(g4717),.A(g2429));
  NOT NOT1_442(.VSS(VSS),.VDD(VDD),.Y(g4720),.A(g2498));
  NOT NOT1_443(.VSS(VSS),.VDD(VDD),.Y(g4721),.A(g2501));
  NOT NOT1_444(.VSS(VSS),.VDD(VDD),.Y(g4724),.A(g2504));
  NOT NOT1_445(.VSS(VSS),.VDD(VDD),.Y(g4725),.A(g2775));
  NOT NOT1_446(.VSS(VSS),.VDD(VDD),.Y(g4728),.A(g2780));
  NOT NOT1_447(.VSS(VSS),.VDD(VDD),.Y(g4731),.A(g2782));
  NOT NOT1_448(.VSS(VSS),.VDD(VDD),.Y(g4734),.A(g11));
  NOT NOT1_449(.VSS(VSS),.VDD(VDD),.Y(I13601),.A(g121));
  NOT NOT1_450(.VSS(VSS),.VDD(VDD),.Y(g4735),.A(I13601));
  NOT NOT1_451(.VSS(VSS),.VDD(VDD),.Y(I13604),.A(g125));
  NOT NOT1_452(.VSS(VSS),.VDD(VDD),.Y(g4736),.A(I13604));
  NOT NOT1_453(.VSS(VSS),.VDD(VDD),.Y(g4737),.A(g376));
  NOT NOT1_454(.VSS(VSS),.VDD(VDD),.Y(g4740),.A(g388));
  NOT NOT1_455(.VSS(VSS),.VDD(VDD),.Y(g4743),.A(g575));
  NOT NOT1_456(.VSS(VSS),.VDD(VDD),.Y(g4746),.A(g580));
  NOT NOT1_457(.VSS(VSS),.VDD(VDD),.Y(g4749),.A(g582));
  NOT NOT1_458(.VSS(VSS),.VDD(VDD),.Y(g4752),.A(g593));
  NOT NOT1_459(.VSS(VSS),.VDD(VDD),.Y(g4753),.A(g599));
  NOT NOT1_460(.VSS(VSS),.VDD(VDD),.Y(g4754),.A(g713));
  NOT NOT1_461(.VSS(VSS),.VDD(VDD),.Y(g4757),.A(g718));
  NOT NOT1_462(.VSS(VSS),.VDD(VDD),.Y(g4760),.A(g720));
  NOT NOT1_463(.VSS(VSS),.VDD(VDD),.Y(g4763),.A(g731));
  NOT NOT1_464(.VSS(VSS),.VDD(VDD),.Y(g4766),.A(g736));
  NOT NOT1_465(.VSS(VSS),.VDD(VDD),.Y(g4769),.A(g1048));
  NOT NOT1_466(.VSS(VSS),.VDD(VDD),.Y(g4772),.A(g1060));
  NOT NOT1_467(.VSS(VSS),.VDD(VDD),.Y(g4775),.A(g1085));
  NOT NOT1_468(.VSS(VSS),.VDD(VDD),.Y(g4778),.A(g1131));
  NOT NOT1_469(.VSS(VSS),.VDD(VDD),.Y(g4779),.A(g1211));
  NOT NOT1_470(.VSS(VSS),.VDD(VDD),.Y(g4780),.A(g1263));
  NOT NOT1_471(.VSS(VSS),.VDD(VDD),.Y(g4783),.A(g1265));
  NOT NOT1_472(.VSS(VSS),.VDD(VDD),.Y(g4786),.A(g1276));
  NOT NOT1_473(.VSS(VSS),.VDD(VDD),.Y(g4787),.A(g1282));
  NOT NOT1_474(.VSS(VSS),.VDD(VDD),.Y(g4788),.A(g1396));
  NOT NOT1_475(.VSS(VSS),.VDD(VDD),.Y(g4791),.A(g1401));
  NOT NOT1_476(.VSS(VSS),.VDD(VDD),.Y(g4794),.A(g1403));
  NOT NOT1_477(.VSS(VSS),.VDD(VDD),.Y(g4797),.A(g1414));
  NOT NOT1_478(.VSS(VSS),.VDD(VDD),.Y(g4800),.A(g1419));
  NOT NOT1_479(.VSS(VSS),.VDD(VDD),.Y(g4803),.A(g1421));
  NOT NOT1_480(.VSS(VSS),.VDD(VDD),.Y(g4806),.A(g1514));
  NOT NOT1_481(.VSS(VSS),.VDD(VDD),.Y(g4809),.A(g1690));
  NOT NOT1_482(.VSS(VSS),.VDD(VDD),.Y(g4818),.A(g1727));
  NOT NOT1_483(.VSS(VSS),.VDD(VDD),.Y(g4821),.A(g1739));
  NOT NOT1_484(.VSS(VSS),.VDD(VDD),.Y(g4824),.A(g1765));
  NOT NOT1_485(.VSS(VSS),.VDD(VDD),.Y(g4827),.A(g1816));
  NOT NOT1_486(.VSS(VSS),.VDD(VDD),.Y(g4828),.A(g1822));
  NOT NOT1_487(.VSS(VSS),.VDD(VDD),.Y(g4829),.A(g1956));
  NOT NOT1_488(.VSS(VSS),.VDD(VDD),.Y(g4832),.A(g1967));
  NOT NOT1_489(.VSS(VSS),.VDD(VDD),.Y(g4833),.A(g2087));
  NOT NOT1_490(.VSS(VSS),.VDD(VDD),.Y(g4836),.A(g2092));
  NOT NOT1_491(.VSS(VSS),.VDD(VDD),.Y(g4839),.A(g2094));
  NOT NOT1_492(.VSS(VSS),.VDD(VDD),.Y(g4842),.A(g2110));
  NOT NOT1_493(.VSS(VSS),.VDD(VDD),.Y(g4845),.A(g2112));
  NOT NOT1_494(.VSS(VSS),.VDD(VDD),.Y(g4848),.A(g2257));
  NOT NOT1_495(.VSS(VSS),.VDD(VDD),.Y(g4851),.A(g2205));
  NOT NOT1_496(.VSS(VSS),.VDD(VDD),.Y(g4854),.A(g2210));
  NOT NOT1_497(.VSS(VSS),.VDD(VDD),.Y(g4857),.A(g2238));
  NOT NOT1_498(.VSS(VSS),.VDD(VDD),.Y(I13652),.A(g2170));
  NOT NOT1_499(.VSS(VSS),.VDD(VDD),.Y(g4860),.A(I13652));
  NOT NOT1_500(.VSS(VSS),.VDD(VDD),.Y(I13655),.A(g2175));
  NOT NOT1_501(.VSS(VSS),.VDD(VDD),.Y(g4861),.A(I13655));
  NOT NOT1_502(.VSS(VSS),.VDD(VDD),.Y(g4862),.A(g2418));
  NOT NOT1_503(.VSS(VSS),.VDD(VDD),.Y(g4865),.A(g2444));
  NOT NOT1_504(.VSS(VSS),.VDD(VDD),.Y(g4868),.A(g2507));
  NOT NOT1_505(.VSS(VSS),.VDD(VDD),.Y(g4869),.A(g2513));
  NOT NOT1_506(.VSS(VSS),.VDD(VDD),.Y(g4870),.A(g2778));
  NOT NOT1_507(.VSS(VSS),.VDD(VDD),.Y(g4873),.A(g2783));
  NOT NOT1_508(.VSS(VSS),.VDD(VDD),.Y(g4876),.A(g2785));
  NOT NOT1_509(.VSS(VSS),.VDD(VDD),.Y(g4879),.A(g2803));
  NOT NOT1_510(.VSS(VSS),.VDD(VDD),.Y(g4882),.A(g391));
  NOT NOT1_511(.VSS(VSS),.VDD(VDD),.Y(g4885),.A(g448));
  NOT NOT1_512(.VSS(VSS),.VDD(VDD),.Y(g4888),.A(g578));
  NOT NOT1_513(.VSS(VSS),.VDD(VDD),.Y(g4891),.A(g583));
  NOT NOT1_514(.VSS(VSS),.VDD(VDD),.Y(g4894),.A(g585));
  NOT NOT1_515(.VSS(VSS),.VDD(VDD),.Y(g4897),.A(g602));
  NOT NOT1_516(.VSS(VSS),.VDD(VDD),.Y(g4898),.A(g605));
  NOT NOT1_517(.VSS(VSS),.VDD(VDD),.Y(g4899),.A(g716));
  NOT NOT1_518(.VSS(VSS),.VDD(VDD),.Y(g4902),.A(g721));
  NOT NOT1_519(.VSS(VSS),.VDD(VDD),.Y(g4905),.A(g723));
  NOT NOT1_520(.VSS(VSS),.VDD(VDD),.Y(g4908),.A(g734));
  NOT NOT1_521(.VSS(VSS),.VDD(VDD),.Y(I13677),.A(g809));
  NOT NOT1_522(.VSS(VSS),.VDD(VDD),.Y(g4911),.A(I13677));
  NOT NOT1_523(.VSS(VSS),.VDD(VDD),.Y(I13680),.A(g813));
  NOT NOT1_524(.VSS(VSS),.VDD(VDD),.Y(g4912),.A(I13680));
  NOT NOT1_525(.VSS(VSS),.VDD(VDD),.Y(g4913),.A(g1063));
  NOT NOT1_526(.VSS(VSS),.VDD(VDD),.Y(g4916),.A(g1075));
  NOT NOT1_527(.VSS(VSS),.VDD(VDD),.Y(g4919),.A(g1261));
  NOT NOT1_528(.VSS(VSS),.VDD(VDD),.Y(g4922),.A(g1266));
  NOT NOT1_529(.VSS(VSS),.VDD(VDD),.Y(g4925),.A(g1268));
  NOT NOT1_530(.VSS(VSS),.VDD(VDD),.Y(g4928),.A(g1279));
  NOT NOT1_531(.VSS(VSS),.VDD(VDD),.Y(g4929),.A(g1285));
  NOT NOT1_532(.VSS(VSS),.VDD(VDD),.Y(g4930),.A(g1399));
  NOT NOT1_533(.VSS(VSS),.VDD(VDD),.Y(g4933),.A(g1404));
  NOT NOT1_534(.VSS(VSS),.VDD(VDD),.Y(g4936),.A(g1406));
  NOT NOT1_535(.VSS(VSS),.VDD(VDD),.Y(g4939),.A(g1417));
  NOT NOT1_536(.VSS(VSS),.VDD(VDD),.Y(g4942),.A(g1422));
  NOT NOT1_537(.VSS(VSS),.VDD(VDD),.Y(g4945),.A(g1742));
  NOT NOT1_538(.VSS(VSS),.VDD(VDD),.Y(g4948),.A(g1754));
  NOT NOT1_539(.VSS(VSS),.VDD(VDD),.Y(g4951),.A(g1779));
  NOT NOT1_540(.VSS(VSS),.VDD(VDD),.Y(g4954),.A(g1825));
  NOT NOT1_541(.VSS(VSS),.VDD(VDD),.Y(g4955),.A(g1905));
  NOT NOT1_542(.VSS(VSS),.VDD(VDD),.Y(g4956),.A(g1957));
  NOT NOT1_543(.VSS(VSS),.VDD(VDD),.Y(g4959),.A(g1959));
  NOT NOT1_544(.VSS(VSS),.VDD(VDD),.Y(g4962),.A(g1970));
  NOT NOT1_545(.VSS(VSS),.VDD(VDD),.Y(g4963),.A(g1976));
  NOT NOT1_546(.VSS(VSS),.VDD(VDD),.Y(g4964),.A(g2090));
  NOT NOT1_547(.VSS(VSS),.VDD(VDD),.Y(g4967),.A(g2095));
  NOT NOT1_548(.VSS(VSS),.VDD(VDD),.Y(g4970),.A(g2097));
  NOT NOT1_549(.VSS(VSS),.VDD(VDD),.Y(g4973),.A(g2108));
  NOT NOT1_550(.VSS(VSS),.VDD(VDD),.Y(g4976),.A(g2113));
  NOT NOT1_551(.VSS(VSS),.VDD(VDD),.Y(g4979),.A(g2115));
  NOT NOT1_552(.VSS(VSS),.VDD(VDD),.Y(g4982),.A(g2208));
  NOT NOT1_553(.VSS(VSS),.VDD(VDD),.Y(g4985),.A(g2384));
  NOT NOT1_554(.VSS(VSS),.VDD(VDD),.Y(g4994),.A(g2421));
  NOT NOT1_555(.VSS(VSS),.VDD(VDD),.Y(g4997),.A(g2433));
  NOT NOT1_556(.VSS(VSS),.VDD(VDD),.Y(g5000),.A(g2459));
  NOT NOT1_557(.VSS(VSS),.VDD(VDD),.Y(g5003),.A(g2510));
  NOT NOT1_558(.VSS(VSS),.VDD(VDD),.Y(g5004),.A(g2516));
  NOT NOT1_559(.VSS(VSS),.VDD(VDD),.Y(g5005),.A(g2650));
  NOT NOT1_560(.VSS(VSS),.VDD(VDD),.Y(g5008),.A(g2661));
  NOT NOT1_561(.VSS(VSS),.VDD(VDD),.Y(g5009),.A(g2781));
  NOT NOT1_562(.VSS(VSS),.VDD(VDD),.Y(g5012),.A(g2786));
  NOT NOT1_563(.VSS(VSS),.VDD(VDD),.Y(g5015),.A(g2788));
  NOT NOT1_564(.VSS(VSS),.VDD(VDD),.Y(g5018),.A(g2804));
  NOT NOT1_565(.VSS(VSS),.VDD(VDD),.Y(g5021),.A(g2806));
  NOT NOT1_566(.VSS(VSS),.VDD(VDD),.Y(g5024),.A(g449));
  NOT NOT1_567(.VSS(VSS),.VDD(VDD),.Y(g5027),.A(g581));
  NOT NOT1_568(.VSS(VSS),.VDD(VDD),.Y(g5030),.A(g586));
  NOT NOT1_569(.VSS(VSS),.VDD(VDD),.Y(g5033),.A(g608));
  NOT NOT1_570(.VSS(VSS),.VDD(VDD),.Y(g5034),.A(g614));
  NOT NOT1_571(.VSS(VSS),.VDD(VDD),.Y(g5035),.A(g719));
  NOT NOT1_572(.VSS(VSS),.VDD(VDD),.Y(g5038),.A(g724));
  NOT NOT1_573(.VSS(VSS),.VDD(VDD),.Y(g5041),.A(g1078));
  NOT NOT1_574(.VSS(VSS),.VDD(VDD),.Y(g5044),.A(g1135));
  NOT NOT1_575(.VSS(VSS),.VDD(VDD),.Y(g5047),.A(g1264));
  NOT NOT1_576(.VSS(VSS),.VDD(VDD),.Y(g5050),.A(g1269));
  NOT NOT1_577(.VSS(VSS),.VDD(VDD),.Y(g5053),.A(g1271));
  NOT NOT1_578(.VSS(VSS),.VDD(VDD),.Y(g5056),.A(g1288));
  NOT NOT1_579(.VSS(VSS),.VDD(VDD),.Y(g5057),.A(g1291));
  NOT NOT1_580(.VSS(VSS),.VDD(VDD),.Y(g5058),.A(g1402));
  NOT NOT1_581(.VSS(VSS),.VDD(VDD),.Y(g5061),.A(g1407));
  NOT NOT1_582(.VSS(VSS),.VDD(VDD),.Y(g5064),.A(g1409));
  NOT NOT1_583(.VSS(VSS),.VDD(VDD),.Y(g5067),.A(g1420));
  NOT NOT1_584(.VSS(VSS),.VDD(VDD),.Y(I13742),.A(g1501));
  NOT NOT1_585(.VSS(VSS),.VDD(VDD),.Y(g5070),.A(I13742));
  NOT NOT1_586(.VSS(VSS),.VDD(VDD),.Y(I13745),.A(g1506));
  NOT NOT1_587(.VSS(VSS),.VDD(VDD),.Y(g5071),.A(I13745));
  NOT NOT1_588(.VSS(VSS),.VDD(VDD),.Y(g5072),.A(g1757));
  NOT NOT1_589(.VSS(VSS),.VDD(VDD),.Y(g5075),.A(g1769));
  NOT NOT1_590(.VSS(VSS),.VDD(VDD),.Y(g5078),.A(g1955));
  NOT NOT1_591(.VSS(VSS),.VDD(VDD),.Y(g5081),.A(g1960));
  NOT NOT1_592(.VSS(VSS),.VDD(VDD),.Y(g5084),.A(g1962));
  NOT NOT1_593(.VSS(VSS),.VDD(VDD),.Y(g5087),.A(g1973));
  NOT NOT1_594(.VSS(VSS),.VDD(VDD),.Y(g5088),.A(g1979));
  NOT NOT1_595(.VSS(VSS),.VDD(VDD),.Y(g5089),.A(g2093));
  NOT NOT1_596(.VSS(VSS),.VDD(VDD),.Y(g5092),.A(g2098));
  NOT NOT1_597(.VSS(VSS),.VDD(VDD),.Y(g5095),.A(g2100));
  NOT NOT1_598(.VSS(VSS),.VDD(VDD),.Y(g5098),.A(g2111));
  NOT NOT1_599(.VSS(VSS),.VDD(VDD),.Y(g5101),.A(g2116));
  NOT NOT1_600(.VSS(VSS),.VDD(VDD),.Y(g5104),.A(g2436));
  NOT NOT1_601(.VSS(VSS),.VDD(VDD),.Y(g5107),.A(g2448));
  NOT NOT1_602(.VSS(VSS),.VDD(VDD),.Y(g5110),.A(g2473));
  NOT NOT1_603(.VSS(VSS),.VDD(VDD),.Y(g5113),.A(g2519));
  NOT NOT1_604(.VSS(VSS),.VDD(VDD),.Y(g5114),.A(g2599));
  NOT NOT1_605(.VSS(VSS),.VDD(VDD),.Y(g5115),.A(g2651));
  NOT NOT1_606(.VSS(VSS),.VDD(VDD),.Y(g5118),.A(g2653));
  NOT NOT1_607(.VSS(VSS),.VDD(VDD),.Y(g5121),.A(g2664));
  NOT NOT1_608(.VSS(VSS),.VDD(VDD),.Y(g5122),.A(g2670));
  NOT NOT1_609(.VSS(VSS),.VDD(VDD),.Y(g5123),.A(g2784));
  NOT NOT1_610(.VSS(VSS),.VDD(VDD),.Y(g5126),.A(g2789));
  NOT NOT1_611(.VSS(VSS),.VDD(VDD),.Y(g5129),.A(g2791));
  NOT NOT1_612(.VSS(VSS),.VDD(VDD),.Y(g5132),.A(g2802));
  NOT NOT1_613(.VSS(VSS),.VDD(VDD),.Y(g5135),.A(g2807));
  NOT NOT1_614(.VSS(VSS),.VDD(VDD),.Y(g5138),.A(g2809));
  NOT NOT1_615(.VSS(VSS),.VDD(VDD),.Y(I13775),.A(g109));
  NOT NOT1_616(.VSS(VSS),.VDD(VDD),.Y(g5141),.A(I13775));
  NOT NOT1_617(.VSS(VSS),.VDD(VDD),.Y(g5142),.A(g447));
  NOT NOT1_618(.VSS(VSS),.VDD(VDD),.Y(g5145),.A(g584));
  NOT NOT1_619(.VSS(VSS),.VDD(VDD),.Y(g5148),.A(g611));
  NOT NOT1_620(.VSS(VSS),.VDD(VDD),.Y(g5149),.A(g617));
  NOT NOT1_621(.VSS(VSS),.VDD(VDD),.Y(g5150),.A(g722));
  NOT NOT1_622(.VSS(VSS),.VDD(VDD),.Y(g5153),.A(g1136));
  NOT NOT1_623(.VSS(VSS),.VDD(VDD),.Y(g5156),.A(g1267));
  NOT NOT1_624(.VSS(VSS),.VDD(VDD),.Y(g5159),.A(g1272));
  NOT NOT1_625(.VSS(VSS),.VDD(VDD),.Y(g5162),.A(g1294));
  NOT NOT1_626(.VSS(VSS),.VDD(VDD),.Y(g5163),.A(g1300));
  NOT NOT1_627(.VSS(VSS),.VDD(VDD),.Y(g5164),.A(g1405));
  NOT NOT1_628(.VSS(VSS),.VDD(VDD),.Y(g5167),.A(g1410));
  NOT NOT1_629(.VSS(VSS),.VDD(VDD),.Y(g5170),.A(g1772));
  NOT NOT1_630(.VSS(VSS),.VDD(VDD),.Y(g5173),.A(g1829));
  NOT NOT1_631(.VSS(VSS),.VDD(VDD),.Y(g5176),.A(g1958));
  NOT NOT1_632(.VSS(VSS),.VDD(VDD),.Y(g5179),.A(g1963));
  NOT NOT1_633(.VSS(VSS),.VDD(VDD),.Y(g5182),.A(g1965));
  NOT NOT1_634(.VSS(VSS),.VDD(VDD),.Y(g5185),.A(g1982));
  NOT NOT1_635(.VSS(VSS),.VDD(VDD),.Y(g5186),.A(g1985));
  NOT NOT1_636(.VSS(VSS),.VDD(VDD),.Y(g5187),.A(g2096));
  NOT NOT1_637(.VSS(VSS),.VDD(VDD),.Y(g5190),.A(g2101));
  NOT NOT1_638(.VSS(VSS),.VDD(VDD),.Y(g5193),.A(g2103));
  NOT NOT1_639(.VSS(VSS),.VDD(VDD),.Y(g5196),.A(g2114));
  NOT NOT1_640(.VSS(VSS),.VDD(VDD),.Y(I13801),.A(g2195));
  NOT NOT1_641(.VSS(VSS),.VDD(VDD),.Y(g5199),.A(I13801));
  NOT NOT1_642(.VSS(VSS),.VDD(VDD),.Y(I13804),.A(g2200));
  NOT NOT1_643(.VSS(VSS),.VDD(VDD),.Y(g5200),.A(I13804));
  NOT NOT1_644(.VSS(VSS),.VDD(VDD),.Y(g5201),.A(g2451));
  NOT NOT1_645(.VSS(VSS),.VDD(VDD),.Y(g5204),.A(g2463));
  NOT NOT1_646(.VSS(VSS),.VDD(VDD),.Y(g5207),.A(g2649));
  NOT NOT1_647(.VSS(VSS),.VDD(VDD),.Y(g5210),.A(g2654));
  NOT NOT1_648(.VSS(VSS),.VDD(VDD),.Y(g5213),.A(g2656));
  NOT NOT1_649(.VSS(VSS),.VDD(VDD),.Y(g5216),.A(g2667));
  NOT NOT1_650(.VSS(VSS),.VDD(VDD),.Y(g5217),.A(g2673));
  NOT NOT1_651(.VSS(VSS),.VDD(VDD),.Y(g5218),.A(g2787));
  NOT NOT1_652(.VSS(VSS),.VDD(VDD),.Y(g5221),.A(g2792));
  NOT NOT1_653(.VSS(VSS),.VDD(VDD),.Y(g5224),.A(g2794));
  NOT NOT1_654(.VSS(VSS),.VDD(VDD),.Y(g5227),.A(g2805));
  NOT NOT1_655(.VSS(VSS),.VDD(VDD),.Y(g5230),.A(g2810));
  NOT NOT1_656(.VSS(VSS),.VDD(VDD),.Y(g5233),.A(g620));
  NOT NOT1_657(.VSS(VSS),.VDD(VDD),.Y(I13820),.A(g797));
  NOT NOT1_658(.VSS(VSS),.VDD(VDD),.Y(g5234),.A(I13820));
  NOT NOT1_659(.VSS(VSS),.VDD(VDD),.Y(g5235),.A(g1134));
  NOT NOT1_660(.VSS(VSS),.VDD(VDD),.Y(g5238),.A(g1270));
  NOT NOT1_661(.VSS(VSS),.VDD(VDD),.Y(g5241),.A(g1297));
  NOT NOT1_662(.VSS(VSS),.VDD(VDD),.Y(g5242),.A(g1303));
  NOT NOT1_663(.VSS(VSS),.VDD(VDD),.Y(g5243),.A(g1408));
  NOT NOT1_664(.VSS(VSS),.VDD(VDD),.Y(g5246),.A(g1830));
  NOT NOT1_665(.VSS(VSS),.VDD(VDD),.Y(g5249),.A(g1961));
  NOT NOT1_666(.VSS(VSS),.VDD(VDD),.Y(g5252),.A(g1966));
  NOT NOT1_667(.VSS(VSS),.VDD(VDD),.Y(g5255),.A(g1988));
  NOT NOT1_668(.VSS(VSS),.VDD(VDD),.Y(g5256),.A(g1994));
  NOT NOT1_669(.VSS(VSS),.VDD(VDD),.Y(g5257),.A(g2099));
  NOT NOT1_670(.VSS(VSS),.VDD(VDD),.Y(g5260),.A(g2104));
  NOT NOT1_671(.VSS(VSS),.VDD(VDD),.Y(g5263),.A(g2466));
  NOT NOT1_672(.VSS(VSS),.VDD(VDD),.Y(g5266),.A(g2523));
  NOT NOT1_673(.VSS(VSS),.VDD(VDD),.Y(g5269),.A(g2652));
  NOT NOT1_674(.VSS(VSS),.VDD(VDD),.Y(g5272),.A(g2657));
  NOT NOT1_675(.VSS(VSS),.VDD(VDD),.Y(g5275),.A(g2659));
  NOT NOT1_676(.VSS(VSS),.VDD(VDD),.Y(g5278),.A(g2676));
  NOT NOT1_677(.VSS(VSS),.VDD(VDD),.Y(g5279),.A(g2679));
  NOT NOT1_678(.VSS(VSS),.VDD(VDD),.Y(g5280),.A(g2790));
  NOT NOT1_679(.VSS(VSS),.VDD(VDD),.Y(g5283),.A(g2795));
  NOT NOT1_680(.VSS(VSS),.VDD(VDD),.Y(g5286),.A(g2797));
  NOT NOT1_681(.VSS(VSS),.VDD(VDD),.Y(g5289),.A(g2808));
  NOT NOT1_682(.VSS(VSS),.VDD(VDD),.Y(g5292),.A(g2857));
  NOT NOT1_683(.VSS(VSS),.VDD(VDD),.Y(g5293),.A(g738));
  NOT NOT1_684(.VSS(VSS),.VDD(VDD),.Y(g5296),.A(g1306));
  NOT NOT1_685(.VSS(VSS),.VDD(VDD),.Y(I13849),.A(g1486));
  NOT NOT1_686(.VSS(VSS),.VDD(VDD),.Y(g5297),.A(I13849));
  NOT NOT1_687(.VSS(VSS),.VDD(VDD),.Y(g5298),.A(g1828));
  NOT NOT1_688(.VSS(VSS),.VDD(VDD),.Y(g5301),.A(g1964));
  NOT NOT1_689(.VSS(VSS),.VDD(VDD),.Y(g5304),.A(g1991));
  NOT NOT1_690(.VSS(VSS),.VDD(VDD),.Y(g5305),.A(g1997));
  NOT NOT1_691(.VSS(VSS),.VDD(VDD),.Y(g5306),.A(g2102));
  NOT NOT1_692(.VSS(VSS),.VDD(VDD),.Y(g5309),.A(g2524));
  NOT NOT1_693(.VSS(VSS),.VDD(VDD),.Y(g5312),.A(g2655));
  NOT NOT1_694(.VSS(VSS),.VDD(VDD),.Y(g5315),.A(g2660));
  NOT NOT1_695(.VSS(VSS),.VDD(VDD),.Y(g5318),.A(g2682));
  NOT NOT1_696(.VSS(VSS),.VDD(VDD),.Y(g5319),.A(g2688));
  NOT NOT1_697(.VSS(VSS),.VDD(VDD),.Y(g5320),.A(g2793));
  NOT NOT1_698(.VSS(VSS),.VDD(VDD),.Y(g5323),.A(g2798));
  NOT NOT1_699(.VSS(VSS),.VDD(VDD),.Y(g5326),.A(g2873));
  NOT NOT1_700(.VSS(VSS),.VDD(VDD),.Y(g5327),.A(g739));
  NOT NOT1_701(.VSS(VSS),.VDD(VDD),.Y(g5330),.A(g1424));
  NOT NOT1_702(.VSS(VSS),.VDD(VDD),.Y(g5333),.A(g2000));
  NOT NOT1_703(.VSS(VSS),.VDD(VDD),.Y(I13868),.A(g2180));
  NOT NOT1_704(.VSS(VSS),.VDD(VDD),.Y(g5334),.A(I13868));
  NOT NOT1_705(.VSS(VSS),.VDD(VDD),.Y(g5335),.A(g2522));
  NOT NOT1_706(.VSS(VSS),.VDD(VDD),.Y(g5338),.A(g2658));
  NOT NOT1_707(.VSS(VSS),.VDD(VDD),.Y(g5341),.A(g2685));
  NOT NOT1_708(.VSS(VSS),.VDD(VDD),.Y(g5342),.A(g2691));
  NOT NOT1_709(.VSS(VSS),.VDD(VDD),.Y(g5343),.A(g2796));
  NOT NOT1_710(.VSS(VSS),.VDD(VDD),.Y(g5346),.A(g3106));
  NOT NOT1_711(.VSS(VSS),.VDD(VDD),.Y(g5349),.A(g2877));
  NOT NOT1_712(.VSS(VSS),.VDD(VDD),.Y(g5352),.A(g737));
  NOT NOT1_713(.VSS(VSS),.VDD(VDD),.Y(g5355),.A(g1425));
  NOT NOT1_714(.VSS(VSS),.VDD(VDD),.Y(g5358),.A(g2118));
  NOT NOT1_715(.VSS(VSS),.VDD(VDD),.Y(g5361),.A(g2694));
  NOT NOT1_716(.VSS(VSS),.VDD(VDD),.Y(g5362),.A(g2817));
  NOT NOT1_717(.VSS(VSS),.VDD(VDD),.Y(g5363),.A(g3107));
  NOT NOT1_718(.VSS(VSS),.VDD(VDD),.Y(g5366),.A(g2878));
  NOT NOT1_719(.VSS(VSS),.VDD(VDD),.Y(g5369),.A(g1423));
  NOT NOT1_720(.VSS(VSS),.VDD(VDD),.Y(g5372),.A(g2119));
  NOT NOT1_721(.VSS(VSS),.VDD(VDD),.Y(g5375),.A(g2812));
  NOT NOT1_722(.VSS(VSS),.VDD(VDD),.Y(g5378),.A(g2933));
  NOT NOT1_723(.VSS(VSS),.VDD(VDD),.Y(g5379),.A(g3108));
  NOT NOT1_724(.VSS(VSS),.VDD(VDD),.Y(g5382),.A(g2117));
  NOT NOT1_725(.VSS(VSS),.VDD(VDD),.Y(g5385),.A(g2813));
  NOT NOT1_726(.VSS(VSS),.VDD(VDD),.Y(I13892),.A(g3040));
  NOT NOT1_727(.VSS(VSS),.VDD(VDD),.Y(g5388),.A(I13892));
  NOT NOT1_728(.VSS(VSS),.VDD(VDD),.Y(g5389),.A(g3040));
  NOT NOT1_729(.VSS(VSS),.VDD(VDD),.Y(I13896),.A(g343));
  NOT NOT1_730(.VSS(VSS),.VDD(VDD),.Y(g5390),.A(I13896));
  NOT NOT1_731(.VSS(VSS),.VDD(VDD),.Y(g5391),.A(g2811));
  NOT NOT1_732(.VSS(VSS),.VDD(VDD),.Y(g5394),.A(g3054));
  NOT NOT1_733(.VSS(VSS),.VDD(VDD),.Y(I13901),.A(g346));
  NOT NOT1_734(.VSS(VSS),.VDD(VDD),.Y(g5395),.A(I13901));
  NOT NOT1_735(.VSS(VSS),.VDD(VDD),.Y(I13904),.A(g358));
  NOT NOT1_736(.VSS(VSS),.VDD(VDD),.Y(g5396),.A(I13904));
  NOT NOT1_737(.VSS(VSS),.VDD(VDD),.Y(I13907),.A(g1030));
  NOT NOT1_738(.VSS(VSS),.VDD(VDD),.Y(g5397),.A(I13907));
  NOT NOT1_739(.VSS(VSS),.VDD(VDD),.Y(I13910),.A(g361));
  NOT NOT1_740(.VSS(VSS),.VDD(VDD),.Y(g5398),.A(I13910));
  NOT NOT1_741(.VSS(VSS),.VDD(VDD),.Y(I13913),.A(g373));
  NOT NOT1_742(.VSS(VSS),.VDD(VDD),.Y(g5399),.A(I13913));
  NOT NOT1_743(.VSS(VSS),.VDD(VDD),.Y(I13916),.A(g1033));
  NOT NOT1_744(.VSS(VSS),.VDD(VDD),.Y(g5400),.A(I13916));
  NOT NOT1_745(.VSS(VSS),.VDD(VDD),.Y(I13919),.A(g1045));
  NOT NOT1_746(.VSS(VSS),.VDD(VDD),.Y(g5401),.A(I13919));
  NOT NOT1_747(.VSS(VSS),.VDD(VDD),.Y(I13922),.A(g1724));
  NOT NOT1_748(.VSS(VSS),.VDD(VDD),.Y(g5402),.A(I13922));
  NOT NOT1_749(.VSS(VSS),.VDD(VDD),.Y(I13925),.A(g376));
  NOT NOT1_750(.VSS(VSS),.VDD(VDD),.Y(g5403),.A(I13925));
  NOT NOT1_751(.VSS(VSS),.VDD(VDD),.Y(I13928),.A(g388));
  NOT NOT1_752(.VSS(VSS),.VDD(VDD),.Y(g5404),.A(I13928));
  NOT NOT1_753(.VSS(VSS),.VDD(VDD),.Y(I13931),.A(g1048));
  NOT NOT1_754(.VSS(VSS),.VDD(VDD),.Y(g5405),.A(I13931));
  NOT NOT1_755(.VSS(VSS),.VDD(VDD),.Y(I13934),.A(g1060));
  NOT NOT1_756(.VSS(VSS),.VDD(VDD),.Y(g5406),.A(I13934));
  NOT NOT1_757(.VSS(VSS),.VDD(VDD),.Y(I13937),.A(g1727));
  NOT NOT1_758(.VSS(VSS),.VDD(VDD),.Y(g5407),.A(I13937));
  NOT NOT1_759(.VSS(VSS),.VDD(VDD),.Y(I13940),.A(g1739));
  NOT NOT1_760(.VSS(VSS),.VDD(VDD),.Y(g5408),.A(I13940));
  NOT NOT1_761(.VSS(VSS),.VDD(VDD),.Y(I13943),.A(g2418));
  NOT NOT1_762(.VSS(VSS),.VDD(VDD),.Y(g5409),.A(I13943));
  NOT NOT1_763(.VSS(VSS),.VDD(VDD),.Y(g5410),.A(g3079));
  NOT NOT1_764(.VSS(VSS),.VDD(VDD),.Y(I13947),.A(g391));
  NOT NOT1_765(.VSS(VSS),.VDD(VDD),.Y(g5411),.A(I13947));
  NOT NOT1_766(.VSS(VSS),.VDD(VDD),.Y(I13950),.A(g1063));
  NOT NOT1_767(.VSS(VSS),.VDD(VDD),.Y(g5412),.A(I13950));
  NOT NOT1_768(.VSS(VSS),.VDD(VDD),.Y(I13953),.A(g1075));
  NOT NOT1_769(.VSS(VSS),.VDD(VDD),.Y(g5413),.A(I13953));
  NOT NOT1_770(.VSS(VSS),.VDD(VDD),.Y(I13956),.A(g1742));
  NOT NOT1_771(.VSS(VSS),.VDD(VDD),.Y(g5414),.A(I13956));
  NOT NOT1_772(.VSS(VSS),.VDD(VDD),.Y(I13959),.A(g1754));
  NOT NOT1_773(.VSS(VSS),.VDD(VDD),.Y(g5415),.A(I13959));
  NOT NOT1_774(.VSS(VSS),.VDD(VDD),.Y(I13962),.A(g2421));
  NOT NOT1_775(.VSS(VSS),.VDD(VDD),.Y(g5416),.A(I13962));
  NOT NOT1_776(.VSS(VSS),.VDD(VDD),.Y(I13965),.A(g2433));
  NOT NOT1_777(.VSS(VSS),.VDD(VDD),.Y(g5417),.A(I13965));
  NOT NOT1_778(.VSS(VSS),.VDD(VDD),.Y(I13968),.A(g1078));
  NOT NOT1_779(.VSS(VSS),.VDD(VDD),.Y(g5418),.A(I13968));
  NOT NOT1_780(.VSS(VSS),.VDD(VDD),.Y(I13971),.A(g1757));
  NOT NOT1_781(.VSS(VSS),.VDD(VDD),.Y(g5419),.A(I13971));
  NOT NOT1_782(.VSS(VSS),.VDD(VDD),.Y(I13974),.A(g1769));
  NOT NOT1_783(.VSS(VSS),.VDD(VDD),.Y(g5420),.A(I13974));
  NOT NOT1_784(.VSS(VSS),.VDD(VDD),.Y(I13977),.A(g2436));
  NOT NOT1_785(.VSS(VSS),.VDD(VDD),.Y(g5421),.A(I13977));
  NOT NOT1_786(.VSS(VSS),.VDD(VDD),.Y(I13980),.A(g2448));
  NOT NOT1_787(.VSS(VSS),.VDD(VDD),.Y(g5422),.A(I13980));
  NOT NOT1_788(.VSS(VSS),.VDD(VDD),.Y(g5423),.A(g2879));
  NOT NOT1_789(.VSS(VSS),.VDD(VDD),.Y(I13984),.A(g1772));
  NOT NOT1_790(.VSS(VSS),.VDD(VDD),.Y(g5424),.A(I13984));
  NOT NOT1_791(.VSS(VSS),.VDD(VDD),.Y(I13987),.A(g2451));
  NOT NOT1_792(.VSS(VSS),.VDD(VDD),.Y(g5425),.A(I13987));
  NOT NOT1_793(.VSS(VSS),.VDD(VDD),.Y(I13990),.A(g2463));
  NOT NOT1_794(.VSS(VSS),.VDD(VDD),.Y(g5426),.A(I13990));
  NOT NOT1_795(.VSS(VSS),.VDD(VDD),.Y(I13993),.A(g2466));
  NOT NOT1_796(.VSS(VSS),.VDD(VDD),.Y(g5427),.A(I13993));
  NOT NOT1_797(.VSS(VSS),.VDD(VDD),.Y(g5428),.A(g3210));
  NOT NOT1_798(.VSS(VSS),.VDD(VDD),.Y(g5431),.A(g3211));
  NOT NOT1_799(.VSS(VSS),.VDD(VDD),.Y(g5434),.A(g3084));
  NOT NOT1_800(.VSS(VSS),.VDD(VDD),.Y(I13999),.A(g276));
  NOT NOT1_801(.VSS(VSS),.VDD(VDD),.Y(g5437),.A(I13999));
  NOT NOT1_802(.VSS(VSS),.VDD(VDD),.Y(I14002),.A(g276));
  NOT NOT1_803(.VSS(VSS),.VDD(VDD),.Y(g5438),.A(I14002));
  NOT NOT1_804(.VSS(VSS),.VDD(VDD),.Y(g5469),.A(g3085));
  NOT NOT1_805(.VSS(VSS),.VDD(VDD),.Y(I14006),.A(g963));
  NOT NOT1_806(.VSS(VSS),.VDD(VDD),.Y(g5472),.A(I14006));
  NOT NOT1_807(.VSS(VSS),.VDD(VDD),.Y(I14009),.A(g963));
  NOT NOT1_808(.VSS(VSS),.VDD(VDD),.Y(g5473),.A(I14009));
  NOT NOT1_809(.VSS(VSS),.VDD(VDD),.Y(g5504),.A(g3086));
  NOT NOT1_810(.VSS(VSS),.VDD(VDD),.Y(g5507),.A(g3155));
  NOT NOT1_811(.VSS(VSS),.VDD(VDD),.Y(I14014),.A(g499));
  NOT NOT1_812(.VSS(VSS),.VDD(VDD),.Y(g5508),.A(I14014));
  NOT NOT1_813(.VSS(VSS),.VDD(VDD),.Y(I14017),.A(g1657));
  NOT NOT1_814(.VSS(VSS),.VDD(VDD),.Y(g5511),.A(I14017));
  NOT NOT1_815(.VSS(VSS),.VDD(VDD),.Y(I14020),.A(g1657));
  NOT NOT1_816(.VSS(VSS),.VDD(VDD),.Y(g5512),.A(I14020));
  NOT NOT1_817(.VSS(VSS),.VDD(VDD),.Y(g5543),.A(g3087));
  NOT NOT1_818(.VSS(VSS),.VDD(VDD),.Y(g5546),.A(g3164));
  NOT NOT1_819(.VSS(VSS),.VDD(VDD),.Y(g5547),.A(g101));
  NOT NOT1_820(.VSS(VSS),.VDD(VDD),.Y(g5548),.A(g105));
  NOT NOT1_821(.VSS(VSS),.VDD(VDD),.Y(I14027),.A(g182));
  NOT NOT1_822(.VSS(VSS),.VDD(VDD),.Y(g5549),.A(I14027));
  NOT NOT1_823(.VSS(VSS),.VDD(VDD),.Y(I14030),.A(g182));
  NOT NOT1_824(.VSS(VSS),.VDD(VDD),.Y(g5550),.A(I14030));
  NOT NOT1_825(.VSS(VSS),.VDD(VDD),.Y(g5551),.A(g514));
  NOT NOT1_826(.VSS(VSS),.VDD(VDD),.Y(I14034),.A(g1186));
  NOT NOT1_827(.VSS(VSS),.VDD(VDD),.Y(g5552),.A(I14034));
  NOT NOT1_828(.VSS(VSS),.VDD(VDD),.Y(I14037),.A(g2351));
  NOT NOT1_829(.VSS(VSS),.VDD(VDD),.Y(g5555),.A(I14037));
  NOT NOT1_830(.VSS(VSS),.VDD(VDD),.Y(I14040),.A(g2351));
  NOT NOT1_831(.VSS(VSS),.VDD(VDD),.Y(g5556),.A(I14040));
  NOT NOT1_832(.VSS(VSS),.VDD(VDD),.Y(g5587),.A(g3091));
  NOT NOT1_833(.VSS(VSS),.VDD(VDD),.Y(g5590),.A(g3158));
  NOT NOT1_834(.VSS(VSS),.VDD(VDD),.Y(g5591),.A(g3173));
  NOT NOT1_835(.VSS(VSS),.VDD(VDD),.Y(g5592),.A(g515));
  NOT NOT1_836(.VSS(VSS),.VDD(VDD),.Y(g5593),.A(g789));
  NOT NOT1_837(.VSS(VSS),.VDD(VDD),.Y(g5594),.A(g793));
  NOT NOT1_838(.VSS(VSS),.VDD(VDD),.Y(I14049),.A(g870));
  NOT NOT1_839(.VSS(VSS),.VDD(VDD),.Y(g5595),.A(I14049));
  NOT NOT1_840(.VSS(VSS),.VDD(VDD),.Y(I14052),.A(g870));
  NOT NOT1_841(.VSS(VSS),.VDD(VDD),.Y(g5596),.A(I14052));
  NOT NOT1_842(.VSS(VSS),.VDD(VDD),.Y(g5597),.A(g1200));
  NOT NOT1_843(.VSS(VSS),.VDD(VDD),.Y(I14056),.A(g1880));
  NOT NOT1_844(.VSS(VSS),.VDD(VDD),.Y(g5598),.A(I14056));
  NOT NOT1_845(.VSS(VSS),.VDD(VDD),.Y(g5601),.A(g3092));
  NOT NOT1_846(.VSS(VSS),.VDD(VDD),.Y(g5604),.A(g3167));
  NOT NOT1_847(.VSS(VSS),.VDD(VDD),.Y(g5605),.A(g3182));
  NOT NOT1_848(.VSS(VSS),.VDD(VDD),.Y(g5606),.A(g79));
  NOT NOT1_849(.VSS(VSS),.VDD(VDD),.Y(g5609),.A(g1201));
  NOT NOT1_850(.VSS(VSS),.VDD(VDD),.Y(g5610),.A(g1476));
  NOT NOT1_851(.VSS(VSS),.VDD(VDD),.Y(g5611),.A(g1481));
  NOT NOT1_852(.VSS(VSS),.VDD(VDD),.Y(I14066),.A(g1564));
  NOT NOT1_853(.VSS(VSS),.VDD(VDD),.Y(g5612),.A(I14066));
  NOT NOT1_854(.VSS(VSS),.VDD(VDD),.Y(I14069),.A(g1564));
  NOT NOT1_855(.VSS(VSS),.VDD(VDD),.Y(g5613),.A(I14069));
  NOT NOT1_856(.VSS(VSS),.VDD(VDD),.Y(g5614),.A(g1894));
  NOT NOT1_857(.VSS(VSS),.VDD(VDD),.Y(I14073),.A(g2574));
  NOT NOT1_858(.VSS(VSS),.VDD(VDD),.Y(g5615),.A(I14073));
  NOT NOT1_859(.VSS(VSS),.VDD(VDD),.Y(g5618),.A(g3093));
  NOT NOT1_860(.VSS(VSS),.VDD(VDD),.Y(g5621),.A(g3161));
  NOT NOT1_861(.VSS(VSS),.VDD(VDD),.Y(g5622),.A(g3176));
  NOT NOT1_862(.VSS(VSS),.VDD(VDD),.Y(g5623),.A(g70));
  NOT NOT1_863(.VSS(VSS),.VDD(VDD),.Y(g5626),.A(g121));
  NOT NOT1_864(.VSS(VSS),.VDD(VDD),.Y(g5627),.A(g125));
  NOT NOT1_865(.VSS(VSS),.VDD(VDD),.Y(g5628),.A(g300));
  NOT NOT1_866(.VSS(VSS),.VDD(VDD),.Y(I14083),.A(g325));
  NOT NOT1_867(.VSS(VSS),.VDD(VDD),.Y(g5629),.A(I14083));
  NOT NOT1_868(.VSS(VSS),.VDD(VDD),.Y(g5631),.A(g767));
  NOT NOT1_869(.VSS(VSS),.VDD(VDD),.Y(g5634),.A(g1895));
  NOT NOT1_870(.VSS(VSS),.VDD(VDD),.Y(g5635),.A(g2170));
  NOT NOT1_871(.VSS(VSS),.VDD(VDD),.Y(g5636),.A(g2175));
  NOT NOT1_872(.VSS(VSS),.VDD(VDD),.Y(I14091),.A(g2258));
  NOT NOT1_873(.VSS(VSS),.VDD(VDD),.Y(g5637),.A(I14091));
  NOT NOT1_874(.VSS(VSS),.VDD(VDD),.Y(I14094),.A(g2258));
  NOT NOT1_875(.VSS(VSS),.VDD(VDD),.Y(g5638),.A(I14094));
  NOT NOT1_876(.VSS(VSS),.VDD(VDD),.Y(g5639),.A(g2588));
  NOT NOT1_877(.VSS(VSS),.VDD(VDD),.Y(g5640),.A(g3170));
  NOT NOT1_878(.VSS(VSS),.VDD(VDD),.Y(g5641),.A(g3185));
  NOT NOT1_879(.VSS(VSS),.VDD(VDD),.Y(g5642),.A(g61));
  NOT NOT1_880(.VSS(VSS),.VDD(VDD),.Y(g5645),.A(g101));
  NOT NOT1_881(.VSS(VSS),.VDD(VDD),.Y(g5646),.A(g213));
  NOT NOT1_882(.VSS(VSS),.VDD(VDD),.Y(g5647),.A(g301));
  NOT NOT1_883(.VSS(VSS),.VDD(VDD),.Y(I14104),.A(g331));
  NOT NOT1_884(.VSS(VSS),.VDD(VDD),.Y(g5648),.A(I14104));
  NOT NOT1_885(.VSS(VSS),.VDD(VDD),.Y(g5651),.A(g758));
  NOT NOT1_886(.VSS(VSS),.VDD(VDD),.Y(g5654),.A(g809));
  NOT NOT1_887(.VSS(VSS),.VDD(VDD),.Y(g5655),.A(g813));
  NOT NOT1_888(.VSS(VSS),.VDD(VDD),.Y(g5656),.A(g987));
  NOT NOT1_889(.VSS(VSS),.VDD(VDD),.Y(I14113),.A(g1012));
  NOT NOT1_890(.VSS(VSS),.VDD(VDD),.Y(g5657),.A(I14113));
  NOT NOT1_891(.VSS(VSS),.VDD(VDD),.Y(g5659),.A(g1453));
  NOT NOT1_892(.VSS(VSS),.VDD(VDD),.Y(g5662),.A(g2589));
  NOT NOT1_893(.VSS(VSS),.VDD(VDD),.Y(g5663),.A(g3179));
  NOT NOT1_894(.VSS(VSS),.VDD(VDD),.Y(g5664),.A(g65));
  NOT NOT1_895(.VSS(VSS),.VDD(VDD),.Y(g5665),.A(g105));
  NOT NOT1_896(.VSS(VSS),.VDD(VDD),.Y(g5666),.A(g216));
  NOT NOT1_897(.VSS(VSS),.VDD(VDD),.Y(g5667),.A(g222));
  NOT NOT1_898(.VSS(VSS),.VDD(VDD),.Y(g5668),.A(g299));
  NOT NOT1_899(.VSS(VSS),.VDD(VDD),.Y(g5675),.A(g302));
  NOT NOT1_900(.VSS(VSS),.VDD(VDD),.Y(g5679),.A(g506));
  NOT NOT1_901(.VSS(VSS),.VDD(VDD),.Y(g5680),.A(g749));
  NOT NOT1_902(.VSS(VSS),.VDD(VDD),.Y(g5683),.A(g789));
  NOT NOT1_903(.VSS(VSS),.VDD(VDD),.Y(g5684),.A(g900));
  NOT NOT1_904(.VSS(VSS),.VDD(VDD),.Y(g5685),.A(g988));
  NOT NOT1_905(.VSS(VSS),.VDD(VDD),.Y(I14134),.A(g1018));
  NOT NOT1_906(.VSS(VSS),.VDD(VDD),.Y(g5686),.A(I14134));
  NOT NOT1_907(.VSS(VSS),.VDD(VDD),.Y(g5689),.A(g1444));
  NOT NOT1_908(.VSS(VSS),.VDD(VDD),.Y(g5692),.A(g1501));
  NOT NOT1_909(.VSS(VSS),.VDD(VDD),.Y(g5693),.A(g1506));
  NOT NOT1_910(.VSS(VSS),.VDD(VDD),.Y(g5694),.A(g1681));
  NOT NOT1_911(.VSS(VSS),.VDD(VDD),.Y(I14143),.A(g1706));
  NOT NOT1_912(.VSS(VSS),.VDD(VDD),.Y(g5695),.A(I14143));
  NOT NOT1_913(.VSS(VSS),.VDD(VDD),.Y(g5697),.A(g2147));
  NOT NOT1_914(.VSS(VSS),.VDD(VDD),.Y(g5700),.A(g3088));
  NOT NOT1_915(.VSS(VSS),.VDD(VDD),.Y(I14149),.A(g3231));
  NOT NOT1_916(.VSS(VSS),.VDD(VDD),.Y(g5701),.A(I14149));
  NOT NOT1_917(.VSS(VSS),.VDD(VDD),.Y(g5702),.A(g56));
  NOT NOT1_918(.VSS(VSS),.VDD(VDD),.Y(g5703),.A(g109));
  NOT NOT1_919(.VSS(VSS),.VDD(VDD),.Y(g5704),.A(g219));
  NOT NOT1_920(.VSS(VSS),.VDD(VDD),.Y(g5705),.A(g225));
  NOT NOT1_921(.VSS(VSS),.VDD(VDD),.Y(g5706),.A(g231));
  NOT NOT1_922(.VSS(VSS),.VDD(VDD),.Y(g5707),.A(g109));
  NOT NOT1_923(.VSS(VSS),.VDD(VDD),.Y(g5708),.A(g303));
  NOT NOT1_924(.VSS(VSS),.VDD(VDD),.Y(g5712),.A(g305));
  NOT NOT1_925(.VSS(VSS),.VDD(VDD),.Y(I14163),.A(g113));
  NOT NOT1_926(.VSS(VSS),.VDD(VDD),.Y(g5713),.A(I14163));
  NOT NOT1_927(.VSS(VSS),.VDD(VDD),.Y(g5714),.A(g507));
  NOT NOT1_928(.VSS(VSS),.VDD(VDD),.Y(g5715),.A(g541));
  NOT NOT1_929(.VSS(VSS),.VDD(VDD),.Y(g5716),.A(g753));
  NOT NOT1_930(.VSS(VSS),.VDD(VDD),.Y(g5717),.A(g793));
  NOT NOT1_931(.VSS(VSS),.VDD(VDD),.Y(g5718),.A(g903));
  NOT NOT1_932(.VSS(VSS),.VDD(VDD),.Y(g5719),.A(g909));
  NOT NOT1_933(.VSS(VSS),.VDD(VDD),.Y(g5720),.A(g986));
  NOT NOT1_934(.VSS(VSS),.VDD(VDD),.Y(g5727),.A(g989));
  NOT NOT1_935(.VSS(VSS),.VDD(VDD),.Y(g5731),.A(g1192));
  NOT NOT1_936(.VSS(VSS),.VDD(VDD),.Y(g5732),.A(g1435));
  NOT NOT1_937(.VSS(VSS),.VDD(VDD),.Y(g5735),.A(g1476));
  NOT NOT1_938(.VSS(VSS),.VDD(VDD),.Y(g5736),.A(g1594));
  NOT NOT1_939(.VSS(VSS),.VDD(VDD),.Y(g5737),.A(g1682));
  NOT NOT1_940(.VSS(VSS),.VDD(VDD),.Y(I14182),.A(g1712));
  NOT NOT1_941(.VSS(VSS),.VDD(VDD),.Y(g5738),.A(I14182));
  NOT NOT1_942(.VSS(VSS),.VDD(VDD),.Y(g5741),.A(g2138));
  NOT NOT1_943(.VSS(VSS),.VDD(VDD),.Y(g5744),.A(g2195));
  NOT NOT1_944(.VSS(VSS),.VDD(VDD),.Y(g5745),.A(g2200));
  NOT NOT1_945(.VSS(VSS),.VDD(VDD),.Y(g5746),.A(g2375));
  NOT NOT1_946(.VSS(VSS),.VDD(VDD),.Y(I14191),.A(g2400));
  NOT NOT1_947(.VSS(VSS),.VDD(VDD),.Y(g5747),.A(I14191));
  NOT NOT1_948(.VSS(VSS),.VDD(VDD),.Y(I14195),.A(g3212));
  NOT NOT1_949(.VSS(VSS),.VDD(VDD),.Y(g5749),.A(I14195));
  NOT NOT1_950(.VSS(VSS),.VDD(VDD),.Y(g5750),.A(g92));
  NOT NOT1_951(.VSS(VSS),.VDD(VDD),.Y(g5751),.A(g52));
  NOT NOT1_952(.VSS(VSS),.VDD(VDD),.Y(g5752),.A(g113));
  NOT NOT1_953(.VSS(VSS),.VDD(VDD),.Y(g5753),.A(g228));
  NOT NOT1_954(.VSS(VSS),.VDD(VDD),.Y(g5754),.A(g234));
  NOT NOT1_955(.VSS(VSS),.VDD(VDD),.Y(g5755),.A(g240));
  NOT NOT1_956(.VSS(VSS),.VDD(VDD),.Y(g5756),.A(g304));
  NOT NOT1_957(.VSS(VSS),.VDD(VDD),.Y(g5759),.A(g508));
  NOT NOT1_958(.VSS(VSS),.VDD(VDD),.Y(g5760),.A(g744));
  NOT NOT1_959(.VSS(VSS),.VDD(VDD),.Y(g5761),.A(g797));
  NOT NOT1_960(.VSS(VSS),.VDD(VDD),.Y(g5762),.A(g906));
  NOT NOT1_961(.VSS(VSS),.VDD(VDD),.Y(g5763),.A(g912));
  NOT NOT1_962(.VSS(VSS),.VDD(VDD),.Y(g5764),.A(g918));
  NOT NOT1_963(.VSS(VSS),.VDD(VDD),.Y(g5765),.A(g797));
  NOT NOT1_964(.VSS(VSS),.VDD(VDD),.Y(g5766),.A(g990));
  NOT NOT1_965(.VSS(VSS),.VDD(VDD),.Y(g5770),.A(g992));
  NOT NOT1_966(.VSS(VSS),.VDD(VDD),.Y(I14219),.A(g801));
  NOT NOT1_967(.VSS(VSS),.VDD(VDD),.Y(g5771),.A(I14219));
  NOT NOT1_968(.VSS(VSS),.VDD(VDD),.Y(g5772),.A(g1193));
  NOT NOT1_969(.VSS(VSS),.VDD(VDD),.Y(g5773),.A(g1227));
  NOT NOT1_970(.VSS(VSS),.VDD(VDD),.Y(g5774),.A(g1439));
  NOT NOT1_971(.VSS(VSS),.VDD(VDD),.Y(g5775),.A(g1481));
  NOT NOT1_972(.VSS(VSS),.VDD(VDD),.Y(g5776),.A(g1597));
  NOT NOT1_973(.VSS(VSS),.VDD(VDD),.Y(g5777),.A(g1603));
  NOT NOT1_974(.VSS(VSS),.VDD(VDD),.Y(g5778),.A(g1680));
  NOT NOT1_975(.VSS(VSS),.VDD(VDD),.Y(g5785),.A(g1683));
  NOT NOT1_976(.VSS(VSS),.VDD(VDD),.Y(g5789),.A(g1886));
  NOT NOT1_977(.VSS(VSS),.VDD(VDD),.Y(g5790),.A(g2129));
  NOT NOT1_978(.VSS(VSS),.VDD(VDD),.Y(g5793),.A(g2170));
  NOT NOT1_979(.VSS(VSS),.VDD(VDD),.Y(g5794),.A(g2288));
  NOT NOT1_980(.VSS(VSS),.VDD(VDD),.Y(g5795),.A(g2376));
  NOT NOT1_981(.VSS(VSS),.VDD(VDD),.Y(I14238),.A(g2406));
  NOT NOT1_982(.VSS(VSS),.VDD(VDD),.Y(g5796),.A(I14238));
  NOT NOT1_983(.VSS(VSS),.VDD(VDD),.Y(I14243),.A(g3221));
  NOT NOT1_984(.VSS(VSS),.VDD(VDD),.Y(g5799),.A(I14243));
  NOT NOT1_985(.VSS(VSS),.VDD(VDD),.Y(I14246),.A(g3227));
  NOT NOT1_986(.VSS(VSS),.VDD(VDD),.Y(g5800),.A(I14246));
  NOT NOT1_987(.VSS(VSS),.VDD(VDD),.Y(I14249),.A(g3216));
  NOT NOT1_988(.VSS(VSS),.VDD(VDD),.Y(g5801),.A(I14249));
  NOT NOT1_989(.VSS(VSS),.VDD(VDD),.Y(g5802),.A(g83));
  NOT NOT1_990(.VSS(VSS),.VDD(VDD),.Y(g5803),.A(g117));
  NOT NOT1_991(.VSS(VSS),.VDD(VDD),.Y(g5804),.A(g237));
  NOT NOT1_992(.VSS(VSS),.VDD(VDD),.Y(g5805),.A(g243));
  NOT NOT1_993(.VSS(VSS),.VDD(VDD),.Y(g5806),.A(g249));
  NOT NOT1_994(.VSS(VSS),.VDD(VDD),.Y(g5808),.A(g509));
  NOT NOT1_995(.VSS(VSS),.VDD(VDD),.Y(g5809),.A(g780));
  NOT NOT1_996(.VSS(VSS),.VDD(VDD),.Y(g5810),.A(g740));
  NOT NOT1_997(.VSS(VSS),.VDD(VDD),.Y(g5811),.A(g801));
  NOT NOT1_998(.VSS(VSS),.VDD(VDD),.Y(g5812),.A(g915));
  NOT NOT1_999(.VSS(VSS),.VDD(VDD),.Y(g5813),.A(g921));
  NOT NOT1_1000(.VSS(VSS),.VDD(VDD),.Y(g5814),.A(g927));
  NOT NOT1_1001(.VSS(VSS),.VDD(VDD),.Y(g5815),.A(g991));
  NOT NOT1_1002(.VSS(VSS),.VDD(VDD),.Y(g5818),.A(g1194));
  NOT NOT1_1003(.VSS(VSS),.VDD(VDD),.Y(g5819),.A(g1430));
  NOT NOT1_1004(.VSS(VSS),.VDD(VDD),.Y(g5820),.A(g1486));
  NOT NOT1_1005(.VSS(VSS),.VDD(VDD),.Y(g5821),.A(g1600));
  NOT NOT1_1006(.VSS(VSS),.VDD(VDD),.Y(g5822),.A(g1606));
  NOT NOT1_1007(.VSS(VSS),.VDD(VDD),.Y(g5823),.A(g1612));
  NOT NOT1_1008(.VSS(VSS),.VDD(VDD),.Y(g5824),.A(g1486));
  NOT NOT1_1009(.VSS(VSS),.VDD(VDD),.Y(g5825),.A(g1684));
  NOT NOT1_1010(.VSS(VSS),.VDD(VDD),.Y(g5829),.A(g1686));
  NOT NOT1_1011(.VSS(VSS),.VDD(VDD),.Y(I14280),.A(g1491));
  NOT NOT1_1012(.VSS(VSS),.VDD(VDD),.Y(g5830),.A(I14280));
  NOT NOT1_1013(.VSS(VSS),.VDD(VDD),.Y(g5831),.A(g1887));
  NOT NOT1_1014(.VSS(VSS),.VDD(VDD),.Y(g5832),.A(g1921));
  NOT NOT1_1015(.VSS(VSS),.VDD(VDD),.Y(g5833),.A(g2133));
  NOT NOT1_1016(.VSS(VSS),.VDD(VDD),.Y(g5834),.A(g2175));
  NOT NOT1_1017(.VSS(VSS),.VDD(VDD),.Y(g5835),.A(g2291));
  NOT NOT1_1018(.VSS(VSS),.VDD(VDD),.Y(g5836),.A(g2297));
  NOT NOT1_1019(.VSS(VSS),.VDD(VDD),.Y(g5837),.A(g2374));
  NOT NOT1_1020(.VSS(VSS),.VDD(VDD),.Y(g5844),.A(g2377));
  NOT NOT1_1021(.VSS(VSS),.VDD(VDD),.Y(g5848),.A(g2580));
  NOT NOT1_1022(.VSS(VSS),.VDD(VDD),.Y(I14295),.A(g3228));
  NOT NOT1_1023(.VSS(VSS),.VDD(VDD),.Y(g5849),.A(I14295));
  NOT NOT1_1024(.VSS(VSS),.VDD(VDD),.Y(I14298),.A(g3217));
  NOT NOT1_1025(.VSS(VSS),.VDD(VDD),.Y(g5850),.A(I14298));
  NOT NOT1_1026(.VSS(VSS),.VDD(VDD),.Y(g5851),.A(g74));
  NOT NOT1_1027(.VSS(VSS),.VDD(VDD),.Y(g5852),.A(g121));
  NOT NOT1_1028(.VSS(VSS),.VDD(VDD),.Y(g5853),.A(g246));
  NOT NOT1_1029(.VSS(VSS),.VDD(VDD),.Y(g5854),.A(g252));
  NOT NOT1_1030(.VSS(VSS),.VDD(VDD),.Y(g5855),.A(g258));
  NOT NOT1_1031(.VSS(VSS),.VDD(VDD),.Y(I14306),.A(g97));
  NOT NOT1_1032(.VSS(VSS),.VDD(VDD),.Y(g5856),.A(I14306));
  NOT NOT1_1033(.VSS(VSS),.VDD(VDD),.Y(g5857),.A(g538));
  NOT NOT1_1034(.VSS(VSS),.VDD(VDD),.Y(g5858),.A(g771));
  NOT NOT1_1035(.VSS(VSS),.VDD(VDD),.Y(g5859),.A(g805));
  NOT NOT1_1036(.VSS(VSS),.VDD(VDD),.Y(g5860),.A(g924));
  NOT NOT1_1037(.VSS(VSS),.VDD(VDD),.Y(g5861),.A(g930));
  NOT NOT1_1038(.VSS(VSS),.VDD(VDD),.Y(g5862),.A(g936));
  NOT NOT1_1039(.VSS(VSS),.VDD(VDD),.Y(g5864),.A(g1195));
  NOT NOT1_1040(.VSS(VSS),.VDD(VDD),.Y(g5865),.A(g1466));
  NOT NOT1_1041(.VSS(VSS),.VDD(VDD),.Y(g5866),.A(g1426));
  NOT NOT1_1042(.VSS(VSS),.VDD(VDD),.Y(g5867),.A(g1491));
  NOT NOT1_1043(.VSS(VSS),.VDD(VDD),.Y(g5868),.A(g1609));
  NOT NOT1_1044(.VSS(VSS),.VDD(VDD),.Y(g5869),.A(g1615));
  NOT NOT1_1045(.VSS(VSS),.VDD(VDD),.Y(g5870),.A(g1621));
  NOT NOT1_1046(.VSS(VSS),.VDD(VDD),.Y(g5871),.A(g1685));
  NOT NOT1_1047(.VSS(VSS),.VDD(VDD),.Y(g5874),.A(g1888));
  NOT NOT1_1048(.VSS(VSS),.VDD(VDD),.Y(g5875),.A(g2124));
  NOT NOT1_1049(.VSS(VSS),.VDD(VDD),.Y(g5876),.A(g2180));
  NOT NOT1_1050(.VSS(VSS),.VDD(VDD),.Y(g5877),.A(g2294));
  NOT NOT1_1051(.VSS(VSS),.VDD(VDD),.Y(g5878),.A(g2300));
  NOT NOT1_1052(.VSS(VSS),.VDD(VDD),.Y(g5879),.A(g2306));
  NOT NOT1_1053(.VSS(VSS),.VDD(VDD),.Y(g5880),.A(g2180));
  NOT NOT1_1054(.VSS(VSS),.VDD(VDD),.Y(g5881),.A(g2378));
  NOT NOT1_1055(.VSS(VSS),.VDD(VDD),.Y(g5885),.A(g2380));
  NOT NOT1_1056(.VSS(VSS),.VDD(VDD),.Y(I14338),.A(g2185));
  NOT NOT1_1057(.VSS(VSS),.VDD(VDD),.Y(g5886),.A(I14338));
  NOT NOT1_1058(.VSS(VSS),.VDD(VDD),.Y(g5887),.A(g2581));
  NOT NOT1_1059(.VSS(VSS),.VDD(VDD),.Y(g5888),.A(g2615));
  NOT NOT1_1060(.VSS(VSS),.VDD(VDD),.Y(I14343),.A(g3219));
  NOT NOT1_1061(.VSS(VSS),.VDD(VDD),.Y(g5889),.A(I14343));
  NOT NOT1_1062(.VSS(VSS),.VDD(VDD),.Y(g5890),.A(g88));
  NOT NOT1_1063(.VSS(VSS),.VDD(VDD),.Y(g5893),.A(g125));
  NOT NOT1_1064(.VSS(VSS),.VDD(VDD),.Y(g5894),.A(g186));
  NOT NOT1_1065(.VSS(VSS),.VDD(VDD),.Y(g5895),.A(g255));
  NOT NOT1_1066(.VSS(VSS),.VDD(VDD),.Y(g5896),.A(g261));
  NOT NOT1_1067(.VSS(VSS),.VDD(VDD),.Y(g5897),.A(g267));
  NOT NOT1_1068(.VSS(VSS),.VDD(VDD),.Y(g5898),.A(g762));
  NOT NOT1_1069(.VSS(VSS),.VDD(VDD),.Y(g5899),.A(g809));
  NOT NOT1_1070(.VSS(VSS),.VDD(VDD),.Y(g5900),.A(g933));
  NOT NOT1_1071(.VSS(VSS),.VDD(VDD),.Y(g5901),.A(g939));
  NOT NOT1_1072(.VSS(VSS),.VDD(VDD),.Y(g5902),.A(g945));
  NOT NOT1_1073(.VSS(VSS),.VDD(VDD),.Y(I14357),.A(g785));
  NOT NOT1_1074(.VSS(VSS),.VDD(VDD),.Y(g5903),.A(I14357));
  NOT NOT1_1075(.VSS(VSS),.VDD(VDD),.Y(g5904),.A(g1224));
  NOT NOT1_1076(.VSS(VSS),.VDD(VDD),.Y(g5905),.A(g1457));
  NOT NOT1_1077(.VSS(VSS),.VDD(VDD),.Y(g5906),.A(g1496));
  NOT NOT1_1078(.VSS(VSS),.VDD(VDD),.Y(g5907),.A(g1618));
  NOT NOT1_1079(.VSS(VSS),.VDD(VDD),.Y(g5908),.A(g1624));
  NOT NOT1_1080(.VSS(VSS),.VDD(VDD),.Y(g5909),.A(g1630));
  NOT NOT1_1081(.VSS(VSS),.VDD(VDD),.Y(g5911),.A(g1889));
  NOT NOT1_1082(.VSS(VSS),.VDD(VDD),.Y(g5912),.A(g2160));
  NOT NOT1_1083(.VSS(VSS),.VDD(VDD),.Y(g5913),.A(g2120));
  NOT NOT1_1084(.VSS(VSS),.VDD(VDD),.Y(g5914),.A(g2185));
  NOT NOT1_1085(.VSS(VSS),.VDD(VDD),.Y(g5915),.A(g2303));
  NOT NOT1_1086(.VSS(VSS),.VDD(VDD),.Y(g5916),.A(g2309));
  NOT NOT1_1087(.VSS(VSS),.VDD(VDD),.Y(g5917),.A(g2315));
  NOT NOT1_1088(.VSS(VSS),.VDD(VDD),.Y(g5918),.A(g2379));
  NOT NOT1_1089(.VSS(VSS),.VDD(VDD),.Y(g5921),.A(g2582));
  NOT NOT1_1090(.VSS(VSS),.VDD(VDD),.Y(I14378),.A(g3234));
  NOT NOT1_1091(.VSS(VSS),.VDD(VDD),.Y(g5922),.A(I14378));
  NOT NOT1_1092(.VSS(VSS),.VDD(VDD),.Y(I14381),.A(g3223));
  NOT NOT1_1093(.VSS(VSS),.VDD(VDD),.Y(g5923),.A(I14381));
  NOT NOT1_1094(.VSS(VSS),.VDD(VDD),.Y(I14384),.A(g3218));
  NOT NOT1_1095(.VSS(VSS),.VDD(VDD),.Y(g5924),.A(I14384));
  NOT NOT1_1096(.VSS(VSS),.VDD(VDD),.Y(g5925),.A(g189));
  NOT NOT1_1097(.VSS(VSS),.VDD(VDD),.Y(g5926),.A(g195));
  NOT NOT1_1098(.VSS(VSS),.VDD(VDD),.Y(g5927),.A(g264));
  NOT NOT1_1099(.VSS(VSS),.VDD(VDD),.Y(g5928),.A(g270));
  NOT NOT1_1100(.VSS(VSS),.VDD(VDD),.Y(g5929),.A(g776));
  NOT NOT1_1101(.VSS(VSS),.VDD(VDD),.Y(g5932),.A(g813));
  NOT NOT1_1102(.VSS(VSS),.VDD(VDD),.Y(g5933),.A(g873));
  NOT NOT1_1103(.VSS(VSS),.VDD(VDD),.Y(g5934),.A(g942));
  NOT NOT1_1104(.VSS(VSS),.VDD(VDD),.Y(g5935),.A(g948));
  NOT NOT1_1105(.VSS(VSS),.VDD(VDD),.Y(g5936),.A(g954));
  NOT NOT1_1106(.VSS(VSS),.VDD(VDD),.Y(g5937),.A(g1448));
  NOT NOT1_1107(.VSS(VSS),.VDD(VDD),.Y(g5938),.A(g1501));
  NOT NOT1_1108(.VSS(VSS),.VDD(VDD),.Y(g5939),.A(g1627));
  NOT NOT1_1109(.VSS(VSS),.VDD(VDD),.Y(g5940),.A(g1633));
  NOT NOT1_1110(.VSS(VSS),.VDD(VDD),.Y(g5941),.A(g1639));
  NOT NOT1_1111(.VSS(VSS),.VDD(VDD),.Y(I14402),.A(g1471));
  NOT NOT1_1112(.VSS(VSS),.VDD(VDD),.Y(g5942),.A(I14402));
  NOT NOT1_1113(.VSS(VSS),.VDD(VDD),.Y(g5943),.A(g1918));
  NOT NOT1_1114(.VSS(VSS),.VDD(VDD),.Y(g5944),.A(g2151));
  NOT NOT1_1115(.VSS(VSS),.VDD(VDD),.Y(g5945),.A(g2190));
  NOT NOT1_1116(.VSS(VSS),.VDD(VDD),.Y(g5946),.A(g2312));
  NOT NOT1_1117(.VSS(VSS),.VDD(VDD),.Y(g5947),.A(g2318));
  NOT NOT1_1118(.VSS(VSS),.VDD(VDD),.Y(g5948),.A(g2324));
  NOT NOT1_1119(.VSS(VSS),.VDD(VDD),.Y(g5950),.A(g2583));
  NOT NOT1_1120(.VSS(VSS),.VDD(VDD),.Y(I14413),.A(g3233));
  NOT NOT1_1121(.VSS(VSS),.VDD(VDD),.Y(g5951),.A(I14413));
  NOT NOT1_1122(.VSS(VSS),.VDD(VDD),.Y(I14416),.A(g3222));
  NOT NOT1_1123(.VSS(VSS),.VDD(VDD),.Y(g5952),.A(I14416));
  NOT NOT1_1124(.VSS(VSS),.VDD(VDD),.Y(g5953),.A(g97));
  NOT NOT1_1125(.VSS(VSS),.VDD(VDD),.Y(g5954),.A(g192));
  NOT NOT1_1126(.VSS(VSS),.VDD(VDD),.Y(g5955),.A(g198));
  NOT NOT1_1127(.VSS(VSS),.VDD(VDD),.Y(g5956),.A(g204));
  NOT NOT1_1128(.VSS(VSS),.VDD(VDD),.Y(g5957),.A(g273));
  NOT NOT1_1129(.VSS(VSS),.VDD(VDD),.Y(I14424),.A(g117));
  NOT NOT1_1130(.VSS(VSS),.VDD(VDD),.Y(g5958),.A(I14424));
  NOT NOT1_1131(.VSS(VSS),.VDD(VDD),.Y(g5959),.A(g876));
  NOT NOT1_1132(.VSS(VSS),.VDD(VDD),.Y(g5960),.A(g882));
  NOT NOT1_1133(.VSS(VSS),.VDD(VDD),.Y(g5961),.A(g951));
  NOT NOT1_1134(.VSS(VSS),.VDD(VDD),.Y(g5962),.A(g957));
  NOT NOT1_1135(.VSS(VSS),.VDD(VDD),.Y(g5963),.A(g1462));
  NOT NOT1_1136(.VSS(VSS),.VDD(VDD),.Y(g5966),.A(g1506));
  NOT NOT1_1137(.VSS(VSS),.VDD(VDD),.Y(g5967),.A(g1567));
  NOT NOT1_1138(.VSS(VSS),.VDD(VDD),.Y(g5968),.A(g1636));
  NOT NOT1_1139(.VSS(VSS),.VDD(VDD),.Y(g5969),.A(g1642));
  NOT NOT1_1140(.VSS(VSS),.VDD(VDD),.Y(g5970),.A(g1648));
  NOT NOT1_1141(.VSS(VSS),.VDD(VDD),.Y(g5971),.A(g2142));
  NOT NOT1_1142(.VSS(VSS),.VDD(VDD),.Y(g5972),.A(g2195));
  NOT NOT1_1143(.VSS(VSS),.VDD(VDD),.Y(g5973),.A(g2321));
  NOT NOT1_1144(.VSS(VSS),.VDD(VDD),.Y(g5974),.A(g2327));
  NOT NOT1_1145(.VSS(VSS),.VDD(VDD),.Y(g5975),.A(g2333));
  NOT NOT1_1146(.VSS(VSS),.VDD(VDD),.Y(I14442),.A(g2165));
  NOT NOT1_1147(.VSS(VSS),.VDD(VDD),.Y(g5976),.A(I14442));
  NOT NOT1_1148(.VSS(VSS),.VDD(VDD),.Y(g5977),.A(g2612));
  NOT NOT1_1149(.VSS(VSS),.VDD(VDD),.Y(I14446),.A(g3230));
  NOT NOT1_1150(.VSS(VSS),.VDD(VDD),.Y(g5978),.A(I14446));
  NOT NOT1_1151(.VSS(VSS),.VDD(VDD),.Y(I14449),.A(g3224));
  NOT NOT1_1152(.VSS(VSS),.VDD(VDD),.Y(g5979),.A(I14449));
  NOT NOT1_1153(.VSS(VSS),.VDD(VDD),.Y(g5980),.A(g201));
  NOT NOT1_1154(.VSS(VSS),.VDD(VDD),.Y(g5981),.A(g207));
  NOT NOT1_1155(.VSS(VSS),.VDD(VDD),.Y(g5982),.A(g785));
  NOT NOT1_1156(.VSS(VSS),.VDD(VDD),.Y(g5983),.A(g879));
  NOT NOT1_1157(.VSS(VSS),.VDD(VDD),.Y(g5984),.A(g885));
  NOT NOT1_1158(.VSS(VSS),.VDD(VDD),.Y(g5985),.A(g891));
  NOT NOT1_1159(.VSS(VSS),.VDD(VDD),.Y(g5986),.A(g960));
  NOT NOT1_1160(.VSS(VSS),.VDD(VDD),.Y(I14459),.A(g805));
  NOT NOT1_1161(.VSS(VSS),.VDD(VDD),.Y(g5987),.A(I14459));
  NOT NOT1_1162(.VSS(VSS),.VDD(VDD),.Y(g5988),.A(g1570));
  NOT NOT1_1163(.VSS(VSS),.VDD(VDD),.Y(g5989),.A(g1576));
  NOT NOT1_1164(.VSS(VSS),.VDD(VDD),.Y(g5990),.A(g1645));
  NOT NOT1_1165(.VSS(VSS),.VDD(VDD),.Y(g5991),.A(g1651));
  NOT NOT1_1166(.VSS(VSS),.VDD(VDD),.Y(g5992),.A(g2156));
  NOT NOT1_1167(.VSS(VSS),.VDD(VDD),.Y(g5995),.A(g2200));
  NOT NOT1_1168(.VSS(VSS),.VDD(VDD),.Y(g5996),.A(g2261));
  NOT NOT1_1169(.VSS(VSS),.VDD(VDD),.Y(g5997),.A(g2330));
  NOT NOT1_1170(.VSS(VSS),.VDD(VDD),.Y(g5998),.A(g2336));
  NOT NOT1_1171(.VSS(VSS),.VDD(VDD),.Y(g5999),.A(g2342));
  NOT NOT1_1172(.VSS(VSS),.VDD(VDD),.Y(I14472),.A(g3080));
  NOT NOT1_1173(.VSS(VSS),.VDD(VDD),.Y(g6000),.A(I14472));
  NOT NOT1_1174(.VSS(VSS),.VDD(VDD),.Y(I14475),.A(g3225));
  NOT NOT1_1175(.VSS(VSS),.VDD(VDD),.Y(g6014),.A(I14475));
  NOT NOT1_1176(.VSS(VSS),.VDD(VDD),.Y(I14478),.A(g3213));
  NOT NOT1_1177(.VSS(VSS),.VDD(VDD),.Y(g6015),.A(I14478));
  NOT NOT1_1178(.VSS(VSS),.VDD(VDD),.Y(g6016),.A(g210));
  NOT NOT1_1179(.VSS(VSS),.VDD(VDD),.Y(g6017),.A(g888));
  NOT NOT1_1180(.VSS(VSS),.VDD(VDD),.Y(g6018),.A(g894));
  NOT NOT1_1181(.VSS(VSS),.VDD(VDD),.Y(g6019),.A(g1471));
  NOT NOT1_1182(.VSS(VSS),.VDD(VDD),.Y(g6020),.A(g1573));
  NOT NOT1_1183(.VSS(VSS),.VDD(VDD),.Y(g6021),.A(g1579));
  NOT NOT1_1184(.VSS(VSS),.VDD(VDD),.Y(g6022),.A(g1585));
  NOT NOT1_1185(.VSS(VSS),.VDD(VDD),.Y(g6023),.A(g1654));
  NOT NOT1_1186(.VSS(VSS),.VDD(VDD),.Y(I14489),.A(g1496));
  NOT NOT1_1187(.VSS(VSS),.VDD(VDD),.Y(g6024),.A(I14489));
  NOT NOT1_1188(.VSS(VSS),.VDD(VDD),.Y(g6025),.A(g2264));
  NOT NOT1_1189(.VSS(VSS),.VDD(VDD),.Y(g6026),.A(g2270));
  NOT NOT1_1190(.VSS(VSS),.VDD(VDD),.Y(g6027),.A(g2339));
  NOT NOT1_1191(.VSS(VSS),.VDD(VDD),.Y(g6028),.A(g2345));
  NOT NOT1_1192(.VSS(VSS),.VDD(VDD),.Y(I14496),.A(g3226));
  NOT NOT1_1193(.VSS(VSS),.VDD(VDD),.Y(g6029),.A(I14496));
  NOT NOT1_1194(.VSS(VSS),.VDD(VDD),.Y(I14499),.A(g3214));
  NOT NOT1_1195(.VSS(VSS),.VDD(VDD),.Y(g6030),.A(I14499));
  NOT NOT1_1196(.VSS(VSS),.VDD(VDD),.Y(I14502),.A(g471));
  NOT NOT1_1197(.VSS(VSS),.VDD(VDD),.Y(g6031),.A(I14502));
  NOT NOT1_1198(.VSS(VSS),.VDD(VDD),.Y(g6032),.A(g897));
  NOT NOT1_1199(.VSS(VSS),.VDD(VDD),.Y(g6033),.A(g1582));
  NOT NOT1_1200(.VSS(VSS),.VDD(VDD),.Y(g6034),.A(g1588));
  NOT NOT1_1201(.VSS(VSS),.VDD(VDD),.Y(g6035),.A(g2165));
  NOT NOT1_1202(.VSS(VSS),.VDD(VDD),.Y(g6036),.A(g2267));
  NOT NOT1_1203(.VSS(VSS),.VDD(VDD),.Y(g6037),.A(g2273));
  NOT NOT1_1204(.VSS(VSS),.VDD(VDD),.Y(g6038),.A(g2279));
  NOT NOT1_1205(.VSS(VSS),.VDD(VDD),.Y(g6039),.A(g2348));
  NOT NOT1_1206(.VSS(VSS),.VDD(VDD),.Y(I14513),.A(g2190));
  NOT NOT1_1207(.VSS(VSS),.VDD(VDD),.Y(g6040),.A(I14513));
  NOT NOT1_1208(.VSS(VSS),.VDD(VDD),.Y(I14516),.A(g3215));
  NOT NOT1_1209(.VSS(VSS),.VDD(VDD),.Y(g6041),.A(I14516));
  NOT NOT1_1210(.VSS(VSS),.VDD(VDD),.Y(I14519),.A(g1158));
  NOT NOT1_1211(.VSS(VSS),.VDD(VDD),.Y(g6042),.A(I14519));
  NOT NOT1_1212(.VSS(VSS),.VDD(VDD),.Y(g6043),.A(g1591));
  NOT NOT1_1213(.VSS(VSS),.VDD(VDD),.Y(g6044),.A(g2276));
  NOT NOT1_1214(.VSS(VSS),.VDD(VDD),.Y(g6045),.A(g2282));
  NOT NOT1_1215(.VSS(VSS),.VDD(VDD),.Y(I14525),.A(g1852));
  NOT NOT1_1216(.VSS(VSS),.VDD(VDD),.Y(g6046),.A(I14525));
  NOT NOT1_1217(.VSS(VSS),.VDD(VDD),.Y(g6047),.A(g2285));
  NOT NOT1_1218(.VSS(VSS),.VDD(VDD),.Y(I14529),.A(g3142));
  NOT NOT1_1219(.VSS(VSS),.VDD(VDD),.Y(g6048),.A(I14529));
  NOT NOT1_1220(.VSS(VSS),.VDD(VDD),.Y(I14532),.A(g354));
  NOT NOT1_1221(.VSS(VSS),.VDD(VDD),.Y(g6051),.A(I14532));
  NOT NOT1_1222(.VSS(VSS),.VDD(VDD),.Y(I14535),.A(g2546));
  NOT NOT1_1223(.VSS(VSS),.VDD(VDD),.Y(g6052),.A(I14535));
  NOT NOT1_1224(.VSS(VSS),.VDD(VDD),.Y(I14538),.A(g369));
  NOT NOT1_1225(.VSS(VSS),.VDD(VDD),.Y(g6053),.A(I14538));
  NOT NOT1_1226(.VSS(VSS),.VDD(VDD),.Y(I14541),.A(g455));
  NOT NOT1_1227(.VSS(VSS),.VDD(VDD),.Y(g6054),.A(I14541));
  NOT NOT1_1228(.VSS(VSS),.VDD(VDD),.Y(I14544),.A(g1041));
  NOT NOT1_1229(.VSS(VSS),.VDD(VDD),.Y(g6055),.A(I14544));
  NOT NOT1_1230(.VSS(VSS),.VDD(VDD),.Y(I14547),.A(g384));
  NOT NOT1_1231(.VSS(VSS),.VDD(VDD),.Y(g6056),.A(I14547));
  NOT NOT1_1232(.VSS(VSS),.VDD(VDD),.Y(I14550),.A(g458));
  NOT NOT1_1233(.VSS(VSS),.VDD(VDD),.Y(g6057),.A(I14550));
  NOT NOT1_1234(.VSS(VSS),.VDD(VDD),.Y(I14553),.A(g1056));
  NOT NOT1_1235(.VSS(VSS),.VDD(VDD),.Y(g6058),.A(I14553));
  NOT NOT1_1236(.VSS(VSS),.VDD(VDD),.Y(I14556),.A(g1142));
  NOT NOT1_1237(.VSS(VSS),.VDD(VDD),.Y(g6059),.A(I14556));
  NOT NOT1_1238(.VSS(VSS),.VDD(VDD),.Y(I14559),.A(g1735));
  NOT NOT1_1239(.VSS(VSS),.VDD(VDD),.Y(g6060),.A(I14559));
  NOT NOT1_1240(.VSS(VSS),.VDD(VDD),.Y(I14562),.A(g398));
  NOT NOT1_1241(.VSS(VSS),.VDD(VDD),.Y(g6061),.A(I14562));
  NOT NOT1_1242(.VSS(VSS),.VDD(VDD),.Y(I14565),.A(g461));
  NOT NOT1_1243(.VSS(VSS),.VDD(VDD),.Y(g6062),.A(I14565));
  NOT NOT1_1244(.VSS(VSS),.VDD(VDD),.Y(I14568),.A(g1071));
  NOT NOT1_1245(.VSS(VSS),.VDD(VDD),.Y(g6063),.A(I14568));
  NOT NOT1_1246(.VSS(VSS),.VDD(VDD),.Y(I14571),.A(g1145));
  NOT NOT1_1247(.VSS(VSS),.VDD(VDD),.Y(g6064),.A(I14571));
  NOT NOT1_1248(.VSS(VSS),.VDD(VDD),.Y(I14574),.A(g1750));
  NOT NOT1_1249(.VSS(VSS),.VDD(VDD),.Y(g6065),.A(I14574));
  NOT NOT1_1250(.VSS(VSS),.VDD(VDD),.Y(I14577),.A(g1836));
  NOT NOT1_1251(.VSS(VSS),.VDD(VDD),.Y(g6066),.A(I14577));
  NOT NOT1_1252(.VSS(VSS),.VDD(VDD),.Y(I14580),.A(g2429));
  NOT NOT1_1253(.VSS(VSS),.VDD(VDD),.Y(g6067),.A(I14580));
  NOT NOT1_1254(.VSS(VSS),.VDD(VDD),.Y(g6068),.A(g499));
  NOT NOT1_1255(.VSS(VSS),.VDD(VDD),.Y(I14584),.A(g465));
  NOT NOT1_1256(.VSS(VSS),.VDD(VDD),.Y(g6079),.A(I14584));
  NOT NOT1_1257(.VSS(VSS),.VDD(VDD),.Y(I14587),.A(g1085));
  NOT NOT1_1258(.VSS(VSS),.VDD(VDD),.Y(g6080),.A(I14587));
  NOT NOT1_1259(.VSS(VSS),.VDD(VDD),.Y(I14590),.A(g1148));
  NOT NOT1_1260(.VSS(VSS),.VDD(VDD),.Y(g6081),.A(I14590));
  NOT NOT1_1261(.VSS(VSS),.VDD(VDD),.Y(I14593),.A(g1765));
  NOT NOT1_1262(.VSS(VSS),.VDD(VDD),.Y(g6082),.A(I14593));
  NOT NOT1_1263(.VSS(VSS),.VDD(VDD),.Y(I14596),.A(g1839));
  NOT NOT1_1264(.VSS(VSS),.VDD(VDD),.Y(g6083),.A(I14596));
  NOT NOT1_1265(.VSS(VSS),.VDD(VDD),.Y(I14599),.A(g2444));
  NOT NOT1_1266(.VSS(VSS),.VDD(VDD),.Y(g6084),.A(I14599));
  NOT NOT1_1267(.VSS(VSS),.VDD(VDD),.Y(I14602),.A(g2530));
  NOT NOT1_1268(.VSS(VSS),.VDD(VDD),.Y(g6085),.A(I14602));
  NOT NOT1_1269(.VSS(VSS),.VDD(VDD),.Y(I14605),.A(g468));
  NOT NOT1_1270(.VSS(VSS),.VDD(VDD),.Y(g6086),.A(I14605));
  NOT NOT1_1271(.VSS(VSS),.VDD(VDD),.Y(g6087),.A(g1186));
  NOT NOT1_1272(.VSS(VSS),.VDD(VDD),.Y(I14609),.A(g1152));
  NOT NOT1_1273(.VSS(VSS),.VDD(VDD),.Y(g6098),.A(I14609));
  NOT NOT1_1274(.VSS(VSS),.VDD(VDD),.Y(I14612),.A(g1779));
  NOT NOT1_1275(.VSS(VSS),.VDD(VDD),.Y(g6099),.A(I14612));
  NOT NOT1_1276(.VSS(VSS),.VDD(VDD),.Y(I14615),.A(g1842));
  NOT NOT1_1277(.VSS(VSS),.VDD(VDD),.Y(g6100),.A(I14615));
  NOT NOT1_1278(.VSS(VSS),.VDD(VDD),.Y(I14618),.A(g2459));
  NOT NOT1_1279(.VSS(VSS),.VDD(VDD),.Y(g6101),.A(I14618));
  NOT NOT1_1280(.VSS(VSS),.VDD(VDD),.Y(I14621),.A(g2533));
  NOT NOT1_1281(.VSS(VSS),.VDD(VDD),.Y(g6102),.A(I14621));
  NOT NOT1_1282(.VSS(VSS),.VDD(VDD),.Y(I14624),.A(g1155));
  NOT NOT1_1283(.VSS(VSS),.VDD(VDD),.Y(g6103),.A(I14624));
  NOT NOT1_1284(.VSS(VSS),.VDD(VDD),.Y(g6104),.A(g1880));
  NOT NOT1_1285(.VSS(VSS),.VDD(VDD),.Y(I14628),.A(g1846));
  NOT NOT1_1286(.VSS(VSS),.VDD(VDD),.Y(g6115),.A(I14628));
  NOT NOT1_1287(.VSS(VSS),.VDD(VDD),.Y(I14631),.A(g2473));
  NOT NOT1_1288(.VSS(VSS),.VDD(VDD),.Y(g6116),.A(I14631));
  NOT NOT1_1289(.VSS(VSS),.VDD(VDD),.Y(I14634),.A(g2536));
  NOT NOT1_1290(.VSS(VSS),.VDD(VDD),.Y(g6117),.A(I14634));
  NOT NOT1_1291(.VSS(VSS),.VDD(VDD),.Y(I14637),.A(g1849));
  NOT NOT1_1292(.VSS(VSS),.VDD(VDD),.Y(g6118),.A(I14637));
  NOT NOT1_1293(.VSS(VSS),.VDD(VDD),.Y(g6119),.A(g2574));
  NOT NOT1_1294(.VSS(VSS),.VDD(VDD),.Y(I14641),.A(g2540));
  NOT NOT1_1295(.VSS(VSS),.VDD(VDD),.Y(g6130),.A(I14641));
  NOT NOT1_1296(.VSS(VSS),.VDD(VDD),.Y(I14644),.A(g3142));
  NOT NOT1_1297(.VSS(VSS),.VDD(VDD),.Y(g6131),.A(I14644));
  NOT NOT1_1298(.VSS(VSS),.VDD(VDD),.Y(I14647),.A(g2543));
  NOT NOT1_1299(.VSS(VSS),.VDD(VDD),.Y(g6134),.A(I14647));
  NOT NOT1_1300(.VSS(VSS),.VDD(VDD),.Y(I14650),.A(g525));
  NOT NOT1_1301(.VSS(VSS),.VDD(VDD),.Y(g6135),.A(I14650));
  NOT NOT1_1302(.VSS(VSS),.VDD(VDD),.Y(g6136),.A(g672));
  NOT NOT1_1303(.VSS(VSS),.VDD(VDD),.Y(I14654),.A(g3220));
  NOT NOT1_1304(.VSS(VSS),.VDD(VDD),.Y(g6139),.A(I14654));
  NOT NOT1_1305(.VSS(VSS),.VDD(VDD),.Y(g6140),.A(g524));
  NOT NOT1_1306(.VSS(VSS),.VDD(VDD),.Y(g6141),.A(g554));
  NOT NOT1_1307(.VSS(VSS),.VDD(VDD),.Y(g6142),.A(g679));
  NOT NOT1_1308(.VSS(VSS),.VDD(VDD),.Y(I14660),.A(g1211));
  NOT NOT1_1309(.VSS(VSS),.VDD(VDD),.Y(g6145),.A(I14660));
  NOT NOT1_1310(.VSS(VSS),.VDD(VDD),.Y(g6146),.A(g1358));
  NOT NOT1_1311(.VSS(VSS),.VDD(VDD),.Y(g6149),.A(g3097));
  NOT NOT1_1312(.VSS(VSS),.VDD(VDD),.Y(I14665),.A(g3147));
  NOT NOT1_1313(.VSS(VSS),.VDD(VDD),.Y(g6153),.A(I14665));
  NOT NOT1_1314(.VSS(VSS),.VDD(VDD),.Y(I14668),.A(g3232));
  NOT NOT1_1315(.VSS(VSS),.VDD(VDD),.Y(g6156),.A(I14668));
  NOT NOT1_1316(.VSS(VSS),.VDD(VDD),.Y(g6157),.A(g686));
  NOT NOT1_1317(.VSS(VSS),.VDD(VDD),.Y(g6161),.A(g1210));
  NOT NOT1_1318(.VSS(VSS),.VDD(VDD),.Y(g6162),.A(g1240));
  NOT NOT1_1319(.VSS(VSS),.VDD(VDD),.Y(g6163),.A(g1365));
  NOT NOT1_1320(.VSS(VSS),.VDD(VDD),.Y(I14675),.A(g1905));
  NOT NOT1_1321(.VSS(VSS),.VDD(VDD),.Y(g6166),.A(I14675));
  NOT NOT1_1322(.VSS(VSS),.VDD(VDD),.Y(g6167),.A(g2052));
  NOT NOT1_1323(.VSS(VSS),.VDD(VDD),.Y(g6170),.A(g3098));
  NOT NOT1_1324(.VSS(VSS),.VDD(VDD),.Y(g6173),.A(g557));
  NOT NOT1_1325(.VSS(VSS),.VDD(VDD),.Y(g6177),.A(g633));
  NOT NOT1_1326(.VSS(VSS),.VDD(VDD),.Y(g6180),.A(g692));
  NOT NOT1_1327(.VSS(VSS),.VDD(VDD),.Y(g6183),.A(g291));
  NOT NOT1_1328(.VSS(VSS),.VDD(VDD),.Y(g6184),.A(g1372));
  NOT NOT1_1329(.VSS(VSS),.VDD(VDD),.Y(g6188),.A(g1904));
  NOT NOT1_1330(.VSS(VSS),.VDD(VDD),.Y(g6189),.A(g1934));
  NOT NOT1_1331(.VSS(VSS),.VDD(VDD),.Y(g6190),.A(g2059));
  NOT NOT1_1332(.VSS(VSS),.VDD(VDD),.Y(I14688),.A(g2599));
  NOT NOT1_1333(.VSS(VSS),.VDD(VDD),.Y(g6193),.A(I14688));
  NOT NOT1_1334(.VSS(VSS),.VDD(VDD),.Y(g6194),.A(g2746));
  NOT NOT1_1335(.VSS(VSS),.VDD(VDD),.Y(g6197),.A(g3099));
  NOT NOT1_1336(.VSS(VSS),.VDD(VDD),.Y(g6200),.A(g542));
  NOT NOT1_1337(.VSS(VSS),.VDD(VDD),.Y(g6201),.A(g646));
  NOT NOT1_1338(.VSS(VSS),.VDD(VDD),.Y(g6204),.A(g289));
  NOT NOT1_1339(.VSS(VSS),.VDD(VDD),.Y(g6205),.A(g1243));
  NOT NOT1_1340(.VSS(VSS),.VDD(VDD),.Y(g6209),.A(g1319));
  NOT NOT1_1341(.VSS(VSS),.VDD(VDD),.Y(g6212),.A(g1378));
  NOT NOT1_1342(.VSS(VSS),.VDD(VDD),.Y(g6215),.A(g978));
  NOT NOT1_1343(.VSS(VSS),.VDD(VDD),.Y(g6216),.A(g2066));
  NOT NOT1_1344(.VSS(VSS),.VDD(VDD),.Y(g6220),.A(g2598));
  NOT NOT1_1345(.VSS(VSS),.VDD(VDD),.Y(g6221),.A(g2628));
  NOT NOT1_1346(.VSS(VSS),.VDD(VDD),.Y(g6222),.A(g2753));
  NOT NOT1_1347(.VSS(VSS),.VDD(VDD),.Y(I14704),.A(g2818));
  NOT NOT1_1348(.VSS(VSS),.VDD(VDD),.Y(g6225),.A(I14704));
  NOT NOT1_1349(.VSS(VSS),.VDD(VDD),.Y(g6226),.A(g2818));
  NOT NOT1_1350(.VSS(VSS),.VDD(VDD),.Y(g6227),.A(g3100));
  NOT NOT1_1351(.VSS(VSS),.VDD(VDD),.Y(I14709),.A(g3229));
  NOT NOT1_1352(.VSS(VSS),.VDD(VDD),.Y(g6230),.A(I14709));
  NOT NOT1_1353(.VSS(VSS),.VDD(VDD),.Y(I14712),.A(g138));
  NOT NOT1_1354(.VSS(VSS),.VDD(VDD),.Y(g6231),.A(I14712));
  NOT NOT1_1355(.VSS(VSS),.VDD(VDD),.Y(I14715),.A(g138));
  NOT NOT1_1356(.VSS(VSS),.VDD(VDD),.Y(g6232),.A(I14715));
  NOT NOT1_1357(.VSS(VSS),.VDD(VDD),.Y(g6281),.A(g510));
  NOT NOT1_1358(.VSS(VSS),.VDD(VDD),.Y(g6284),.A(g640));
  NOT NOT1_1359(.VSS(VSS),.VDD(VDD),.Y(g6288),.A(g287));
  NOT NOT1_1360(.VSS(VSS),.VDD(VDD),.Y(g6289),.A(g1228));
  NOT NOT1_1361(.VSS(VSS),.VDD(VDD),.Y(g6290),.A(g1332));
  NOT NOT1_1362(.VSS(VSS),.VDD(VDD),.Y(g6293),.A(g976));
  NOT NOT1_1363(.VSS(VSS),.VDD(VDD),.Y(g6294),.A(g1937));
  NOT NOT1_1364(.VSS(VSS),.VDD(VDD),.Y(g6298),.A(g2013));
  NOT NOT1_1365(.VSS(VSS),.VDD(VDD),.Y(g6301),.A(g2072));
  NOT NOT1_1366(.VSS(VSS),.VDD(VDD),.Y(g6304),.A(g1672));
  NOT NOT1_1367(.VSS(VSS),.VDD(VDD),.Y(g6305),.A(g2760));
  NOT NOT1_1368(.VSS(VSS),.VDD(VDD),.Y(g6309),.A(g14));
  NOT NOT1_1369(.VSS(VSS),.VDD(VDD),.Y(g6310),.A(g3101));
  NOT NOT1_1370(.VSS(VSS),.VDD(VDD),.Y(I14731),.A(g135));
  NOT NOT1_1371(.VSS(VSS),.VDD(VDD),.Y(g6313),.A(I14731));
  NOT NOT1_1372(.VSS(VSS),.VDD(VDD),.Y(I14734),.A(g135));
  NOT NOT1_1373(.VSS(VSS),.VDD(VDD),.Y(g6314),.A(I14734));
  NOT NOT1_1374(.VSS(VSS),.VDD(VDD),.Y(g6363),.A(g653));
  NOT NOT1_1375(.VSS(VSS),.VDD(VDD),.Y(g6367),.A(g285));
  NOT NOT1_1376(.VSS(VSS),.VDD(VDD),.Y(I14739),.A(g826));
  NOT NOT1_1377(.VSS(VSS),.VDD(VDD),.Y(g6368),.A(I14739));
  NOT NOT1_1378(.VSS(VSS),.VDD(VDD),.Y(I14742),.A(g826));
  NOT NOT1_1379(.VSS(VSS),.VDD(VDD),.Y(g6369),.A(I14742));
  NOT NOT1_1380(.VSS(VSS),.VDD(VDD),.Y(g6418),.A(g1196));
  NOT NOT1_1381(.VSS(VSS),.VDD(VDD),.Y(g6421),.A(g1326));
  NOT NOT1_1382(.VSS(VSS),.VDD(VDD),.Y(g6425),.A(g974));
  NOT NOT1_1383(.VSS(VSS),.VDD(VDD),.Y(g6426),.A(g1922));
  NOT NOT1_1384(.VSS(VSS),.VDD(VDD),.Y(g6427),.A(g2026));
  NOT NOT1_1385(.VSS(VSS),.VDD(VDD),.Y(g6430),.A(g1670));
  NOT NOT1_1386(.VSS(VSS),.VDD(VDD),.Y(g6431),.A(g2631));
  NOT NOT1_1387(.VSS(VSS),.VDD(VDD),.Y(g6435),.A(g2707));
  NOT NOT1_1388(.VSS(VSS),.VDD(VDD),.Y(g6438),.A(g2766));
  NOT NOT1_1389(.VSS(VSS),.VDD(VDD),.Y(g6441),.A(g2366));
  NOT NOT1_1390(.VSS(VSS),.VDD(VDD),.Y(I14755),.A(g2821));
  NOT NOT1_1391(.VSS(VSS),.VDD(VDD),.Y(g6442),.A(I14755));
  NOT NOT1_1392(.VSS(VSS),.VDD(VDD),.Y(g6443),.A(g2821));
  NOT NOT1_1393(.VSS(VSS),.VDD(VDD),.Y(g6444),.A(g3102));
  NOT NOT1_1394(.VSS(VSS),.VDD(VDD),.Y(I14760),.A(g405));
  NOT NOT1_1395(.VSS(VSS),.VDD(VDD),.Y(g6447),.A(I14760));
  NOT NOT1_1396(.VSS(VSS),.VDD(VDD),.Y(I14763),.A(g405));
  NOT NOT1_1397(.VSS(VSS),.VDD(VDD),.Y(g6448),.A(I14763));
  NOT NOT1_1398(.VSS(VSS),.VDD(VDD),.Y(I14766),.A(g545));
  NOT NOT1_1399(.VSS(VSS),.VDD(VDD),.Y(g6485),.A(I14766));
  NOT NOT1_1400(.VSS(VSS),.VDD(VDD),.Y(I14769),.A(g545));
  NOT NOT1_1401(.VSS(VSS),.VDD(VDD),.Y(g6486),.A(I14769));
  NOT NOT1_1402(.VSS(VSS),.VDD(VDD),.Y(g6512),.A(g544));
  NOT NOT1_1403(.VSS(VSS),.VDD(VDD),.Y(g6513),.A(g660));
  NOT NOT1_1404(.VSS(VSS),.VDD(VDD),.Y(g6517),.A(g283));
  NOT NOT1_1405(.VSS(VSS),.VDD(VDD),.Y(I14775),.A(g823));
  NOT NOT1_1406(.VSS(VSS),.VDD(VDD),.Y(g6518),.A(I14775));
  NOT NOT1_1407(.VSS(VSS),.VDD(VDD),.Y(I14778),.A(g823));
  NOT NOT1_1408(.VSS(VSS),.VDD(VDD),.Y(g6519),.A(I14778));
  NOT NOT1_1409(.VSS(VSS),.VDD(VDD),.Y(g6568),.A(g1339));
  NOT NOT1_1410(.VSS(VSS),.VDD(VDD),.Y(g6572),.A(g972));
  NOT NOT1_1411(.VSS(VSS),.VDD(VDD),.Y(I14783),.A(g1520));
  NOT NOT1_1412(.VSS(VSS),.VDD(VDD),.Y(g6573),.A(I14783));
  NOT NOT1_1413(.VSS(VSS),.VDD(VDD),.Y(I14786),.A(g1520));
  NOT NOT1_1414(.VSS(VSS),.VDD(VDD),.Y(g6574),.A(I14786));
  NOT NOT1_1415(.VSS(VSS),.VDD(VDD),.Y(g6623),.A(g1890));
  NOT NOT1_1416(.VSS(VSS),.VDD(VDD),.Y(g6626),.A(g2020));
  NOT NOT1_1417(.VSS(VSS),.VDD(VDD),.Y(g6630),.A(g1668));
  NOT NOT1_1418(.VSS(VSS),.VDD(VDD),.Y(g6631),.A(g2616));
  NOT NOT1_1419(.VSS(VSS),.VDD(VDD),.Y(g6632),.A(g2720));
  NOT NOT1_1420(.VSS(VSS),.VDD(VDD),.Y(g6635),.A(g2364));
  NOT NOT1_1421(.VSS(VSS),.VDD(VDD),.Y(g6636),.A(g1491));
  NOT NOT1_1422(.VSS(VSS),.VDD(VDD),.Y(g6637),.A(g5));
  NOT NOT1_1423(.VSS(VSS),.VDD(VDD),.Y(g6638),.A(g3103));
  NOT NOT1_1424(.VSS(VSS),.VDD(VDD),.Y(g6641),.A(g113));
  NOT NOT1_1425(.VSS(VSS),.VDD(VDD),.Y(I14799),.A(g551));
  NOT NOT1_1426(.VSS(VSS),.VDD(VDD),.Y(g6642),.A(I14799));
  NOT NOT1_1427(.VSS(VSS),.VDD(VDD),.Y(I14802),.A(g551));
  NOT NOT1_1428(.VSS(VSS),.VDD(VDD),.Y(g6643),.A(I14802));
  NOT NOT1_1429(.VSS(VSS),.VDD(VDD),.Y(g6672),.A(g464));
  NOT NOT1_1430(.VSS(VSS),.VDD(VDD),.Y(g6675),.A(g458));
  NOT NOT1_1431(.VSS(VSS),.VDD(VDD),.Y(g6676),.A(g559));
  NOT NOT1_1432(.VSS(VSS),.VDD(VDD),.Y(I14808),.A(g623));
  NOT NOT1_1433(.VSS(VSS),.VDD(VDD),.Y(g6677),.A(I14808));
  NOT NOT1_1434(.VSS(VSS),.VDD(VDD),.Y(I14811),.A(g623));
  NOT NOT1_1435(.VSS(VSS),.VDD(VDD),.Y(g6678),.A(I14811));
  NOT NOT1_1436(.VSS(VSS),.VDD(VDD),.Y(g6707),.A(g666));
  NOT NOT1_1437(.VSS(VSS),.VDD(VDD),.Y(g6711),.A(g281));
  NOT NOT1_1438(.VSS(VSS),.VDD(VDD),.Y(I14816),.A(g1092));
  NOT NOT1_1439(.VSS(VSS),.VDD(VDD),.Y(g6712),.A(I14816));
  NOT NOT1_1440(.VSS(VSS),.VDD(VDD),.Y(I14819),.A(g1092));
  NOT NOT1_1441(.VSS(VSS),.VDD(VDD),.Y(g6713),.A(I14819));
  NOT NOT1_1442(.VSS(VSS),.VDD(VDD),.Y(I14822),.A(g1231));
  NOT NOT1_1443(.VSS(VSS),.VDD(VDD),.Y(g6750),.A(I14822));
  NOT NOT1_1444(.VSS(VSS),.VDD(VDD),.Y(I14825),.A(g1231));
  NOT NOT1_1445(.VSS(VSS),.VDD(VDD),.Y(g6751),.A(I14825));
  NOT NOT1_1446(.VSS(VSS),.VDD(VDD),.Y(g6776),.A(g1230));
  NOT NOT1_1447(.VSS(VSS),.VDD(VDD),.Y(g6777),.A(g1346));
  NOT NOT1_1448(.VSS(VSS),.VDD(VDD),.Y(g6781),.A(g970));
  NOT NOT1_1449(.VSS(VSS),.VDD(VDD),.Y(I14831),.A(g1517));
  NOT NOT1_1450(.VSS(VSS),.VDD(VDD),.Y(g6782),.A(I14831));
  NOT NOT1_1451(.VSS(VSS),.VDD(VDD),.Y(I14834),.A(g1517));
  NOT NOT1_1452(.VSS(VSS),.VDD(VDD),.Y(g6783),.A(I14834));
  NOT NOT1_1453(.VSS(VSS),.VDD(VDD),.Y(g6832),.A(g2033));
  NOT NOT1_1454(.VSS(VSS),.VDD(VDD),.Y(g6836),.A(g1666));
  NOT NOT1_1455(.VSS(VSS),.VDD(VDD),.Y(I14839),.A(g2214));
  NOT NOT1_1456(.VSS(VSS),.VDD(VDD),.Y(g6837),.A(I14839));
  NOT NOT1_1457(.VSS(VSS),.VDD(VDD),.Y(I14842),.A(g2214));
  NOT NOT1_1458(.VSS(VSS),.VDD(VDD),.Y(g6838),.A(I14842));
  NOT NOT1_1459(.VSS(VSS),.VDD(VDD),.Y(g6887),.A(g2584));
  NOT NOT1_1460(.VSS(VSS),.VDD(VDD),.Y(g6890),.A(g2714));
  NOT NOT1_1461(.VSS(VSS),.VDD(VDD),.Y(g6894),.A(g2362));
  NOT NOT1_1462(.VSS(VSS),.VDD(VDD),.Y(I14848),.A(g2824));
  NOT NOT1_1463(.VSS(VSS),.VDD(VDD),.Y(g6895),.A(I14848));
  NOT NOT1_1464(.VSS(VSS),.VDD(VDD),.Y(g6896),.A(g2824));
  NOT NOT1_1465(.VSS(VSS),.VDD(VDD),.Y(g6897),.A(g1486));
  NOT NOT1_1466(.VSS(VSS),.VDD(VDD),.Y(g6898),.A(g2993));
  NOT NOT1_1467(.VSS(VSS),.VDD(VDD),.Y(g6901),.A(g3006));
  NOT NOT1_1468(.VSS(VSS),.VDD(VDD),.Y(g6905),.A(g3104));
  NOT NOT1_1469(.VSS(VSS),.VDD(VDD),.Y(g6908),.A(g484));
  NOT NOT1_1470(.VSS(VSS),.VDD(VDD),.Y(I14857),.A(g626));
  NOT NOT1_1471(.VSS(VSS),.VDD(VDD),.Y(g6911),.A(I14857));
  NOT NOT1_1472(.VSS(VSS),.VDD(VDD),.Y(I14860),.A(g626));
  NOT NOT1_1473(.VSS(VSS),.VDD(VDD),.Y(g6912),.A(I14860));
  NOT NOT1_1474(.VSS(VSS),.VDD(VDD),.Y(g6942),.A(g279));
  NOT NOT1_1475(.VSS(VSS),.VDD(VDD),.Y(g6943),.A(g801));
  NOT NOT1_1476(.VSS(VSS),.VDD(VDD),.Y(I14865),.A(g1237));
  NOT NOT1_1477(.VSS(VSS),.VDD(VDD),.Y(g6944),.A(I14865));
  NOT NOT1_1478(.VSS(VSS),.VDD(VDD),.Y(I14868),.A(g1237));
  NOT NOT1_1479(.VSS(VSS),.VDD(VDD),.Y(g6945),.A(I14868));
  NOT NOT1_1480(.VSS(VSS),.VDD(VDD),.Y(g6974),.A(g1151));
  NOT NOT1_1481(.VSS(VSS),.VDD(VDD),.Y(g6977),.A(g1145));
  NOT NOT1_1482(.VSS(VSS),.VDD(VDD),.Y(g6978),.A(g1245));
  NOT NOT1_1483(.VSS(VSS),.VDD(VDD),.Y(I14874),.A(g1309));
  NOT NOT1_1484(.VSS(VSS),.VDD(VDD),.Y(g6979),.A(I14874));
  NOT NOT1_1485(.VSS(VSS),.VDD(VDD),.Y(I14877),.A(g1309));
  NOT NOT1_1486(.VSS(VSS),.VDD(VDD),.Y(g6980),.A(I14877));
  NOT NOT1_1487(.VSS(VSS),.VDD(VDD),.Y(g7009),.A(g1352));
  NOT NOT1_1488(.VSS(VSS),.VDD(VDD),.Y(g7013),.A(g968));
  NOT NOT1_1489(.VSS(VSS),.VDD(VDD),.Y(I14882),.A(g1786));
  NOT NOT1_1490(.VSS(VSS),.VDD(VDD),.Y(g7014),.A(I14882));
  NOT NOT1_1491(.VSS(VSS),.VDD(VDD),.Y(I14885),.A(g1786));
  NOT NOT1_1492(.VSS(VSS),.VDD(VDD),.Y(g7015),.A(I14885));
  NOT NOT1_1493(.VSS(VSS),.VDD(VDD),.Y(I14888),.A(g1925));
  NOT NOT1_1494(.VSS(VSS),.VDD(VDD),.Y(g7052),.A(I14888));
  NOT NOT1_1495(.VSS(VSS),.VDD(VDD),.Y(I14891),.A(g1925));
  NOT NOT1_1496(.VSS(VSS),.VDD(VDD),.Y(g7053),.A(I14891));
  NOT NOT1_1497(.VSS(VSS),.VDD(VDD),.Y(g7078),.A(g1924));
  NOT NOT1_1498(.VSS(VSS),.VDD(VDD),.Y(g7079),.A(g2040));
  NOT NOT1_1499(.VSS(VSS),.VDD(VDD),.Y(g7083),.A(g1664));
  NOT NOT1_1500(.VSS(VSS),.VDD(VDD),.Y(I14897),.A(g2211));
  NOT NOT1_1501(.VSS(VSS),.VDD(VDD),.Y(g7084),.A(I14897));
  NOT NOT1_1502(.VSS(VSS),.VDD(VDD),.Y(I14900),.A(g2211));
  NOT NOT1_1503(.VSS(VSS),.VDD(VDD),.Y(g7085),.A(I14900));
  NOT NOT1_1504(.VSS(VSS),.VDD(VDD),.Y(g7134),.A(g2727));
  NOT NOT1_1505(.VSS(VSS),.VDD(VDD),.Y(g7138),.A(g2360));
  NOT NOT1_1506(.VSS(VSS),.VDD(VDD),.Y(g7139),.A(g1481));
  NOT NOT1_1507(.VSS(VSS),.VDD(VDD),.Y(g7140),.A(g2170));
  NOT NOT1_1508(.VSS(VSS),.VDD(VDD),.Y(g7141),.A(g2195));
  NOT NOT1_1509(.VSS(VSS),.VDD(VDD),.Y(g7142),.A(g8));
  NOT NOT1_1510(.VSS(VSS),.VDD(VDD),.Y(g7143),.A(g2998));
  NOT NOT1_1511(.VSS(VSS),.VDD(VDD),.Y(g7146),.A(g3013));
  NOT NOT1_1512(.VSS(VSS),.VDD(VDD),.Y(g7149),.A(g3105));
  NOT NOT1_1513(.VSS(VSS),.VDD(VDD),.Y(g7152),.A(g3136));
  NOT NOT1_1514(.VSS(VSS),.VDD(VDD),.Y(g7153),.A(g480));
  NOT NOT1_1515(.VSS(VSS),.VDD(VDD),.Y(g7156),.A(g461));
  NOT NOT1_1516(.VSS(VSS),.VDD(VDD),.Y(g7157),.A(g453));
  NOT NOT1_1517(.VSS(VSS),.VDD(VDD),.Y(g7158),.A(g1171));
  NOT NOT1_1518(.VSS(VSS),.VDD(VDD),.Y(I14917),.A(g1312));
  NOT NOT1_1519(.VSS(VSS),.VDD(VDD),.Y(g7161),.A(I14917));
  NOT NOT1_1520(.VSS(VSS),.VDD(VDD),.Y(I14920),.A(g1312));
  NOT NOT1_1521(.VSS(VSS),.VDD(VDD),.Y(g7162),.A(I14920));
  NOT NOT1_1522(.VSS(VSS),.VDD(VDD),.Y(g7192),.A(g966));
  NOT NOT1_1523(.VSS(VSS),.VDD(VDD),.Y(g7193),.A(g1491));
  NOT NOT1_1524(.VSS(VSS),.VDD(VDD),.Y(I14925),.A(g1931));
  NOT NOT1_1525(.VSS(VSS),.VDD(VDD),.Y(g7194),.A(I14925));
  NOT NOT1_1526(.VSS(VSS),.VDD(VDD),.Y(I14928),.A(g1931));
  NOT NOT1_1527(.VSS(VSS),.VDD(VDD),.Y(g7195),.A(I14928));
  NOT NOT1_1528(.VSS(VSS),.VDD(VDD),.Y(g7224),.A(g1845));
  NOT NOT1_1529(.VSS(VSS),.VDD(VDD),.Y(g7227),.A(g1839));
  NOT NOT1_1530(.VSS(VSS),.VDD(VDD),.Y(g7228),.A(g1939));
  NOT NOT1_1531(.VSS(VSS),.VDD(VDD),.Y(I14934),.A(g2003));
  NOT NOT1_1532(.VSS(VSS),.VDD(VDD),.Y(g7229),.A(I14934));
  NOT NOT1_1533(.VSS(VSS),.VDD(VDD),.Y(I14937),.A(g2003));
  NOT NOT1_1534(.VSS(VSS),.VDD(VDD),.Y(g7230),.A(I14937));
  NOT NOT1_1535(.VSS(VSS),.VDD(VDD),.Y(g7259),.A(g2046));
  NOT NOT1_1536(.VSS(VSS),.VDD(VDD),.Y(g7263),.A(g1662));
  NOT NOT1_1537(.VSS(VSS),.VDD(VDD),.Y(I14942),.A(g2480));
  NOT NOT1_1538(.VSS(VSS),.VDD(VDD),.Y(g7264),.A(I14942));
  NOT NOT1_1539(.VSS(VSS),.VDD(VDD),.Y(I14945),.A(g2480));
  NOT NOT1_1540(.VSS(VSS),.VDD(VDD),.Y(g7265),.A(I14945));
  NOT NOT1_1541(.VSS(VSS),.VDD(VDD),.Y(I14948),.A(g2619));
  NOT NOT1_1542(.VSS(VSS),.VDD(VDD),.Y(g7302),.A(I14948));
  NOT NOT1_1543(.VSS(VSS),.VDD(VDD),.Y(I14951),.A(g2619));
  NOT NOT1_1544(.VSS(VSS),.VDD(VDD),.Y(g7303),.A(I14951));
  NOT NOT1_1545(.VSS(VSS),.VDD(VDD),.Y(g7328),.A(g2618));
  NOT NOT1_1546(.VSS(VSS),.VDD(VDD),.Y(g7329),.A(g2734));
  NOT NOT1_1547(.VSS(VSS),.VDD(VDD),.Y(g7333),.A(g2358));
  NOT NOT1_1548(.VSS(VSS),.VDD(VDD),.Y(I14957),.A(g2827));
  NOT NOT1_1549(.VSS(VSS),.VDD(VDD),.Y(g7334),.A(I14957));
  NOT NOT1_1550(.VSS(VSS),.VDD(VDD),.Y(g7335),.A(g2827));
  NOT NOT1_1551(.VSS(VSS),.VDD(VDD),.Y(g7336),.A(g1476));
  NOT NOT1_1552(.VSS(VSS),.VDD(VDD),.Y(g7337),.A(g2190));
  NOT NOT1_1553(.VSS(VSS),.VDD(VDD),.Y(g7338),.A(g3002));
  NOT NOT1_1554(.VSS(VSS),.VDD(VDD),.Y(g7342),.A(g3024));
  NOT NOT1_1555(.VSS(VSS),.VDD(VDD),.Y(g7345),.A(g3139));
  NOT NOT1_1556(.VSS(VSS),.VDD(VDD),.Y(g7346),.A(g97));
  NOT NOT1_1557(.VSS(VSS),.VDD(VDD),.Y(g7347),.A(g490));
  NOT NOT1_1558(.VSS(VSS),.VDD(VDD),.Y(g7348),.A(g451));
  NOT NOT1_1559(.VSS(VSS),.VDD(VDD),.Y(g7349),.A(g1167));
  NOT NOT1_1560(.VSS(VSS),.VDD(VDD),.Y(g7352),.A(g1148));
  NOT NOT1_1561(.VSS(VSS),.VDD(VDD),.Y(g7353),.A(g1140));
  NOT NOT1_1562(.VSS(VSS),.VDD(VDD),.Y(g7354),.A(g1865));
  NOT NOT1_1563(.VSS(VSS),.VDD(VDD),.Y(I14973),.A(g2006));
  NOT NOT1_1564(.VSS(VSS),.VDD(VDD),.Y(g7357),.A(I14973));
  NOT NOT1_1565(.VSS(VSS),.VDD(VDD),.Y(I14976),.A(g2006));
  NOT NOT1_1566(.VSS(VSS),.VDD(VDD),.Y(g7358),.A(I14976));
  NOT NOT1_1567(.VSS(VSS),.VDD(VDD),.Y(g7388),.A(g1660));
  NOT NOT1_1568(.VSS(VSS),.VDD(VDD),.Y(g7389),.A(g2185));
  NOT NOT1_1569(.VSS(VSS),.VDD(VDD),.Y(I14981),.A(g2625));
  NOT NOT1_1570(.VSS(VSS),.VDD(VDD),.Y(g7390),.A(I14981));
  NOT NOT1_1571(.VSS(VSS),.VDD(VDD),.Y(I14984),.A(g2625));
  NOT NOT1_1572(.VSS(VSS),.VDD(VDD),.Y(g7391),.A(I14984));
  NOT NOT1_1573(.VSS(VSS),.VDD(VDD),.Y(g7420),.A(g2539));
  NOT NOT1_1574(.VSS(VSS),.VDD(VDD),.Y(g7423),.A(g2533));
  NOT NOT1_1575(.VSS(VSS),.VDD(VDD),.Y(g7424),.A(g2633));
  NOT NOT1_1576(.VSS(VSS),.VDD(VDD),.Y(I14990),.A(g2697));
  NOT NOT1_1577(.VSS(VSS),.VDD(VDD),.Y(g7425),.A(I14990));
  NOT NOT1_1578(.VSS(VSS),.VDD(VDD),.Y(I14993),.A(g2697));
  NOT NOT1_1579(.VSS(VSS),.VDD(VDD),.Y(g7426),.A(I14993));
  NOT NOT1_1580(.VSS(VSS),.VDD(VDD),.Y(g7455),.A(g2740));
  NOT NOT1_1581(.VSS(VSS),.VDD(VDD),.Y(g7459),.A(g2356));
  NOT NOT1_1582(.VSS(VSS),.VDD(VDD),.Y(g7460),.A(g1471));
  NOT NOT1_1583(.VSS(VSS),.VDD(VDD),.Y(g7461),.A(g2175));
  NOT NOT1_1584(.VSS(VSS),.VDD(VDD),.Y(g7462),.A(g2912));
  NOT NOT1_1585(.VSS(VSS),.VDD(VDD),.Y(g7465),.A(g2));
  NOT NOT1_1586(.VSS(VSS),.VDD(VDD),.Y(g7466),.A(g3010));
  NOT NOT1_1587(.VSS(VSS),.VDD(VDD),.Y(g7471),.A(g3036));
  NOT NOT1_1588(.VSS(VSS),.VDD(VDD),.Y(g7475),.A(g493));
  NOT NOT1_1589(.VSS(VSS),.VDD(VDD),.Y(g7476),.A(g785));
  NOT NOT1_1590(.VSS(VSS),.VDD(VDD),.Y(g7477),.A(g1177));
  NOT NOT1_1591(.VSS(VSS),.VDD(VDD),.Y(g7478),.A(g1138));
  NOT NOT1_1592(.VSS(VSS),.VDD(VDD),.Y(g7479),.A(g1861));
  NOT NOT1_1593(.VSS(VSS),.VDD(VDD),.Y(g7482),.A(g1842));
  NOT NOT1_1594(.VSS(VSS),.VDD(VDD),.Y(g7483),.A(g1834));
  NOT NOT1_1595(.VSS(VSS),.VDD(VDD),.Y(g7484),.A(g2559));
  NOT NOT1_1596(.VSS(VSS),.VDD(VDD),.Y(I15012),.A(g2700));
  NOT NOT1_1597(.VSS(VSS),.VDD(VDD),.Y(g7487),.A(I15012));
  NOT NOT1_1598(.VSS(VSS),.VDD(VDD),.Y(I15015),.A(g2700));
  NOT NOT1_1599(.VSS(VSS),.VDD(VDD),.Y(g7488),.A(I15015));
  NOT NOT1_1600(.VSS(VSS),.VDD(VDD),.Y(g7518),.A(g2354));
  NOT NOT1_1601(.VSS(VSS),.VDD(VDD),.Y(I15019),.A(g2830));
  NOT NOT1_1602(.VSS(VSS),.VDD(VDD),.Y(g7519),.A(I15019));
  NOT NOT1_1603(.VSS(VSS),.VDD(VDD),.Y(g7520),.A(g2830));
  NOT NOT1_1604(.VSS(VSS),.VDD(VDD),.Y(g7521),.A(g2200));
  NOT NOT1_1605(.VSS(VSS),.VDD(VDD),.Y(g7522),.A(g2917));
  NOT NOT1_1606(.VSS(VSS),.VDD(VDD),.Y(g7527),.A(g3018));
  NOT NOT1_1607(.VSS(VSS),.VDD(VDD),.Y(g7529),.A(g465));
  NOT NOT1_1608(.VSS(VSS),.VDD(VDD),.Y(g7530),.A(g496));
  NOT NOT1_1609(.VSS(VSS),.VDD(VDD),.Y(g7531),.A(g1180));
  NOT NOT1_1610(.VSS(VSS),.VDD(VDD),.Y(g7532),.A(g1471));
  NOT NOT1_1611(.VSS(VSS),.VDD(VDD),.Y(g7533),.A(g1871));
  NOT NOT1_1612(.VSS(VSS),.VDD(VDD),.Y(g7534),.A(g1832));
  NOT NOT1_1613(.VSS(VSS),.VDD(VDD),.Y(g7535),.A(g2555));
  NOT NOT1_1614(.VSS(VSS),.VDD(VDD),.Y(g7538),.A(g2536));
  NOT NOT1_1615(.VSS(VSS),.VDD(VDD),.Y(g7539),.A(g2528));
  NOT NOT1_1616(.VSS(VSS),.VDD(VDD),.Y(g7540),.A(g1506));
  NOT NOT1_1617(.VSS(VSS),.VDD(VDD),.Y(g7541),.A(g2180));
  NOT NOT1_1618(.VSS(VSS),.VDD(VDD),.Y(g7542),.A(g2883));
  NOT NOT1_1619(.VSS(VSS),.VDD(VDD),.Y(g7545),.A(g2920));
  NOT NOT1_1620(.VSS(VSS),.VDD(VDD),.Y(g7548),.A(g2990));
  NOT NOT1_1621(.VSS(VSS),.VDD(VDD),.Y(g7549),.A(g3028));
  NOT NOT1_1622(.VSS(VSS),.VDD(VDD),.Y(g7553),.A(g3114));
  NOT NOT1_1623(.VSS(VSS),.VDD(VDD),.Y(g7554),.A(g117));
  NOT NOT1_1624(.VSS(VSS),.VDD(VDD),.Y(g7555),.A(g1152));
  NOT NOT1_1625(.VSS(VSS),.VDD(VDD),.Y(g7556),.A(g1183));
  NOT NOT1_1626(.VSS(VSS),.VDD(VDD),.Y(g7557),.A(g1874));
  NOT NOT1_1627(.VSS(VSS),.VDD(VDD),.Y(g7558),.A(g2165));
  NOT NOT1_1628(.VSS(VSS),.VDD(VDD),.Y(g7559),.A(g2565));
  NOT NOT1_1629(.VSS(VSS),.VDD(VDD),.Y(g7560),.A(g2526));
  NOT NOT1_1630(.VSS(VSS),.VDD(VDD),.Y(g7561),.A(g1501));
  NOT NOT1_1631(.VSS(VSS),.VDD(VDD),.Y(g7562),.A(g2888));
  NOT NOT1_1632(.VSS(VSS),.VDD(VDD),.Y(g7566),.A(g2896));
  NOT NOT1_1633(.VSS(VSS),.VDD(VDD),.Y(g7570),.A(g3032));
  NOT NOT1_1634(.VSS(VSS),.VDD(VDD),.Y(g7573),.A(g3120));
  NOT NOT1_1635(.VSS(VSS),.VDD(VDD),.Y(g7574),.A(g3128));
  NOT NOT1_1636(.VSS(VSS),.VDD(VDD),.Y(g7576),.A(g468));
  NOT NOT1_1637(.VSS(VSS),.VDD(VDD),.Y(g7577),.A(g805));
  NOT NOT1_1638(.VSS(VSS),.VDD(VDD),.Y(g7578),.A(g1846));
  NOT NOT1_1639(.VSS(VSS),.VDD(VDD),.Y(g7579),.A(g1877));
  NOT NOT1_1640(.VSS(VSS),.VDD(VDD),.Y(g7580),.A(g2568));
  NOT NOT1_1641(.VSS(VSS),.VDD(VDD),.Y(g7581),.A(g1496));
  NOT NOT1_1642(.VSS(VSS),.VDD(VDD),.Y(g7582),.A(g2185));
  NOT NOT1_1643(.VSS(VSS),.VDD(VDD),.Y(g7583),.A(g2892));
  NOT NOT1_1644(.VSS(VSS),.VDD(VDD),.Y(g7587),.A(g2903));
  NOT NOT1_1645(.VSS(VSS),.VDD(VDD),.Y(g7590),.A(g1155));
  NOT NOT1_1646(.VSS(VSS),.VDD(VDD),.Y(g7591),.A(g1496));
  NOT NOT1_1647(.VSS(VSS),.VDD(VDD),.Y(g7592),.A(g2540));
  NOT NOT1_1648(.VSS(VSS),.VDD(VDD),.Y(g7593),.A(g2571));
  NOT NOT1_1649(.VSS(VSS),.VDD(VDD),.Y(g7594),.A(g2165));
  NOT NOT1_1650(.VSS(VSS),.VDD(VDD),.Y(g7595),.A(g2900));
  NOT NOT1_1651(.VSS(VSS),.VDD(VDD),.Y(g7600),.A(g2908));
  NOT NOT1_1652(.VSS(VSS),.VDD(VDD),.Y(g7603),.A(g3133));
  NOT NOT1_1653(.VSS(VSS),.VDD(VDD),.Y(g7604),.A(g471));
  NOT NOT1_1654(.VSS(VSS),.VDD(VDD),.Y(g7605),.A(g1849));
  NOT NOT1_1655(.VSS(VSS),.VDD(VDD),.Y(g7606),.A(g2190));
  NOT NOT1_1656(.VSS(VSS),.VDD(VDD),.Y(g7607),.A(g2924));
  NOT NOT1_1657(.VSS(VSS),.VDD(VDD),.Y(g7610),.A(g312));
  NOT NOT1_1658(.VSS(VSS),.VDD(VDD),.Y(g7613),.A(g1158));
  NOT NOT1_1659(.VSS(VSS),.VDD(VDD),.Y(g7614),.A(g2543));
  NOT NOT1_1660(.VSS(VSS),.VDD(VDD),.Y(g7615),.A(g3123));
  NOT NOT1_1661(.VSS(VSS),.VDD(VDD),.Y(g7616),.A(g313));
  NOT NOT1_1662(.VSS(VSS),.VDD(VDD),.Y(g7619),.A(g999));
  NOT NOT1_1663(.VSS(VSS),.VDD(VDD),.Y(g7622),.A(g1852));
  NOT NOT1_1664(.VSS(VSS),.VDD(VDD),.Y(g7623),.A(g314));
  NOT NOT1_1665(.VSS(VSS),.VDD(VDD),.Y(g7626),.A(g315));
  NOT NOT1_1666(.VSS(VSS),.VDD(VDD),.Y(g7629),.A(g403));
  NOT NOT1_1667(.VSS(VSS),.VDD(VDD),.Y(g7632),.A(g1000));
  NOT NOT1_1668(.VSS(VSS),.VDD(VDD),.Y(g7635),.A(g1693));
  NOT NOT1_1669(.VSS(VSS),.VDD(VDD),.Y(g7638),.A(g2546));
  NOT NOT1_1670(.VSS(VSS),.VDD(VDD),.Y(g7639),.A(g3094));
  NOT NOT1_1671(.VSS(VSS),.VDD(VDD),.Y(g7642),.A(g3125));
  NOT NOT1_1672(.VSS(VSS),.VDD(VDD),.Y(g7643),.A(g316));
  NOT NOT1_1673(.VSS(VSS),.VDD(VDD),.Y(g7646),.A(g318));
  NOT NOT1_1674(.VSS(VSS),.VDD(VDD),.Y(g7649),.A(g404));
  NOT NOT1_1675(.VSS(VSS),.VDD(VDD),.Y(g7652),.A(g1001));
  NOT NOT1_1676(.VSS(VSS),.VDD(VDD),.Y(g7655),.A(g1002));
  NOT NOT1_1677(.VSS(VSS),.VDD(VDD),.Y(g7658),.A(g1090));
  NOT NOT1_1678(.VSS(VSS),.VDD(VDD),.Y(g7661),.A(g1694));
  NOT NOT1_1679(.VSS(VSS),.VDD(VDD),.Y(g7664),.A(g2387));
  NOT NOT1_1680(.VSS(VSS),.VDD(VDD),.Y(g7667),.A(g3095));
  NOT NOT1_1681(.VSS(VSS),.VDD(VDD),.Y(g7670),.A(g317));
  NOT NOT1_1682(.VSS(VSS),.VDD(VDD),.Y(g7673),.A(g319));
  NOT NOT1_1683(.VSS(VSS),.VDD(VDD),.Y(g7676),.A(g402));
  NOT NOT1_1684(.VSS(VSS),.VDD(VDD),.Y(g7679),.A(g1003));
  NOT NOT1_1685(.VSS(VSS),.VDD(VDD),.Y(g7682),.A(g1005));
  NOT NOT1_1686(.VSS(VSS),.VDD(VDD),.Y(g7685),.A(g1091));
  NOT NOT1_1687(.VSS(VSS),.VDD(VDD),.Y(g7688),.A(g1695));
  NOT NOT1_1688(.VSS(VSS),.VDD(VDD),.Y(g7691),.A(g1696));
  NOT NOT1_1689(.VSS(VSS),.VDD(VDD),.Y(g7694),.A(g1784));
  NOT NOT1_1690(.VSS(VSS),.VDD(VDD),.Y(g7697),.A(g2388));
  NOT NOT1_1691(.VSS(VSS),.VDD(VDD),.Y(g7700),.A(g3096));
  NOT NOT1_1692(.VSS(VSS),.VDD(VDD),.Y(g7703),.A(g320));
  NOT NOT1_1693(.VSS(VSS),.VDD(VDD),.Y(g7706),.A(g1004));
  NOT NOT1_1694(.VSS(VSS),.VDD(VDD),.Y(g7709),.A(g1006));
  NOT NOT1_1695(.VSS(VSS),.VDD(VDD),.Y(g7712),.A(g1089));
  NOT NOT1_1696(.VSS(VSS),.VDD(VDD),.Y(g7715),.A(g1697));
  NOT NOT1_1697(.VSS(VSS),.VDD(VDD),.Y(g7718),.A(g1699));
  NOT NOT1_1698(.VSS(VSS),.VDD(VDD),.Y(g7721),.A(g1785));
  NOT NOT1_1699(.VSS(VSS),.VDD(VDD),.Y(g7724),.A(g2389));
  NOT NOT1_1700(.VSS(VSS),.VDD(VDD),.Y(g7727),.A(g2390));
  NOT NOT1_1701(.VSS(VSS),.VDD(VDD),.Y(g7730),.A(g2478));
  NOT NOT1_1702(.VSS(VSS),.VDD(VDD),.Y(g7733),.A(g1007));
  NOT NOT1_1703(.VSS(VSS),.VDD(VDD),.Y(g7736),.A(g1698));
  NOT NOT1_1704(.VSS(VSS),.VDD(VDD),.Y(g7739),.A(g1700));
  NOT NOT1_1705(.VSS(VSS),.VDD(VDD),.Y(g7742),.A(g1783));
  NOT NOT1_1706(.VSS(VSS),.VDD(VDD),.Y(g7745),.A(g2391));
  NOT NOT1_1707(.VSS(VSS),.VDD(VDD),.Y(g7748),.A(g2393));
  NOT NOT1_1708(.VSS(VSS),.VDD(VDD),.Y(g7751),.A(g2479));
  NOT NOT1_1709(.VSS(VSS),.VDD(VDD),.Y(g7754),.A(g322));
  NOT NOT1_1710(.VSS(VSS),.VDD(VDD),.Y(g7757),.A(g1701));
  NOT NOT1_1711(.VSS(VSS),.VDD(VDD),.Y(g7760),.A(g2392));
  NOT NOT1_1712(.VSS(VSS),.VDD(VDD),.Y(g7763),.A(g2394));
  NOT NOT1_1713(.VSS(VSS),.VDD(VDD),.Y(g7766),.A(g2477));
  NOT NOT1_1714(.VSS(VSS),.VDD(VDD),.Y(g7769),.A(g323));
  NOT NOT1_1715(.VSS(VSS),.VDD(VDD),.Y(g7772),.A(g659));
  NOT NOT1_1716(.VSS(VSS),.VDD(VDD),.Y(g7776),.A(g1009));
  NOT NOT1_1717(.VSS(VSS),.VDD(VDD),.Y(g7779),.A(g2395));
  NOT NOT1_1718(.VSS(VSS),.VDD(VDD),.Y(g7782),.A(g321));
  NOT NOT1_1719(.VSS(VSS),.VDD(VDD),.Y(g7785),.A(g1010));
  NOT NOT1_1720(.VSS(VSS),.VDD(VDD),.Y(g7788),.A(g1345));
  NOT NOT1_1721(.VSS(VSS),.VDD(VDD),.Y(g7792),.A(g1703));
  NOT NOT1_1722(.VSS(VSS),.VDD(VDD),.Y(g7796),.A(g1008));
  NOT NOT1_1723(.VSS(VSS),.VDD(VDD),.Y(g7799),.A(g1704));
  NOT NOT1_1724(.VSS(VSS),.VDD(VDD),.Y(g7802),.A(g2039));
  NOT NOT1_1725(.VSS(VSS),.VDD(VDD),.Y(g7806),.A(g2397));
  NOT NOT1_1726(.VSS(VSS),.VDD(VDD),.Y(g7809),.A(g1702));
  NOT NOT1_1727(.VSS(VSS),.VDD(VDD),.Y(g7812),.A(g2398));
  NOT NOT1_1728(.VSS(VSS),.VDD(VDD),.Y(g7815),.A(g2733));
  NOT NOT1_1729(.VSS(VSS),.VDD(VDD),.Y(g7819),.A(g479));
  NOT NOT1_1730(.VSS(VSS),.VDD(VDD),.Y(g7822),.A(g510));
  NOT NOT1_1731(.VSS(VSS),.VDD(VDD),.Y(g7823),.A(g2396));
  NOT NOT1_1732(.VSS(VSS),.VDD(VDD),.Y(g7826),.A(g2987));
  NOT NOT1_1733(.VSS(VSS),.VDD(VDD),.Y(g7827),.A(g478));
  NOT NOT1_1734(.VSS(VSS),.VDD(VDD),.Y(g7830),.A(g1166));
  NOT NOT1_1735(.VSS(VSS),.VDD(VDD),.Y(g7833),.A(g1196));
  NOT NOT1_1736(.VSS(VSS),.VDD(VDD),.Y(g7834),.A(g2953));
  NOT NOT1_1737(.VSS(VSS),.VDD(VDD),.Y(g7837),.A(g3044));
  NOT NOT1_1738(.VSS(VSS),.VDD(VDD),.Y(g7838),.A(g477));
  NOT NOT1_1739(.VSS(VSS),.VDD(VDD),.Y(g7841),.A(g630));
  NOT NOT1_1740(.VSS(VSS),.VDD(VDD),.Y(g7842),.A(g1165));
  NOT NOT1_1741(.VSS(VSS),.VDD(VDD),.Y(g7845),.A(g1860));
  NOT NOT1_1742(.VSS(VSS),.VDD(VDD),.Y(g7848),.A(g1890));
  NOT NOT1_1743(.VSS(VSS),.VDD(VDD),.Y(g7849),.A(g2956));
  NOT NOT1_1744(.VSS(VSS),.VDD(VDD),.Y(g7852),.A(g2981));
  NOT NOT1_1745(.VSS(VSS),.VDD(VDD),.Y(g7856),.A(g3045));
  NOT NOT1_1746(.VSS(VSS),.VDD(VDD),.Y(g7857),.A(g3055));
  NOT NOT1_1747(.VSS(VSS),.VDD(VDD),.Y(g7858),.A(g1164));
  NOT NOT1_1748(.VSS(VSS),.VDD(VDD),.Y(g7861),.A(g1316));
  NOT NOT1_1749(.VSS(VSS),.VDD(VDD),.Y(g7862),.A(g1859));
  NOT NOT1_1750(.VSS(VSS),.VDD(VDD),.Y(g7865),.A(g2554));
  NOT NOT1_1751(.VSS(VSS),.VDD(VDD),.Y(g7868),.A(g2584));
  NOT NOT1_1752(.VSS(VSS),.VDD(VDD),.Y(g7869),.A(g2959));
  NOT NOT1_1753(.VSS(VSS),.VDD(VDD),.Y(g7872),.A(g2874));
  NOT NOT1_1754(.VSS(VSS),.VDD(VDD),.Y(g7877),.A(g3046));
  NOT NOT1_1755(.VSS(VSS),.VDD(VDD),.Y(g7878),.A(g3056));
  NOT NOT1_1756(.VSS(VSS),.VDD(VDD),.Y(g7879),.A(g3065));
  NOT NOT1_1757(.VSS(VSS),.VDD(VDD),.Y(g7880),.A(g3201));
  NOT NOT1_1758(.VSS(VSS),.VDD(VDD),.Y(g7888),.A(g1858));
  NOT NOT1_1759(.VSS(VSS),.VDD(VDD),.Y(g7891),.A(g2010));
  NOT NOT1_1760(.VSS(VSS),.VDD(VDD),.Y(g7892),.A(g2553));
  NOT NOT1_1761(.VSS(VSS),.VDD(VDD),.Y(g7897),.A(g3047));
  NOT NOT1_1762(.VSS(VSS),.VDD(VDD),.Y(g7898),.A(g3057));
  NOT NOT1_1763(.VSS(VSS),.VDD(VDD),.Y(g7899),.A(g3066));
  NOT NOT1_1764(.VSS(VSS),.VDD(VDD),.Y(g7900),.A(g3075));
  NOT NOT1_1765(.VSS(VSS),.VDD(VDD),.Y(I15222),.A(g3151));
  NOT NOT1_1766(.VSS(VSS),.VDD(VDD),.Y(g7901),.A(I15222));
  NOT NOT1_1767(.VSS(VSS),.VDD(VDD),.Y(g7906),.A(g488));
  NOT NOT1_1768(.VSS(VSS),.VDD(VDD),.Y(I15226),.A(g474));
  NOT NOT1_1769(.VSS(VSS),.VDD(VDD),.Y(g7909),.A(I15226));
  NOT NOT1_1770(.VSS(VSS),.VDD(VDD),.Y(g7910),.A(g474));
  NOT NOT1_1771(.VSS(VSS),.VDD(VDD),.Y(I15230),.A(g499));
  NOT NOT1_1772(.VSS(VSS),.VDD(VDD),.Y(g7911),.A(I15230));
  NOT NOT1_1773(.VSS(VSS),.VDD(VDD),.Y(g7912),.A(g2552));
  NOT NOT1_1774(.VSS(VSS),.VDD(VDD),.Y(g7915),.A(g2704));
  NOT NOT1_1775(.VSS(VSS),.VDD(VDD),.Y(g7916),.A(g2935));
  NOT NOT1_1776(.VSS(VSS),.VDD(VDD),.Y(g7919),.A(g2963));
  NOT NOT1_1777(.VSS(VSS),.VDD(VDD),.Y(g7924),.A(g3048));
  NOT NOT1_1778(.VSS(VSS),.VDD(VDD),.Y(g7925),.A(g3058));
  NOT NOT1_1779(.VSS(VSS),.VDD(VDD),.Y(g7926),.A(g3067));
  NOT NOT1_1780(.VSS(VSS),.VDD(VDD),.Y(g7927),.A(g3076));
  NOT NOT1_1781(.VSS(VSS),.VDD(VDD),.Y(g7928),.A(g3204));
  NOT NOT1_1782(.VSS(VSS),.VDD(VDD),.Y(I15256),.A(g2950));
  NOT NOT1_1783(.VSS(VSS),.VDD(VDD),.Y(g7936),.A(I15256));
  NOT NOT1_1784(.VSS(VSS),.VDD(VDD),.Y(g7949),.A(g165));
  NOT NOT1_1785(.VSS(VSS),.VDD(VDD),.Y(g7950),.A(g142));
  NOT NOT1_1786(.VSS(VSS),.VDD(VDD),.Y(g7953),.A(g487));
  NOT NOT1_1787(.VSS(VSS),.VDD(VDD),.Y(I15262),.A(g481));
  NOT NOT1_1788(.VSS(VSS),.VDD(VDD),.Y(g7956),.A(I15262));
  NOT NOT1_1789(.VSS(VSS),.VDD(VDD),.Y(g7957),.A(g481));
  NOT NOT1_1790(.VSS(VSS),.VDD(VDD),.Y(g7958),.A(g1175));
  NOT NOT1_1791(.VSS(VSS),.VDD(VDD),.Y(I15267),.A(g1161));
  NOT NOT1_1792(.VSS(VSS),.VDD(VDD),.Y(g7961),.A(I15267));
  NOT NOT1_1793(.VSS(VSS),.VDD(VDD),.Y(g7962),.A(g1161));
  NOT NOT1_1794(.VSS(VSS),.VDD(VDD),.Y(I15271),.A(g1186));
  NOT NOT1_1795(.VSS(VSS),.VDD(VDD),.Y(g7963),.A(I15271));
  NOT NOT1_1796(.VSS(VSS),.VDD(VDD),.Y(g7964),.A(g2938));
  NOT NOT1_1797(.VSS(VSS),.VDD(VDD),.Y(g7967),.A(g2966));
  NOT NOT1_1798(.VSS(VSS),.VDD(VDD),.Y(g7971),.A(g3049));
  NOT NOT1_1799(.VSS(VSS),.VDD(VDD),.Y(g7972),.A(g3059));
  NOT NOT1_1800(.VSS(VSS),.VDD(VDD),.Y(g7973),.A(g3068));
  NOT NOT1_1801(.VSS(VSS),.VDD(VDD),.Y(g7974),.A(g3077));
  NOT NOT1_1802(.VSS(VSS),.VDD(VDD),.Y(g7975),.A(g39));
  NOT NOT1_1803(.VSS(VSS),.VDD(VDD),.Y(I15288),.A(g3109));
  NOT NOT1_1804(.VSS(VSS),.VDD(VDD),.Y(g7976),.A(I15288));
  NOT NOT1_1805(.VSS(VSS),.VDD(VDD),.Y(g7989),.A(g3191));
  NOT NOT1_1806(.VSS(VSS),.VDD(VDD),.Y(g7990),.A(g143));
  NOT NOT1_1807(.VSS(VSS),.VDD(VDD),.Y(g7993),.A(g145));
  NOT NOT1_1808(.VSS(VSS),.VDD(VDD),.Y(g7996),.A(g486));
  NOT NOT1_1809(.VSS(VSS),.VDD(VDD),.Y(g7999),.A(g485));
  NOT NOT1_1810(.VSS(VSS),.VDD(VDD),.Y(g8000),.A(g853));
  NOT NOT1_1811(.VSS(VSS),.VDD(VDD),.Y(g8001),.A(g830));
  NOT NOT1_1812(.VSS(VSS),.VDD(VDD),.Y(g8004),.A(g1174));
  NOT NOT1_1813(.VSS(VSS),.VDD(VDD),.Y(I15299),.A(g1168));
  NOT NOT1_1814(.VSS(VSS),.VDD(VDD),.Y(g8007),.A(I15299));
  NOT NOT1_1815(.VSS(VSS),.VDD(VDD),.Y(g8008),.A(g1168));
  NOT NOT1_1816(.VSS(VSS),.VDD(VDD),.Y(g8009),.A(g1869));
  NOT NOT1_1817(.VSS(VSS),.VDD(VDD),.Y(I15304),.A(g1855));
  NOT NOT1_1818(.VSS(VSS),.VDD(VDD),.Y(g8012),.A(I15304));
  NOT NOT1_1819(.VSS(VSS),.VDD(VDD),.Y(g8013),.A(g1855));
  NOT NOT1_1820(.VSS(VSS),.VDD(VDD),.Y(I15308),.A(g1880));
  NOT NOT1_1821(.VSS(VSS),.VDD(VDD),.Y(g8014),.A(I15308));
  NOT NOT1_1822(.VSS(VSS),.VDD(VDD),.Y(g8015),.A(g2941));
  NOT NOT1_1823(.VSS(VSS),.VDD(VDD),.Y(g8018),.A(g2969));
  NOT NOT1_1824(.VSS(VSS),.VDD(VDD),.Y(I15313),.A(g2930));
  NOT NOT1_1825(.VSS(VSS),.VDD(VDD),.Y(g8021),.A(I15313));
  NOT NOT1_1826(.VSS(VSS),.VDD(VDD),.Y(g8022),.A(g2930));
  NOT NOT1_1827(.VSS(VSS),.VDD(VDD),.Y(I15317),.A(g2842));
  NOT NOT1_1828(.VSS(VSS),.VDD(VDD),.Y(g8023),.A(I15317));
  NOT NOT1_1829(.VSS(VSS),.VDD(VDD),.Y(g8024),.A(g2842));
  NOT NOT1_1830(.VSS(VSS),.VDD(VDD),.Y(g8025),.A(g3050));
  NOT NOT1_1831(.VSS(VSS),.VDD(VDD),.Y(g8026),.A(g3060));
  NOT NOT1_1832(.VSS(VSS),.VDD(VDD),.Y(g8027),.A(g3069));
  NOT NOT1_1833(.VSS(VSS),.VDD(VDD),.Y(g8028),.A(g3078));
  NOT NOT1_1834(.VSS(VSS),.VDD(VDD),.Y(g8029),.A(g3083));
  NOT NOT1_1835(.VSS(VSS),.VDD(VDD),.Y(I15326),.A(g3117));
  NOT NOT1_1836(.VSS(VSS),.VDD(VDD),.Y(g8030),.A(I15326));
  NOT NOT1_1837(.VSS(VSS),.VDD(VDD),.Y(I15329),.A(g3117));
  NOT NOT1_1838(.VSS(VSS),.VDD(VDD),.Y(g8031),.A(I15329));
  NOT NOT1_1839(.VSS(VSS),.VDD(VDD),.Y(g8044),.A(g3194));
  NOT NOT1_1840(.VSS(VSS),.VDD(VDD),.Y(g8045),.A(g3207));
  NOT NOT1_1841(.VSS(VSS),.VDD(VDD),.Y(g8053),.A(g141));
  NOT NOT1_1842(.VSS(VSS),.VDD(VDD),.Y(g8056),.A(g146));
  NOT NOT1_1843(.VSS(VSS),.VDD(VDD),.Y(g8059),.A(g148));
  NOT NOT1_1844(.VSS(VSS),.VDD(VDD),.Y(g8062),.A(g169));
  NOT NOT1_1845(.VSS(VSS),.VDD(VDD),.Y(g8065),.A(g831));
  NOT NOT1_1846(.VSS(VSS),.VDD(VDD),.Y(g8068),.A(g833));
  NOT NOT1_1847(.VSS(VSS),.VDD(VDD),.Y(g8071),.A(g1173));
  NOT NOT1_1848(.VSS(VSS),.VDD(VDD),.Y(g8074),.A(g1172));
  NOT NOT1_1849(.VSS(VSS),.VDD(VDD),.Y(g8075),.A(g1547));
  NOT NOT1_1850(.VSS(VSS),.VDD(VDD),.Y(g8076),.A(g1524));
  NOT NOT1_1851(.VSS(VSS),.VDD(VDD),.Y(g8079),.A(g1868));
  NOT NOT1_1852(.VSS(VSS),.VDD(VDD),.Y(I15345),.A(g1862));
  NOT NOT1_1853(.VSS(VSS),.VDD(VDD),.Y(g8082),.A(I15345));
  NOT NOT1_1854(.VSS(VSS),.VDD(VDD),.Y(g8083),.A(g1862));
  NOT NOT1_1855(.VSS(VSS),.VDD(VDD),.Y(g8084),.A(g2563));
  NOT NOT1_1856(.VSS(VSS),.VDD(VDD),.Y(I15350),.A(g2549));
  NOT NOT1_1857(.VSS(VSS),.VDD(VDD),.Y(g8087),.A(I15350));
  NOT NOT1_1858(.VSS(VSS),.VDD(VDD),.Y(g8088),.A(g2549));
  NOT NOT1_1859(.VSS(VSS),.VDD(VDD),.Y(I15354),.A(g2574));
  NOT NOT1_1860(.VSS(VSS),.VDD(VDD),.Y(g8089),.A(I15354));
  NOT NOT1_1861(.VSS(VSS),.VDD(VDD),.Y(g8090),.A(g2944));
  NOT NOT1_1862(.VSS(VSS),.VDD(VDD),.Y(g8093),.A(g2972));
  NOT NOT1_1863(.VSS(VSS),.VDD(VDD),.Y(I15359),.A(g2858));
  NOT NOT1_1864(.VSS(VSS),.VDD(VDD),.Y(g8096),.A(I15359));
  NOT NOT1_1865(.VSS(VSS),.VDD(VDD),.Y(g8097),.A(g2858));
  NOT NOT1_1866(.VSS(VSS),.VDD(VDD),.Y(g8098),.A(g3051));
  NOT NOT1_1867(.VSS(VSS),.VDD(VDD),.Y(g8099),.A(g3061));
  NOT NOT1_1868(.VSS(VSS),.VDD(VDD),.Y(g8100),.A(g3070));
  NOT NOT1_1869(.VSS(VSS),.VDD(VDD),.Y(g8101),.A(g2997));
  NOT NOT1_1870(.VSS(VSS),.VDD(VDD),.Y(g8102),.A(g27));
  NOT NOT1_1871(.VSS(VSS),.VDD(VDD),.Y(g8103),.A(g185));
  NOT NOT1_1872(.VSS(VSS),.VDD(VDD),.Y(I15369),.A(g3129));
  NOT NOT1_1873(.VSS(VSS),.VDD(VDD),.Y(g8106),.A(I15369));
  NOT NOT1_1874(.VSS(VSS),.VDD(VDD),.Y(I15372),.A(g3129));
  NOT NOT1_1875(.VSS(VSS),.VDD(VDD),.Y(g8107),.A(I15372));
  NOT NOT1_1876(.VSS(VSS),.VDD(VDD),.Y(g8120),.A(g3197));
  NOT NOT1_1877(.VSS(VSS),.VDD(VDD),.Y(g8123),.A(g144));
  NOT NOT1_1878(.VSS(VSS),.VDD(VDD),.Y(g8126),.A(g149));
  NOT NOT1_1879(.VSS(VSS),.VDD(VDD),.Y(g8129),.A(g151));
  NOT NOT1_1880(.VSS(VSS),.VDD(VDD),.Y(g8132),.A(g170));
  NOT NOT1_1881(.VSS(VSS),.VDD(VDD),.Y(g8135),.A(g172));
  NOT NOT1_1882(.VSS(VSS),.VDD(VDD),.Y(g8138),.A(g829));
  NOT NOT1_1883(.VSS(VSS),.VDD(VDD),.Y(g8141),.A(g834));
  NOT NOT1_1884(.VSS(VSS),.VDD(VDD),.Y(g8144),.A(g836));
  NOT NOT1_1885(.VSS(VSS),.VDD(VDD),.Y(g8147),.A(g857));
  NOT NOT1_1886(.VSS(VSS),.VDD(VDD),.Y(g8150),.A(g1525));
  NOT NOT1_1887(.VSS(VSS),.VDD(VDD),.Y(g8153),.A(g1527));
  NOT NOT1_1888(.VSS(VSS),.VDD(VDD),.Y(g8156),.A(g1867));
  NOT NOT1_1889(.VSS(VSS),.VDD(VDD),.Y(g8159),.A(g1866));
  NOT NOT1_1890(.VSS(VSS),.VDD(VDD),.Y(g8160),.A(g2241));
  NOT NOT1_1891(.VSS(VSS),.VDD(VDD),.Y(g8161),.A(g2218));
  NOT NOT1_1892(.VSS(VSS),.VDD(VDD),.Y(g8164),.A(g2562));
  NOT NOT1_1893(.VSS(VSS),.VDD(VDD),.Y(I15392),.A(g2556));
  NOT NOT1_1894(.VSS(VSS),.VDD(VDD),.Y(g8167),.A(I15392));
  NOT NOT1_1895(.VSS(VSS),.VDD(VDD),.Y(g8168),.A(g2556));
  NOT NOT1_1896(.VSS(VSS),.VDD(VDD),.Y(g8169),.A(g2947));
  NOT NOT1_1897(.VSS(VSS),.VDD(VDD),.Y(g8172),.A(g2975));
  NOT NOT1_1898(.VSS(VSS),.VDD(VDD),.Y(I15398),.A(g2845));
  NOT NOT1_1899(.VSS(VSS),.VDD(VDD),.Y(g8175),.A(I15398));
  NOT NOT1_1900(.VSS(VSS),.VDD(VDD),.Y(g8176),.A(g2845));
  NOT NOT1_1901(.VSS(VSS),.VDD(VDD),.Y(g8177),.A(g3043));
  NOT NOT1_1902(.VSS(VSS),.VDD(VDD),.Y(g8178),.A(g3052));
  NOT NOT1_1903(.VSS(VSS),.VDD(VDD),.Y(g8179),.A(g3062));
  NOT NOT1_1904(.VSS(VSS),.VDD(VDD),.Y(g8180),.A(g3071));
  NOT NOT1_1905(.VSS(VSS),.VDD(VDD),.Y(g8181),.A(g48));
  NOT NOT1_1906(.VSS(VSS),.VDD(VDD),.Y(g8182),.A(g3198));
  NOT NOT1_1907(.VSS(VSS),.VDD(VDD),.Y(g8183),.A(g3188));
  NOT NOT1_1908(.VSS(VSS),.VDD(VDD),.Y(g8191),.A(g147));
  NOT NOT1_1909(.VSS(VSS),.VDD(VDD),.Y(g8194),.A(g152));
  NOT NOT1_1910(.VSS(VSS),.VDD(VDD),.Y(g8197),.A(g154));
  NOT NOT1_1911(.VSS(VSS),.VDD(VDD),.Y(g8200),.A(g168));
  NOT NOT1_1912(.VSS(VSS),.VDD(VDD),.Y(g8203),.A(g173));
  NOT NOT1_1913(.VSS(VSS),.VDD(VDD),.Y(g8206),.A(g175));
  NOT NOT1_1914(.VSS(VSS),.VDD(VDD),.Y(g8209),.A(g832));
  NOT NOT1_1915(.VSS(VSS),.VDD(VDD),.Y(g8212),.A(g837));
  NOT NOT1_1916(.VSS(VSS),.VDD(VDD),.Y(g8215),.A(g839));
  NOT NOT1_1917(.VSS(VSS),.VDD(VDD),.Y(g8218),.A(g858));
  NOT NOT1_1918(.VSS(VSS),.VDD(VDD),.Y(g8221),.A(g860));
  NOT NOT1_1919(.VSS(VSS),.VDD(VDD),.Y(g8224),.A(g1523));
  NOT NOT1_1920(.VSS(VSS),.VDD(VDD),.Y(g8227),.A(g1528));
  NOT NOT1_1921(.VSS(VSS),.VDD(VDD),.Y(g8230),.A(g1530));
  NOT NOT1_1922(.VSS(VSS),.VDD(VDD),.Y(g8233),.A(g1551));
  NOT NOT1_1923(.VSS(VSS),.VDD(VDD),.Y(g8236),.A(g2219));
  NOT NOT1_1924(.VSS(VSS),.VDD(VDD),.Y(g8239),.A(g2221));
  NOT NOT1_1925(.VSS(VSS),.VDD(VDD),.Y(g8242),.A(g2561));
  NOT NOT1_1926(.VSS(VSS),.VDD(VDD),.Y(g8245),.A(g2560));
  NOT NOT1_1927(.VSS(VSS),.VDD(VDD),.Y(g8246),.A(g2978));
  NOT NOT1_1928(.VSS(VSS),.VDD(VDD),.Y(I15429),.A(g2833));
  NOT NOT1_1929(.VSS(VSS),.VDD(VDD),.Y(g8249),.A(I15429));
  NOT NOT1_1930(.VSS(VSS),.VDD(VDD),.Y(g8250),.A(g2833));
  NOT NOT1_1931(.VSS(VSS),.VDD(VDD),.Y(I15433),.A(g2861));
  NOT NOT1_1932(.VSS(VSS),.VDD(VDD),.Y(g8251),.A(I15433));
  NOT NOT1_1933(.VSS(VSS),.VDD(VDD),.Y(g8252),.A(g2861));
  NOT NOT1_1934(.VSS(VSS),.VDD(VDD),.Y(g8253),.A(g3053));
  NOT NOT1_1935(.VSS(VSS),.VDD(VDD),.Y(g8254),.A(g3063));
  NOT NOT1_1936(.VSS(VSS),.VDD(VDD),.Y(g8255),.A(g3072));
  NOT NOT1_1937(.VSS(VSS),.VDD(VDD),.Y(g8256),.A(g30));
  NOT NOT1_1938(.VSS(VSS),.VDD(VDD),.Y(g8257),.A(g3201));
  NOT NOT1_1939(.VSS(VSS),.VDD(VDD),.Y(I15442),.A(g3235));
  NOT NOT1_1940(.VSS(VSS),.VDD(VDD),.Y(g8258),.A(I15442));
  NOT NOT1_1941(.VSS(VSS),.VDD(VDD),.Y(I15445),.A(g3236));
  NOT NOT1_1942(.VSS(VSS),.VDD(VDD),.Y(g8259),.A(I15445));
  NOT NOT1_1943(.VSS(VSS),.VDD(VDD),.Y(I15448),.A(g3237));
  NOT NOT1_1944(.VSS(VSS),.VDD(VDD),.Y(g8260),.A(I15448));
  NOT NOT1_1945(.VSS(VSS),.VDD(VDD),.Y(I15451),.A(g3238));
  NOT NOT1_1946(.VSS(VSS),.VDD(VDD),.Y(g8261),.A(I15451));
  NOT NOT1_1947(.VSS(VSS),.VDD(VDD),.Y(I15454),.A(g3239));
  NOT NOT1_1948(.VSS(VSS),.VDD(VDD),.Y(g8262),.A(I15454));
  NOT NOT1_1949(.VSS(VSS),.VDD(VDD),.Y(I15457),.A(g3240));
  NOT NOT1_1950(.VSS(VSS),.VDD(VDD),.Y(g8263),.A(I15457));
  NOT NOT1_1951(.VSS(VSS),.VDD(VDD),.Y(I15460),.A(g3241));
  NOT NOT1_1952(.VSS(VSS),.VDD(VDD),.Y(g8264),.A(I15460));
  NOT NOT1_1953(.VSS(VSS),.VDD(VDD),.Y(I15463),.A(g3242));
  NOT NOT1_1954(.VSS(VSS),.VDD(VDD),.Y(g8265),.A(I15463));
  NOT NOT1_1955(.VSS(VSS),.VDD(VDD),.Y(I15466),.A(g3243));
  NOT NOT1_1956(.VSS(VSS),.VDD(VDD),.Y(g8266),.A(I15466));
  NOT NOT1_1957(.VSS(VSS),.VDD(VDD),.Y(I15469),.A(g3244));
  NOT NOT1_1958(.VSS(VSS),.VDD(VDD),.Y(g8267),.A(I15469));
  NOT NOT1_1959(.VSS(VSS),.VDD(VDD),.Y(I15472),.A(g3245));
  NOT NOT1_1960(.VSS(VSS),.VDD(VDD),.Y(g8268),.A(I15472));
  NOT NOT1_1961(.VSS(VSS),.VDD(VDD),.Y(I15475),.A(g3246));
  NOT NOT1_1962(.VSS(VSS),.VDD(VDD),.Y(g8269),.A(I15475));
  NOT NOT1_1963(.VSS(VSS),.VDD(VDD),.Y(I15478),.A(g3247));
  NOT NOT1_1964(.VSS(VSS),.VDD(VDD),.Y(g8270),.A(I15478));
  NOT NOT1_1965(.VSS(VSS),.VDD(VDD),.Y(I15481),.A(g3248));
  NOT NOT1_1966(.VSS(VSS),.VDD(VDD),.Y(g8271),.A(I15481));
  NOT NOT1_1967(.VSS(VSS),.VDD(VDD),.Y(I15484),.A(g3249));
  NOT NOT1_1968(.VSS(VSS),.VDD(VDD),.Y(g8272),.A(I15484));
  NOT NOT1_1969(.VSS(VSS),.VDD(VDD),.Y(I15487),.A(g3250));
  NOT NOT1_1970(.VSS(VSS),.VDD(VDD),.Y(g8273),.A(I15487));
  NOT NOT1_1971(.VSS(VSS),.VDD(VDD),.Y(I15490),.A(g3251));
  NOT NOT1_1972(.VSS(VSS),.VDD(VDD),.Y(g8274),.A(I15490));
  NOT NOT1_1973(.VSS(VSS),.VDD(VDD),.Y(I15493),.A(g3252));
  NOT NOT1_1974(.VSS(VSS),.VDD(VDD),.Y(g8275),.A(I15493));
  NOT NOT1_1975(.VSS(VSS),.VDD(VDD),.Y(g8276),.A(g3253));
  NOT NOT1_1976(.VSS(VSS),.VDD(VDD),.Y(g8277),.A(g3305));
  NOT NOT1_1977(.VSS(VSS),.VDD(VDD),.Y(g8278),.A(g3337));
  NOT NOT1_1978(.VSS(VSS),.VDD(VDD),.Y(I15499),.A(g7911));
  NOT NOT1_1979(.VSS(VSS),.VDD(VDD),.Y(g8284),.A(I15499));
  NOT NOT1_1980(.VSS(VSS),.VDD(VDD),.Y(g8285),.A(g3365));
  NOT NOT1_1981(.VSS(VSS),.VDD(VDD),.Y(g8286),.A(g3461));
  NOT NOT1_1982(.VSS(VSS),.VDD(VDD),.Y(g8287),.A(g3493));
  NOT NOT1_1983(.VSS(VSS),.VDD(VDD),.Y(I15505),.A(g7963));
  NOT NOT1_1984(.VSS(VSS),.VDD(VDD),.Y(g8293),.A(I15505));
  NOT NOT1_1985(.VSS(VSS),.VDD(VDD),.Y(g8294),.A(g3521));
  NOT NOT1_1986(.VSS(VSS),.VDD(VDD),.Y(g8295),.A(g3617));
  NOT NOT1_1987(.VSS(VSS),.VDD(VDD),.Y(g8296),.A(g3649));
  NOT NOT1_1988(.VSS(VSS),.VDD(VDD),.Y(I15511),.A(g8014));
  NOT NOT1_1989(.VSS(VSS),.VDD(VDD),.Y(g8302),.A(I15511));
  NOT NOT1_1990(.VSS(VSS),.VDD(VDD),.Y(g8303),.A(g3677));
  NOT NOT1_1991(.VSS(VSS),.VDD(VDD),.Y(g8304),.A(g3773));
  NOT NOT1_1992(.VSS(VSS),.VDD(VDD),.Y(g8305),.A(g3805));
  NOT NOT1_1993(.VSS(VSS),.VDD(VDD),.Y(I15517),.A(g8089));
  NOT NOT1_1994(.VSS(VSS),.VDD(VDD),.Y(g8311),.A(I15517));
  NOT NOT1_1995(.VSS(VSS),.VDD(VDD),.Y(g8312),.A(g3833));
  NOT NOT1_1996(.VSS(VSS),.VDD(VDD),.Y(g8313),.A(g3897));
  NOT NOT1_1997(.VSS(VSS),.VDD(VDD),.Y(g8317),.A(g3919));
  NOT NOT1_1998(.VSS(VSS),.VDD(VDD),.Y(I15523),.A(g3254));
  NOT NOT1_1999(.VSS(VSS),.VDD(VDD),.Y(g8321),.A(I15523));
  NOT NOT1_2000(.VSS(VSS),.VDD(VDD),.Y(I15526),.A(g6314));
  NOT NOT1_2001(.VSS(VSS),.VDD(VDD),.Y(g8324),.A(I15526));
  NOT NOT1_2002(.VSS(VSS),.VDD(VDD),.Y(I15532),.A(g3410));
  NOT NOT1_2003(.VSS(VSS),.VDD(VDD),.Y(g8330),.A(I15532));
  NOT NOT1_2004(.VSS(VSS),.VDD(VDD),.Y(I15535),.A(g6519));
  NOT NOT1_2005(.VSS(VSS),.VDD(VDD),.Y(g8333),.A(I15535));
  NOT NOT1_2006(.VSS(VSS),.VDD(VDD),.Y(I15538),.A(g6369));
  NOT NOT1_2007(.VSS(VSS),.VDD(VDD),.Y(g8336),.A(I15538));
  NOT NOT1_2008(.VSS(VSS),.VDD(VDD),.Y(I15543),.A(g3410));
  NOT NOT1_2009(.VSS(VSS),.VDD(VDD),.Y(g8341),.A(I15543));
  NOT NOT1_2010(.VSS(VSS),.VDD(VDD),.Y(I15546),.A(g6783));
  NOT NOT1_2011(.VSS(VSS),.VDD(VDD),.Y(g8344),.A(I15546));
  NOT NOT1_2012(.VSS(VSS),.VDD(VDD),.Y(I15549),.A(g6574));
  NOT NOT1_2013(.VSS(VSS),.VDD(VDD),.Y(g8347),.A(I15549));
  NOT NOT1_2014(.VSS(VSS),.VDD(VDD),.Y(I15553),.A(g3566));
  NOT NOT1_2015(.VSS(VSS),.VDD(VDD),.Y(g8351),.A(I15553));
  NOT NOT1_2016(.VSS(VSS),.VDD(VDD),.Y(I15556),.A(g6783));
  NOT NOT1_2017(.VSS(VSS),.VDD(VDD),.Y(g8354),.A(I15556));
  NOT NOT1_2018(.VSS(VSS),.VDD(VDD),.Y(I15559),.A(g7015));
  NOT NOT1_2019(.VSS(VSS),.VDD(VDD),.Y(g8357),.A(I15559));
  NOT NOT1_2020(.VSS(VSS),.VDD(VDD),.Y(I15562),.A(g5778));
  NOT NOT1_2021(.VSS(VSS),.VDD(VDD),.Y(g8360),.A(I15562));
  NOT NOT1_2022(.VSS(VSS),.VDD(VDD),.Y(I15565),.A(g6838));
  NOT NOT1_2023(.VSS(VSS),.VDD(VDD),.Y(g8363),.A(I15565));
  NOT NOT1_2024(.VSS(VSS),.VDD(VDD),.Y(I15568),.A(g3722));
  NOT NOT1_2025(.VSS(VSS),.VDD(VDD),.Y(g8366),.A(I15568));
  NOT NOT1_2026(.VSS(VSS),.VDD(VDD),.Y(I15571),.A(g7085));
  NOT NOT1_2027(.VSS(VSS),.VDD(VDD),.Y(g8369),.A(I15571));
  NOT NOT1_2028(.VSS(VSS),.VDD(VDD),.Y(I15574),.A(g6838));
  NOT NOT1_2029(.VSS(VSS),.VDD(VDD),.Y(g8372),.A(I15574));
  NOT NOT1_2030(.VSS(VSS),.VDD(VDD),.Y(I15577),.A(g7265));
  NOT NOT1_2031(.VSS(VSS),.VDD(VDD),.Y(g8375),.A(I15577));
  NOT NOT1_2032(.VSS(VSS),.VDD(VDD),.Y(I15580),.A(g5837));
  NOT NOT1_2033(.VSS(VSS),.VDD(VDD),.Y(g8378),.A(I15580));
  NOT NOT1_2034(.VSS(VSS),.VDD(VDD),.Y(I15584),.A(g3254));
  NOT NOT1_2035(.VSS(VSS),.VDD(VDD),.Y(g8382),.A(I15584));
  NOT NOT1_2036(.VSS(VSS),.VDD(VDD),.Y(I15590),.A(g3410));
  NOT NOT1_2037(.VSS(VSS),.VDD(VDD),.Y(g8388),.A(I15590));
  NOT NOT1_2038(.VSS(VSS),.VDD(VDD),.Y(I15593),.A(g6519));
  NOT NOT1_2039(.VSS(VSS),.VDD(VDD),.Y(g8391),.A(I15593));
  NOT NOT1_2040(.VSS(VSS),.VDD(VDD),.Y(I15599),.A(g3566));
  NOT NOT1_2041(.VSS(VSS),.VDD(VDD),.Y(g8397),.A(I15599));
  NOT NOT1_2042(.VSS(VSS),.VDD(VDD),.Y(I15602),.A(g6783));
  NOT NOT1_2043(.VSS(VSS),.VDD(VDD),.Y(g8400),.A(I15602));
  NOT NOT1_2044(.VSS(VSS),.VDD(VDD),.Y(I15605),.A(g6574));
  NOT NOT1_2045(.VSS(VSS),.VDD(VDD),.Y(g8403),.A(I15605));
  NOT NOT1_2046(.VSS(VSS),.VDD(VDD),.Y(I15610),.A(g3566));
  NOT NOT1_2047(.VSS(VSS),.VDD(VDD),.Y(g8408),.A(I15610));
  NOT NOT1_2048(.VSS(VSS),.VDD(VDD),.Y(I15613),.A(g7085));
  NOT NOT1_2049(.VSS(VSS),.VDD(VDD),.Y(g8411),.A(I15613));
  NOT NOT1_2050(.VSS(VSS),.VDD(VDD),.Y(I15616),.A(g6838));
  NOT NOT1_2051(.VSS(VSS),.VDD(VDD),.Y(g8414),.A(I15616));
  NOT NOT1_2052(.VSS(VSS),.VDD(VDD),.Y(I15620),.A(g3722));
  NOT NOT1_2053(.VSS(VSS),.VDD(VDD),.Y(g8418),.A(I15620));
  NOT NOT1_2054(.VSS(VSS),.VDD(VDD),.Y(I15623),.A(g7085));
  NOT NOT1_2055(.VSS(VSS),.VDD(VDD),.Y(g8421),.A(I15623));
  NOT NOT1_2056(.VSS(VSS),.VDD(VDD),.Y(I15626),.A(g7265));
  NOT NOT1_2057(.VSS(VSS),.VDD(VDD),.Y(g8424),.A(I15626));
  NOT NOT1_2058(.VSS(VSS),.VDD(VDD),.Y(I15629),.A(g5837));
  NOT NOT1_2059(.VSS(VSS),.VDD(VDD),.Y(g8427),.A(I15629));
  NOT NOT1_2060(.VSS(VSS),.VDD(VDD),.Y(I15636),.A(g3410));
  NOT NOT1_2061(.VSS(VSS),.VDD(VDD),.Y(g8434),.A(I15636));
  NOT NOT1_2062(.VSS(VSS),.VDD(VDD),.Y(I15642),.A(g3566));
  NOT NOT1_2063(.VSS(VSS),.VDD(VDD),.Y(g8440),.A(I15642));
  NOT NOT1_2064(.VSS(VSS),.VDD(VDD),.Y(I15645),.A(g6783));
  NOT NOT1_2065(.VSS(VSS),.VDD(VDD),.Y(g8443),.A(I15645));
  NOT NOT1_2066(.VSS(VSS),.VDD(VDD),.Y(I15651),.A(g3722));
  NOT NOT1_2067(.VSS(VSS),.VDD(VDD),.Y(g8449),.A(I15651));
  NOT NOT1_2068(.VSS(VSS),.VDD(VDD),.Y(I15654),.A(g7085));
  NOT NOT1_2069(.VSS(VSS),.VDD(VDD),.Y(g8452),.A(I15654));
  NOT NOT1_2070(.VSS(VSS),.VDD(VDD),.Y(I15657),.A(g6838));
  NOT NOT1_2071(.VSS(VSS),.VDD(VDD),.Y(g8455),.A(I15657));
  NOT NOT1_2072(.VSS(VSS),.VDD(VDD),.Y(I15662),.A(g3722));
  NOT NOT1_2073(.VSS(VSS),.VDD(VDD),.Y(g8460),.A(I15662));
  NOT NOT1_2074(.VSS(VSS),.VDD(VDD),.Y(I15671),.A(g3566));
  NOT NOT1_2075(.VSS(VSS),.VDD(VDD),.Y(g8469),.A(I15671));
  NOT NOT1_2076(.VSS(VSS),.VDD(VDD),.Y(I15677),.A(g3722));
  NOT NOT1_2077(.VSS(VSS),.VDD(VDD),.Y(g8475),.A(I15677));
  NOT NOT1_2078(.VSS(VSS),.VDD(VDD),.Y(I15680),.A(g7085));
  NOT NOT1_2079(.VSS(VSS),.VDD(VDD),.Y(g8478),.A(I15680));
  NOT NOT1_2080(.VSS(VSS),.VDD(VDD),.Y(I15696),.A(g3722));
  NOT NOT1_2081(.VSS(VSS),.VDD(VDD),.Y(g8494),.A(I15696));
  NOT NOT1_2082(.VSS(VSS),.VDD(VDD),.Y(g8514),.A(g6139));
  NOT NOT1_2083(.VSS(VSS),.VDD(VDD),.Y(g8530),.A(g6156));
  NOT NOT1_2084(.VSS(VSS),.VDD(VDD),.Y(g8568),.A(g6230));
  NOT NOT1_2085(.VSS(VSS),.VDD(VDD),.Y(I15771),.A(g6000));
  NOT NOT1_2086(.VSS(VSS),.VDD(VDD),.Y(g8569),.A(I15771));
  NOT NOT1_2087(.VSS(VSS),.VDD(VDD),.Y(I15779),.A(g6000));
  NOT NOT1_2088(.VSS(VSS),.VDD(VDD),.Y(g8575),.A(I15779));
  NOT NOT1_2089(.VSS(VSS),.VDD(VDD),.Y(I15784),.A(g6000));
  NOT NOT1_2090(.VSS(VSS),.VDD(VDD),.Y(g8578),.A(I15784));
  NOT NOT1_2091(.VSS(VSS),.VDD(VDD),.Y(I15787),.A(g6000));
  NOT NOT1_2092(.VSS(VSS),.VDD(VDD),.Y(g8579),.A(I15787));
  NOT NOT1_2093(.VSS(VSS),.VDD(VDD),.Y(g8580),.A(g6281));
  NOT NOT1_2094(.VSS(VSS),.VDD(VDD),.Y(g8587),.A(g6418));
  NOT NOT1_2095(.VSS(VSS),.VDD(VDD),.Y(g8594),.A(g6623));
  NOT NOT1_2096(.VSS(VSS),.VDD(VDD),.Y(I15794),.A(g3338));
  NOT NOT1_2097(.VSS(VSS),.VDD(VDD),.Y(g8602),.A(I15794));
  NOT NOT1_2098(.VSS(VSS),.VDD(VDD),.Y(g8605),.A(g6887));
  NOT NOT1_2099(.VSS(VSS),.VDD(VDD),.Y(I15800),.A(g3494));
  NOT NOT1_2100(.VSS(VSS),.VDD(VDD),.Y(g8614),.A(I15800));
  NOT NOT1_2101(.VSS(VSS),.VDD(VDD),.Y(I15803),.A(g8107));
  NOT NOT1_2102(.VSS(VSS),.VDD(VDD),.Y(g8617),.A(I15803));
  NOT NOT1_2103(.VSS(VSS),.VDD(VDD),.Y(I15806),.A(g5550));
  NOT NOT1_2104(.VSS(VSS),.VDD(VDD),.Y(g8620),.A(I15806));
  NOT NOT1_2105(.VSS(VSS),.VDD(VDD),.Y(I15810),.A(g3338));
  NOT NOT1_2106(.VSS(VSS),.VDD(VDD),.Y(g8622),.A(I15810));
  NOT NOT1_2107(.VSS(VSS),.VDD(VDD),.Y(I15815),.A(g3650));
  NOT NOT1_2108(.VSS(VSS),.VDD(VDD),.Y(g8627),.A(I15815));
  NOT NOT1_2109(.VSS(VSS),.VDD(VDD),.Y(I15818),.A(g5596));
  NOT NOT1_2110(.VSS(VSS),.VDD(VDD),.Y(g8630),.A(I15818));
  NOT NOT1_2111(.VSS(VSS),.VDD(VDD),.Y(I15822),.A(g3494));
  NOT NOT1_2112(.VSS(VSS),.VDD(VDD),.Y(g8632),.A(I15822));
  NOT NOT1_2113(.VSS(VSS),.VDD(VDD),.Y(I15827),.A(g3806));
  NOT NOT1_2114(.VSS(VSS),.VDD(VDD),.Y(g8637),.A(I15827));
  NOT NOT1_2115(.VSS(VSS),.VDD(VDD),.Y(I15830),.A(g8031));
  NOT NOT1_2116(.VSS(VSS),.VDD(VDD),.Y(g8640),.A(I15830));
  NOT NOT1_2117(.VSS(VSS),.VDD(VDD),.Y(I15833),.A(g3338));
  NOT NOT1_2118(.VSS(VSS),.VDD(VDD),.Y(g8643),.A(I15833));
  NOT NOT1_2119(.VSS(VSS),.VDD(VDD),.Y(I15836),.A(g3366));
  NOT NOT1_2120(.VSS(VSS),.VDD(VDD),.Y(g8646),.A(I15836));
  NOT NOT1_2121(.VSS(VSS),.VDD(VDD),.Y(I15839),.A(g5613));
  NOT NOT1_2122(.VSS(VSS),.VDD(VDD),.Y(g8649),.A(I15839));
  NOT NOT1_2123(.VSS(VSS),.VDD(VDD),.Y(I15843),.A(g3650));
  NOT NOT1_2124(.VSS(VSS),.VDD(VDD),.Y(g8651),.A(I15843));
  NOT NOT1_2125(.VSS(VSS),.VDD(VDD),.Y(I15847),.A(g3878));
  NOT NOT1_2126(.VSS(VSS),.VDD(VDD),.Y(g8655),.A(I15847));
  NOT NOT1_2127(.VSS(VSS),.VDD(VDD),.Y(I15850),.A(g5627));
  NOT NOT1_2128(.VSS(VSS),.VDD(VDD),.Y(g8658),.A(I15850));
  NOT NOT1_2129(.VSS(VSS),.VDD(VDD),.Y(I15853),.A(g3494));
  NOT NOT1_2130(.VSS(VSS),.VDD(VDD),.Y(g8659),.A(I15853));
  NOT NOT1_2131(.VSS(VSS),.VDD(VDD),.Y(I15856),.A(g3522));
  NOT NOT1_2132(.VSS(VSS),.VDD(VDD),.Y(g8662),.A(I15856));
  NOT NOT1_2133(.VSS(VSS),.VDD(VDD),.Y(I15859),.A(g5638));
  NOT NOT1_2134(.VSS(VSS),.VDD(VDD),.Y(g8665),.A(I15859));
  NOT NOT1_2135(.VSS(VSS),.VDD(VDD),.Y(I15863),.A(g3806));
  NOT NOT1_2136(.VSS(VSS),.VDD(VDD),.Y(g8667),.A(I15863));
  NOT NOT1_2137(.VSS(VSS),.VDD(VDD),.Y(I15866),.A(g3878));
  NOT NOT1_2138(.VSS(VSS),.VDD(VDD),.Y(g8670),.A(I15866));
  NOT NOT1_2139(.VSS(VSS),.VDD(VDD),.Y(I15869),.A(g7976));
  NOT NOT1_2140(.VSS(VSS),.VDD(VDD),.Y(g8673),.A(I15869));
  NOT NOT1_2141(.VSS(VSS),.VDD(VDD),.Y(I15873),.A(g5655));
  NOT NOT1_2142(.VSS(VSS),.VDD(VDD),.Y(g8677),.A(I15873));
  NOT NOT1_2143(.VSS(VSS),.VDD(VDD),.Y(I15876),.A(g3650));
  NOT NOT1_2144(.VSS(VSS),.VDD(VDD),.Y(g8678),.A(I15876));
  NOT NOT1_2145(.VSS(VSS),.VDD(VDD),.Y(I15879),.A(g3678));
  NOT NOT1_2146(.VSS(VSS),.VDD(VDD),.Y(g8681),.A(I15879));
  NOT NOT1_2147(.VSS(VSS),.VDD(VDD),.Y(I15882),.A(g3878));
  NOT NOT1_2148(.VSS(VSS),.VDD(VDD),.Y(g8684),.A(I15882));
  NOT NOT1_2149(.VSS(VSS),.VDD(VDD),.Y(I15887),.A(g5693));
  NOT NOT1_2150(.VSS(VSS),.VDD(VDD),.Y(g8689),.A(I15887));
  NOT NOT1_2151(.VSS(VSS),.VDD(VDD),.Y(I15890),.A(g3806));
  NOT NOT1_2152(.VSS(VSS),.VDD(VDD),.Y(g8690),.A(I15890));
  NOT NOT1_2153(.VSS(VSS),.VDD(VDD),.Y(I15893),.A(g3834));
  NOT NOT1_2154(.VSS(VSS),.VDD(VDD),.Y(g8693),.A(I15893));
  NOT NOT1_2155(.VSS(VSS),.VDD(VDD),.Y(I15896),.A(g3878));
  NOT NOT1_2156(.VSS(VSS),.VDD(VDD),.Y(g8696),.A(I15896));
  NOT NOT1_2157(.VSS(VSS),.VDD(VDD),.Y(I15899),.A(g5626));
  NOT NOT1_2158(.VSS(VSS),.VDD(VDD),.Y(g8699),.A(I15899));
  NOT NOT1_2159(.VSS(VSS),.VDD(VDD),.Y(I15902),.A(g6486));
  NOT NOT1_2160(.VSS(VSS),.VDD(VDD),.Y(g8700),.A(I15902));
  NOT NOT1_2161(.VSS(VSS),.VDD(VDD),.Y(I15909),.A(g5745));
  NOT NOT1_2162(.VSS(VSS),.VDD(VDD),.Y(g8707),.A(I15909));
  NOT NOT1_2163(.VSS(VSS),.VDD(VDD),.Y(I15912),.A(g3878));
  NOT NOT1_2164(.VSS(VSS),.VDD(VDD),.Y(g8708),.A(I15912));
  NOT NOT1_2165(.VSS(VSS),.VDD(VDD),.Y(I15915),.A(g3878));
  NOT NOT1_2166(.VSS(VSS),.VDD(VDD),.Y(g8711),.A(I15915));
  NOT NOT1_2167(.VSS(VSS),.VDD(VDD),.Y(I15918),.A(g6643));
  NOT NOT1_2168(.VSS(VSS),.VDD(VDD),.Y(g8714),.A(I15918));
  NOT NOT1_2169(.VSS(VSS),.VDD(VDD),.Y(I15922),.A(g5654));
  NOT NOT1_2170(.VSS(VSS),.VDD(VDD),.Y(g8718),.A(I15922));
  NOT NOT1_2171(.VSS(VSS),.VDD(VDD),.Y(I15925),.A(g6751));
  NOT NOT1_2172(.VSS(VSS),.VDD(VDD),.Y(g8719),.A(I15925));
  NOT NOT1_2173(.VSS(VSS),.VDD(VDD),.Y(I15932),.A(g5423));
  NOT NOT1_2174(.VSS(VSS),.VDD(VDD),.Y(g8726),.A(I15932));
  NOT NOT1_2175(.VSS(VSS),.VDD(VDD),.Y(I15935),.A(g3878));
  NOT NOT1_2176(.VSS(VSS),.VDD(VDD),.Y(g8745),.A(I15935));
  NOT NOT1_2177(.VSS(VSS),.VDD(VDD),.Y(I15938),.A(g3338));
  NOT NOT1_2178(.VSS(VSS),.VDD(VDD),.Y(g8748),.A(I15938));
  NOT NOT1_2179(.VSS(VSS),.VDD(VDD),.Y(I15942),.A(g6945));
  NOT NOT1_2180(.VSS(VSS),.VDD(VDD),.Y(g8752),.A(I15942));
  NOT NOT1_2181(.VSS(VSS),.VDD(VDD),.Y(I15946),.A(g5692));
  NOT NOT1_2182(.VSS(VSS),.VDD(VDD),.Y(g8756),.A(I15946));
  NOT NOT1_2183(.VSS(VSS),.VDD(VDD),.Y(I15949),.A(g7053));
  NOT NOT1_2184(.VSS(VSS),.VDD(VDD),.Y(g8757),.A(I15949));
  NOT NOT1_2185(.VSS(VSS),.VDD(VDD),.Y(I15955),.A(g3878));
  NOT NOT1_2186(.VSS(VSS),.VDD(VDD),.Y(g8763),.A(I15955));
  NOT NOT1_2187(.VSS(VSS),.VDD(VDD),.Y(I15958),.A(g3878));
  NOT NOT1_2188(.VSS(VSS),.VDD(VDD),.Y(g8766),.A(I15958));
  NOT NOT1_2189(.VSS(VSS),.VDD(VDD),.Y(I15961),.A(g6051));
  NOT NOT1_2190(.VSS(VSS),.VDD(VDD),.Y(g8769),.A(I15961));
  NOT NOT1_2191(.VSS(VSS),.VDD(VDD),.Y(I15964),.A(g7554));
  NOT NOT1_2192(.VSS(VSS),.VDD(VDD),.Y(g8770),.A(I15964));
  NOT NOT1_2193(.VSS(VSS),.VDD(VDD),.Y(I15967),.A(g3494));
  NOT NOT1_2194(.VSS(VSS),.VDD(VDD),.Y(g8771),.A(I15967));
  NOT NOT1_2195(.VSS(VSS),.VDD(VDD),.Y(I15971),.A(g7195));
  NOT NOT1_2196(.VSS(VSS),.VDD(VDD),.Y(g8775),.A(I15971));
  NOT NOT1_2197(.VSS(VSS),.VDD(VDD),.Y(I15975),.A(g5744));
  NOT NOT1_2198(.VSS(VSS),.VDD(VDD),.Y(g8779),.A(I15975));
  NOT NOT1_2199(.VSS(VSS),.VDD(VDD),.Y(I15978),.A(g7303));
  NOT NOT1_2200(.VSS(VSS),.VDD(VDD),.Y(g8780),.A(I15978));
  NOT NOT1_2201(.VSS(VSS),.VDD(VDD),.Y(I15983),.A(g3878));
  NOT NOT1_2202(.VSS(VSS),.VDD(VDD),.Y(g8785),.A(I15983));
  NOT NOT1_2203(.VSS(VSS),.VDD(VDD),.Y(I15986),.A(g3878));
  NOT NOT1_2204(.VSS(VSS),.VDD(VDD),.Y(g8788),.A(I15986));
  NOT NOT1_2205(.VSS(VSS),.VDD(VDD),.Y(I15989),.A(g6053));
  NOT NOT1_2206(.VSS(VSS),.VDD(VDD),.Y(g8791),.A(I15989));
  NOT NOT1_2207(.VSS(VSS),.VDD(VDD),.Y(I15992),.A(g6055));
  NOT NOT1_2208(.VSS(VSS),.VDD(VDD),.Y(g8792),.A(I15992));
  NOT NOT1_2209(.VSS(VSS),.VDD(VDD),.Y(I15995),.A(g7577));
  NOT NOT1_2210(.VSS(VSS),.VDD(VDD),.Y(g8793),.A(I15995));
  NOT NOT1_2211(.VSS(VSS),.VDD(VDD),.Y(I15998),.A(g3650));
  NOT NOT1_2212(.VSS(VSS),.VDD(VDD),.Y(g8794),.A(I15998));
  NOT NOT1_2213(.VSS(VSS),.VDD(VDD),.Y(I16002),.A(g7391));
  NOT NOT1_2214(.VSS(VSS),.VDD(VDD),.Y(g8798),.A(I16002));
  NOT NOT1_2215(.VSS(VSS),.VDD(VDD),.Y(I16006),.A(g3878));
  NOT NOT1_2216(.VSS(VSS),.VDD(VDD),.Y(g8802),.A(I16006));
  NOT NOT1_2217(.VSS(VSS),.VDD(VDD),.Y(I16009),.A(g3878));
  NOT NOT1_2218(.VSS(VSS),.VDD(VDD),.Y(g8805),.A(I16009));
  NOT NOT1_2219(.VSS(VSS),.VDD(VDD),.Y(I16012),.A(g5390));
  NOT NOT1_2220(.VSS(VSS),.VDD(VDD),.Y(g8808),.A(I16012));
  NOT NOT1_2221(.VSS(VSS),.VDD(VDD),.Y(I16015),.A(g6056));
  NOT NOT1_2222(.VSS(VSS),.VDD(VDD),.Y(g8809),.A(I16015));
  NOT NOT1_2223(.VSS(VSS),.VDD(VDD),.Y(I16018),.A(g6058));
  NOT NOT1_2224(.VSS(VSS),.VDD(VDD),.Y(g8810),.A(I16018));
  NOT NOT1_2225(.VSS(VSS),.VDD(VDD),.Y(I16021),.A(g6060));
  NOT NOT1_2226(.VSS(VSS),.VDD(VDD),.Y(g8811),.A(I16021));
  NOT NOT1_2227(.VSS(VSS),.VDD(VDD),.Y(I16024),.A(g7591));
  NOT NOT1_2228(.VSS(VSS),.VDD(VDD),.Y(g8812),.A(I16024));
  NOT NOT1_2229(.VSS(VSS),.VDD(VDD),.Y(I16027),.A(g3806));
  NOT NOT1_2230(.VSS(VSS),.VDD(VDD),.Y(g8813),.A(I16027));
  NOT NOT1_2231(.VSS(VSS),.VDD(VDD),.Y(I16031),.A(g3878));
  NOT NOT1_2232(.VSS(VSS),.VDD(VDD),.Y(g8817),.A(I16031));
  NOT NOT1_2233(.VSS(VSS),.VDD(VDD),.Y(I16034),.A(g5396));
  NOT NOT1_2234(.VSS(VSS),.VDD(VDD),.Y(g8820),.A(I16034));
  NOT NOT1_2235(.VSS(VSS),.VDD(VDD),.Y(I16037),.A(g6061));
  NOT NOT1_2236(.VSS(VSS),.VDD(VDD),.Y(g8821),.A(I16037));
  NOT NOT1_2237(.VSS(VSS),.VDD(VDD),.Y(g8822),.A(g4602));
  NOT NOT1_2238(.VSS(VSS),.VDD(VDD),.Y(I16041),.A(g6486));
  NOT NOT1_2239(.VSS(VSS),.VDD(VDD),.Y(g8823),.A(I16041));
  NOT NOT1_2240(.VSS(VSS),.VDD(VDD),.Y(I16044),.A(g5397));
  NOT NOT1_2241(.VSS(VSS),.VDD(VDD),.Y(g8824),.A(I16044));
  NOT NOT1_2242(.VSS(VSS),.VDD(VDD),.Y(I16047),.A(g6063));
  NOT NOT1_2243(.VSS(VSS),.VDD(VDD),.Y(g8825),.A(I16047));
  NOT NOT1_2244(.VSS(VSS),.VDD(VDD),.Y(I16050),.A(g6065));
  NOT NOT1_2245(.VSS(VSS),.VDD(VDD),.Y(g8826),.A(I16050));
  NOT NOT1_2246(.VSS(VSS),.VDD(VDD),.Y(I16053),.A(g6067));
  NOT NOT1_2247(.VSS(VSS),.VDD(VDD),.Y(g8827),.A(I16053));
  NOT NOT1_2248(.VSS(VSS),.VDD(VDD),.Y(I16056),.A(g7606));
  NOT NOT1_2249(.VSS(VSS),.VDD(VDD),.Y(g8828),.A(I16056));
  NOT NOT1_2250(.VSS(VSS),.VDD(VDD),.Y(I16059),.A(g3878));
  NOT NOT1_2251(.VSS(VSS),.VDD(VDD),.Y(g8829),.A(I16059));
  NOT NOT1_2252(.VSS(VSS),.VDD(VDD),.Y(I16062),.A(g3900));
  NOT NOT1_2253(.VSS(VSS),.VDD(VDD),.Y(g8832),.A(I16062));
  NOT NOT1_2254(.VSS(VSS),.VDD(VDD),.Y(I16065),.A(g7936));
  NOT NOT1_2255(.VSS(VSS),.VDD(VDD),.Y(g8835),.A(I16065));
  NOT NOT1_2256(.VSS(VSS),.VDD(VDD),.Y(I16068),.A(g5438));
  NOT NOT1_2257(.VSS(VSS),.VDD(VDD),.Y(g8836),.A(I16068));
  NOT NOT1_2258(.VSS(VSS),.VDD(VDD),.Y(I16071),.A(g5395));
  NOT NOT1_2259(.VSS(VSS),.VDD(VDD),.Y(g8839),.A(I16071));
  NOT NOT1_2260(.VSS(VSS),.VDD(VDD),.Y(I16074),.A(g5399));
  NOT NOT1_2261(.VSS(VSS),.VDD(VDD),.Y(g8840),.A(I16074));
  NOT NOT1_2262(.VSS(VSS),.VDD(VDD),.Y(I16079),.A(g6086));
  NOT NOT1_2263(.VSS(VSS),.VDD(VDD),.Y(g8843),.A(I16079));
  NOT NOT1_2264(.VSS(VSS),.VDD(VDD),.Y(I16082),.A(g5401));
  NOT NOT1_2265(.VSS(VSS),.VDD(VDD),.Y(g8844),.A(I16082));
  NOT NOT1_2266(.VSS(VSS),.VDD(VDD),.Y(I16085),.A(g6080));
  NOT NOT1_2267(.VSS(VSS),.VDD(VDD),.Y(g8845),.A(I16085));
  NOT NOT1_2268(.VSS(VSS),.VDD(VDD),.Y(g8846),.A(g4779));
  NOT NOT1_2269(.VSS(VSS),.VDD(VDD),.Y(I16089),.A(g6751));
  NOT NOT1_2270(.VSS(VSS),.VDD(VDD),.Y(g8847),.A(I16089));
  NOT NOT1_2271(.VSS(VSS),.VDD(VDD),.Y(I16092),.A(g5402));
  NOT NOT1_2272(.VSS(VSS),.VDD(VDD),.Y(g8850),.A(I16092));
  NOT NOT1_2273(.VSS(VSS),.VDD(VDD),.Y(I16095),.A(g6082));
  NOT NOT1_2274(.VSS(VSS),.VDD(VDD),.Y(g8851),.A(I16095));
  NOT NOT1_2275(.VSS(VSS),.VDD(VDD),.Y(I16098),.A(g6084));
  NOT NOT1_2276(.VSS(VSS),.VDD(VDD),.Y(g8852),.A(I16098));
  NOT NOT1_2277(.VSS(VSS),.VDD(VDD),.Y(I16101),.A(g3878));
  NOT NOT1_2278(.VSS(VSS),.VDD(VDD),.Y(g8853),.A(I16101));
  NOT NOT1_2279(.VSS(VSS),.VDD(VDD),.Y(I16104),.A(g6448));
  NOT NOT1_2280(.VSS(VSS),.VDD(VDD),.Y(g8856),.A(I16104));
  NOT NOT1_2281(.VSS(VSS),.VDD(VDD),.Y(I16107),.A(g5398));
  NOT NOT1_2282(.VSS(VSS),.VDD(VDD),.Y(g8859),.A(I16107));
  NOT NOT1_2283(.VSS(VSS),.VDD(VDD),.Y(I16110),.A(g5404));
  NOT NOT1_2284(.VSS(VSS),.VDD(VDD),.Y(g8860),.A(I16110));
  NOT NOT1_2285(.VSS(VSS),.VDD(VDD),.Y(I16114),.A(g7936));
  NOT NOT1_2286(.VSS(VSS),.VDD(VDD),.Y(g8862),.A(I16114));
  NOT NOT1_2287(.VSS(VSS),.VDD(VDD),.Y(I16117),.A(g5473));
  NOT NOT1_2288(.VSS(VSS),.VDD(VDD),.Y(g8863),.A(I16117));
  NOT NOT1_2289(.VSS(VSS),.VDD(VDD),.Y(I16120),.A(g5400));
  NOT NOT1_2290(.VSS(VSS),.VDD(VDD),.Y(g8866),.A(I16120));
  NOT NOT1_2291(.VSS(VSS),.VDD(VDD),.Y(I16123),.A(g5406));
  NOT NOT1_2292(.VSS(VSS),.VDD(VDD),.Y(g8867),.A(I16123));
  NOT NOT1_2293(.VSS(VSS),.VDD(VDD),.Y(I16128),.A(g6103));
  NOT NOT1_2294(.VSS(VSS),.VDD(VDD),.Y(g8870),.A(I16128));
  NOT NOT1_2295(.VSS(VSS),.VDD(VDD),.Y(I16131),.A(g5408));
  NOT NOT1_2296(.VSS(VSS),.VDD(VDD),.Y(g8871),.A(I16131));
  NOT NOT1_2297(.VSS(VSS),.VDD(VDD),.Y(I16134),.A(g6099));
  NOT NOT1_2298(.VSS(VSS),.VDD(VDD),.Y(g8872),.A(I16134));
  NOT NOT1_2299(.VSS(VSS),.VDD(VDD),.Y(g8873),.A(g4955));
  NOT NOT1_2300(.VSS(VSS),.VDD(VDD),.Y(I16138),.A(g7053));
  NOT NOT1_2301(.VSS(VSS),.VDD(VDD),.Y(g8874),.A(I16138));
  NOT NOT1_2302(.VSS(VSS),.VDD(VDD),.Y(I16141),.A(g5409));
  NOT NOT1_2303(.VSS(VSS),.VDD(VDD),.Y(g8877),.A(I16141));
  NOT NOT1_2304(.VSS(VSS),.VDD(VDD),.Y(I16144),.A(g6101));
  NOT NOT1_2305(.VSS(VSS),.VDD(VDD),.Y(g8878),.A(I16144));
  NOT NOT1_2306(.VSS(VSS),.VDD(VDD),.Y(I16147),.A(g3878));
  NOT NOT1_2307(.VSS(VSS),.VDD(VDD),.Y(g8879),.A(I16147));
  NOT NOT1_2308(.VSS(VSS),.VDD(VDD),.Y(I16150),.A(g3900));
  NOT NOT1_2309(.VSS(VSS),.VDD(VDD),.Y(g8882),.A(I16150));
  NOT NOT1_2310(.VSS(VSS),.VDD(VDD),.Y(I16153),.A(g3306));
  NOT NOT1_2311(.VSS(VSS),.VDD(VDD),.Y(g8885),.A(I16153));
  NOT NOT1_2312(.VSS(VSS),.VDD(VDD),.Y(I16156),.A(g5438));
  NOT NOT1_2313(.VSS(VSS),.VDD(VDD),.Y(g8888),.A(I16156));
  NOT NOT1_2314(.VSS(VSS),.VDD(VDD),.Y(I16159),.A(g5403));
  NOT NOT1_2315(.VSS(VSS),.VDD(VDD),.Y(g8891),.A(I16159));
  NOT NOT1_2316(.VSS(VSS),.VDD(VDD),.Y(I16163),.A(g6031));
  NOT NOT1_2317(.VSS(VSS),.VDD(VDD),.Y(g8893),.A(I16163));
  NOT NOT1_2318(.VSS(VSS),.VDD(VDD),.Y(I16166),.A(g6713));
  NOT NOT1_2319(.VSS(VSS),.VDD(VDD),.Y(g8894),.A(I16166));
  NOT NOT1_2320(.VSS(VSS),.VDD(VDD),.Y(I16169),.A(g5405));
  NOT NOT1_2321(.VSS(VSS),.VDD(VDD),.Y(g8897),.A(I16169));
  NOT NOT1_2322(.VSS(VSS),.VDD(VDD),.Y(I16172),.A(g5413));
  NOT NOT1_2323(.VSS(VSS),.VDD(VDD),.Y(g8898),.A(I16172));
  NOT NOT1_2324(.VSS(VSS),.VDD(VDD),.Y(I16176),.A(g7936));
  NOT NOT1_2325(.VSS(VSS),.VDD(VDD),.Y(g8900),.A(I16176));
  NOT NOT1_2326(.VSS(VSS),.VDD(VDD),.Y(I16179),.A(g5512));
  NOT NOT1_2327(.VSS(VSS),.VDD(VDD),.Y(g8901),.A(I16179));
  NOT NOT1_2328(.VSS(VSS),.VDD(VDD),.Y(I16182),.A(g5407));
  NOT NOT1_2329(.VSS(VSS),.VDD(VDD),.Y(g8904),.A(I16182));
  NOT NOT1_2330(.VSS(VSS),.VDD(VDD),.Y(I16185),.A(g5415));
  NOT NOT1_2331(.VSS(VSS),.VDD(VDD),.Y(g8905),.A(I16185));
  NOT NOT1_2332(.VSS(VSS),.VDD(VDD),.Y(I16190),.A(g6118));
  NOT NOT1_2333(.VSS(VSS),.VDD(VDD),.Y(g8908),.A(I16190));
  NOT NOT1_2334(.VSS(VSS),.VDD(VDD),.Y(I16193),.A(g5417));
  NOT NOT1_2335(.VSS(VSS),.VDD(VDD),.Y(g8909),.A(I16193));
  NOT NOT1_2336(.VSS(VSS),.VDD(VDD),.Y(I16196),.A(g6116));
  NOT NOT1_2337(.VSS(VSS),.VDD(VDD),.Y(g8910),.A(I16196));
  NOT NOT1_2338(.VSS(VSS),.VDD(VDD),.Y(g8911),.A(g5114));
  NOT NOT1_2339(.VSS(VSS),.VDD(VDD),.Y(I16200),.A(g7303));
  NOT NOT1_2340(.VSS(VSS),.VDD(VDD),.Y(g8912),.A(I16200));
  NOT NOT1_2341(.VSS(VSS),.VDD(VDD),.Y(I16203),.A(g3878));
  NOT NOT1_2342(.VSS(VSS),.VDD(VDD),.Y(g8915),.A(I16203));
  NOT NOT1_2343(.VSS(VSS),.VDD(VDD),.Y(I16206),.A(g6448));
  NOT NOT1_2344(.VSS(VSS),.VDD(VDD),.Y(g8918),.A(I16206));
  NOT NOT1_2345(.VSS(VSS),.VDD(VDD),.Y(I16209),.A(g5438));
  NOT NOT1_2346(.VSS(VSS),.VDD(VDD),.Y(g8921),.A(I16209));
  NOT NOT1_2347(.VSS(VSS),.VDD(VDD),.Y(I16212),.A(g5411));
  NOT NOT1_2348(.VSS(VSS),.VDD(VDD),.Y(g8924),.A(I16212));
  NOT NOT1_2349(.VSS(VSS),.VDD(VDD),.Y(I16215),.A(g3462));
  NOT NOT1_2350(.VSS(VSS),.VDD(VDD),.Y(g8925),.A(I16215));
  NOT NOT1_2351(.VSS(VSS),.VDD(VDD),.Y(I16218),.A(g5473));
  NOT NOT1_2352(.VSS(VSS),.VDD(VDD),.Y(g8928),.A(I16218));
  NOT NOT1_2353(.VSS(VSS),.VDD(VDD),.Y(I16221),.A(g5412));
  NOT NOT1_2354(.VSS(VSS),.VDD(VDD),.Y(g8931),.A(I16221));
  NOT NOT1_2355(.VSS(VSS),.VDD(VDD),.Y(I16225),.A(g6042));
  NOT NOT1_2356(.VSS(VSS),.VDD(VDD),.Y(g8933),.A(I16225));
  NOT NOT1_2357(.VSS(VSS),.VDD(VDD),.Y(I16228),.A(g7015));
  NOT NOT1_2358(.VSS(VSS),.VDD(VDD),.Y(g8934),.A(I16228));
  NOT NOT1_2359(.VSS(VSS),.VDD(VDD),.Y(I16231),.A(g5414));
  NOT NOT1_2360(.VSS(VSS),.VDD(VDD),.Y(g8937),.A(I16231));
  NOT NOT1_2361(.VSS(VSS),.VDD(VDD),.Y(I16234),.A(g5420));
  NOT NOT1_2362(.VSS(VSS),.VDD(VDD),.Y(g8938),.A(I16234));
  NOT NOT1_2363(.VSS(VSS),.VDD(VDD),.Y(I16238),.A(g7936));
  NOT NOT1_2364(.VSS(VSS),.VDD(VDD),.Y(g8940),.A(I16238));
  NOT NOT1_2365(.VSS(VSS),.VDD(VDD),.Y(I16241),.A(g5556));
  NOT NOT1_2366(.VSS(VSS),.VDD(VDD),.Y(g8941),.A(I16241));
  NOT NOT1_2367(.VSS(VSS),.VDD(VDD),.Y(I16244),.A(g5416));
  NOT NOT1_2368(.VSS(VSS),.VDD(VDD),.Y(g8944),.A(I16244));
  NOT NOT1_2369(.VSS(VSS),.VDD(VDD),.Y(I16247),.A(g5422));
  NOT NOT1_2370(.VSS(VSS),.VDD(VDD),.Y(g8945),.A(I16247));
  NOT NOT1_2371(.VSS(VSS),.VDD(VDD),.Y(I16252),.A(g6134));
  NOT NOT1_2372(.VSS(VSS),.VDD(VDD),.Y(g8948),.A(I16252));
  NOT NOT1_2373(.VSS(VSS),.VDD(VDD),.Y(I16255),.A(g3900));
  NOT NOT1_2374(.VSS(VSS),.VDD(VDD),.Y(g8949),.A(I16255));
  NOT NOT1_2375(.VSS(VSS),.VDD(VDD),.Y(I16258),.A(g3306));
  NOT NOT1_2376(.VSS(VSS),.VDD(VDD),.Y(g8952),.A(I16258));
  NOT NOT1_2377(.VSS(VSS),.VDD(VDD),.Y(I16261),.A(g6448));
  NOT NOT1_2378(.VSS(VSS),.VDD(VDD),.Y(g8955),.A(I16261));
  NOT NOT1_2379(.VSS(VSS),.VDD(VDD),.Y(I16264),.A(g6713));
  NOT NOT1_2380(.VSS(VSS),.VDD(VDD),.Y(g8958),.A(I16264));
  NOT NOT1_2381(.VSS(VSS),.VDD(VDD),.Y(I16267),.A(g5473));
  NOT NOT1_2382(.VSS(VSS),.VDD(VDD),.Y(g8961),.A(I16267));
  NOT NOT1_2383(.VSS(VSS),.VDD(VDD),.Y(I16270),.A(g5418));
  NOT NOT1_2384(.VSS(VSS),.VDD(VDD),.Y(g8964),.A(I16270));
  NOT NOT1_2385(.VSS(VSS),.VDD(VDD),.Y(I16273),.A(g3618));
  NOT NOT1_2386(.VSS(VSS),.VDD(VDD),.Y(g8965),.A(I16273));
  NOT NOT1_2387(.VSS(VSS),.VDD(VDD),.Y(I16276),.A(g5512));
  NOT NOT1_2388(.VSS(VSS),.VDD(VDD),.Y(g8968),.A(I16276));
  NOT NOT1_2389(.VSS(VSS),.VDD(VDD),.Y(I16279),.A(g5419));
  NOT NOT1_2390(.VSS(VSS),.VDD(VDD),.Y(g8971),.A(I16279));
  NOT NOT1_2391(.VSS(VSS),.VDD(VDD),.Y(I16283),.A(g6046));
  NOT NOT1_2392(.VSS(VSS),.VDD(VDD),.Y(g8973),.A(I16283));
  NOT NOT1_2393(.VSS(VSS),.VDD(VDD),.Y(I16286),.A(g7265));
  NOT NOT1_2394(.VSS(VSS),.VDD(VDD),.Y(g8974),.A(I16286));
  NOT NOT1_2395(.VSS(VSS),.VDD(VDD),.Y(I16289),.A(g5421));
  NOT NOT1_2396(.VSS(VSS),.VDD(VDD),.Y(g8977),.A(I16289));
  NOT NOT1_2397(.VSS(VSS),.VDD(VDD),.Y(I16292),.A(g5426));
  NOT NOT1_2398(.VSS(VSS),.VDD(VDD),.Y(g8978),.A(I16292));
  NOT NOT1_2399(.VSS(VSS),.VDD(VDD),.Y(I16296),.A(g3306));
  NOT NOT1_2400(.VSS(VSS),.VDD(VDD),.Y(g8980),.A(I16296));
  NOT NOT1_2401(.VSS(VSS),.VDD(VDD),.Y(g8983),.A(g6486));
  NOT NOT1_2402(.VSS(VSS),.VDD(VDD),.Y(I16300),.A(g3462));
  NOT NOT1_2403(.VSS(VSS),.VDD(VDD),.Y(g8984),.A(I16300));
  NOT NOT1_2404(.VSS(VSS),.VDD(VDD),.Y(I16303),.A(g6713));
  NOT NOT1_2405(.VSS(VSS),.VDD(VDD),.Y(g8987),.A(I16303));
  NOT NOT1_2406(.VSS(VSS),.VDD(VDD),.Y(I16306),.A(g7015));
  NOT NOT1_2407(.VSS(VSS),.VDD(VDD),.Y(g8990),.A(I16306));
  NOT NOT1_2408(.VSS(VSS),.VDD(VDD),.Y(I16309),.A(g5512));
  NOT NOT1_2409(.VSS(VSS),.VDD(VDD),.Y(g8993),.A(I16309));
  NOT NOT1_2410(.VSS(VSS),.VDD(VDD),.Y(I16312),.A(g5424));
  NOT NOT1_2411(.VSS(VSS),.VDD(VDD),.Y(g8996),.A(I16312));
  NOT NOT1_2412(.VSS(VSS),.VDD(VDD),.Y(I16315),.A(g3774));
  NOT NOT1_2413(.VSS(VSS),.VDD(VDD),.Y(g8997),.A(I16315));
  NOT NOT1_2414(.VSS(VSS),.VDD(VDD),.Y(I16318),.A(g5556));
  NOT NOT1_2415(.VSS(VSS),.VDD(VDD),.Y(g9000),.A(I16318));
  NOT NOT1_2416(.VSS(VSS),.VDD(VDD),.Y(I16321),.A(g5425));
  NOT NOT1_2417(.VSS(VSS),.VDD(VDD),.Y(g9003),.A(I16321));
  NOT NOT1_2418(.VSS(VSS),.VDD(VDD),.Y(I16325),.A(g6052));
  NOT NOT1_2419(.VSS(VSS),.VDD(VDD),.Y(g9005),.A(I16325));
  NOT NOT1_2420(.VSS(VSS),.VDD(VDD),.Y(I16328),.A(g3900));
  NOT NOT1_2421(.VSS(VSS),.VDD(VDD),.Y(g9006),.A(I16328));
  NOT NOT1_2422(.VSS(VSS),.VDD(VDD),.Y(I16332),.A(g3462));
  NOT NOT1_2423(.VSS(VSS),.VDD(VDD),.Y(g9010),.A(I16332));
  NOT NOT1_2424(.VSS(VSS),.VDD(VDD),.Y(I16335),.A(g3618));
  NOT NOT1_2425(.VSS(VSS),.VDD(VDD),.Y(g9013),.A(I16335));
  NOT NOT1_2426(.VSS(VSS),.VDD(VDD),.Y(I16338),.A(g7015));
  NOT NOT1_2427(.VSS(VSS),.VDD(VDD),.Y(g9016),.A(I16338));
  NOT NOT1_2428(.VSS(VSS),.VDD(VDD),.Y(I16341),.A(g7265));
  NOT NOT1_2429(.VSS(VSS),.VDD(VDD),.Y(g9019),.A(I16341));
  NOT NOT1_2430(.VSS(VSS),.VDD(VDD),.Y(I16344),.A(g5556));
  NOT NOT1_2431(.VSS(VSS),.VDD(VDD),.Y(g9022),.A(I16344));
  NOT NOT1_2432(.VSS(VSS),.VDD(VDD),.Y(I16347),.A(g5427));
  NOT NOT1_2433(.VSS(VSS),.VDD(VDD),.Y(g9025),.A(I16347));
  NOT NOT1_2434(.VSS(VSS),.VDD(VDD),.Y(g9027),.A(g5679));
  NOT NOT1_2435(.VSS(VSS),.VDD(VDD),.Y(I16354),.A(g3618));
  NOT NOT1_2436(.VSS(VSS),.VDD(VDD),.Y(g9035),.A(I16354));
  NOT NOT1_2437(.VSS(VSS),.VDD(VDD),.Y(I16357),.A(g3774));
  NOT NOT1_2438(.VSS(VSS),.VDD(VDD),.Y(g9038),.A(I16357));
  NOT NOT1_2439(.VSS(VSS),.VDD(VDD),.Y(I16360),.A(g7265));
  NOT NOT1_2440(.VSS(VSS),.VDD(VDD),.Y(g9041),.A(I16360));
  NOT NOT1_2441(.VSS(VSS),.VDD(VDD),.Y(I16363),.A(g3900));
  NOT NOT1_2442(.VSS(VSS),.VDD(VDD),.Y(g9044),.A(I16363));
  NOT NOT1_2443(.VSS(VSS),.VDD(VDD),.Y(g9050),.A(g5731));
  NOT NOT1_2444(.VSS(VSS),.VDD(VDD),.Y(I16372),.A(g3774));
  NOT NOT1_2445(.VSS(VSS),.VDD(VDD),.Y(g9058),.A(I16372));
  NOT NOT1_2446(.VSS(VSS),.VDD(VDD),.Y(g9067),.A(g5789));
  NOT NOT1_2447(.VSS(VSS),.VDD(VDD),.Y(g9084),.A(g5848));
  NOT NOT1_2448(.VSS(VSS),.VDD(VDD),.Y(I16432),.A(g3366));
  NOT NOT1_2449(.VSS(VSS),.VDD(VDD),.Y(g9128),.A(I16432));
  NOT NOT1_2450(.VSS(VSS),.VDD(VDD),.Y(I16438),.A(g3522));
  NOT NOT1_2451(.VSS(VSS),.VDD(VDD),.Y(g9134),.A(I16438));
  NOT NOT1_2452(.VSS(VSS),.VDD(VDD),.Y(I16444),.A(g3678));
  NOT NOT1_2453(.VSS(VSS),.VDD(VDD),.Y(g9140),.A(I16444));
  NOT NOT1_2454(.VSS(VSS),.VDD(VDD),.Y(I16450),.A(g3834));
  NOT NOT1_2455(.VSS(VSS),.VDD(VDD),.Y(g9146),.A(I16450));
  NOT NOT1_2456(.VSS(VSS),.VDD(VDD),.Y(I16453),.A(g7936));
  NOT NOT1_2457(.VSS(VSS),.VDD(VDD),.Y(g9149),.A(I16453));
  NOT NOT1_2458(.VSS(VSS),.VDD(VDD),.Y(g9150),.A(g5893));
  NOT NOT1_2459(.VSS(VSS),.VDD(VDD),.Y(I16457),.A(g7936));
  NOT NOT1_2460(.VSS(VSS),.VDD(VDD),.Y(g9159),.A(I16457));
  NOT NOT1_2461(.VSS(VSS),.VDD(VDD),.Y(g9160),.A(g6170));
  NOT NOT1_2462(.VSS(VSS),.VDD(VDD),.Y(g9161),.A(g5852));
  NOT NOT1_2463(.VSS(VSS),.VDD(VDD),.Y(I16462),.A(g5438));
  NOT NOT1_2464(.VSS(VSS),.VDD(VDD),.Y(g9170),.A(I16462));
  NOT NOT1_2465(.VSS(VSS),.VDD(VDD),.Y(I16465),.A(g6000));
  NOT NOT1_2466(.VSS(VSS),.VDD(VDD),.Y(g9173),.A(I16465));
  NOT NOT1_2467(.VSS(VSS),.VDD(VDD),.Y(g9174),.A(g5932));
  NOT NOT1_2468(.VSS(VSS),.VDD(VDD),.Y(I16469),.A(g7936));
  NOT NOT1_2469(.VSS(VSS),.VDD(VDD),.Y(g9183),.A(I16469));
  NOT NOT1_2470(.VSS(VSS),.VDD(VDD),.Y(I16472),.A(g7901));
  NOT NOT1_2471(.VSS(VSS),.VDD(VDD),.Y(g9184),.A(I16472));
  NOT NOT1_2472(.VSS(VSS),.VDD(VDD),.Y(g9187),.A(g5803));
  NOT NOT1_2473(.VSS(VSS),.VDD(VDD),.Y(I16476),.A(g6448));
  NOT NOT1_2474(.VSS(VSS),.VDD(VDD),.Y(g9196),.A(I16476));
  NOT NOT1_2475(.VSS(VSS),.VDD(VDD),.Y(I16479),.A(g5438));
  NOT NOT1_2476(.VSS(VSS),.VDD(VDD),.Y(g9199),.A(I16479));
  NOT NOT1_2477(.VSS(VSS),.VDD(VDD),.Y(I16482),.A(g6000));
  NOT NOT1_2478(.VSS(VSS),.VDD(VDD),.Y(g9202),.A(I16482));
  NOT NOT1_2479(.VSS(VSS),.VDD(VDD),.Y(g9203),.A(g5899));
  NOT NOT1_2480(.VSS(VSS),.VDD(VDD),.Y(I16486),.A(g5473));
  NOT NOT1_2481(.VSS(VSS),.VDD(VDD),.Y(g9212),.A(I16486));
  NOT NOT1_2482(.VSS(VSS),.VDD(VDD),.Y(I16489),.A(g6000));
  NOT NOT1_2483(.VSS(VSS),.VDD(VDD),.Y(g9215),.A(I16489));
  NOT NOT1_2484(.VSS(VSS),.VDD(VDD),.Y(g9216),.A(g5966));
  NOT NOT1_2485(.VSS(VSS),.VDD(VDD),.Y(I16493),.A(g7936));
  NOT NOT1_2486(.VSS(VSS),.VDD(VDD),.Y(g9225),.A(I16493));
  NOT NOT1_2487(.VSS(VSS),.VDD(VDD),.Y(g9226),.A(g5434));
  NOT NOT1_2488(.VSS(VSS),.VDD(VDD),.Y(g9227),.A(g5587));
  NOT NOT1_2489(.VSS(VSS),.VDD(VDD),.Y(g9228),.A(g7667));
  NOT NOT1_2490(.VSS(VSS),.VDD(VDD),.Y(I16499),.A(g7901));
  NOT NOT1_2491(.VSS(VSS),.VDD(VDD),.Y(g9229),.A(I16499));
  NOT NOT1_2492(.VSS(VSS),.VDD(VDD),.Y(g9232),.A(g5752));
  NOT NOT1_2493(.VSS(VSS),.VDD(VDD),.Y(I16504),.A(g3306));
  NOT NOT1_2494(.VSS(VSS),.VDD(VDD),.Y(g9242),.A(I16504));
  NOT NOT1_2495(.VSS(VSS),.VDD(VDD),.Y(I16507),.A(g6448));
  NOT NOT1_2496(.VSS(VSS),.VDD(VDD),.Y(g9245),.A(I16507));
  NOT NOT1_2497(.VSS(VSS),.VDD(VDD),.Y(g9248),.A(g5859));
  NOT NOT1_2498(.VSS(VSS),.VDD(VDD),.Y(I16511),.A(g6713));
  NOT NOT1_2499(.VSS(VSS),.VDD(VDD),.Y(g9257),.A(I16511));
  NOT NOT1_2500(.VSS(VSS),.VDD(VDD),.Y(I16514),.A(g5473));
  NOT NOT1_2501(.VSS(VSS),.VDD(VDD),.Y(g9260),.A(I16514));
  NOT NOT1_2502(.VSS(VSS),.VDD(VDD),.Y(I16517),.A(g6000));
  NOT NOT1_2503(.VSS(VSS),.VDD(VDD),.Y(g9263),.A(I16517));
  NOT NOT1_2504(.VSS(VSS),.VDD(VDD),.Y(g9264),.A(g5938));
  NOT NOT1_2505(.VSS(VSS),.VDD(VDD),.Y(I16521),.A(g5512));
  NOT NOT1_2506(.VSS(VSS),.VDD(VDD),.Y(g9273),.A(I16521));
  NOT NOT1_2507(.VSS(VSS),.VDD(VDD),.Y(I16524),.A(g6000));
  NOT NOT1_2508(.VSS(VSS),.VDD(VDD),.Y(g9276),.A(I16524));
  NOT NOT1_2509(.VSS(VSS),.VDD(VDD),.Y(g9277),.A(g5995));
  NOT NOT1_2510(.VSS(VSS),.VDD(VDD),.Y(g9286),.A(g6197));
  NOT NOT1_2511(.VSS(VSS),.VDD(VDD),.Y(g9287),.A(g6638));
  NOT NOT1_2512(.VSS(VSS),.VDD(VDD),.Y(g9288),.A(g5363));
  NOT NOT1_2513(.VSS(VSS),.VDD(VDD),.Y(g9289),.A(g5379));
  NOT NOT1_2514(.VSS(VSS),.VDD(VDD),.Y(I16532),.A(g7901));
  NOT NOT1_2515(.VSS(VSS),.VDD(VDD),.Y(g9290),.A(I16532));
  NOT NOT1_2516(.VSS(VSS),.VDD(VDD),.Y(g9293),.A(g5703));
  NOT NOT1_2517(.VSS(VSS),.VDD(VDD),.Y(I16538),.A(g3306));
  NOT NOT1_2518(.VSS(VSS),.VDD(VDD),.Y(g9303),.A(I16538));
  NOT NOT1_2519(.VSS(VSS),.VDD(VDD),.Y(I16541),.A(g5438));
  NOT NOT1_2520(.VSS(VSS),.VDD(VDD),.Y(g9306),.A(I16541));
  NOT NOT1_2521(.VSS(VSS),.VDD(VDD),.Y(I16544),.A(g6054));
  NOT NOT1_2522(.VSS(VSS),.VDD(VDD),.Y(g9309),.A(I16544));
  NOT NOT1_2523(.VSS(VSS),.VDD(VDD),.Y(g9310),.A(g5811));
  NOT NOT1_2524(.VSS(VSS),.VDD(VDD),.Y(I16549),.A(g3462));
  NOT NOT1_2525(.VSS(VSS),.VDD(VDD),.Y(g9320),.A(I16549));
  NOT NOT1_2526(.VSS(VSS),.VDD(VDD),.Y(I16552),.A(g6713));
  NOT NOT1_2527(.VSS(VSS),.VDD(VDD),.Y(g9323),.A(I16552));
  NOT NOT1_2528(.VSS(VSS),.VDD(VDD),.Y(g9326),.A(g5906));
  NOT NOT1_2529(.VSS(VSS),.VDD(VDD),.Y(I16556),.A(g7015));
  NOT NOT1_2530(.VSS(VSS),.VDD(VDD),.Y(g9335),.A(I16556));
  NOT NOT1_2531(.VSS(VSS),.VDD(VDD),.Y(I16559),.A(g5512));
  NOT NOT1_2532(.VSS(VSS),.VDD(VDD),.Y(g9338),.A(I16559));
  NOT NOT1_2533(.VSS(VSS),.VDD(VDD),.Y(I16562),.A(g6000));
  NOT NOT1_2534(.VSS(VSS),.VDD(VDD),.Y(g9341),.A(I16562));
  NOT NOT1_2535(.VSS(VSS),.VDD(VDD),.Y(g9342),.A(g5972));
  NOT NOT1_2536(.VSS(VSS),.VDD(VDD),.Y(I16566),.A(g5556));
  NOT NOT1_2537(.VSS(VSS),.VDD(VDD),.Y(g9351),.A(I16566));
  NOT NOT1_2538(.VSS(VSS),.VDD(VDD),.Y(I16569),.A(g6000));
  NOT NOT1_2539(.VSS(VSS),.VDD(VDD),.Y(g9354),.A(I16569));
  NOT NOT1_2540(.VSS(VSS),.VDD(VDD),.Y(g9355),.A(g7639));
  NOT NOT1_2541(.VSS(VSS),.VDD(VDD),.Y(g9356),.A(g5665));
  NOT NOT1_2542(.VSS(VSS),.VDD(VDD),.Y(I16578),.A(g6448));
  NOT NOT1_2543(.VSS(VSS),.VDD(VDD),.Y(g9368),.A(I16578));
  NOT NOT1_2544(.VSS(VSS),.VDD(VDD),.Y(I16581),.A(g5438));
  NOT NOT1_2545(.VSS(VSS),.VDD(VDD),.Y(g9371),.A(I16581));
  NOT NOT1_2546(.VSS(VSS),.VDD(VDD),.Y(g9374),.A(g5761));
  NOT NOT1_2547(.VSS(VSS),.VDD(VDD),.Y(I16587),.A(g3462));
  NOT NOT1_2548(.VSS(VSS),.VDD(VDD),.Y(g9384),.A(I16587));
  NOT NOT1_2549(.VSS(VSS),.VDD(VDD),.Y(I16590),.A(g5473));
  NOT NOT1_2550(.VSS(VSS),.VDD(VDD),.Y(g9387),.A(I16590));
  NOT NOT1_2551(.VSS(VSS),.VDD(VDD),.Y(I16593),.A(g6059));
  NOT NOT1_2552(.VSS(VSS),.VDD(VDD),.Y(g9390),.A(I16593));
  NOT NOT1_2553(.VSS(VSS),.VDD(VDD),.Y(g9391),.A(g5867));
  NOT NOT1_2554(.VSS(VSS),.VDD(VDD),.Y(I16598),.A(g3618));
  NOT NOT1_2555(.VSS(VSS),.VDD(VDD),.Y(g9401),.A(I16598));
  NOT NOT1_2556(.VSS(VSS),.VDD(VDD),.Y(I16601),.A(g7015));
  NOT NOT1_2557(.VSS(VSS),.VDD(VDD),.Y(g9404),.A(I16601));
  NOT NOT1_2558(.VSS(VSS),.VDD(VDD),.Y(g9407),.A(g5945));
  NOT NOT1_2559(.VSS(VSS),.VDD(VDD),.Y(I16605),.A(g7265));
  NOT NOT1_2560(.VSS(VSS),.VDD(VDD),.Y(g9416),.A(I16605));
  NOT NOT1_2561(.VSS(VSS),.VDD(VDD),.Y(I16608),.A(g5556));
  NOT NOT1_2562(.VSS(VSS),.VDD(VDD),.Y(g9419),.A(I16608));
  NOT NOT1_2563(.VSS(VSS),.VDD(VDD),.Y(I16611),.A(g6000));
  NOT NOT1_2564(.VSS(VSS),.VDD(VDD),.Y(g9422),.A(I16611));
  NOT NOT1_2565(.VSS(VSS),.VDD(VDD),.Y(g9423),.A(g5428));
  NOT NOT1_2566(.VSS(VSS),.VDD(VDD),.Y(g9424),.A(g5469));
  NOT NOT1_2567(.VSS(VSS),.VDD(VDD),.Y(g9425),.A(g5346));
  NOT NOT1_2568(.VSS(VSS),.VDD(VDD),.Y(g9426),.A(g5543));
  NOT NOT1_2569(.VSS(VSS),.VDD(VDD),.Y(g9427),.A(g5645));
  NOT NOT1_2570(.VSS(VSS),.VDD(VDD),.Y(I16624),.A(g3306));
  NOT NOT1_2571(.VSS(VSS),.VDD(VDD),.Y(g9443),.A(I16624));
  NOT NOT1_2572(.VSS(VSS),.VDD(VDD),.Y(I16627),.A(g6448));
  NOT NOT1_2573(.VSS(VSS),.VDD(VDD),.Y(g9446),.A(I16627));
  NOT NOT1_2574(.VSS(VSS),.VDD(VDD),.Y(I16630),.A(g6057));
  NOT NOT1_2575(.VSS(VSS),.VDD(VDD),.Y(g9449),.A(I16630));
  NOT NOT1_2576(.VSS(VSS),.VDD(VDD),.Y(I16633),.A(g6486));
  NOT NOT1_2577(.VSS(VSS),.VDD(VDD),.Y(g9450),.A(I16633));
  NOT NOT1_2578(.VSS(VSS),.VDD(VDD),.Y(g9453),.A(g5717));
  NOT NOT1_2579(.VSS(VSS),.VDD(VDD),.Y(I16641),.A(g6713));
  NOT NOT1_2580(.VSS(VSS),.VDD(VDD),.Y(g9465),.A(I16641));
  NOT NOT1_2581(.VSS(VSS),.VDD(VDD),.Y(I16644),.A(g5473));
  NOT NOT1_2582(.VSS(VSS),.VDD(VDD),.Y(g9468),.A(I16644));
  NOT NOT1_2583(.VSS(VSS),.VDD(VDD),.Y(g9471),.A(g5820));
  NOT NOT1_2584(.VSS(VSS),.VDD(VDD),.Y(I16650),.A(g3618));
  NOT NOT1_2585(.VSS(VSS),.VDD(VDD),.Y(g9481),.A(I16650));
  NOT NOT1_2586(.VSS(VSS),.VDD(VDD),.Y(I16653),.A(g5512));
  NOT NOT1_2587(.VSS(VSS),.VDD(VDD),.Y(g9484),.A(I16653));
  NOT NOT1_2588(.VSS(VSS),.VDD(VDD),.Y(I16656),.A(g6066));
  NOT NOT1_2589(.VSS(VSS),.VDD(VDD),.Y(g9487),.A(I16656));
  NOT NOT1_2590(.VSS(VSS),.VDD(VDD),.Y(g9488),.A(g5914));
  NOT NOT1_2591(.VSS(VSS),.VDD(VDD),.Y(I16661),.A(g3774));
  NOT NOT1_2592(.VSS(VSS),.VDD(VDD),.Y(g9498),.A(I16661));
  NOT NOT1_2593(.VSS(VSS),.VDD(VDD),.Y(I16664),.A(g7265));
  NOT NOT1_2594(.VSS(VSS),.VDD(VDD),.Y(g9501),.A(I16664));
  NOT NOT1_2595(.VSS(VSS),.VDD(VDD),.Y(g9504),.A(g6149));
  NOT NOT1_2596(.VSS(VSS),.VDD(VDD),.Y(g9505),.A(g6227));
  NOT NOT1_2597(.VSS(VSS),.VDD(VDD),.Y(g9506),.A(g6444));
  NOT NOT1_2598(.VSS(VSS),.VDD(VDD),.Y(g9507),.A(g5953));
  NOT NOT1_2599(.VSS(VSS),.VDD(VDD),.Y(I16677),.A(g3306));
  NOT NOT1_2600(.VSS(VSS),.VDD(VDD),.Y(g9524),.A(I16677));
  NOT NOT1_2601(.VSS(VSS),.VDD(VDD),.Y(g9527),.A(g5508));
  NOT NOT1_2602(.VSS(VSS),.VDD(VDD),.Y(I16681),.A(g6643));
  NOT NOT1_2603(.VSS(VSS),.VDD(VDD),.Y(g9528),.A(I16681));
  NOT NOT1_2604(.VSS(VSS),.VDD(VDD),.Y(I16684),.A(g6486));
  NOT NOT1_2605(.VSS(VSS),.VDD(VDD),.Y(g9531),.A(I16684));
  NOT NOT1_2606(.VSS(VSS),.VDD(VDD),.Y(g9569),.A(g5683));
  NOT NOT1_2607(.VSS(VSS),.VDD(VDD),.Y(I16694),.A(g3462));
  NOT NOT1_2608(.VSS(VSS),.VDD(VDD),.Y(g9585),.A(I16694));
  NOT NOT1_2609(.VSS(VSS),.VDD(VDD),.Y(I16697),.A(g6713));
  NOT NOT1_2610(.VSS(VSS),.VDD(VDD),.Y(g9588),.A(I16697));
  NOT NOT1_2611(.VSS(VSS),.VDD(VDD),.Y(I16700),.A(g6064));
  NOT NOT1_2612(.VSS(VSS),.VDD(VDD),.Y(g9591),.A(I16700));
  NOT NOT1_2613(.VSS(VSS),.VDD(VDD),.Y(I16703),.A(g6751));
  NOT NOT1_2614(.VSS(VSS),.VDD(VDD),.Y(g9592),.A(I16703));
  NOT NOT1_2615(.VSS(VSS),.VDD(VDD),.Y(g9595),.A(g5775));
  NOT NOT1_2616(.VSS(VSS),.VDD(VDD),.Y(I16711),.A(g7015));
  NOT NOT1_2617(.VSS(VSS),.VDD(VDD),.Y(g9607),.A(I16711));
  NOT NOT1_2618(.VSS(VSS),.VDD(VDD),.Y(I16714),.A(g5512));
  NOT NOT1_2619(.VSS(VSS),.VDD(VDD),.Y(g9610),.A(I16714));
  NOT NOT1_2620(.VSS(VSS),.VDD(VDD),.Y(g9613),.A(g5876));
  NOT NOT1_2621(.VSS(VSS),.VDD(VDD),.Y(I16720),.A(g3774));
  NOT NOT1_2622(.VSS(VSS),.VDD(VDD),.Y(g9623),.A(I16720));
  NOT NOT1_2623(.VSS(VSS),.VDD(VDD),.Y(I16723),.A(g5556));
  NOT NOT1_2624(.VSS(VSS),.VDD(VDD),.Y(g9626),.A(I16723));
  NOT NOT1_2625(.VSS(VSS),.VDD(VDD),.Y(I16726),.A(g6085));
  NOT NOT1_2626(.VSS(VSS),.VDD(VDD),.Y(g9629),.A(I16726));
  NOT NOT1_2627(.VSS(VSS),.VDD(VDD),.Y(I16741),.A(g6062));
  NOT NOT1_2628(.VSS(VSS),.VDD(VDD),.Y(g9640),.A(I16741));
  NOT NOT1_2629(.VSS(VSS),.VDD(VDD),.Y(I16744),.A(g3338));
  NOT NOT1_2630(.VSS(VSS),.VDD(VDD),.Y(g9641),.A(I16744));
  NOT NOT1_2631(.VSS(VSS),.VDD(VDD),.Y(I16747),.A(g6643));
  NOT NOT1_2632(.VSS(VSS),.VDD(VDD),.Y(g9644),.A(I16747));
  NOT NOT1_2633(.VSS(VSS),.VDD(VDD),.Y(g9649),.A(g5982));
  NOT NOT1_2634(.VSS(VSS),.VDD(VDD),.Y(I16759),.A(g3462));
  NOT NOT1_2635(.VSS(VSS),.VDD(VDD),.Y(g9666),.A(I16759));
  NOT NOT1_2636(.VSS(VSS),.VDD(VDD),.Y(g9669),.A(g5552));
  NOT NOT1_2637(.VSS(VSS),.VDD(VDD),.Y(I16763),.A(g6945));
  NOT NOT1_2638(.VSS(VSS),.VDD(VDD),.Y(g9670),.A(I16763));
  NOT NOT1_2639(.VSS(VSS),.VDD(VDD),.Y(I16766),.A(g6751));
  NOT NOT1_2640(.VSS(VSS),.VDD(VDD),.Y(g9673),.A(I16766));
  NOT NOT1_2641(.VSS(VSS),.VDD(VDD),.Y(g9711),.A(g5735));
  NOT NOT1_2642(.VSS(VSS),.VDD(VDD),.Y(I16776),.A(g3618));
  NOT NOT1_2643(.VSS(VSS),.VDD(VDD),.Y(g9727),.A(I16776));
  NOT NOT1_2644(.VSS(VSS),.VDD(VDD),.Y(I16779),.A(g7015));
  NOT NOT1_2645(.VSS(VSS),.VDD(VDD),.Y(g9730),.A(I16779));
  NOT NOT1_2646(.VSS(VSS),.VDD(VDD),.Y(I16782),.A(g6083));
  NOT NOT1_2647(.VSS(VSS),.VDD(VDD),.Y(g9733),.A(I16782));
  NOT NOT1_2648(.VSS(VSS),.VDD(VDD),.Y(I16785),.A(g7053));
  NOT NOT1_2649(.VSS(VSS),.VDD(VDD),.Y(g9734),.A(I16785));
  NOT NOT1_2650(.VSS(VSS),.VDD(VDD),.Y(g9737),.A(g5834));
  NOT NOT1_2651(.VSS(VSS),.VDD(VDD),.Y(I16793),.A(g7265));
  NOT NOT1_2652(.VSS(VSS),.VDD(VDD),.Y(g9749),.A(I16793));
  NOT NOT1_2653(.VSS(VSS),.VDD(VDD),.Y(I16796),.A(g5556));
  NOT NOT1_2654(.VSS(VSS),.VDD(VDD),.Y(g9752),.A(I16796));
  NOT NOT1_2655(.VSS(VSS),.VDD(VDD),.Y(g9755),.A(g5431));
  NOT NOT1_2656(.VSS(VSS),.VDD(VDD),.Y(g9756),.A(g5504));
  NOT NOT1_2657(.VSS(VSS),.VDD(VDD),.Y(g9757),.A(g5601));
  NOT NOT1_2658(.VSS(VSS),.VDD(VDD),.Y(g9758),.A(g5618));
  NOT NOT1_2659(.VSS(VSS),.VDD(VDD),.Y(I16811),.A(g3338));
  NOT NOT1_2660(.VSS(VSS),.VDD(VDD),.Y(g9767),.A(I16811));
  NOT NOT1_2661(.VSS(VSS),.VDD(VDD),.Y(I16814),.A(g6486));
  NOT NOT1_2662(.VSS(VSS),.VDD(VDD),.Y(g9770),.A(I16814));
  NOT NOT1_2663(.VSS(VSS),.VDD(VDD),.Y(I16832),.A(g6081));
  NOT NOT1_2664(.VSS(VSS),.VDD(VDD),.Y(g9786),.A(I16832));
  NOT NOT1_2665(.VSS(VSS),.VDD(VDD),.Y(I16835),.A(g3494));
  NOT NOT1_2666(.VSS(VSS),.VDD(VDD),.Y(g9787),.A(I16835));
  NOT NOT1_2667(.VSS(VSS),.VDD(VDD),.Y(I16838),.A(g6945));
  NOT NOT1_2668(.VSS(VSS),.VDD(VDD),.Y(g9790),.A(I16838));
  NOT NOT1_2669(.VSS(VSS),.VDD(VDD),.Y(g9795),.A(g6019));
  NOT NOT1_2670(.VSS(VSS),.VDD(VDD),.Y(I16850),.A(g3618));
  NOT NOT1_2671(.VSS(VSS),.VDD(VDD),.Y(g9812),.A(I16850));
  NOT NOT1_2672(.VSS(VSS),.VDD(VDD),.Y(g9815),.A(g5598));
  NOT NOT1_2673(.VSS(VSS),.VDD(VDD),.Y(I16854),.A(g7195));
  NOT NOT1_2674(.VSS(VSS),.VDD(VDD),.Y(g9816),.A(I16854));
  NOT NOT1_2675(.VSS(VSS),.VDD(VDD),.Y(I16857),.A(g7053));
  NOT NOT1_2676(.VSS(VSS),.VDD(VDD),.Y(g9819),.A(I16857));
  NOT NOT1_2677(.VSS(VSS),.VDD(VDD),.Y(g9857),.A(g5793));
  NOT NOT1_2678(.VSS(VSS),.VDD(VDD),.Y(I16867),.A(g3774));
  NOT NOT1_2679(.VSS(VSS),.VDD(VDD),.Y(g9873),.A(I16867));
  NOT NOT1_2680(.VSS(VSS),.VDD(VDD),.Y(I16870),.A(g7265));
  NOT NOT1_2681(.VSS(VSS),.VDD(VDD),.Y(g9876),.A(I16870));
  NOT NOT1_2682(.VSS(VSS),.VDD(VDD),.Y(I16873),.A(g6102));
  NOT NOT1_2683(.VSS(VSS),.VDD(VDD),.Y(g9879),.A(I16873));
  NOT NOT1_2684(.VSS(VSS),.VDD(VDD),.Y(I16876),.A(g7303));
  NOT NOT1_2685(.VSS(VSS),.VDD(VDD),.Y(g9880),.A(I16876));
  NOT NOT1_2686(.VSS(VSS),.VDD(VDD),.Y(g9884),.A(g6310));
  NOT NOT1_2687(.VSS(VSS),.VDD(VDD),.Y(g9885),.A(g6905));
  NOT NOT1_2688(.VSS(VSS),.VDD(VDD),.Y(g9886),.A(g7149));
  NOT NOT1_2689(.VSS(VSS),.VDD(VDD),.Y(I16897),.A(g6643));
  NOT NOT1_2690(.VSS(VSS),.VDD(VDD),.Y(g9895),.A(I16897));
  NOT NOT1_2691(.VSS(VSS),.VDD(VDD),.Y(I16900),.A(g6486));
  NOT NOT1_2692(.VSS(VSS),.VDD(VDD),.Y(g9898),.A(I16900));
  NOT NOT1_2693(.VSS(VSS),.VDD(VDD),.Y(I16915),.A(g3494));
  NOT NOT1_2694(.VSS(VSS),.VDD(VDD),.Y(g9913),.A(I16915));
  NOT NOT1_2695(.VSS(VSS),.VDD(VDD),.Y(I16918),.A(g6751));
  NOT NOT1_2696(.VSS(VSS),.VDD(VDD),.Y(g9916),.A(I16918));
  NOT NOT1_2697(.VSS(VSS),.VDD(VDD),.Y(I16936),.A(g6100));
  NOT NOT1_2698(.VSS(VSS),.VDD(VDD),.Y(g9932),.A(I16936));
  NOT NOT1_2699(.VSS(VSS),.VDD(VDD),.Y(I16939),.A(g3650));
  NOT NOT1_2700(.VSS(VSS),.VDD(VDD),.Y(g9933),.A(I16939));
  NOT NOT1_2701(.VSS(VSS),.VDD(VDD),.Y(I16942),.A(g7195));
  NOT NOT1_2702(.VSS(VSS),.VDD(VDD),.Y(g9936),.A(I16942));
  NOT NOT1_2703(.VSS(VSS),.VDD(VDD),.Y(g9941),.A(g6035));
  NOT NOT1_2704(.VSS(VSS),.VDD(VDD),.Y(I16954),.A(g3774));
  NOT NOT1_2705(.VSS(VSS),.VDD(VDD),.Y(g9958),.A(I16954));
  NOT NOT1_2706(.VSS(VSS),.VDD(VDD),.Y(g9961),.A(g5615));
  NOT NOT1_2707(.VSS(VSS),.VDD(VDD),.Y(I16958),.A(g7391));
  NOT NOT1_2708(.VSS(VSS),.VDD(VDD),.Y(g9962),.A(I16958));
  NOT NOT1_2709(.VSS(VSS),.VDD(VDD),.Y(I16961),.A(g7303));
  NOT NOT1_2710(.VSS(VSS),.VDD(VDD),.Y(g9965),.A(I16961));
  NOT NOT1_2711(.VSS(VSS),.VDD(VDD),.Y(I16972),.A(g3900));
  NOT NOT1_2712(.VSS(VSS),.VDD(VDD),.Y(g10004),.A(I16972));
  NOT NOT1_2713(.VSS(VSS),.VDD(VDD),.Y(g10015),.A(g5292));
  NOT NOT1_2714(.VSS(VSS),.VDD(VDD),.Y(I16984),.A(g7936));
  NOT NOT1_2715(.VSS(VSS),.VDD(VDD),.Y(g10016),.A(I16984));
  NOT NOT1_2716(.VSS(VSS),.VDD(VDD),.Y(I16987),.A(g6079));
  NOT NOT1_2717(.VSS(VSS),.VDD(VDD),.Y(g10017),.A(I16987));
  NOT NOT1_2718(.VSS(VSS),.VDD(VDD),.Y(I16990),.A(g3338));
  NOT NOT1_2719(.VSS(VSS),.VDD(VDD),.Y(g10018),.A(I16990));
  NOT NOT1_2720(.VSS(VSS),.VDD(VDD),.Y(I16993),.A(g6643));
  NOT NOT1_2721(.VSS(VSS),.VDD(VDD),.Y(g10021),.A(I16993));
  NOT NOT1_2722(.VSS(VSS),.VDD(VDD),.Y(I17009),.A(g6945));
  NOT NOT1_2723(.VSS(VSS),.VDD(VDD),.Y(g10049),.A(I17009));
  NOT NOT1_2724(.VSS(VSS),.VDD(VDD),.Y(I17012),.A(g6751));
  NOT NOT1_2725(.VSS(VSS),.VDD(VDD),.Y(g10052),.A(I17012));
  NOT NOT1_2726(.VSS(VSS),.VDD(VDD),.Y(I17027),.A(g3650));
  NOT NOT1_2727(.VSS(VSS),.VDD(VDD),.Y(g10067),.A(I17027));
  NOT NOT1_2728(.VSS(VSS),.VDD(VDD),.Y(I17030),.A(g7053));
  NOT NOT1_2729(.VSS(VSS),.VDD(VDD),.Y(g10070),.A(I17030));
  NOT NOT1_2730(.VSS(VSS),.VDD(VDD),.Y(I17048),.A(g6117));
  NOT NOT1_2731(.VSS(VSS),.VDD(VDD),.Y(g10086),.A(I17048));
  NOT NOT1_2732(.VSS(VSS),.VDD(VDD),.Y(I17051),.A(g3806));
  NOT NOT1_2733(.VSS(VSS),.VDD(VDD),.Y(g10087),.A(I17051));
  NOT NOT1_2734(.VSS(VSS),.VDD(VDD),.Y(I17054),.A(g7391));
  NOT NOT1_2735(.VSS(VSS),.VDD(VDD),.Y(g10090),.A(I17054));
  NOT NOT1_2736(.VSS(VSS),.VDD(VDD),.Y(I17066),.A(g3900));
  NOT NOT1_2737(.VSS(VSS),.VDD(VDD),.Y(g10096),.A(I17066));
  NOT NOT1_2738(.VSS(VSS),.VDD(VDD),.Y(g10099),.A(g7700));
  NOT NOT1_2739(.VSS(VSS),.VDD(VDD),.Y(I17070),.A(g7528));
  NOT NOT1_2740(.VSS(VSS),.VDD(VDD),.Y(g10100),.A(I17070));
  NOT NOT1_2741(.VSS(VSS),.VDD(VDD),.Y(I17081),.A(g3338));
  NOT NOT1_2742(.VSS(VSS),.VDD(VDD),.Y(g10109),.A(I17081));
  NOT NOT1_2743(.VSS(VSS),.VDD(VDD),.Y(g10124),.A(g5326));
  NOT NOT1_2744(.VSS(VSS),.VDD(VDD),.Y(I17097),.A(g7936));
  NOT NOT1_2745(.VSS(VSS),.VDD(VDD),.Y(g10125),.A(I17097));
  NOT NOT1_2746(.VSS(VSS),.VDD(VDD),.Y(I17100),.A(g6098));
  NOT NOT1_2747(.VSS(VSS),.VDD(VDD),.Y(g10126),.A(I17100));
  NOT NOT1_2748(.VSS(VSS),.VDD(VDD),.Y(I17103),.A(g3494));
  NOT NOT1_2749(.VSS(VSS),.VDD(VDD),.Y(g10127),.A(I17103));
  NOT NOT1_2750(.VSS(VSS),.VDD(VDD),.Y(I17106),.A(g6945));
  NOT NOT1_2751(.VSS(VSS),.VDD(VDD),.Y(g10130),.A(I17106));
  NOT NOT1_2752(.VSS(VSS),.VDD(VDD),.Y(I17122),.A(g7195));
  NOT NOT1_2753(.VSS(VSS),.VDD(VDD),.Y(g10158),.A(I17122));
  NOT NOT1_2754(.VSS(VSS),.VDD(VDD),.Y(I17125),.A(g7053));
  NOT NOT1_2755(.VSS(VSS),.VDD(VDD),.Y(g10161),.A(I17125));
  NOT NOT1_2756(.VSS(VSS),.VDD(VDD),.Y(I17140),.A(g3806));
  NOT NOT1_2757(.VSS(VSS),.VDD(VDD),.Y(g10176),.A(I17140));
  NOT NOT1_2758(.VSS(VSS),.VDD(VDD),.Y(I17143),.A(g7303));
  NOT NOT1_2759(.VSS(VSS),.VDD(VDD),.Y(g10179),.A(I17143));
  NOT NOT1_2760(.VSS(VSS),.VDD(VDD),.Y(I17159),.A(g3900));
  NOT NOT1_2761(.VSS(VSS),.VDD(VDD),.Y(g10189),.A(I17159));
  NOT NOT1_2762(.VSS(VSS),.VDD(VDD),.Y(I17184),.A(g3494));
  NOT NOT1_2763(.VSS(VSS),.VDD(VDD),.Y(g10214),.A(I17184));
  NOT NOT1_2764(.VSS(VSS),.VDD(VDD),.Y(g10229),.A(g5349));
  NOT NOT1_2765(.VSS(VSS),.VDD(VDD),.Y(I17200),.A(g7936));
  NOT NOT1_2766(.VSS(VSS),.VDD(VDD),.Y(g10230),.A(I17200));
  NOT NOT1_2767(.VSS(VSS),.VDD(VDD),.Y(I17203),.A(g6115));
  NOT NOT1_2768(.VSS(VSS),.VDD(VDD),.Y(g10231),.A(I17203));
  NOT NOT1_2769(.VSS(VSS),.VDD(VDD),.Y(I17206),.A(g3650));
  NOT NOT1_2770(.VSS(VSS),.VDD(VDD),.Y(g10232),.A(I17206));
  NOT NOT1_2771(.VSS(VSS),.VDD(VDD),.Y(I17209),.A(g7195));
  NOT NOT1_2772(.VSS(VSS),.VDD(VDD),.Y(g10235),.A(I17209));
  NOT NOT1_2773(.VSS(VSS),.VDD(VDD),.Y(I17225),.A(g7391));
  NOT NOT1_2774(.VSS(VSS),.VDD(VDD),.Y(g10263),.A(I17225));
  NOT NOT1_2775(.VSS(VSS),.VDD(VDD),.Y(I17228),.A(g7303));
  NOT NOT1_2776(.VSS(VSS),.VDD(VDD),.Y(g10266),.A(I17228));
  NOT NOT1_2777(.VSS(VSS),.VDD(VDD),.Y(I17235),.A(g3900));
  NOT NOT1_2778(.VSS(VSS),.VDD(VDD),.Y(g10273),.A(I17235));
  NOT NOT1_2779(.VSS(VSS),.VDD(VDD),.Y(I17238),.A(g3900));
  NOT NOT1_2780(.VSS(VSS),.VDD(VDD),.Y(g10276),.A(I17238));
  NOT NOT1_2781(.VSS(VSS),.VDD(VDD),.Y(I17278),.A(g3650));
  NOT NOT1_2782(.VSS(VSS),.VDD(VDD),.Y(g10316),.A(I17278));
  NOT NOT1_2783(.VSS(VSS),.VDD(VDD),.Y(g10331),.A(g5366));
  NOT NOT1_2784(.VSS(VSS),.VDD(VDD),.Y(I17294),.A(g7936));
  NOT NOT1_2785(.VSS(VSS),.VDD(VDD),.Y(g10332),.A(I17294));
  NOT NOT1_2786(.VSS(VSS),.VDD(VDD),.Y(I17297),.A(g6130));
  NOT NOT1_2787(.VSS(VSS),.VDD(VDD),.Y(g10333),.A(I17297));
  NOT NOT1_2788(.VSS(VSS),.VDD(VDD),.Y(I17300),.A(g3806));
  NOT NOT1_2789(.VSS(VSS),.VDD(VDD),.Y(g10334),.A(I17300));
  NOT NOT1_2790(.VSS(VSS),.VDD(VDD),.Y(I17303),.A(g7391));
  NOT NOT1_2791(.VSS(VSS),.VDD(VDD),.Y(g10337),.A(I17303));
  NOT NOT1_2792(.VSS(VSS),.VDD(VDD),.Y(I17311),.A(g3900));
  NOT NOT1_2793(.VSS(VSS),.VDD(VDD),.Y(g10357),.A(I17311));
  NOT NOT1_2794(.VSS(VSS),.VDD(VDD),.Y(I17363),.A(g3806));
  NOT NOT1_2795(.VSS(VSS),.VDD(VDD),.Y(g10409),.A(I17363));
  NOT NOT1_2796(.VSS(VSS),.VDD(VDD),.Y(I17370),.A(g3900));
  NOT NOT1_2797(.VSS(VSS),.VDD(VDD),.Y(g10416),.A(I17370));
  NOT NOT1_2798(.VSS(VSS),.VDD(VDD),.Y(I17373),.A(g3900));
  NOT NOT1_2799(.VSS(VSS),.VDD(VDD),.Y(g10419),.A(I17373));
  NOT NOT1_2800(.VSS(VSS),.VDD(VDD),.Y(g10424),.A(g7910));
  NOT NOT1_2801(.VSS(VSS),.VDD(VDD),.Y(g10481),.A(g7826));
  NOT NOT1_2802(.VSS(VSS),.VDD(VDD),.Y(I17433),.A(g3900));
  NOT NOT1_2803(.VSS(VSS),.VDD(VDD),.Y(g10482),.A(I17433));
  NOT NOT1_2804(.VSS(VSS),.VDD(VDD),.Y(g10486),.A(g7957));
  NOT NOT1_2805(.VSS(VSS),.VDD(VDD),.Y(g10500),.A(g7962));
  NOT NOT1_2806(.VSS(VSS),.VDD(VDD),.Y(I17483),.A(g3900));
  NOT NOT1_2807(.VSS(VSS),.VDD(VDD),.Y(g10542),.A(I17483));
  NOT NOT1_2808(.VSS(VSS),.VDD(VDD),.Y(I17486),.A(g3900));
  NOT NOT1_2809(.VSS(VSS),.VDD(VDD),.Y(g10545),.A(I17486));
  NOT NOT1_2810(.VSS(VSS),.VDD(VDD),.Y(g10549),.A(g7999));
  NOT NOT1_2811(.VSS(VSS),.VDD(VDD),.Y(g10560),.A(g8008));
  NOT NOT1_2812(.VSS(VSS),.VDD(VDD),.Y(g10574),.A(g8013));
  NOT NOT1_2813(.VSS(VSS),.VDD(VDD),.Y(I17527),.A(g3900));
  NOT NOT1_2814(.VSS(VSS),.VDD(VDD),.Y(g10601),.A(I17527));
  NOT NOT1_2815(.VSS(VSS),.VDD(VDD),.Y(g10606),.A(g8074));
  NOT NOT1_2816(.VSS(VSS),.VDD(VDD),.Y(g10617),.A(g8083));
  NOT NOT1_2817(.VSS(VSS),.VDD(VDD),.Y(g10631),.A(g8088));
  NOT NOT1_2818(.VSS(VSS),.VDD(VDD),.Y(I17557),.A(g3900));
  NOT NOT1_2819(.VSS(VSS),.VDD(VDD),.Y(g10646),.A(I17557));
  NOT NOT1_2820(.VSS(VSS),.VDD(VDD),.Y(g10653),.A(g8159));
  NOT NOT1_2821(.VSS(VSS),.VDD(VDD),.Y(g10664),.A(g8168));
  NOT NOT1_2822(.VSS(VSS),.VDD(VDD),.Y(g10683),.A(g8245));
  NOT NOT1_2823(.VSS(VSS),.VDD(VDD),.Y(g10694),.A(g4326));
  NOT NOT1_2824(.VSS(VSS),.VDD(VDD),.Y(g10714),.A(g4495));
  NOT NOT1_2825(.VSS(VSS),.VDD(VDD),.Y(g10730),.A(g6173));
  NOT NOT1_2826(.VSS(VSS),.VDD(VDD),.Y(g10735),.A(g4671));
  NOT NOT1_2827(.VSS(VSS),.VDD(VDD),.Y(g10749),.A(g6205));
  NOT NOT1_2828(.VSS(VSS),.VDD(VDD),.Y(g10754),.A(g4848));
  NOT NOT1_2829(.VSS(VSS),.VDD(VDD),.Y(g10765),.A(g6048));
  NOT NOT1_2830(.VSS(VSS),.VDD(VDD),.Y(g10766),.A(g6676));
  NOT NOT1_2831(.VSS(VSS),.VDD(VDD),.Y(g10767),.A(g6294));
  NOT NOT1_2832(.VSS(VSS),.VDD(VDD),.Y(g10772),.A(g6978));
  NOT NOT1_2833(.VSS(VSS),.VDD(VDD),.Y(g10773),.A(g6431));
  NOT NOT1_2834(.VSS(VSS),.VDD(VDD),.Y(I17627),.A(g7575));
  NOT NOT1_2835(.VSS(VSS),.VDD(VDD),.Y(g10779),.A(I17627));
  NOT NOT1_2836(.VSS(VSS),.VDD(VDD),.Y(g10783),.A(g7228));
  NOT NOT1_2837(.VSS(VSS),.VDD(VDD),.Y(I17632),.A(g6183));
  NOT NOT1_2838(.VSS(VSS),.VDD(VDD),.Y(g10787),.A(I17632));
  NOT NOT1_2839(.VSS(VSS),.VDD(VDD),.Y(g10788),.A(g7424));
  NOT NOT1_2840(.VSS(VSS),.VDD(VDD),.Y(I17637),.A(g6204));
  NOT NOT1_2841(.VSS(VSS),.VDD(VDD),.Y(g10792),.A(I17637));
  NOT NOT1_2842(.VSS(VSS),.VDD(VDD),.Y(I17641),.A(g6215));
  NOT NOT1_2843(.VSS(VSS),.VDD(VDD),.Y(g10796),.A(I17641));
  NOT NOT1_2844(.VSS(VSS),.VDD(VDD),.Y(I17645),.A(g6288));
  NOT NOT1_2845(.VSS(VSS),.VDD(VDD),.Y(g10800),.A(I17645));
  NOT NOT1_2846(.VSS(VSS),.VDD(VDD),.Y(I17649),.A(g6293));
  NOT NOT1_2847(.VSS(VSS),.VDD(VDD),.Y(g10804),.A(I17649));
  NOT NOT1_2848(.VSS(VSS),.VDD(VDD),.Y(I17653),.A(g6304));
  NOT NOT1_2849(.VSS(VSS),.VDD(VDD),.Y(g10808),.A(I17653));
  NOT NOT1_2850(.VSS(VSS),.VDD(VDD),.Y(g10809),.A(g5701));
  NOT NOT1_2851(.VSS(VSS),.VDD(VDD),.Y(I17658),.A(g6367));
  NOT NOT1_2852(.VSS(VSS),.VDD(VDD),.Y(g10813),.A(I17658));
  NOT NOT1_2853(.VSS(VSS),.VDD(VDD),.Y(I17662),.A(g6425));
  NOT NOT1_2854(.VSS(VSS),.VDD(VDD),.Y(g10817),.A(I17662));
  NOT NOT1_2855(.VSS(VSS),.VDD(VDD),.Y(I17666),.A(g6430));
  NOT NOT1_2856(.VSS(VSS),.VDD(VDD),.Y(g10821),.A(I17666));
  NOT NOT1_2857(.VSS(VSS),.VDD(VDD),.Y(I17670),.A(g6441));
  NOT NOT1_2858(.VSS(VSS),.VDD(VDD),.Y(g10825),.A(I17670));
  NOT NOT1_2859(.VSS(VSS),.VDD(VDD),.Y(I17673),.A(g8107));
  NOT NOT1_2860(.VSS(VSS),.VDD(VDD),.Y(g10826),.A(I17673));
  NOT NOT1_2861(.VSS(VSS),.VDD(VDD),.Y(g10829),.A(g5749));
  NOT NOT1_2862(.VSS(VSS),.VDD(VDD),.Y(I17677),.A(g6517));
  NOT NOT1_2863(.VSS(VSS),.VDD(VDD),.Y(g10830),.A(I17677));
  NOT NOT1_2864(.VSS(VSS),.VDD(VDD),.Y(I17681),.A(g6572));
  NOT NOT1_2865(.VSS(VSS),.VDD(VDD),.Y(g10834),.A(I17681));
  NOT NOT1_2866(.VSS(VSS),.VDD(VDD),.Y(I17685),.A(g6630));
  NOT NOT1_2867(.VSS(VSS),.VDD(VDD),.Y(g10838),.A(I17685));
  NOT NOT1_2868(.VSS(VSS),.VDD(VDD),.Y(I17689),.A(g6635));
  NOT NOT1_2869(.VSS(VSS),.VDD(VDD),.Y(g10842),.A(I17689));
  NOT NOT1_2870(.VSS(VSS),.VDD(VDD),.Y(I17692),.A(g8107));
  NOT NOT1_2871(.VSS(VSS),.VDD(VDD),.Y(g10843),.A(I17692));
  NOT NOT1_2872(.VSS(VSS),.VDD(VDD),.Y(g10846),.A(g5799));
  NOT NOT1_2873(.VSS(VSS),.VDD(VDD),.Y(g10847),.A(g5800));
  NOT NOT1_2874(.VSS(VSS),.VDD(VDD),.Y(g10848),.A(g5801));
  NOT NOT1_2875(.VSS(VSS),.VDD(VDD),.Y(I17698),.A(g6711));
  NOT NOT1_2876(.VSS(VSS),.VDD(VDD),.Y(g10849),.A(I17698));
  NOT NOT1_2877(.VSS(VSS),.VDD(VDD),.Y(I17701),.A(g6781));
  NOT NOT1_2878(.VSS(VSS),.VDD(VDD),.Y(g10850),.A(I17701));
  NOT NOT1_2879(.VSS(VSS),.VDD(VDD),.Y(I17705),.A(g6836));
  NOT NOT1_2880(.VSS(VSS),.VDD(VDD),.Y(g10854),.A(I17705));
  NOT NOT1_2881(.VSS(VSS),.VDD(VDD),.Y(I17709),.A(g6894));
  NOT NOT1_2882(.VSS(VSS),.VDD(VDD),.Y(g10858),.A(I17709));
  NOT NOT1_2883(.VSS(VSS),.VDD(VDD),.Y(I17712),.A(g8031));
  NOT NOT1_2884(.VSS(VSS),.VDD(VDD),.Y(g10859),.A(I17712));
  NOT NOT1_2885(.VSS(VSS),.VDD(VDD),.Y(I17715),.A(g8107));
  NOT NOT1_2886(.VSS(VSS),.VDD(VDD),.Y(g10862),.A(I17715));
  NOT NOT1_2887(.VSS(VSS),.VDD(VDD),.Y(g10865),.A(g6131));
  NOT NOT1_2888(.VSS(VSS),.VDD(VDD),.Y(g10866),.A(g5849));
  NOT NOT1_2889(.VSS(VSS),.VDD(VDD),.Y(g10867),.A(g5850));
  NOT NOT1_2890(.VSS(VSS),.VDD(VDD),.Y(I17721),.A(g6641));
  NOT NOT1_2891(.VSS(VSS),.VDD(VDD),.Y(g10868),.A(I17721));
  NOT NOT1_2892(.VSS(VSS),.VDD(VDD),.Y(I17724),.A(g6942));
  NOT NOT1_2893(.VSS(VSS),.VDD(VDD),.Y(g10869),.A(I17724));
  NOT NOT1_2894(.VSS(VSS),.VDD(VDD),.Y(I17727),.A(g7013));
  NOT NOT1_2895(.VSS(VSS),.VDD(VDD),.Y(g10870),.A(I17727));
  NOT NOT1_2896(.VSS(VSS),.VDD(VDD),.Y(I17730),.A(g7083));
  NOT NOT1_2897(.VSS(VSS),.VDD(VDD),.Y(g10871),.A(I17730));
  NOT NOT1_2898(.VSS(VSS),.VDD(VDD),.Y(I17734),.A(g7138));
  NOT NOT1_2899(.VSS(VSS),.VDD(VDD),.Y(g10875),.A(I17734));
  NOT NOT1_2900(.VSS(VSS),.VDD(VDD),.Y(I17737),.A(g6000));
  NOT NOT1_2901(.VSS(VSS),.VDD(VDD),.Y(g10876),.A(I17737));
  NOT NOT1_2902(.VSS(VSS),.VDD(VDD),.Y(I17740),.A(g8031));
  NOT NOT1_2903(.VSS(VSS),.VDD(VDD),.Y(g10877),.A(I17740));
  NOT NOT1_2904(.VSS(VSS),.VDD(VDD),.Y(I17743),.A(g8107));
  NOT NOT1_2905(.VSS(VSS),.VDD(VDD),.Y(g10880),.A(I17743));
  NOT NOT1_2906(.VSS(VSS),.VDD(VDD),.Y(I17746),.A(g8107));
  NOT NOT1_2907(.VSS(VSS),.VDD(VDD),.Y(g10883),.A(I17746));
  NOT NOT1_2908(.VSS(VSS),.VDD(VDD),.Y(g10886),.A(g5889));
  NOT NOT1_2909(.VSS(VSS),.VDD(VDD),.Y(I17750),.A(g7157));
  NOT NOT1_2910(.VSS(VSS),.VDD(VDD),.Y(g10887),.A(I17750));
  NOT NOT1_2911(.VSS(VSS),.VDD(VDD),.Y(I17753),.A(g6943));
  NOT NOT1_2912(.VSS(VSS),.VDD(VDD),.Y(g10888),.A(I17753));
  NOT NOT1_2913(.VSS(VSS),.VDD(VDD),.Y(I17756),.A(g7192));
  NOT NOT1_2914(.VSS(VSS),.VDD(VDD),.Y(g10889),.A(I17756));
  NOT NOT1_2915(.VSS(VSS),.VDD(VDD),.Y(I17759),.A(g7263));
  NOT NOT1_2916(.VSS(VSS),.VDD(VDD),.Y(g10890),.A(I17759));
  NOT NOT1_2917(.VSS(VSS),.VDD(VDD),.Y(I17762),.A(g7333));
  NOT NOT1_2918(.VSS(VSS),.VDD(VDD),.Y(g10891),.A(I17762));
  NOT NOT1_2919(.VSS(VSS),.VDD(VDD),.Y(I17765),.A(g7976));
  NOT NOT1_2920(.VSS(VSS),.VDD(VDD),.Y(g10892),.A(I17765));
  NOT NOT1_2921(.VSS(VSS),.VDD(VDD),.Y(I17768),.A(g8031));
  NOT NOT1_2922(.VSS(VSS),.VDD(VDD),.Y(g10895),.A(I17768));
  NOT NOT1_2923(.VSS(VSS),.VDD(VDD),.Y(I17771),.A(g8107));
  NOT NOT1_2924(.VSS(VSS),.VDD(VDD),.Y(g10898),.A(I17771));
  NOT NOT1_2925(.VSS(VSS),.VDD(VDD),.Y(I17774),.A(g8107));
  NOT NOT1_2926(.VSS(VSS),.VDD(VDD),.Y(g10901),.A(I17774));
  NOT NOT1_2927(.VSS(VSS),.VDD(VDD),.Y(g10904),.A(g5922));
  NOT NOT1_2928(.VSS(VSS),.VDD(VDD),.Y(g10905),.A(g5923));
  NOT NOT1_2929(.VSS(VSS),.VDD(VDD),.Y(g10906),.A(g5924));
  NOT NOT1_2930(.VSS(VSS),.VDD(VDD),.Y(I17780),.A(g7348));
  NOT NOT1_2931(.VSS(VSS),.VDD(VDD),.Y(g10907),.A(I17780));
  NOT NOT1_2932(.VSS(VSS),.VDD(VDD),.Y(I17783),.A(g7353));
  NOT NOT1_2933(.VSS(VSS),.VDD(VDD),.Y(g10908),.A(I17783));
  NOT NOT1_2934(.VSS(VSS),.VDD(VDD),.Y(I17786),.A(g7193));
  NOT NOT1_2935(.VSS(VSS),.VDD(VDD),.Y(g10909),.A(I17786));
  NOT NOT1_2936(.VSS(VSS),.VDD(VDD),.Y(I17789),.A(g7388));
  NOT NOT1_2937(.VSS(VSS),.VDD(VDD),.Y(g10910),.A(I17789));
  NOT NOT1_2938(.VSS(VSS),.VDD(VDD),.Y(I17792),.A(g7459));
  NOT NOT1_2939(.VSS(VSS),.VDD(VDD),.Y(g10911),.A(I17792));
  NOT NOT1_2940(.VSS(VSS),.VDD(VDD),.Y(I17795),.A(g7976));
  NOT NOT1_2941(.VSS(VSS),.VDD(VDD),.Y(g10912),.A(I17795));
  NOT NOT1_2942(.VSS(VSS),.VDD(VDD),.Y(I17798),.A(g8031));
  NOT NOT1_2943(.VSS(VSS),.VDD(VDD),.Y(g10915),.A(I17798));
  NOT NOT1_2944(.VSS(VSS),.VDD(VDD),.Y(I17801),.A(g8107));
  NOT NOT1_2945(.VSS(VSS),.VDD(VDD),.Y(g10918),.A(I17801));
  NOT NOT1_2946(.VSS(VSS),.VDD(VDD),.Y(I17804),.A(g8031));
  NOT NOT1_2947(.VSS(VSS),.VDD(VDD),.Y(g10921),.A(I17804));
  NOT NOT1_2948(.VSS(VSS),.VDD(VDD),.Y(I17807),.A(g8107));
  NOT NOT1_2949(.VSS(VSS),.VDD(VDD),.Y(g10924),.A(I17807));
  NOT NOT1_2950(.VSS(VSS),.VDD(VDD),.Y(g10927),.A(g6153));
  NOT NOT1_2951(.VSS(VSS),.VDD(VDD),.Y(g10928),.A(g5951));
  NOT NOT1_2952(.VSS(VSS),.VDD(VDD),.Y(g10929),.A(g5952));
  NOT NOT1_2953(.VSS(VSS),.VDD(VDD),.Y(I17813),.A(g5707));
  NOT NOT1_2954(.VSS(VSS),.VDD(VDD),.Y(g10930),.A(I17813));
  NOT NOT1_2955(.VSS(VSS),.VDD(VDD),.Y(I17816),.A(g7346));
  NOT NOT1_2956(.VSS(VSS),.VDD(VDD),.Y(g10931),.A(I17816));
  NOT NOT1_2957(.VSS(VSS),.VDD(VDD),.Y(I17819),.A(g6448));
  NOT NOT1_2958(.VSS(VSS),.VDD(VDD),.Y(g10932),.A(I17819));
  NOT NOT1_2959(.VSS(VSS),.VDD(VDD),.Y(I17822),.A(g7478));
  NOT NOT1_2960(.VSS(VSS),.VDD(VDD),.Y(g10933),.A(I17822));
  NOT NOT1_2961(.VSS(VSS),.VDD(VDD),.Y(I17825),.A(g7483));
  NOT NOT1_2962(.VSS(VSS),.VDD(VDD),.Y(g10934),.A(I17825));
  NOT NOT1_2963(.VSS(VSS),.VDD(VDD),.Y(I17828),.A(g7389));
  NOT NOT1_2964(.VSS(VSS),.VDD(VDD),.Y(g10935),.A(I17828));
  NOT NOT1_2965(.VSS(VSS),.VDD(VDD),.Y(I17831),.A(g7518));
  NOT NOT1_2966(.VSS(VSS),.VDD(VDD),.Y(g10936),.A(I17831));
  NOT NOT1_2967(.VSS(VSS),.VDD(VDD),.Y(I17834),.A(g7976));
  NOT NOT1_2968(.VSS(VSS),.VDD(VDD),.Y(g10937),.A(I17834));
  NOT NOT1_2969(.VSS(VSS),.VDD(VDD),.Y(I17837),.A(g8031));
  NOT NOT1_2970(.VSS(VSS),.VDD(VDD),.Y(g10940),.A(I17837));
  NOT NOT1_2971(.VSS(VSS),.VDD(VDD),.Y(I17840),.A(g8107));
  NOT NOT1_2972(.VSS(VSS),.VDD(VDD),.Y(g10943),.A(I17840));
  NOT NOT1_2973(.VSS(VSS),.VDD(VDD),.Y(I17843),.A(g8031));
  NOT NOT1_2974(.VSS(VSS),.VDD(VDD),.Y(g10946),.A(I17843));
  NOT NOT1_2975(.VSS(VSS),.VDD(VDD),.Y(I17846),.A(g8107));
  NOT NOT1_2976(.VSS(VSS),.VDD(VDD),.Y(g10949),.A(I17846));
  NOT NOT1_2977(.VSS(VSS),.VDD(VDD),.Y(I17849),.A(g8103));
  NOT NOT1_2978(.VSS(VSS),.VDD(VDD),.Y(g10952),.A(I17849));
  NOT NOT1_2979(.VSS(VSS),.VDD(VDD),.Y(g10961),.A(g5978));
  NOT NOT1_2980(.VSS(VSS),.VDD(VDD),.Y(g10962),.A(g5979));
  NOT NOT1_2981(.VSS(VSS),.VDD(VDD),.Y(I17854),.A(g6232));
  NOT NOT1_2982(.VSS(VSS),.VDD(VDD),.Y(g10963),.A(I17854));
  NOT NOT1_2983(.VSS(VSS),.VDD(VDD),.Y(I17857),.A(g6448));
  NOT NOT1_2984(.VSS(VSS),.VDD(VDD),.Y(g10966),.A(I17857));
  NOT NOT1_2985(.VSS(VSS),.VDD(VDD),.Y(I17860),.A(g5765));
  NOT NOT1_2986(.VSS(VSS),.VDD(VDD),.Y(g10967),.A(I17860));
  NOT NOT1_2987(.VSS(VSS),.VDD(VDD),.Y(I17863),.A(g7476));
  NOT NOT1_2988(.VSS(VSS),.VDD(VDD),.Y(g10968),.A(I17863));
  NOT NOT1_2989(.VSS(VSS),.VDD(VDD),.Y(I17866),.A(g6713));
  NOT NOT1_2990(.VSS(VSS),.VDD(VDD),.Y(g10969),.A(I17866));
  NOT NOT1_2991(.VSS(VSS),.VDD(VDD),.Y(I17869),.A(g7534));
  NOT NOT1_2992(.VSS(VSS),.VDD(VDD),.Y(g10972),.A(I17869));
  NOT NOT1_2993(.VSS(VSS),.VDD(VDD),.Y(I17872),.A(g7539));
  NOT NOT1_2994(.VSS(VSS),.VDD(VDD),.Y(g10973),.A(I17872));
  NOT NOT1_2995(.VSS(VSS),.VDD(VDD),.Y(I17875),.A(g7976));
  NOT NOT1_2996(.VSS(VSS),.VDD(VDD),.Y(g10974),.A(I17875));
  NOT NOT1_2997(.VSS(VSS),.VDD(VDD),.Y(I17878),.A(g8031));
  NOT NOT1_2998(.VSS(VSS),.VDD(VDD),.Y(g10977),.A(I17878));
  NOT NOT1_2999(.VSS(VSS),.VDD(VDD),.Y(I17881),.A(g7976));
  NOT NOT1_3000(.VSS(VSS),.VDD(VDD),.Y(g10980),.A(I17881));
  NOT NOT1_3001(.VSS(VSS),.VDD(VDD),.Y(I17884),.A(g8031));
  NOT NOT1_3002(.VSS(VSS),.VDD(VDD),.Y(g10983),.A(I17884));
  NOT NOT1_3003(.VSS(VSS),.VDD(VDD),.Y(g10986),.A(g6014));
  NOT NOT1_3004(.VSS(VSS),.VDD(VDD),.Y(g10987),.A(g6015));
  NOT NOT1_3005(.VSS(VSS),.VDD(VDD),.Y(I17889),.A(g6314));
  NOT NOT1_3006(.VSS(VSS),.VDD(VDD),.Y(g10988),.A(I17889));
  NOT NOT1_3007(.VSS(VSS),.VDD(VDD),.Y(I17892),.A(g6232));
  NOT NOT1_3008(.VSS(VSS),.VDD(VDD),.Y(g10991),.A(I17892));
  NOT NOT1_3009(.VSS(VSS),.VDD(VDD),.Y(I17895),.A(g6448));
  NOT NOT1_3010(.VSS(VSS),.VDD(VDD),.Y(g10994),.A(I17895));
  NOT NOT1_3011(.VSS(VSS),.VDD(VDD),.Y(I17898),.A(g6643));
  NOT NOT1_3012(.VSS(VSS),.VDD(VDD),.Y(g10995),.A(I17898));
  NOT NOT1_3013(.VSS(VSS),.VDD(VDD),.Y(I17901),.A(g6369));
  NOT NOT1_3014(.VSS(VSS),.VDD(VDD),.Y(g10996),.A(I17901));
  NOT NOT1_3015(.VSS(VSS),.VDD(VDD),.Y(I17904),.A(g6713));
  NOT NOT1_3016(.VSS(VSS),.VDD(VDD),.Y(g10999),.A(I17904));
  NOT NOT1_3017(.VSS(VSS),.VDD(VDD),.Y(I17907),.A(g5824));
  NOT NOT1_3018(.VSS(VSS),.VDD(VDD),.Y(g11002),.A(I17907));
  NOT NOT1_3019(.VSS(VSS),.VDD(VDD),.Y(I17910),.A(g7532));
  NOT NOT1_3020(.VSS(VSS),.VDD(VDD),.Y(g11003),.A(I17910));
  NOT NOT1_3021(.VSS(VSS),.VDD(VDD),.Y(I17913),.A(g7015));
  NOT NOT1_3022(.VSS(VSS),.VDD(VDD),.Y(g11004),.A(I17913));
  NOT NOT1_3023(.VSS(VSS),.VDD(VDD),.Y(I17916),.A(g7560));
  NOT NOT1_3024(.VSS(VSS),.VDD(VDD),.Y(g11007),.A(I17916));
  NOT NOT1_3025(.VSS(VSS),.VDD(VDD),.Y(I17919),.A(g7976));
  NOT NOT1_3026(.VSS(VSS),.VDD(VDD),.Y(g11008),.A(I17919));
  NOT NOT1_3027(.VSS(VSS),.VDD(VDD),.Y(I17922),.A(g8031));
  NOT NOT1_3028(.VSS(VSS),.VDD(VDD),.Y(g11011),.A(I17922));
  NOT NOT1_3029(.VSS(VSS),.VDD(VDD),.Y(I17925),.A(g7976));
  NOT NOT1_3030(.VSS(VSS),.VDD(VDD),.Y(g11014),.A(I17925));
  NOT NOT1_3031(.VSS(VSS),.VDD(VDD),.Y(I17928),.A(g8031));
  NOT NOT1_3032(.VSS(VSS),.VDD(VDD),.Y(g11017),.A(I17928));
  NOT NOT1_3033(.VSS(VSS),.VDD(VDD),.Y(g11020),.A(g6029));
  NOT NOT1_3034(.VSS(VSS),.VDD(VDD),.Y(g11021),.A(g6030));
  NOT NOT1_3035(.VSS(VSS),.VDD(VDD),.Y(I17933),.A(g3254));
  NOT NOT1_3036(.VSS(VSS),.VDD(VDD),.Y(g11022),.A(I17933));
  NOT NOT1_3037(.VSS(VSS),.VDD(VDD),.Y(I17936),.A(g6314));
  NOT NOT1_3038(.VSS(VSS),.VDD(VDD),.Y(g11025),.A(I17936));
  NOT NOT1_3039(.VSS(VSS),.VDD(VDD),.Y(I17939),.A(g6232));
  NOT NOT1_3040(.VSS(VSS),.VDD(VDD),.Y(g11028),.A(I17939));
  NOT NOT1_3041(.VSS(VSS),.VDD(VDD),.Y(I17942),.A(g5548));
  NOT NOT1_3042(.VSS(VSS),.VDD(VDD),.Y(g11031),.A(I17942));
  NOT NOT1_3043(.VSS(VSS),.VDD(VDD),.Y(I17945),.A(g5668));
  NOT NOT1_3044(.VSS(VSS),.VDD(VDD),.Y(g11032),.A(I17945));
  NOT NOT1_3045(.VSS(VSS),.VDD(VDD),.Y(I17948),.A(g6643));
  NOT NOT1_3046(.VSS(VSS),.VDD(VDD),.Y(g11035),.A(I17948));
  NOT NOT1_3047(.VSS(VSS),.VDD(VDD),.Y(I17951),.A(g6519));
  NOT NOT1_3048(.VSS(VSS),.VDD(VDD),.Y(g11036),.A(I17951));
  NOT NOT1_3049(.VSS(VSS),.VDD(VDD),.Y(I17954),.A(g6369));
  NOT NOT1_3050(.VSS(VSS),.VDD(VDD),.Y(g11039),.A(I17954));
  NOT NOT1_3051(.VSS(VSS),.VDD(VDD),.Y(I17957),.A(g6713));
  NOT NOT1_3052(.VSS(VSS),.VDD(VDD),.Y(g11042),.A(I17957));
  NOT NOT1_3053(.VSS(VSS),.VDD(VDD),.Y(I17960),.A(g6945));
  NOT NOT1_3054(.VSS(VSS),.VDD(VDD),.Y(g11045),.A(I17960));
  NOT NOT1_3055(.VSS(VSS),.VDD(VDD),.Y(I17963),.A(g6574));
  NOT NOT1_3056(.VSS(VSS),.VDD(VDD),.Y(g11048),.A(I17963));
  NOT NOT1_3057(.VSS(VSS),.VDD(VDD),.Y(I17966),.A(g7015));
  NOT NOT1_3058(.VSS(VSS),.VDD(VDD),.Y(g11051),.A(I17966));
  NOT NOT1_3059(.VSS(VSS),.VDD(VDD),.Y(I17969),.A(g5880));
  NOT NOT1_3060(.VSS(VSS),.VDD(VDD),.Y(g11054),.A(I17969));
  NOT NOT1_3061(.VSS(VSS),.VDD(VDD),.Y(I17972),.A(g7558));
  NOT NOT1_3062(.VSS(VSS),.VDD(VDD),.Y(g11055),.A(I17972));
  NOT NOT1_3063(.VSS(VSS),.VDD(VDD),.Y(I17975),.A(g7265));
  NOT NOT1_3064(.VSS(VSS),.VDD(VDD),.Y(g11056),.A(I17975));
  NOT NOT1_3065(.VSS(VSS),.VDD(VDD),.Y(I17978),.A(g7795));
  NOT NOT1_3066(.VSS(VSS),.VDD(VDD),.Y(g11059),.A(I17978));
  NOT NOT1_3067(.VSS(VSS),.VDD(VDD),.Y(I17981),.A(g7976));
  NOT NOT1_3068(.VSS(VSS),.VDD(VDD),.Y(g11063),.A(I17981));
  NOT NOT1_3069(.VSS(VSS),.VDD(VDD),.Y(I17984),.A(g7976));
  NOT NOT1_3070(.VSS(VSS),.VDD(VDD),.Y(g11066),.A(I17984));
  NOT NOT1_3071(.VSS(VSS),.VDD(VDD),.Y(g11069),.A(g8257));
  NOT NOT1_3072(.VSS(VSS),.VDD(VDD),.Y(g11078),.A(g6041));
  NOT NOT1_3073(.VSS(VSS),.VDD(VDD),.Y(I17989),.A(g3254));
  NOT NOT1_3074(.VSS(VSS),.VDD(VDD),.Y(g11079),.A(I17989));
  NOT NOT1_3075(.VSS(VSS),.VDD(VDD),.Y(I17992),.A(g6314));
  NOT NOT1_3076(.VSS(VSS),.VDD(VDD),.Y(g11082),.A(I17992));
  NOT NOT1_3077(.VSS(VSS),.VDD(VDD),.Y(I17995),.A(g6232));
  NOT NOT1_3078(.VSS(VSS),.VDD(VDD),.Y(g11085),.A(I17995));
  NOT NOT1_3079(.VSS(VSS),.VDD(VDD),.Y(I17998),.A(g5668));
  NOT NOT1_3080(.VSS(VSS),.VDD(VDD),.Y(g11088),.A(I17998));
  NOT NOT1_3081(.VSS(VSS),.VDD(VDD),.Y(I18001),.A(g6643));
  NOT NOT1_3082(.VSS(VSS),.VDD(VDD),.Y(g11091),.A(I18001));
  NOT NOT1_3083(.VSS(VSS),.VDD(VDD),.Y(I18004),.A(g3410));
  NOT NOT1_3084(.VSS(VSS),.VDD(VDD),.Y(g11092),.A(I18004));
  NOT NOT1_3085(.VSS(VSS),.VDD(VDD),.Y(I18007),.A(g6519));
  NOT NOT1_3086(.VSS(VSS),.VDD(VDD),.Y(g11095),.A(I18007));
  NOT NOT1_3087(.VSS(VSS),.VDD(VDD),.Y(I18010),.A(g6369));
  NOT NOT1_3088(.VSS(VSS),.VDD(VDD),.Y(g11098),.A(I18010));
  NOT NOT1_3089(.VSS(VSS),.VDD(VDD),.Y(I18013),.A(g5594));
  NOT NOT1_3090(.VSS(VSS),.VDD(VDD),.Y(g11101),.A(I18013));
  NOT NOT1_3091(.VSS(VSS),.VDD(VDD),.Y(I18016),.A(g5720));
  NOT NOT1_3092(.VSS(VSS),.VDD(VDD),.Y(g11102),.A(I18016));
  NOT NOT1_3093(.VSS(VSS),.VDD(VDD),.Y(I18019),.A(g6945));
  NOT NOT1_3094(.VSS(VSS),.VDD(VDD),.Y(g11105),.A(I18019));
  NOT NOT1_3095(.VSS(VSS),.VDD(VDD),.Y(I18022),.A(g6783));
  NOT NOT1_3096(.VSS(VSS),.VDD(VDD),.Y(g11108),.A(I18022));
  NOT NOT1_3097(.VSS(VSS),.VDD(VDD),.Y(I18025),.A(g6574));
  NOT NOT1_3098(.VSS(VSS),.VDD(VDD),.Y(g11111),.A(I18025));
  NOT NOT1_3099(.VSS(VSS),.VDD(VDD),.Y(I18028),.A(g7015));
  NOT NOT1_3100(.VSS(VSS),.VDD(VDD),.Y(g11114),.A(I18028));
  NOT NOT1_3101(.VSS(VSS),.VDD(VDD),.Y(I18031),.A(g7195));
  NOT NOT1_3102(.VSS(VSS),.VDD(VDD),.Y(g11117),.A(I18031));
  NOT NOT1_3103(.VSS(VSS),.VDD(VDD),.Y(I18034),.A(g6838));
  NOT NOT1_3104(.VSS(VSS),.VDD(VDD),.Y(g11120),.A(I18034));
  NOT NOT1_3105(.VSS(VSS),.VDD(VDD),.Y(I18037),.A(g7265));
  NOT NOT1_3106(.VSS(VSS),.VDD(VDD),.Y(g11123),.A(I18037));
  NOT NOT1_3107(.VSS(VSS),.VDD(VDD),.Y(I18040),.A(g7976));
  NOT NOT1_3108(.VSS(VSS),.VDD(VDD),.Y(g11126),.A(I18040));
  NOT NOT1_3109(.VSS(VSS),.VDD(VDD),.Y(I18043),.A(g7976));
  NOT NOT1_3110(.VSS(VSS),.VDD(VDD),.Y(g11129),.A(I18043));
  NOT NOT1_3111(.VSS(VSS),.VDD(VDD),.Y(I18046),.A(g3254));
  NOT NOT1_3112(.VSS(VSS),.VDD(VDD),.Y(g11132),.A(I18046));
  NOT NOT1_3113(.VSS(VSS),.VDD(VDD),.Y(I18049),.A(g6314));
  NOT NOT1_3114(.VSS(VSS),.VDD(VDD),.Y(g11135),.A(I18049));
  NOT NOT1_3115(.VSS(VSS),.VDD(VDD),.Y(I18052),.A(g6232));
  NOT NOT1_3116(.VSS(VSS),.VDD(VDD),.Y(g11138),.A(I18052));
  NOT NOT1_3117(.VSS(VSS),.VDD(VDD),.Y(I18055),.A(g5668));
  NOT NOT1_3118(.VSS(VSS),.VDD(VDD),.Y(g11141),.A(I18055));
  NOT NOT1_3119(.VSS(VSS),.VDD(VDD),.Y(I18058),.A(g6643));
  NOT NOT1_3120(.VSS(VSS),.VDD(VDD),.Y(g11144),.A(I18058));
  NOT NOT1_3121(.VSS(VSS),.VDD(VDD),.Y(I18061),.A(g3410));
  NOT NOT1_3122(.VSS(VSS),.VDD(VDD),.Y(g11145),.A(I18061));
  NOT NOT1_3123(.VSS(VSS),.VDD(VDD),.Y(I18064),.A(g6519));
  NOT NOT1_3124(.VSS(VSS),.VDD(VDD),.Y(g11148),.A(I18064));
  NOT NOT1_3125(.VSS(VSS),.VDD(VDD),.Y(I18067),.A(g6369));
  NOT NOT1_3126(.VSS(VSS),.VDD(VDD),.Y(g11151),.A(I18067));
  NOT NOT1_3127(.VSS(VSS),.VDD(VDD),.Y(I18070),.A(g5720));
  NOT NOT1_3128(.VSS(VSS),.VDD(VDD),.Y(g11154),.A(I18070));
  NOT NOT1_3129(.VSS(VSS),.VDD(VDD),.Y(I18073),.A(g6945));
  NOT NOT1_3130(.VSS(VSS),.VDD(VDD),.Y(g11157),.A(I18073));
  NOT NOT1_3131(.VSS(VSS),.VDD(VDD),.Y(I18076),.A(g3566));
  NOT NOT1_3132(.VSS(VSS),.VDD(VDD),.Y(g11160),.A(I18076));
  NOT NOT1_3133(.VSS(VSS),.VDD(VDD),.Y(I18079),.A(g6783));
  NOT NOT1_3134(.VSS(VSS),.VDD(VDD),.Y(g11163),.A(I18079));
  NOT NOT1_3135(.VSS(VSS),.VDD(VDD),.Y(I18082),.A(g6574));
  NOT NOT1_3136(.VSS(VSS),.VDD(VDD),.Y(g11166),.A(I18082));
  NOT NOT1_3137(.VSS(VSS),.VDD(VDD),.Y(I18085),.A(g5611));
  NOT NOT1_3138(.VSS(VSS),.VDD(VDD),.Y(g11169),.A(I18085));
  NOT NOT1_3139(.VSS(VSS),.VDD(VDD),.Y(I18088),.A(g5778));
  NOT NOT1_3140(.VSS(VSS),.VDD(VDD),.Y(g11170),.A(I18088));
  NOT NOT1_3141(.VSS(VSS),.VDD(VDD),.Y(I18091),.A(g7195));
  NOT NOT1_3142(.VSS(VSS),.VDD(VDD),.Y(g11173),.A(I18091));
  NOT NOT1_3143(.VSS(VSS),.VDD(VDD),.Y(I18094),.A(g7085));
  NOT NOT1_3144(.VSS(VSS),.VDD(VDD),.Y(g11176),.A(I18094));
  NOT NOT1_3145(.VSS(VSS),.VDD(VDD),.Y(I18097),.A(g6838));
  NOT NOT1_3146(.VSS(VSS),.VDD(VDD),.Y(g11179),.A(I18097));
  NOT NOT1_3147(.VSS(VSS),.VDD(VDD),.Y(I18100),.A(g7265));
  NOT NOT1_3148(.VSS(VSS),.VDD(VDD),.Y(g11182),.A(I18100));
  NOT NOT1_3149(.VSS(VSS),.VDD(VDD),.Y(I18103),.A(g7391));
  NOT NOT1_3150(.VSS(VSS),.VDD(VDD),.Y(g11185),.A(I18103));
  NOT NOT1_3151(.VSS(VSS),.VDD(VDD),.Y(g11190),.A(g3999));
  NOT NOT1_3152(.VSS(VSS),.VDD(VDD),.Y(I18121),.A(g3254));
  NOT NOT1_3153(.VSS(VSS),.VDD(VDD),.Y(g11199),.A(I18121));
  NOT NOT1_3154(.VSS(VSS),.VDD(VDD),.Y(I18124),.A(g6314));
  NOT NOT1_3155(.VSS(VSS),.VDD(VDD),.Y(g11202),.A(I18124));
  NOT NOT1_3156(.VSS(VSS),.VDD(VDD),.Y(I18127),.A(g6232));
  NOT NOT1_3157(.VSS(VSS),.VDD(VDD),.Y(g11205),.A(I18127));
  NOT NOT1_3158(.VSS(VSS),.VDD(VDD),.Y(I18130),.A(g5547));
  NOT NOT1_3159(.VSS(VSS),.VDD(VDD),.Y(g11208),.A(I18130));
  NOT NOT1_3160(.VSS(VSS),.VDD(VDD),.Y(I18133),.A(g6448));
  NOT NOT1_3161(.VSS(VSS),.VDD(VDD),.Y(g11209),.A(I18133));
  NOT NOT1_3162(.VSS(VSS),.VDD(VDD),.Y(I18136),.A(g5668));
  NOT NOT1_3163(.VSS(VSS),.VDD(VDD),.Y(g11210),.A(I18136));
  NOT NOT1_3164(.VSS(VSS),.VDD(VDD),.Y(I18139),.A(g6643));
  NOT NOT1_3165(.VSS(VSS),.VDD(VDD),.Y(g11213),.A(I18139));
  NOT NOT1_3166(.VSS(VSS),.VDD(VDD),.Y(I18142),.A(g3410));
  NOT NOT1_3167(.VSS(VSS),.VDD(VDD),.Y(g11216),.A(I18142));
  NOT NOT1_3168(.VSS(VSS),.VDD(VDD),.Y(I18145),.A(g6519));
  NOT NOT1_3169(.VSS(VSS),.VDD(VDD),.Y(g11219),.A(I18145));
  NOT NOT1_3170(.VSS(VSS),.VDD(VDD),.Y(I18148),.A(g6369));
  NOT NOT1_3171(.VSS(VSS),.VDD(VDD),.Y(g11222),.A(I18148));
  NOT NOT1_3172(.VSS(VSS),.VDD(VDD),.Y(I18151),.A(g5720));
  NOT NOT1_3173(.VSS(VSS),.VDD(VDD),.Y(g11225),.A(I18151));
  NOT NOT1_3174(.VSS(VSS),.VDD(VDD),.Y(I18154),.A(g6945));
  NOT NOT1_3175(.VSS(VSS),.VDD(VDD),.Y(g11228),.A(I18154));
  NOT NOT1_3176(.VSS(VSS),.VDD(VDD),.Y(I18157),.A(g3566));
  NOT NOT1_3177(.VSS(VSS),.VDD(VDD),.Y(g11231),.A(I18157));
  NOT NOT1_3178(.VSS(VSS),.VDD(VDD),.Y(I18160),.A(g6783));
  NOT NOT1_3179(.VSS(VSS),.VDD(VDD),.Y(g11234),.A(I18160));
  NOT NOT1_3180(.VSS(VSS),.VDD(VDD),.Y(I18163),.A(g6574));
  NOT NOT1_3181(.VSS(VSS),.VDD(VDD),.Y(g11237),.A(I18163));
  NOT NOT1_3182(.VSS(VSS),.VDD(VDD),.Y(I18166),.A(g5778));
  NOT NOT1_3183(.VSS(VSS),.VDD(VDD),.Y(g11240),.A(I18166));
  NOT NOT1_3184(.VSS(VSS),.VDD(VDD),.Y(I18169),.A(g7195));
  NOT NOT1_3185(.VSS(VSS),.VDD(VDD),.Y(g11243),.A(I18169));
  NOT NOT1_3186(.VSS(VSS),.VDD(VDD),.Y(I18172),.A(g3722));
  NOT NOT1_3187(.VSS(VSS),.VDD(VDD),.Y(g11246),.A(I18172));
  NOT NOT1_3188(.VSS(VSS),.VDD(VDD),.Y(I18175),.A(g7085));
  NOT NOT1_3189(.VSS(VSS),.VDD(VDD),.Y(g11249),.A(I18175));
  NOT NOT1_3190(.VSS(VSS),.VDD(VDD),.Y(I18178),.A(g6838));
  NOT NOT1_3191(.VSS(VSS),.VDD(VDD),.Y(g11252),.A(I18178));
  NOT NOT1_3192(.VSS(VSS),.VDD(VDD),.Y(I18181),.A(g5636));
  NOT NOT1_3193(.VSS(VSS),.VDD(VDD),.Y(g11255),.A(I18181));
  NOT NOT1_3194(.VSS(VSS),.VDD(VDD),.Y(I18184),.A(g5837));
  NOT NOT1_3195(.VSS(VSS),.VDD(VDD),.Y(g11256),.A(I18184));
  NOT NOT1_3196(.VSS(VSS),.VDD(VDD),.Y(I18187),.A(g7391));
  NOT NOT1_3197(.VSS(VSS),.VDD(VDD),.Y(g11259),.A(I18187));
  NOT NOT1_3198(.VSS(VSS),.VDD(VDD),.Y(I18211),.A(g6232));
  NOT NOT1_3199(.VSS(VSS),.VDD(VDD),.Y(g11265),.A(I18211));
  NOT NOT1_3200(.VSS(VSS),.VDD(VDD),.Y(I18214),.A(g3254));
  NOT NOT1_3201(.VSS(VSS),.VDD(VDD),.Y(g11268),.A(I18214));
  NOT NOT1_3202(.VSS(VSS),.VDD(VDD),.Y(I18217),.A(g6314));
  NOT NOT1_3203(.VSS(VSS),.VDD(VDD),.Y(g11271),.A(I18217));
  NOT NOT1_3204(.VSS(VSS),.VDD(VDD),.Y(I18220),.A(g6232));
  NOT NOT1_3205(.VSS(VSS),.VDD(VDD),.Y(g11274),.A(I18220));
  NOT NOT1_3206(.VSS(VSS),.VDD(VDD),.Y(I18223),.A(g6448));
  NOT NOT1_3207(.VSS(VSS),.VDD(VDD),.Y(g11277),.A(I18223));
  NOT NOT1_3208(.VSS(VSS),.VDD(VDD),.Y(I18226),.A(g5668));
  NOT NOT1_3209(.VSS(VSS),.VDD(VDD),.Y(g11278),.A(I18226));
  NOT NOT1_3210(.VSS(VSS),.VDD(VDD),.Y(I18229),.A(g3410));
  NOT NOT1_3211(.VSS(VSS),.VDD(VDD),.Y(g11281),.A(I18229));
  NOT NOT1_3212(.VSS(VSS),.VDD(VDD),.Y(I18232),.A(g6519));
  NOT NOT1_3213(.VSS(VSS),.VDD(VDD),.Y(g11284),.A(I18232));
  NOT NOT1_3214(.VSS(VSS),.VDD(VDD),.Y(I18235),.A(g6369));
  NOT NOT1_3215(.VSS(VSS),.VDD(VDD),.Y(g11287),.A(I18235));
  NOT NOT1_3216(.VSS(VSS),.VDD(VDD),.Y(I18238),.A(g5593));
  NOT NOT1_3217(.VSS(VSS),.VDD(VDD),.Y(g11290),.A(I18238));
  NOT NOT1_3218(.VSS(VSS),.VDD(VDD),.Y(I18241),.A(g6713));
  NOT NOT1_3219(.VSS(VSS),.VDD(VDD),.Y(g11291),.A(I18241));
  NOT NOT1_3220(.VSS(VSS),.VDD(VDD),.Y(I18244),.A(g5720));
  NOT NOT1_3221(.VSS(VSS),.VDD(VDD),.Y(g11294),.A(I18244));
  NOT NOT1_3222(.VSS(VSS),.VDD(VDD),.Y(I18247),.A(g6945));
  NOT NOT1_3223(.VSS(VSS),.VDD(VDD),.Y(g11297),.A(I18247));
  NOT NOT1_3224(.VSS(VSS),.VDD(VDD),.Y(I18250),.A(g3566));
  NOT NOT1_3225(.VSS(VSS),.VDD(VDD),.Y(g11300),.A(I18250));
  NOT NOT1_3226(.VSS(VSS),.VDD(VDD),.Y(I18253),.A(g6783));
  NOT NOT1_3227(.VSS(VSS),.VDD(VDD),.Y(g11303),.A(I18253));
  NOT NOT1_3228(.VSS(VSS),.VDD(VDD),.Y(I18256),.A(g6574));
  NOT NOT1_3229(.VSS(VSS),.VDD(VDD),.Y(g11306),.A(I18256));
  NOT NOT1_3230(.VSS(VSS),.VDD(VDD),.Y(I18259),.A(g5778));
  NOT NOT1_3231(.VSS(VSS),.VDD(VDD),.Y(g11309),.A(I18259));
  NOT NOT1_3232(.VSS(VSS),.VDD(VDD),.Y(I18262),.A(g7195));
  NOT NOT1_3233(.VSS(VSS),.VDD(VDD),.Y(g11312),.A(I18262));
  NOT NOT1_3234(.VSS(VSS),.VDD(VDD),.Y(I18265),.A(g3722));
  NOT NOT1_3235(.VSS(VSS),.VDD(VDD),.Y(g11315),.A(I18265));
  NOT NOT1_3236(.VSS(VSS),.VDD(VDD),.Y(I18268),.A(g7085));
  NOT NOT1_3237(.VSS(VSS),.VDD(VDD),.Y(g11318),.A(I18268));
  NOT NOT1_3238(.VSS(VSS),.VDD(VDD),.Y(I18271),.A(g6838));
  NOT NOT1_3239(.VSS(VSS),.VDD(VDD),.Y(g11321),.A(I18271));
  NOT NOT1_3240(.VSS(VSS),.VDD(VDD),.Y(I18274),.A(g5837));
  NOT NOT1_3241(.VSS(VSS),.VDD(VDD),.Y(g11324),.A(I18274));
  NOT NOT1_3242(.VSS(VSS),.VDD(VDD),.Y(I18277),.A(g7391));
  NOT NOT1_3243(.VSS(VSS),.VDD(VDD),.Y(g11327),.A(I18277));
  NOT NOT1_3244(.VSS(VSS),.VDD(VDD),.Y(g11332),.A(g4094));
  NOT NOT1_3245(.VSS(VSS),.VDD(VDD),.Y(I18295),.A(g6314));
  NOT NOT1_3246(.VSS(VSS),.VDD(VDD),.Y(g11341),.A(I18295));
  NOT NOT1_3247(.VSS(VSS),.VDD(VDD),.Y(I18298),.A(g6232));
  NOT NOT1_3248(.VSS(VSS),.VDD(VDD),.Y(g11344),.A(I18298));
  NOT NOT1_3249(.VSS(VSS),.VDD(VDD),.Y(I18302),.A(g3254));
  NOT NOT1_3250(.VSS(VSS),.VDD(VDD),.Y(g11348),.A(I18302));
  NOT NOT1_3251(.VSS(VSS),.VDD(VDD),.Y(I18305),.A(g6314));
  NOT NOT1_3252(.VSS(VSS),.VDD(VDD),.Y(g11351),.A(I18305));
  NOT NOT1_3253(.VSS(VSS),.VDD(VDD),.Y(I18308),.A(g6448));
  NOT NOT1_3254(.VSS(VSS),.VDD(VDD),.Y(g11354),.A(I18308));
  NOT NOT1_3255(.VSS(VSS),.VDD(VDD),.Y(I18311),.A(g5668));
  NOT NOT1_3256(.VSS(VSS),.VDD(VDD),.Y(g11355),.A(I18311));
  NOT NOT1_3257(.VSS(VSS),.VDD(VDD),.Y(I18314),.A(g6369));
  NOT NOT1_3258(.VSS(VSS),.VDD(VDD),.Y(g11358),.A(I18314));
  NOT NOT1_3259(.VSS(VSS),.VDD(VDD),.Y(I18317),.A(g3410));
  NOT NOT1_3260(.VSS(VSS),.VDD(VDD),.Y(g11361),.A(I18317));
  NOT NOT1_3261(.VSS(VSS),.VDD(VDD),.Y(I18320),.A(g6519));
  NOT NOT1_3262(.VSS(VSS),.VDD(VDD),.Y(g11364),.A(I18320));
  NOT NOT1_3263(.VSS(VSS),.VDD(VDD),.Y(I18323),.A(g6369));
  NOT NOT1_3264(.VSS(VSS),.VDD(VDD),.Y(g11367),.A(I18323));
  NOT NOT1_3265(.VSS(VSS),.VDD(VDD),.Y(I18326),.A(g6713));
  NOT NOT1_3266(.VSS(VSS),.VDD(VDD),.Y(g11370),.A(I18326));
  NOT NOT1_3267(.VSS(VSS),.VDD(VDD),.Y(I18329),.A(g5720));
  NOT NOT1_3268(.VSS(VSS),.VDD(VDD),.Y(g11373),.A(I18329));
  NOT NOT1_3269(.VSS(VSS),.VDD(VDD),.Y(I18332),.A(g3566));
  NOT NOT1_3270(.VSS(VSS),.VDD(VDD),.Y(g11376),.A(I18332));
  NOT NOT1_3271(.VSS(VSS),.VDD(VDD),.Y(I18335),.A(g6783));
  NOT NOT1_3272(.VSS(VSS),.VDD(VDD),.Y(g11379),.A(I18335));
  NOT NOT1_3273(.VSS(VSS),.VDD(VDD),.Y(I18338),.A(g6574));
  NOT NOT1_3274(.VSS(VSS),.VDD(VDD),.Y(g11382),.A(I18338));
  NOT NOT1_3275(.VSS(VSS),.VDD(VDD),.Y(I18341),.A(g5610));
  NOT NOT1_3276(.VSS(VSS),.VDD(VDD),.Y(g11385),.A(I18341));
  NOT NOT1_3277(.VSS(VSS),.VDD(VDD),.Y(I18344),.A(g7015));
  NOT NOT1_3278(.VSS(VSS),.VDD(VDD),.Y(g11386),.A(I18344));
  NOT NOT1_3279(.VSS(VSS),.VDD(VDD),.Y(I18347),.A(g5778));
  NOT NOT1_3280(.VSS(VSS),.VDD(VDD),.Y(g11389),.A(I18347));
  NOT NOT1_3281(.VSS(VSS),.VDD(VDD),.Y(I18350),.A(g7195));
  NOT NOT1_3282(.VSS(VSS),.VDD(VDD),.Y(g11392),.A(I18350));
  NOT NOT1_3283(.VSS(VSS),.VDD(VDD),.Y(I18353),.A(g3722));
  NOT NOT1_3284(.VSS(VSS),.VDD(VDD),.Y(g11395),.A(I18353));
  NOT NOT1_3285(.VSS(VSS),.VDD(VDD),.Y(I18356),.A(g7085));
  NOT NOT1_3286(.VSS(VSS),.VDD(VDD),.Y(g11398),.A(I18356));
  NOT NOT1_3287(.VSS(VSS),.VDD(VDD),.Y(I18359),.A(g6838));
  NOT NOT1_3288(.VSS(VSS),.VDD(VDD),.Y(g11401),.A(I18359));
  NOT NOT1_3289(.VSS(VSS),.VDD(VDD),.Y(I18362),.A(g5837));
  NOT NOT1_3290(.VSS(VSS),.VDD(VDD),.Y(g11404),.A(I18362));
  NOT NOT1_3291(.VSS(VSS),.VDD(VDD),.Y(I18365),.A(g7391));
  NOT NOT1_3292(.VSS(VSS),.VDD(VDD),.Y(g11407),.A(I18365));
  NOT NOT1_3293(.VSS(VSS),.VDD(VDD),.Y(I18375),.A(g3254));
  NOT NOT1_3294(.VSS(VSS),.VDD(VDD),.Y(g11411),.A(I18375));
  NOT NOT1_3295(.VSS(VSS),.VDD(VDD),.Y(I18378),.A(g6314));
  NOT NOT1_3296(.VSS(VSS),.VDD(VDD),.Y(g11414),.A(I18378));
  NOT NOT1_3297(.VSS(VSS),.VDD(VDD),.Y(I18381),.A(g6232));
  NOT NOT1_3298(.VSS(VSS),.VDD(VDD),.Y(g11417),.A(I18381));
  NOT NOT1_3299(.VSS(VSS),.VDD(VDD),.Y(I18386),.A(g3254));
  NOT NOT1_3300(.VSS(VSS),.VDD(VDD),.Y(g11422),.A(I18386));
  NOT NOT1_3301(.VSS(VSS),.VDD(VDD),.Y(I18389),.A(g6519));
  NOT NOT1_3302(.VSS(VSS),.VDD(VDD),.Y(g11425),.A(I18389));
  NOT NOT1_3303(.VSS(VSS),.VDD(VDD),.Y(I18392),.A(g6369));
  NOT NOT1_3304(.VSS(VSS),.VDD(VDD),.Y(g11428),.A(I18392));
  NOT NOT1_3305(.VSS(VSS),.VDD(VDD),.Y(I18396),.A(g3410));
  NOT NOT1_3306(.VSS(VSS),.VDD(VDD),.Y(g11432),.A(I18396));
  NOT NOT1_3307(.VSS(VSS),.VDD(VDD),.Y(I18399),.A(g6519));
  NOT NOT1_3308(.VSS(VSS),.VDD(VDD),.Y(g11435),.A(I18399));
  NOT NOT1_3309(.VSS(VSS),.VDD(VDD),.Y(I18402),.A(g6713));
  NOT NOT1_3310(.VSS(VSS),.VDD(VDD),.Y(g11438),.A(I18402));
  NOT NOT1_3311(.VSS(VSS),.VDD(VDD),.Y(I18405),.A(g5720));
  NOT NOT1_3312(.VSS(VSS),.VDD(VDD),.Y(g11441),.A(I18405));
  NOT NOT1_3313(.VSS(VSS),.VDD(VDD),.Y(I18408),.A(g6574));
  NOT NOT1_3314(.VSS(VSS),.VDD(VDD),.Y(g11444),.A(I18408));
  NOT NOT1_3315(.VSS(VSS),.VDD(VDD),.Y(I18411),.A(g3566));
  NOT NOT1_3316(.VSS(VSS),.VDD(VDD),.Y(g11447),.A(I18411));
  NOT NOT1_3317(.VSS(VSS),.VDD(VDD),.Y(I18414),.A(g6783));
  NOT NOT1_3318(.VSS(VSS),.VDD(VDD),.Y(g11450),.A(I18414));
  NOT NOT1_3319(.VSS(VSS),.VDD(VDD),.Y(I18417),.A(g6574));
  NOT NOT1_3320(.VSS(VSS),.VDD(VDD),.Y(g11453),.A(I18417));
  NOT NOT1_3321(.VSS(VSS),.VDD(VDD),.Y(I18420),.A(g7015));
  NOT NOT1_3322(.VSS(VSS),.VDD(VDD),.Y(g11456),.A(I18420));
  NOT NOT1_3323(.VSS(VSS),.VDD(VDD),.Y(I18423),.A(g5778));
  NOT NOT1_3324(.VSS(VSS),.VDD(VDD),.Y(g11459),.A(I18423));
  NOT NOT1_3325(.VSS(VSS),.VDD(VDD),.Y(I18426),.A(g3722));
  NOT NOT1_3326(.VSS(VSS),.VDD(VDD),.Y(g11462),.A(I18426));
  NOT NOT1_3327(.VSS(VSS),.VDD(VDD),.Y(I18429),.A(g7085));
  NOT NOT1_3328(.VSS(VSS),.VDD(VDD),.Y(g11465),.A(I18429));
  NOT NOT1_3329(.VSS(VSS),.VDD(VDD),.Y(I18432),.A(g6838));
  NOT NOT1_3330(.VSS(VSS),.VDD(VDD),.Y(g11468),.A(I18432));
  NOT NOT1_3331(.VSS(VSS),.VDD(VDD),.Y(I18435),.A(g5635));
  NOT NOT1_3332(.VSS(VSS),.VDD(VDD),.Y(g11471),.A(I18435));
  NOT NOT1_3333(.VSS(VSS),.VDD(VDD),.Y(I18438),.A(g7265));
  NOT NOT1_3334(.VSS(VSS),.VDD(VDD),.Y(g11472),.A(I18438));
  NOT NOT1_3335(.VSS(VSS),.VDD(VDD),.Y(I18441),.A(g5837));
  NOT NOT1_3336(.VSS(VSS),.VDD(VDD),.Y(g11475),.A(I18441));
  NOT NOT1_3337(.VSS(VSS),.VDD(VDD),.Y(I18444),.A(g7391));
  NOT NOT1_3338(.VSS(VSS),.VDD(VDD),.Y(g11478),.A(I18444));
  NOT NOT1_3339(.VSS(VSS),.VDD(VDD),.Y(g11481),.A(g4204));
  NOT NOT1_3340(.VSS(VSS),.VDD(VDD),.Y(g11490),.A(g8276));
  NOT NOT1_3341(.VSS(VSS),.VDD(VDD),.Y(I18449),.A(g10868));
  NOT NOT1_3342(.VSS(VSS),.VDD(VDD),.Y(g11491),.A(I18449));
  NOT NOT1_3343(.VSS(VSS),.VDD(VDD),.Y(I18452),.A(g10930));
  NOT NOT1_3344(.VSS(VSS),.VDD(VDD),.Y(g11492),.A(I18452));
  NOT NOT1_3345(.VSS(VSS),.VDD(VDD),.Y(I18455),.A(g11031));
  NOT NOT1_3346(.VSS(VSS),.VDD(VDD),.Y(g11493),.A(I18455));
  NOT NOT1_3347(.VSS(VSS),.VDD(VDD),.Y(I18458),.A(g11208));
  NOT NOT1_3348(.VSS(VSS),.VDD(VDD),.Y(g11494),.A(I18458));
  NOT NOT1_3349(.VSS(VSS),.VDD(VDD),.Y(I18461),.A(g10931));
  NOT NOT1_3350(.VSS(VSS),.VDD(VDD),.Y(g11495),.A(I18461));
  NOT NOT1_3351(.VSS(VSS),.VDD(VDD),.Y(I18464),.A(g8620));
  NOT NOT1_3352(.VSS(VSS),.VDD(VDD),.Y(g11496),.A(I18464));
  NOT NOT1_3353(.VSS(VSS),.VDD(VDD),.Y(I18467),.A(g8769));
  NOT NOT1_3354(.VSS(VSS),.VDD(VDD),.Y(g11497),.A(I18467));
  NOT NOT1_3355(.VSS(VSS),.VDD(VDD),.Y(I18470),.A(g8808));
  NOT NOT1_3356(.VSS(VSS),.VDD(VDD),.Y(g11498),.A(I18470));
  NOT NOT1_3357(.VSS(VSS),.VDD(VDD),.Y(I18473),.A(g8839));
  NOT NOT1_3358(.VSS(VSS),.VDD(VDD),.Y(g11499),.A(I18473));
  NOT NOT1_3359(.VSS(VSS),.VDD(VDD),.Y(I18476),.A(g8791));
  NOT NOT1_3360(.VSS(VSS),.VDD(VDD),.Y(g11500),.A(I18476));
  NOT NOT1_3361(.VSS(VSS),.VDD(VDD),.Y(I18479),.A(g8820));
  NOT NOT1_3362(.VSS(VSS),.VDD(VDD),.Y(g11501),.A(I18479));
  NOT NOT1_3363(.VSS(VSS),.VDD(VDD),.Y(I18482),.A(g8859));
  NOT NOT1_3364(.VSS(VSS),.VDD(VDD),.Y(g11502),.A(I18482));
  NOT NOT1_3365(.VSS(VSS),.VDD(VDD),.Y(I18485),.A(g8809));
  NOT NOT1_3366(.VSS(VSS),.VDD(VDD),.Y(g11503),.A(I18485));
  NOT NOT1_3367(.VSS(VSS),.VDD(VDD),.Y(I18488),.A(g8840));
  NOT NOT1_3368(.VSS(VSS),.VDD(VDD),.Y(g11504),.A(I18488));
  NOT NOT1_3369(.VSS(VSS),.VDD(VDD),.Y(I18491),.A(g8891));
  NOT NOT1_3370(.VSS(VSS),.VDD(VDD),.Y(g11505),.A(I18491));
  NOT NOT1_3371(.VSS(VSS),.VDD(VDD),.Y(I18494),.A(g8821));
  NOT NOT1_3372(.VSS(VSS),.VDD(VDD),.Y(g11506),.A(I18494));
  NOT NOT1_3373(.VSS(VSS),.VDD(VDD),.Y(I18497),.A(g8860));
  NOT NOT1_3374(.VSS(VSS),.VDD(VDD),.Y(g11507),.A(I18497));
  NOT NOT1_3375(.VSS(VSS),.VDD(VDD),.Y(I18500),.A(g8924));
  NOT NOT1_3376(.VSS(VSS),.VDD(VDD),.Y(g11508),.A(I18500));
  NOT NOT1_3377(.VSS(VSS),.VDD(VDD),.Y(I18503),.A(g8658));
  NOT NOT1_3378(.VSS(VSS),.VDD(VDD),.Y(g11509),.A(I18503));
  NOT NOT1_3379(.VSS(VSS),.VDD(VDD),.Y(I18506),.A(g8699));
  NOT NOT1_3380(.VSS(VSS),.VDD(VDD),.Y(g11510),.A(I18506));
  NOT NOT1_3381(.VSS(VSS),.VDD(VDD),.Y(I18509),.A(g8770));
  NOT NOT1_3382(.VSS(VSS),.VDD(VDD),.Y(g11511),.A(I18509));
  NOT NOT1_3383(.VSS(VSS),.VDD(VDD),.Y(I18512),.A(g9309));
  NOT NOT1_3384(.VSS(VSS),.VDD(VDD),.Y(g11512),.A(I18512));
  NOT NOT1_3385(.VSS(VSS),.VDD(VDD),.Y(I18515),.A(g8843));
  NOT NOT1_3386(.VSS(VSS),.VDD(VDD),.Y(g11513),.A(I18515));
  NOT NOT1_3387(.VSS(VSS),.VDD(VDD),.Y(I18518),.A(g8893));
  NOT NOT1_3388(.VSS(VSS),.VDD(VDD),.Y(g11514),.A(I18518));
  NOT NOT1_3389(.VSS(VSS),.VDD(VDD),.Y(I18521),.A(g9449));
  NOT NOT1_3390(.VSS(VSS),.VDD(VDD),.Y(g11515),.A(I18521));
  NOT NOT1_3391(.VSS(VSS),.VDD(VDD),.Y(I18524),.A(g9640));
  NOT NOT1_3392(.VSS(VSS),.VDD(VDD),.Y(g11516),.A(I18524));
  NOT NOT1_3393(.VSS(VSS),.VDD(VDD),.Y(I18527),.A(g10017));
  NOT NOT1_3394(.VSS(VSS),.VDD(VDD),.Y(g11517),.A(I18527));
  NOT NOT1_3395(.VSS(VSS),.VDD(VDD),.Y(I18530),.A(g10888));
  NOT NOT1_3396(.VSS(VSS),.VDD(VDD),.Y(g11518),.A(I18530));
  NOT NOT1_3397(.VSS(VSS),.VDD(VDD),.Y(I18533),.A(g10967));
  NOT NOT1_3398(.VSS(VSS),.VDD(VDD),.Y(g11519),.A(I18533));
  NOT NOT1_3399(.VSS(VSS),.VDD(VDD),.Y(I18536),.A(g11101));
  NOT NOT1_3400(.VSS(VSS),.VDD(VDD),.Y(g11520),.A(I18536));
  NOT NOT1_3401(.VSS(VSS),.VDD(VDD),.Y(I18539),.A(g11290));
  NOT NOT1_3402(.VSS(VSS),.VDD(VDD),.Y(g11521),.A(I18539));
  NOT NOT1_3403(.VSS(VSS),.VDD(VDD),.Y(I18542),.A(g10968));
  NOT NOT1_3404(.VSS(VSS),.VDD(VDD),.Y(g11522),.A(I18542));
  NOT NOT1_3405(.VSS(VSS),.VDD(VDD),.Y(I18545),.A(g8630));
  NOT NOT1_3406(.VSS(VSS),.VDD(VDD),.Y(g11523),.A(I18545));
  NOT NOT1_3407(.VSS(VSS),.VDD(VDD),.Y(I18548),.A(g8792));
  NOT NOT1_3408(.VSS(VSS),.VDD(VDD),.Y(g11524),.A(I18548));
  NOT NOT1_3409(.VSS(VSS),.VDD(VDD),.Y(I18551),.A(g8824));
  NOT NOT1_3410(.VSS(VSS),.VDD(VDD),.Y(g11525),.A(I18551));
  NOT NOT1_3411(.VSS(VSS),.VDD(VDD),.Y(I18554),.A(g8866));
  NOT NOT1_3412(.VSS(VSS),.VDD(VDD),.Y(g11526),.A(I18554));
  NOT NOT1_3413(.VSS(VSS),.VDD(VDD),.Y(I18557),.A(g8810));
  NOT NOT1_3414(.VSS(VSS),.VDD(VDD),.Y(g11527),.A(I18557));
  NOT NOT1_3415(.VSS(VSS),.VDD(VDD),.Y(I18560),.A(g8844));
  NOT NOT1_3416(.VSS(VSS),.VDD(VDD),.Y(g11528),.A(I18560));
  NOT NOT1_3417(.VSS(VSS),.VDD(VDD),.Y(I18563),.A(g8897));
  NOT NOT1_3418(.VSS(VSS),.VDD(VDD),.Y(g11529),.A(I18563));
  NOT NOT1_3419(.VSS(VSS),.VDD(VDD),.Y(I18566),.A(g8825));
  NOT NOT1_3420(.VSS(VSS),.VDD(VDD),.Y(g11530),.A(I18566));
  NOT NOT1_3421(.VSS(VSS),.VDD(VDD),.Y(I18569),.A(g8867));
  NOT NOT1_3422(.VSS(VSS),.VDD(VDD),.Y(g11531),.A(I18569));
  NOT NOT1_3423(.VSS(VSS),.VDD(VDD),.Y(I18572),.A(g8931));
  NOT NOT1_3424(.VSS(VSS),.VDD(VDD),.Y(g11532),.A(I18572));
  NOT NOT1_3425(.VSS(VSS),.VDD(VDD),.Y(I18575),.A(g8845));
  NOT NOT1_3426(.VSS(VSS),.VDD(VDD),.Y(g11533),.A(I18575));
  NOT NOT1_3427(.VSS(VSS),.VDD(VDD),.Y(I18578),.A(g8898));
  NOT NOT1_3428(.VSS(VSS),.VDD(VDD),.Y(g11534),.A(I18578));
  NOT NOT1_3429(.VSS(VSS),.VDD(VDD),.Y(I18581),.A(g8964));
  NOT NOT1_3430(.VSS(VSS),.VDD(VDD),.Y(g11535),.A(I18581));
  NOT NOT1_3431(.VSS(VSS),.VDD(VDD),.Y(I18584),.A(g8677));
  NOT NOT1_3432(.VSS(VSS),.VDD(VDD),.Y(g11536),.A(I18584));
  NOT NOT1_3433(.VSS(VSS),.VDD(VDD),.Y(I18587),.A(g8718));
  NOT NOT1_3434(.VSS(VSS),.VDD(VDD),.Y(g11537),.A(I18587));
  NOT NOT1_3435(.VSS(VSS),.VDD(VDD),.Y(I18590),.A(g8793));
  NOT NOT1_3436(.VSS(VSS),.VDD(VDD),.Y(g11538),.A(I18590));
  NOT NOT1_3437(.VSS(VSS),.VDD(VDD),.Y(I18593),.A(g9390));
  NOT NOT1_3438(.VSS(VSS),.VDD(VDD),.Y(g11539),.A(I18593));
  NOT NOT1_3439(.VSS(VSS),.VDD(VDD),.Y(I18596),.A(g8870));
  NOT NOT1_3440(.VSS(VSS),.VDD(VDD),.Y(g11540),.A(I18596));
  NOT NOT1_3441(.VSS(VSS),.VDD(VDD),.Y(I18599),.A(g8933));
  NOT NOT1_3442(.VSS(VSS),.VDD(VDD),.Y(g11541),.A(I18599));
  NOT NOT1_3443(.VSS(VSS),.VDD(VDD),.Y(I18602),.A(g9591));
  NOT NOT1_3444(.VSS(VSS),.VDD(VDD),.Y(g11542),.A(I18602));
  NOT NOT1_3445(.VSS(VSS),.VDD(VDD),.Y(I18605),.A(g9786));
  NOT NOT1_3446(.VSS(VSS),.VDD(VDD),.Y(g11543),.A(I18605));
  NOT NOT1_3447(.VSS(VSS),.VDD(VDD),.Y(I18608),.A(g10126));
  NOT NOT1_3448(.VSS(VSS),.VDD(VDD),.Y(g11544),.A(I18608));
  NOT NOT1_3449(.VSS(VSS),.VDD(VDD),.Y(I18611),.A(g10909));
  NOT NOT1_3450(.VSS(VSS),.VDD(VDD),.Y(g11545),.A(I18611));
  NOT NOT1_3451(.VSS(VSS),.VDD(VDD),.Y(I18614),.A(g11002));
  NOT NOT1_3452(.VSS(VSS),.VDD(VDD),.Y(g11546),.A(I18614));
  NOT NOT1_3453(.VSS(VSS),.VDD(VDD),.Y(I18617),.A(g11169));
  NOT NOT1_3454(.VSS(VSS),.VDD(VDD),.Y(g11547),.A(I18617));
  NOT NOT1_3455(.VSS(VSS),.VDD(VDD),.Y(I18620),.A(g11385));
  NOT NOT1_3456(.VSS(VSS),.VDD(VDD),.Y(g11548),.A(I18620));
  NOT NOT1_3457(.VSS(VSS),.VDD(VDD),.Y(I18623),.A(g11003));
  NOT NOT1_3458(.VSS(VSS),.VDD(VDD),.Y(g11549),.A(I18623));
  NOT NOT1_3459(.VSS(VSS),.VDD(VDD),.Y(I18626),.A(g8649));
  NOT NOT1_3460(.VSS(VSS),.VDD(VDD),.Y(g11550),.A(I18626));
  NOT NOT1_3461(.VSS(VSS),.VDD(VDD),.Y(I18629),.A(g8811));
  NOT NOT1_3462(.VSS(VSS),.VDD(VDD),.Y(g11551),.A(I18629));
  NOT NOT1_3463(.VSS(VSS),.VDD(VDD),.Y(I18632),.A(g8850));
  NOT NOT1_3464(.VSS(VSS),.VDD(VDD),.Y(g11552),.A(I18632));
  NOT NOT1_3465(.VSS(VSS),.VDD(VDD),.Y(I18635),.A(g8904));
  NOT NOT1_3466(.VSS(VSS),.VDD(VDD),.Y(g11553),.A(I18635));
  NOT NOT1_3467(.VSS(VSS),.VDD(VDD),.Y(I18638),.A(g8826));
  NOT NOT1_3468(.VSS(VSS),.VDD(VDD),.Y(g11554),.A(I18638));
  NOT NOT1_3469(.VSS(VSS),.VDD(VDD),.Y(I18641),.A(g8871));
  NOT NOT1_3470(.VSS(VSS),.VDD(VDD),.Y(g11555),.A(I18641));
  NOT NOT1_3471(.VSS(VSS),.VDD(VDD),.Y(I18644),.A(g8937));
  NOT NOT1_3472(.VSS(VSS),.VDD(VDD),.Y(g11556),.A(I18644));
  NOT NOT1_3473(.VSS(VSS),.VDD(VDD),.Y(I18647),.A(g8851));
  NOT NOT1_3474(.VSS(VSS),.VDD(VDD),.Y(g11557),.A(I18647));
  NOT NOT1_3475(.VSS(VSS),.VDD(VDD),.Y(I18650),.A(g8905));
  NOT NOT1_3476(.VSS(VSS),.VDD(VDD),.Y(g11558),.A(I18650));
  NOT NOT1_3477(.VSS(VSS),.VDD(VDD),.Y(I18653),.A(g8971));
  NOT NOT1_3478(.VSS(VSS),.VDD(VDD),.Y(g11559),.A(I18653));
  NOT NOT1_3479(.VSS(VSS),.VDD(VDD),.Y(I18656),.A(g8872));
  NOT NOT1_3480(.VSS(VSS),.VDD(VDD),.Y(g11560),.A(I18656));
  NOT NOT1_3481(.VSS(VSS),.VDD(VDD),.Y(I18659),.A(g8938));
  NOT NOT1_3482(.VSS(VSS),.VDD(VDD),.Y(g11561),.A(I18659));
  NOT NOT1_3483(.VSS(VSS),.VDD(VDD),.Y(I18662),.A(g8996));
  NOT NOT1_3484(.VSS(VSS),.VDD(VDD),.Y(g11562),.A(I18662));
  NOT NOT1_3485(.VSS(VSS),.VDD(VDD),.Y(I18665),.A(g8689));
  NOT NOT1_3486(.VSS(VSS),.VDD(VDD),.Y(g11563),.A(I18665));
  NOT NOT1_3487(.VSS(VSS),.VDD(VDD),.Y(I18668),.A(g8756));
  NOT NOT1_3488(.VSS(VSS),.VDD(VDD),.Y(g11564),.A(I18668));
  NOT NOT1_3489(.VSS(VSS),.VDD(VDD),.Y(I18671),.A(g8812));
  NOT NOT1_3490(.VSS(VSS),.VDD(VDD),.Y(g11565),.A(I18671));
  NOT NOT1_3491(.VSS(VSS),.VDD(VDD),.Y(I18674),.A(g9487));
  NOT NOT1_3492(.VSS(VSS),.VDD(VDD),.Y(g11566),.A(I18674));
  NOT NOT1_3493(.VSS(VSS),.VDD(VDD),.Y(I18677),.A(g8908));
  NOT NOT1_3494(.VSS(VSS),.VDD(VDD),.Y(g11567),.A(I18677));
  NOT NOT1_3495(.VSS(VSS),.VDD(VDD),.Y(I18680),.A(g8973));
  NOT NOT1_3496(.VSS(VSS),.VDD(VDD),.Y(g11568),.A(I18680));
  NOT NOT1_3497(.VSS(VSS),.VDD(VDD),.Y(I18683),.A(g9733));
  NOT NOT1_3498(.VSS(VSS),.VDD(VDD),.Y(g11569),.A(I18683));
  NOT NOT1_3499(.VSS(VSS),.VDD(VDD),.Y(I18686),.A(g9932));
  NOT NOT1_3500(.VSS(VSS),.VDD(VDD),.Y(g11570),.A(I18686));
  NOT NOT1_3501(.VSS(VSS),.VDD(VDD),.Y(I18689),.A(g10231));
  NOT NOT1_3502(.VSS(VSS),.VDD(VDD),.Y(g11571),.A(I18689));
  NOT NOT1_3503(.VSS(VSS),.VDD(VDD),.Y(I18692),.A(g10935));
  NOT NOT1_3504(.VSS(VSS),.VDD(VDD),.Y(g11572),.A(I18692));
  NOT NOT1_3505(.VSS(VSS),.VDD(VDD),.Y(I18695),.A(g11054));
  NOT NOT1_3506(.VSS(VSS),.VDD(VDD),.Y(g11573),.A(I18695));
  NOT NOT1_3507(.VSS(VSS),.VDD(VDD),.Y(I18698),.A(g11255));
  NOT NOT1_3508(.VSS(VSS),.VDD(VDD),.Y(g11574),.A(I18698));
  NOT NOT1_3509(.VSS(VSS),.VDD(VDD),.Y(I18701),.A(g11471));
  NOT NOT1_3510(.VSS(VSS),.VDD(VDD),.Y(g11575),.A(I18701));
  NOT NOT1_3511(.VSS(VSS),.VDD(VDD),.Y(I18704),.A(g11055));
  NOT NOT1_3512(.VSS(VSS),.VDD(VDD),.Y(g11576),.A(I18704));
  NOT NOT1_3513(.VSS(VSS),.VDD(VDD),.Y(I18707),.A(g8665));
  NOT NOT1_3514(.VSS(VSS),.VDD(VDD),.Y(g11577),.A(I18707));
  NOT NOT1_3515(.VSS(VSS),.VDD(VDD),.Y(I18710),.A(g8827));
  NOT NOT1_3516(.VSS(VSS),.VDD(VDD),.Y(g11578),.A(I18710));
  NOT NOT1_3517(.VSS(VSS),.VDD(VDD),.Y(I18713),.A(g8877));
  NOT NOT1_3518(.VSS(VSS),.VDD(VDD),.Y(g11579),.A(I18713));
  NOT NOT1_3519(.VSS(VSS),.VDD(VDD),.Y(I18716),.A(g8944));
  NOT NOT1_3520(.VSS(VSS),.VDD(VDD),.Y(g11580),.A(I18716));
  NOT NOT1_3521(.VSS(VSS),.VDD(VDD),.Y(I18719),.A(g8852));
  NOT NOT1_3522(.VSS(VSS),.VDD(VDD),.Y(g11581),.A(I18719));
  NOT NOT1_3523(.VSS(VSS),.VDD(VDD),.Y(I18722),.A(g8909));
  NOT NOT1_3524(.VSS(VSS),.VDD(VDD),.Y(g11582),.A(I18722));
  NOT NOT1_3525(.VSS(VSS),.VDD(VDD),.Y(I18725),.A(g8977));
  NOT NOT1_3526(.VSS(VSS),.VDD(VDD),.Y(g11583),.A(I18725));
  NOT NOT1_3527(.VSS(VSS),.VDD(VDD),.Y(I18728),.A(g8878));
  NOT NOT1_3528(.VSS(VSS),.VDD(VDD),.Y(g11584),.A(I18728));
  NOT NOT1_3529(.VSS(VSS),.VDD(VDD),.Y(I18731),.A(g8945));
  NOT NOT1_3530(.VSS(VSS),.VDD(VDD),.Y(g11585),.A(I18731));
  NOT NOT1_3531(.VSS(VSS),.VDD(VDD),.Y(I18734),.A(g9003));
  NOT NOT1_3532(.VSS(VSS),.VDD(VDD),.Y(g11586),.A(I18734));
  NOT NOT1_3533(.VSS(VSS),.VDD(VDD),.Y(I18737),.A(g8910));
  NOT NOT1_3534(.VSS(VSS),.VDD(VDD),.Y(g11587),.A(I18737));
  NOT NOT1_3535(.VSS(VSS),.VDD(VDD),.Y(I18740),.A(g8978));
  NOT NOT1_3536(.VSS(VSS),.VDD(VDD),.Y(g11588),.A(I18740));
  NOT NOT1_3537(.VSS(VSS),.VDD(VDD),.Y(I18743),.A(g9025));
  NOT NOT1_3538(.VSS(VSS),.VDD(VDD),.Y(g11589),.A(I18743));
  NOT NOT1_3539(.VSS(VSS),.VDD(VDD),.Y(I18746),.A(g8707));
  NOT NOT1_3540(.VSS(VSS),.VDD(VDD),.Y(g11590),.A(I18746));
  NOT NOT1_3541(.VSS(VSS),.VDD(VDD),.Y(I18749),.A(g8779));
  NOT NOT1_3542(.VSS(VSS),.VDD(VDD),.Y(g11591),.A(I18749));
  NOT NOT1_3543(.VSS(VSS),.VDD(VDD),.Y(I18752),.A(g8828));
  NOT NOT1_3544(.VSS(VSS),.VDD(VDD),.Y(g11592),.A(I18752));
  NOT NOT1_3545(.VSS(VSS),.VDD(VDD),.Y(I18755),.A(g9629));
  NOT NOT1_3546(.VSS(VSS),.VDD(VDD),.Y(g11593),.A(I18755));
  NOT NOT1_3547(.VSS(VSS),.VDD(VDD),.Y(I18758),.A(g8948));
  NOT NOT1_3548(.VSS(VSS),.VDD(VDD),.Y(g11594),.A(I18758));
  NOT NOT1_3549(.VSS(VSS),.VDD(VDD),.Y(I18761),.A(g9005));
  NOT NOT1_3550(.VSS(VSS),.VDD(VDD),.Y(g11595),.A(I18761));
  NOT NOT1_3551(.VSS(VSS),.VDD(VDD),.Y(I18764),.A(g9879));
  NOT NOT1_3552(.VSS(VSS),.VDD(VDD),.Y(g11596),.A(I18764));
  NOT NOT1_3553(.VSS(VSS),.VDD(VDD),.Y(I18767),.A(g10086));
  NOT NOT1_3554(.VSS(VSS),.VDD(VDD),.Y(g11597),.A(I18767));
  NOT NOT1_3555(.VSS(VSS),.VDD(VDD),.Y(I18770),.A(g10333));
  NOT NOT1_3556(.VSS(VSS),.VDD(VDD),.Y(g11598),.A(I18770));
  NOT NOT1_3557(.VSS(VSS),.VDD(VDD),.Y(I18773),.A(g10830));
  NOT NOT1_3558(.VSS(VSS),.VDD(VDD),.Y(g11599),.A(I18773));
  NOT NOT1_3559(.VSS(VSS),.VDD(VDD),.Y(I18777),.A(g9050));
  NOT NOT1_3560(.VSS(VSS),.VDD(VDD),.Y(g11603),.A(I18777));
  NOT NOT1_3561(.VSS(VSS),.VDD(VDD),.Y(I18780),.A(g10870));
  NOT NOT1_3562(.VSS(VSS),.VDD(VDD),.Y(g11606),.A(I18780));
  NOT NOT1_3563(.VSS(VSS),.VDD(VDD),.Y(I18784),.A(g9067));
  NOT NOT1_3564(.VSS(VSS),.VDD(VDD),.Y(g11608),.A(I18784));
  NOT NOT1_3565(.VSS(VSS),.VDD(VDD),.Y(I18787),.A(g10910));
  NOT NOT1_3566(.VSS(VSS),.VDD(VDD),.Y(g11611),.A(I18787));
  NOT NOT1_3567(.VSS(VSS),.VDD(VDD),.Y(I18791),.A(g9084));
  NOT NOT1_3568(.VSS(VSS),.VDD(VDD),.Y(g11613),.A(I18791));
  NOT NOT1_3569(.VSS(VSS),.VDD(VDD),.Y(I18794),.A(g10973));
  NOT NOT1_3570(.VSS(VSS),.VDD(VDD),.Y(g11616),.A(I18794));
  NOT NOT1_3571(.VSS(VSS),.VDD(VDD),.Y(g11620),.A(g10601));
  NOT NOT1_3572(.VSS(VSS),.VDD(VDD),.Y(g11623),.A(g10961));
  NOT NOT1_3573(.VSS(VSS),.VDD(VDD),.Y(I18810),.A(g10813));
  NOT NOT1_3574(.VSS(VSS),.VDD(VDD),.Y(g11628),.A(I18810));
  NOT NOT1_3575(.VSS(VSS),.VDD(VDD),.Y(I18813),.A(g10850));
  NOT NOT1_3576(.VSS(VSS),.VDD(VDD),.Y(g11629),.A(I18813));
  NOT NOT1_3577(.VSS(VSS),.VDD(VDD),.Y(I18817),.A(g9067));
  NOT NOT1_3578(.VSS(VSS),.VDD(VDD),.Y(g11633),.A(I18817));
  NOT NOT1_3579(.VSS(VSS),.VDD(VDD),.Y(I18820),.A(g10890));
  NOT NOT1_3580(.VSS(VSS),.VDD(VDD),.Y(g11636),.A(I18820));
  NOT NOT1_3581(.VSS(VSS),.VDD(VDD),.Y(I18824),.A(g9084));
  NOT NOT1_3582(.VSS(VSS),.VDD(VDD),.Y(g11638),.A(I18824));
  NOT NOT1_3583(.VSS(VSS),.VDD(VDD),.Y(I18827),.A(g10936));
  NOT NOT1_3584(.VSS(VSS),.VDD(VDD),.Y(g11641),.A(I18827));
  NOT NOT1_3585(.VSS(VSS),.VDD(VDD),.Y(g11642),.A(g10646));
  NOT NOT1_3586(.VSS(VSS),.VDD(VDD),.Y(I18835),.A(g10834));
  NOT NOT1_3587(.VSS(VSS),.VDD(VDD),.Y(g11651),.A(I18835));
  NOT NOT1_3588(.VSS(VSS),.VDD(VDD),.Y(I18838),.A(g10871));
  NOT NOT1_3589(.VSS(VSS),.VDD(VDD),.Y(g11652),.A(I18838));
  NOT NOT1_3590(.VSS(VSS),.VDD(VDD),.Y(I18842),.A(g9084));
  NOT NOT1_3591(.VSS(VSS),.VDD(VDD),.Y(g11656),.A(I18842));
  NOT NOT1_3592(.VSS(VSS),.VDD(VDD),.Y(I18845),.A(g10911));
  NOT NOT1_3593(.VSS(VSS),.VDD(VDD),.Y(g11659),.A(I18845));
  NOT NOT1_3594(.VSS(VSS),.VDD(VDD),.Y(I18854),.A(g10854));
  NOT NOT1_3595(.VSS(VSS),.VDD(VDD),.Y(g11670),.A(I18854));
  NOT NOT1_3596(.VSS(VSS),.VDD(VDD),.Y(I18857),.A(g10891));
  NOT NOT1_3597(.VSS(VSS),.VDD(VDD),.Y(g11671),.A(I18857));
  NOT NOT1_3598(.VSS(VSS),.VDD(VDD),.Y(I18866),.A(g10875));
  NOT NOT1_3599(.VSS(VSS),.VDD(VDD),.Y(g11682),.A(I18866));
  NOT NOT1_3600(.VSS(VSS),.VDD(VDD),.Y(g11706),.A(g10928));
  NOT NOT1_3601(.VSS(VSS),.VDD(VDD),.Y(g11732),.A(g10826));
  NOT NOT1_3602(.VSS(VSS),.VDD(VDD),.Y(g11734),.A(g10843));
  NOT NOT1_3603(.VSS(VSS),.VDD(VDD),.Y(g11735),.A(g10859));
  NOT NOT1_3604(.VSS(VSS),.VDD(VDD),.Y(g11736),.A(g10862));
  NOT NOT1_3605(.VSS(VSS),.VDD(VDD),.Y(g11737),.A(g10809));
  NOT NOT1_3606(.VSS(VSS),.VDD(VDD),.Y(g11740),.A(g10877));
  NOT NOT1_3607(.VSS(VSS),.VDD(VDD),.Y(g11741),.A(g10880));
  NOT NOT1_3608(.VSS(VSS),.VDD(VDD),.Y(g11742),.A(g10883));
  NOT NOT1_3609(.VSS(VSS),.VDD(VDD),.Y(g11743),.A(g8530));
  NOT NOT1_3610(.VSS(VSS),.VDD(VDD),.Y(g11745),.A(g10892));
  NOT NOT1_3611(.VSS(VSS),.VDD(VDD),.Y(g11746),.A(g10895));
  NOT NOT1_3612(.VSS(VSS),.VDD(VDD),.Y(g11747),.A(g10898));
  NOT NOT1_3613(.VSS(VSS),.VDD(VDD),.Y(g11748),.A(g10901));
  NOT NOT1_3614(.VSS(VSS),.VDD(VDD),.Y(I18929),.A(g10711));
  NOT NOT1_3615(.VSS(VSS),.VDD(VDD),.Y(g11749),.A(I18929));
  NOT NOT1_3616(.VSS(VSS),.VDD(VDD),.Y(g11758),.A(g8514));
  NOT NOT1_3617(.VSS(VSS),.VDD(VDD),.Y(g11761),.A(g10912));
  NOT NOT1_3618(.VSS(VSS),.VDD(VDD),.Y(g11762),.A(g10915));
  NOT NOT1_3619(.VSS(VSS),.VDD(VDD),.Y(g11763),.A(g10918));
  NOT NOT1_3620(.VSS(VSS),.VDD(VDD),.Y(g11764),.A(g10921));
  NOT NOT1_3621(.VSS(VSS),.VDD(VDD),.Y(g11765),.A(g10924));
  NOT NOT1_3622(.VSS(VSS),.VDD(VDD),.Y(g11766),.A(g10886));
  NOT NOT1_3623(.VSS(VSS),.VDD(VDD),.Y(I18943),.A(g9149));
  NOT NOT1_3624(.VSS(VSS),.VDD(VDD),.Y(g11769),.A(I18943));
  NOT NOT1_3625(.VSS(VSS),.VDD(VDD),.Y(g11770),.A(g10932));
  NOT NOT1_3626(.VSS(VSS),.VDD(VDD),.Y(g11774),.A(g10937));
  NOT NOT1_3627(.VSS(VSS),.VDD(VDD),.Y(g11775),.A(g10940));
  NOT NOT1_3628(.VSS(VSS),.VDD(VDD),.Y(g11776),.A(g10943));
  NOT NOT1_3629(.VSS(VSS),.VDD(VDD),.Y(g11777),.A(g10946));
  NOT NOT1_3630(.VSS(VSS),.VDD(VDD),.Y(g11778),.A(g10949));
  NOT NOT1_3631(.VSS(VSS),.VDD(VDD),.Y(g11779),.A(g10906));
  NOT NOT1_3632(.VSS(VSS),.VDD(VDD),.Y(g11782),.A(g10963));
  NOT NOT1_3633(.VSS(VSS),.VDD(VDD),.Y(g11783),.A(g10966));
  NOT NOT1_3634(.VSS(VSS),.VDD(VDD),.Y(I18962),.A(g9159));
  NOT NOT1_3635(.VSS(VSS),.VDD(VDD),.Y(g11786),.A(I18962));
  NOT NOT1_3636(.VSS(VSS),.VDD(VDD),.Y(g11787),.A(g10969));
  NOT NOT1_3637(.VSS(VSS),.VDD(VDD),.Y(I18969),.A(g8726));
  NOT NOT1_3638(.VSS(VSS),.VDD(VDD),.Y(g11791),.A(I18969));
  NOT NOT1_3639(.VSS(VSS),.VDD(VDD),.Y(g11794),.A(g10974));
  NOT NOT1_3640(.VSS(VSS),.VDD(VDD),.Y(g11795),.A(g10977));
  NOT NOT1_3641(.VSS(VSS),.VDD(VDD),.Y(g11796),.A(g10980));
  NOT NOT1_3642(.VSS(VSS),.VDD(VDD),.Y(g11797),.A(g10983));
  NOT NOT1_3643(.VSS(VSS),.VDD(VDD),.Y(g11798),.A(g10867));
  NOT NOT1_3644(.VSS(VSS),.VDD(VDD),.Y(g11801),.A(g10988));
  NOT NOT1_3645(.VSS(VSS),.VDD(VDD),.Y(g11802),.A(g10991));
  NOT NOT1_3646(.VSS(VSS),.VDD(VDD),.Y(g11803),.A(g10994));
  NOT NOT1_3647(.VSS(VSS),.VDD(VDD),.Y(g11804),.A(g10995));
  NOT NOT1_3648(.VSS(VSS),.VDD(VDD),.Y(g11808),.A(g10996));
  NOT NOT1_3649(.VSS(VSS),.VDD(VDD),.Y(g11809),.A(g10999));
  NOT NOT1_3650(.VSS(VSS),.VDD(VDD),.Y(I18990),.A(g9183));
  NOT NOT1_3651(.VSS(VSS),.VDD(VDD),.Y(g11812),.A(I18990));
  NOT NOT1_3652(.VSS(VSS),.VDD(VDD),.Y(g11813),.A(g11004));
  NOT NOT1_3653(.VSS(VSS),.VDD(VDD),.Y(g11817),.A(g11008));
  NOT NOT1_3654(.VSS(VSS),.VDD(VDD),.Y(g11818),.A(g11011));
  NOT NOT1_3655(.VSS(VSS),.VDD(VDD),.Y(g11819),.A(g11014));
  NOT NOT1_3656(.VSS(VSS),.VDD(VDD),.Y(g11820),.A(g11017));
  NOT NOT1_3657(.VSS(VSS),.VDD(VDD),.Y(g11821),.A(g10848));
  NOT NOT1_3658(.VSS(VSS),.VDD(VDD),.Y(g11824),.A(g11022));
  NOT NOT1_3659(.VSS(VSS),.VDD(VDD),.Y(g11825),.A(g11025));
  NOT NOT1_3660(.VSS(VSS),.VDD(VDD),.Y(g11826),.A(g11028));
  NOT NOT1_3661(.VSS(VSS),.VDD(VDD),.Y(g11827),.A(g11032));
  NOT NOT1_3662(.VSS(VSS),.VDD(VDD),.Y(g11829),.A(g11035));
  NOT NOT1_3663(.VSS(VSS),.VDD(VDD),.Y(g11834),.A(g11036));
  NOT NOT1_3664(.VSS(VSS),.VDD(VDD),.Y(g11835),.A(g11039));
  NOT NOT1_3665(.VSS(VSS),.VDD(VDD),.Y(g11836),.A(g11042));
  NOT NOT1_3666(.VSS(VSS),.VDD(VDD),.Y(g11837),.A(g11045));
  NOT NOT1_3667(.VSS(VSS),.VDD(VDD),.Y(g11841),.A(g11048));
  NOT NOT1_3668(.VSS(VSS),.VDD(VDD),.Y(g11842),.A(g11051));
  NOT NOT1_3669(.VSS(VSS),.VDD(VDD),.Y(I19025),.A(g9225));
  NOT NOT1_3670(.VSS(VSS),.VDD(VDD),.Y(g11845),.A(I19025));
  NOT NOT1_3671(.VSS(VSS),.VDD(VDD),.Y(g11846),.A(g11056));
  NOT NOT1_3672(.VSS(VSS),.VDD(VDD),.Y(I19030),.A(g8726));
  NOT NOT1_3673(.VSS(VSS),.VDD(VDD),.Y(g11848),.A(I19030));
  NOT NOT1_3674(.VSS(VSS),.VDD(VDD),.Y(g11852),.A(g11063));
  NOT NOT1_3675(.VSS(VSS),.VDD(VDD),.Y(g11853),.A(g11066));
  NOT NOT1_3676(.VSS(VSS),.VDD(VDD),.Y(g11854),.A(g11078));
  NOT NOT1_3677(.VSS(VSS),.VDD(VDD),.Y(g11856),.A(g11079));
  NOT NOT1_3678(.VSS(VSS),.VDD(VDD),.Y(g11857),.A(g11082));
  NOT NOT1_3679(.VSS(VSS),.VDD(VDD),.Y(g11858),.A(g11085));
  NOT NOT1_3680(.VSS(VSS),.VDD(VDD),.Y(g11859),.A(g11088));
  NOT NOT1_3681(.VSS(VSS),.VDD(VDD),.Y(g11862),.A(g11091));
  NOT NOT1_3682(.VSS(VSS),.VDD(VDD),.Y(g11866),.A(g11092));
  NOT NOT1_3683(.VSS(VSS),.VDD(VDD),.Y(g11867),.A(g11095));
  NOT NOT1_3684(.VSS(VSS),.VDD(VDD),.Y(g11868),.A(g11098));
  NOT NOT1_3685(.VSS(VSS),.VDD(VDD),.Y(g11869),.A(g11102));
  NOT NOT1_3686(.VSS(VSS),.VDD(VDD),.Y(g11871),.A(g11105));
  NOT NOT1_3687(.VSS(VSS),.VDD(VDD),.Y(g11876),.A(g11108));
  NOT NOT1_3688(.VSS(VSS),.VDD(VDD),.Y(g11877),.A(g11111));
  NOT NOT1_3689(.VSS(VSS),.VDD(VDD),.Y(g11878),.A(g11114));
  NOT NOT1_3690(.VSS(VSS),.VDD(VDD),.Y(g11879),.A(g11117));
  NOT NOT1_3691(.VSS(VSS),.VDD(VDD),.Y(g11883),.A(g11120));
  NOT NOT1_3692(.VSS(VSS),.VDD(VDD),.Y(g11884),.A(g11123));
  NOT NOT1_3693(.VSS(VSS),.VDD(VDD),.Y(g11886),.A(g11126));
  NOT NOT1_3694(.VSS(VSS),.VDD(VDD),.Y(g11887),.A(g11129));
  NOT NOT1_3695(.VSS(VSS),.VDD(VDD),.Y(g11888),.A(g11021));
  NOT NOT1_3696(.VSS(VSS),.VDD(VDD),.Y(g11891),.A(g11132));
  NOT NOT1_3697(.VSS(VSS),.VDD(VDD),.Y(g11892),.A(g11135));
  NOT NOT1_3698(.VSS(VSS),.VDD(VDD),.Y(g11893),.A(g11138));
  NOT NOT1_3699(.VSS(VSS),.VDD(VDD),.Y(g11894),.A(g11141));
  NOT NOT1_3700(.VSS(VSS),.VDD(VDD),.Y(g11895),.A(g11144));
  NOT NOT1_3701(.VSS(VSS),.VDD(VDD),.Y(g11898),.A(g11145));
  NOT NOT1_3702(.VSS(VSS),.VDD(VDD),.Y(g11899),.A(g11148));
  NOT NOT1_3703(.VSS(VSS),.VDD(VDD),.Y(g11900),.A(g11151));
  NOT NOT1_3704(.VSS(VSS),.VDD(VDD),.Y(g11901),.A(g11154));
  NOT NOT1_3705(.VSS(VSS),.VDD(VDD),.Y(g11904),.A(g11157));
  NOT NOT1_3706(.VSS(VSS),.VDD(VDD),.Y(g11908),.A(g11160));
  NOT NOT1_3707(.VSS(VSS),.VDD(VDD),.Y(g11909),.A(g11163));
  NOT NOT1_3708(.VSS(VSS),.VDD(VDD),.Y(g11910),.A(g11166));
  NOT NOT1_3709(.VSS(VSS),.VDD(VDD),.Y(g11911),.A(g11170));
  NOT NOT1_3710(.VSS(VSS),.VDD(VDD),.Y(g11913),.A(g11173));
  NOT NOT1_3711(.VSS(VSS),.VDD(VDD),.Y(g11918),.A(g11176));
  NOT NOT1_3712(.VSS(VSS),.VDD(VDD),.Y(g11919),.A(g11179));
  NOT NOT1_3713(.VSS(VSS),.VDD(VDD),.Y(g11920),.A(g11182));
  NOT NOT1_3714(.VSS(VSS),.VDD(VDD),.Y(g11921),.A(g11185));
  NOT NOT1_3715(.VSS(VSS),.VDD(VDD),.Y(I19105),.A(g8726));
  NOT NOT1_3716(.VSS(VSS),.VDD(VDD),.Y(g11923),.A(I19105));
  NOT NOT1_3717(.VSS(VSS),.VDD(VDD),.Y(g11927),.A(g10987));
  NOT NOT1_3718(.VSS(VSS),.VDD(VDD),.Y(g11929),.A(g11199));
  NOT NOT1_3719(.VSS(VSS),.VDD(VDD),.Y(g11930),.A(g11202));
  NOT NOT1_3720(.VSS(VSS),.VDD(VDD),.Y(g11931),.A(g11205));
  NOT NOT1_3721(.VSS(VSS),.VDD(VDD),.Y(g11932),.A(g11209));
  NOT NOT1_3722(.VSS(VSS),.VDD(VDD),.Y(g11933),.A(g11210));
  NOT NOT1_3723(.VSS(VSS),.VDD(VDD),.Y(g11936),.A(g11213));
  NOT NOT1_3724(.VSS(VSS),.VDD(VDD),.Y(I19119),.A(g9202));
  NOT NOT1_3725(.VSS(VSS),.VDD(VDD),.Y(g11937),.A(I19119));
  NOT NOT1_3726(.VSS(VSS),.VDD(VDD),.Y(g11941),.A(g11216));
  NOT NOT1_3727(.VSS(VSS),.VDD(VDD),.Y(g11942),.A(g11219));
  NOT NOT1_3728(.VSS(VSS),.VDD(VDD),.Y(g11943),.A(g11222));
  NOT NOT1_3729(.VSS(VSS),.VDD(VDD),.Y(g11944),.A(g11225));
  NOT NOT1_3730(.VSS(VSS),.VDD(VDD),.Y(g11945),.A(g11228));
  NOT NOT1_3731(.VSS(VSS),.VDD(VDD),.Y(g11948),.A(g11231));
  NOT NOT1_3732(.VSS(VSS),.VDD(VDD),.Y(g11949),.A(g11234));
  NOT NOT1_3733(.VSS(VSS),.VDD(VDD),.Y(g11950),.A(g11237));
  NOT NOT1_3734(.VSS(VSS),.VDD(VDD),.Y(g11951),.A(g11240));
  NOT NOT1_3735(.VSS(VSS),.VDD(VDD),.Y(g11954),.A(g11243));
  NOT NOT1_3736(.VSS(VSS),.VDD(VDD),.Y(g11958),.A(g11246));
  NOT NOT1_3737(.VSS(VSS),.VDD(VDD),.Y(g11959),.A(g11249));
  NOT NOT1_3738(.VSS(VSS),.VDD(VDD),.Y(g11960),.A(g11252));
  NOT NOT1_3739(.VSS(VSS),.VDD(VDD),.Y(g11961),.A(g11256));
  NOT NOT1_3740(.VSS(VSS),.VDD(VDD),.Y(g11963),.A(g11259));
  NOT NOT1_3741(.VSS(VSS),.VDD(VDD),.Y(g11968),.A(g11265));
  NOT NOT1_3742(.VSS(VSS),.VDD(VDD),.Y(g11969),.A(g11268));
  NOT NOT1_3743(.VSS(VSS),.VDD(VDD),.Y(g11970),.A(g11271));
  NOT NOT1_3744(.VSS(VSS),.VDD(VDD),.Y(g11971),.A(g11274));
  NOT NOT1_3745(.VSS(VSS),.VDD(VDD),.Y(g11972),.A(g11277));
  NOT NOT1_3746(.VSS(VSS),.VDD(VDD),.Y(g11973),.A(g11278));
  NOT NOT1_3747(.VSS(VSS),.VDD(VDD),.Y(I19160),.A(g10549));
  NOT NOT1_3748(.VSS(VSS),.VDD(VDD),.Y(g11976),.A(I19160));
  NOT NOT1_3749(.VSS(VSS),.VDD(VDD),.Y(g11982),.A(g11281));
  NOT NOT1_3750(.VSS(VSS),.VDD(VDD),.Y(g11983),.A(g11284));
  NOT NOT1_3751(.VSS(VSS),.VDD(VDD),.Y(g11984),.A(g11287));
  NOT NOT1_3752(.VSS(VSS),.VDD(VDD),.Y(g11985),.A(g11291));
  NOT NOT1_3753(.VSS(VSS),.VDD(VDD),.Y(g11986),.A(g11294));
  NOT NOT1_3754(.VSS(VSS),.VDD(VDD),.Y(g11989),.A(g11297));
  NOT NOT1_3755(.VSS(VSS),.VDD(VDD),.Y(I19174),.A(g9263));
  NOT NOT1_3756(.VSS(VSS),.VDD(VDD),.Y(g11990),.A(I19174));
  NOT NOT1_3757(.VSS(VSS),.VDD(VDD),.Y(g11994),.A(g11300));
  NOT NOT1_3758(.VSS(VSS),.VDD(VDD),.Y(g11995),.A(g11303));
  NOT NOT1_3759(.VSS(VSS),.VDD(VDD),.Y(g11996),.A(g11306));
  NOT NOT1_3760(.VSS(VSS),.VDD(VDD),.Y(g11997),.A(g11309));
  NOT NOT1_3761(.VSS(VSS),.VDD(VDD),.Y(g11998),.A(g11312));
  NOT NOT1_3762(.VSS(VSS),.VDD(VDD),.Y(g12001),.A(g11315));
  NOT NOT1_3763(.VSS(VSS),.VDD(VDD),.Y(g12002),.A(g11318));
  NOT NOT1_3764(.VSS(VSS),.VDD(VDD),.Y(g12003),.A(g11321));
  NOT NOT1_3765(.VSS(VSS),.VDD(VDD),.Y(g12004),.A(g11324));
  NOT NOT1_3766(.VSS(VSS),.VDD(VDD),.Y(g12007),.A(g11327));
  NOT NOT1_3767(.VSS(VSS),.VDD(VDD),.Y(I19195),.A(g8726));
  NOT NOT1_3768(.VSS(VSS),.VDD(VDD),.Y(g12009),.A(I19195));
  NOT NOT1_3769(.VSS(VSS),.VDD(VDD),.Y(g12013),.A(g10772));
  NOT NOT1_3770(.VSS(VSS),.VDD(VDD),.Y(g12017),.A(g10100));
  NOT NOT1_3771(.VSS(VSS),.VDD(VDD),.Y(g12020),.A(g11341));
  NOT NOT1_3772(.VSS(VSS),.VDD(VDD),.Y(g12021),.A(g11344));
  NOT NOT1_3773(.VSS(VSS),.VDD(VDD),.Y(g12022),.A(g11348));
  NOT NOT1_3774(.VSS(VSS),.VDD(VDD),.Y(g12023),.A(g11351));
  NOT NOT1_3775(.VSS(VSS),.VDD(VDD),.Y(g12024),.A(g11354));
  NOT NOT1_3776(.VSS(VSS),.VDD(VDD),.Y(g12025),.A(g11355));
  NOT NOT1_3777(.VSS(VSS),.VDD(VDD),.Y(I19208),.A(g10424));
  NOT NOT1_3778(.VSS(VSS),.VDD(VDD),.Y(g12027),.A(I19208));
  NOT NOT1_3779(.VSS(VSS),.VDD(VDD),.Y(I19211),.A(g10486));
  NOT NOT1_3780(.VSS(VSS),.VDD(VDD),.Y(g12030),.A(I19211));
  NOT NOT1_3781(.VSS(VSS),.VDD(VDD),.Y(g12037),.A(g11358));
  NOT NOT1_3782(.VSS(VSS),.VDD(VDD),.Y(g12038),.A(g11361));
  NOT NOT1_3783(.VSS(VSS),.VDD(VDD),.Y(g12039),.A(g11364));
  NOT NOT1_3784(.VSS(VSS),.VDD(VDD),.Y(g12040),.A(g11367));
  NOT NOT1_3785(.VSS(VSS),.VDD(VDD),.Y(g12041),.A(g11370));
  NOT NOT1_3786(.VSS(VSS),.VDD(VDD),.Y(g12042),.A(g11373));
  NOT NOT1_3787(.VSS(VSS),.VDD(VDD),.Y(I19226),.A(g10606));
  NOT NOT1_3788(.VSS(VSS),.VDD(VDD),.Y(g12045),.A(I19226));
  NOT NOT1_3789(.VSS(VSS),.VDD(VDD),.Y(g12051),.A(g11376));
  NOT NOT1_3790(.VSS(VSS),.VDD(VDD),.Y(g12052),.A(g11379));
  NOT NOT1_3791(.VSS(VSS),.VDD(VDD),.Y(g12053),.A(g11382));
  NOT NOT1_3792(.VSS(VSS),.VDD(VDD),.Y(g12054),.A(g11386));
  NOT NOT1_3793(.VSS(VSS),.VDD(VDD),.Y(g12055),.A(g11389));
  NOT NOT1_3794(.VSS(VSS),.VDD(VDD),.Y(g12058),.A(g11392));
  NOT NOT1_3795(.VSS(VSS),.VDD(VDD),.Y(I19240),.A(g9341));
  NOT NOT1_3796(.VSS(VSS),.VDD(VDD),.Y(g12059),.A(I19240));
  NOT NOT1_3797(.VSS(VSS),.VDD(VDD),.Y(g12063),.A(g11395));
  NOT NOT1_3798(.VSS(VSS),.VDD(VDD),.Y(g12064),.A(g11398));
  NOT NOT1_3799(.VSS(VSS),.VDD(VDD),.Y(g12065),.A(g11401));
  NOT NOT1_3800(.VSS(VSS),.VDD(VDD),.Y(g12066),.A(g11404));
  NOT NOT1_3801(.VSS(VSS),.VDD(VDD),.Y(g12067),.A(g11407));
  NOT NOT1_3802(.VSS(VSS),.VDD(VDD),.Y(g12071),.A(g10783));
  NOT NOT1_3803(.VSS(VSS),.VDD(VDD),.Y(g12075),.A(g11411));
  NOT NOT1_3804(.VSS(VSS),.VDD(VDD),.Y(g12076),.A(g11414));
  NOT NOT1_3805(.VSS(VSS),.VDD(VDD),.Y(g12077),.A(g11417));
  NOT NOT1_3806(.VSS(VSS),.VDD(VDD),.Y(g12078),.A(g11422));
  NOT NOT1_3807(.VSS(VSS),.VDD(VDD),.Y(g12084),.A(g11425));
  NOT NOT1_3808(.VSS(VSS),.VDD(VDD),.Y(g12085),.A(g11428));
  NOT NOT1_3809(.VSS(VSS),.VDD(VDD),.Y(g12086),.A(g11432));
  NOT NOT1_3810(.VSS(VSS),.VDD(VDD),.Y(g12087),.A(g11435));
  NOT NOT1_3811(.VSS(VSS),.VDD(VDD),.Y(g12088),.A(g11438));
  NOT NOT1_3812(.VSS(VSS),.VDD(VDD),.Y(g12089),.A(g11441));
  NOT NOT1_3813(.VSS(VSS),.VDD(VDD),.Y(I19271),.A(g10500));
  NOT NOT1_3814(.VSS(VSS),.VDD(VDD),.Y(g12091),.A(I19271));
  NOT NOT1_3815(.VSS(VSS),.VDD(VDD),.Y(I19274),.A(g10560));
  NOT NOT1_3816(.VSS(VSS),.VDD(VDD),.Y(g12094),.A(I19274));
  NOT NOT1_3817(.VSS(VSS),.VDD(VDD),.Y(g12101),.A(g11444));
  NOT NOT1_3818(.VSS(VSS),.VDD(VDD),.Y(g12102),.A(g11447));
  NOT NOT1_3819(.VSS(VSS),.VDD(VDD),.Y(g12103),.A(g11450));
  NOT NOT1_3820(.VSS(VSS),.VDD(VDD),.Y(g12104),.A(g11453));
  NOT NOT1_3821(.VSS(VSS),.VDD(VDD),.Y(g12105),.A(g11456));
  NOT NOT1_3822(.VSS(VSS),.VDD(VDD),.Y(g12106),.A(g11459));
  NOT NOT1_3823(.VSS(VSS),.VDD(VDD),.Y(I19289),.A(g10653));
  NOT NOT1_3824(.VSS(VSS),.VDD(VDD),.Y(g12109),.A(I19289));
  NOT NOT1_3825(.VSS(VSS),.VDD(VDD),.Y(g12115),.A(g11462));
  NOT NOT1_3826(.VSS(VSS),.VDD(VDD),.Y(g12116),.A(g11465));
  NOT NOT1_3827(.VSS(VSS),.VDD(VDD),.Y(g12117),.A(g11468));
  NOT NOT1_3828(.VSS(VSS),.VDD(VDD),.Y(g12118),.A(g11472));
  NOT NOT1_3829(.VSS(VSS),.VDD(VDD),.Y(g12119),.A(g11475));
  NOT NOT1_3830(.VSS(VSS),.VDD(VDD),.Y(g12122),.A(g11478));
  NOT NOT1_3831(.VSS(VSS),.VDD(VDD),.Y(I19303),.A(g9422));
  NOT NOT1_3832(.VSS(VSS),.VDD(VDD),.Y(g12123),.A(I19303));
  NOT NOT1_3833(.VSS(VSS),.VDD(VDD),.Y(I19307),.A(g8726));
  NOT NOT1_3834(.VSS(VSS),.VDD(VDD),.Y(g12125),.A(I19307));
  NOT NOT1_3835(.VSS(VSS),.VDD(VDD),.Y(g12130),.A(g10788));
  NOT NOT1_3836(.VSS(VSS),.VDD(VDD),.Y(g12134),.A(g8321));
  NOT NOT1_3837(.VSS(VSS),.VDD(VDD),.Y(g12135),.A(g8324));
  NOT NOT1_3838(.VSS(VSS),.VDD(VDD),.Y(I19315),.A(g10424));
  NOT NOT1_3839(.VSS(VSS),.VDD(VDD),.Y(g12136),.A(I19315));
  NOT NOT1_3840(.VSS(VSS),.VDD(VDD),.Y(I19318),.A(g10486));
  NOT NOT1_3841(.VSS(VSS),.VDD(VDD),.Y(g12139),.A(I19318));
  NOT NOT1_3842(.VSS(VSS),.VDD(VDD),.Y(I19321),.A(g10549));
  NOT NOT1_3843(.VSS(VSS),.VDD(VDD),.Y(g12142),.A(I19321));
  NOT NOT1_3844(.VSS(VSS),.VDD(VDD),.Y(g12147),.A(g8330));
  NOT NOT1_3845(.VSS(VSS),.VDD(VDD),.Y(g12148),.A(g8333));
  NOT NOT1_3846(.VSS(VSS),.VDD(VDD),.Y(g12149),.A(g8336));
  NOT NOT1_3847(.VSS(VSS),.VDD(VDD),.Y(g12150),.A(g8341));
  NOT NOT1_3848(.VSS(VSS),.VDD(VDD),.Y(g12156),.A(g8344));
  NOT NOT1_3849(.VSS(VSS),.VDD(VDD),.Y(g12157),.A(g8347));
  NOT NOT1_3850(.VSS(VSS),.VDD(VDD),.Y(g12158),.A(g8351));
  NOT NOT1_3851(.VSS(VSS),.VDD(VDD),.Y(g12159),.A(g8354));
  NOT NOT1_3852(.VSS(VSS),.VDD(VDD),.Y(g12160),.A(g8357));
  NOT NOT1_3853(.VSS(VSS),.VDD(VDD),.Y(g12161),.A(g8360));
  NOT NOT1_3854(.VSS(VSS),.VDD(VDD),.Y(I19342),.A(g10574));
  NOT NOT1_3855(.VSS(VSS),.VDD(VDD),.Y(g12163),.A(I19342));
  NOT NOT1_3856(.VSS(VSS),.VDD(VDD),.Y(I19345),.A(g10617));
  NOT NOT1_3857(.VSS(VSS),.VDD(VDD),.Y(g12166),.A(I19345));
  NOT NOT1_3858(.VSS(VSS),.VDD(VDD),.Y(g12173),.A(g8363));
  NOT NOT1_3859(.VSS(VSS),.VDD(VDD),.Y(g12174),.A(g8366));
  NOT NOT1_3860(.VSS(VSS),.VDD(VDD),.Y(g12175),.A(g8369));
  NOT NOT1_3861(.VSS(VSS),.VDD(VDD),.Y(g12176),.A(g8372));
  NOT NOT1_3862(.VSS(VSS),.VDD(VDD),.Y(g12177),.A(g8375));
  NOT NOT1_3863(.VSS(VSS),.VDD(VDD),.Y(g12178),.A(g8378));
  NOT NOT1_3864(.VSS(VSS),.VDD(VDD),.Y(I19360),.A(g10683));
  NOT NOT1_3865(.VSS(VSS),.VDD(VDD),.Y(g12181),.A(I19360));
  NOT NOT1_3866(.VSS(VSS),.VDD(VDD),.Y(g12187),.A(g8285));
  NOT NOT1_3867(.VSS(VSS),.VDD(VDD),.Y(g12191),.A(g8382));
  NOT NOT1_3868(.VSS(VSS),.VDD(VDD),.Y(g12196),.A(g8388));
  NOT NOT1_3869(.VSS(VSS),.VDD(VDD),.Y(g12197),.A(g8391));
  NOT NOT1_3870(.VSS(VSS),.VDD(VDD),.Y(I19374),.A(g10500));
  NOT NOT1_3871(.VSS(VSS),.VDD(VDD),.Y(g12198),.A(I19374));
  NOT NOT1_3872(.VSS(VSS),.VDD(VDD),.Y(I19377),.A(g10560));
  NOT NOT1_3873(.VSS(VSS),.VDD(VDD),.Y(g12201),.A(I19377));
  NOT NOT1_3874(.VSS(VSS),.VDD(VDD),.Y(I19380),.A(g10606));
  NOT NOT1_3875(.VSS(VSS),.VDD(VDD),.Y(g12204),.A(I19380));
  NOT NOT1_3876(.VSS(VSS),.VDD(VDD),.Y(g12209),.A(g8397));
  NOT NOT1_3877(.VSS(VSS),.VDD(VDD),.Y(g12210),.A(g8400));
  NOT NOT1_3878(.VSS(VSS),.VDD(VDD),.Y(g12211),.A(g8403));
  NOT NOT1_3879(.VSS(VSS),.VDD(VDD),.Y(g12212),.A(g8408));
  NOT NOT1_3880(.VSS(VSS),.VDD(VDD),.Y(g12218),.A(g8411));
  NOT NOT1_3881(.VSS(VSS),.VDD(VDD),.Y(g12219),.A(g8414));
  NOT NOT1_3882(.VSS(VSS),.VDD(VDD),.Y(g12220),.A(g8418));
  NOT NOT1_3883(.VSS(VSS),.VDD(VDD),.Y(g12221),.A(g8421));
  NOT NOT1_3884(.VSS(VSS),.VDD(VDD),.Y(g12222),.A(g8424));
  NOT NOT1_3885(.VSS(VSS),.VDD(VDD),.Y(g12223),.A(g8427));
  NOT NOT1_3886(.VSS(VSS),.VDD(VDD),.Y(I19401),.A(g10631));
  NOT NOT1_3887(.VSS(VSS),.VDD(VDD),.Y(g12225),.A(I19401));
  NOT NOT1_3888(.VSS(VSS),.VDD(VDD),.Y(I19404),.A(g10664));
  NOT NOT1_3889(.VSS(VSS),.VDD(VDD),.Y(g12228),.A(I19404));
  NOT NOT1_3890(.VSS(VSS),.VDD(VDD),.Y(g12235),.A(g8294));
  NOT NOT1_3891(.VSS(VSS),.VDD(VDD),.Y(I19412),.A(g10486));
  NOT NOT1_3892(.VSS(VSS),.VDD(VDD),.Y(g12239),.A(I19412));
  NOT NOT1_3893(.VSS(VSS),.VDD(VDD),.Y(I19415),.A(g10549));
  NOT NOT1_3894(.VSS(VSS),.VDD(VDD),.Y(g12242),.A(I19415));
  NOT NOT1_3895(.VSS(VSS),.VDD(VDD),.Y(g12246),.A(g8434));
  NOT NOT1_3896(.VSS(VSS),.VDD(VDD),.Y(g12251),.A(g8440));
  NOT NOT1_3897(.VSS(VSS),.VDD(VDD),.Y(g12252),.A(g8443));
  NOT NOT1_3898(.VSS(VSS),.VDD(VDD),.Y(I19426),.A(g10574));
  NOT NOT1_3899(.VSS(VSS),.VDD(VDD),.Y(g12253),.A(I19426));
  NOT NOT1_3900(.VSS(VSS),.VDD(VDD),.Y(I19429),.A(g10617));
  NOT NOT1_3901(.VSS(VSS),.VDD(VDD),.Y(g12256),.A(I19429));
  NOT NOT1_3902(.VSS(VSS),.VDD(VDD),.Y(I19432),.A(g10653));
  NOT NOT1_3903(.VSS(VSS),.VDD(VDD),.Y(g12259),.A(I19432));
  NOT NOT1_3904(.VSS(VSS),.VDD(VDD),.Y(g12264),.A(g8449));
  NOT NOT1_3905(.VSS(VSS),.VDD(VDD),.Y(g12265),.A(g8452));
  NOT NOT1_3906(.VSS(VSS),.VDD(VDD),.Y(g12266),.A(g8455));
  NOT NOT1_3907(.VSS(VSS),.VDD(VDD),.Y(g12267),.A(g8460));
  NOT NOT1_3908(.VSS(VSS),.VDD(VDD),.Y(g12275),.A(g8303));
  NOT NOT1_3909(.VSS(VSS),.VDD(VDD),.Y(I19449),.A(g10424));
  NOT NOT1_3910(.VSS(VSS),.VDD(VDD),.Y(g12279),.A(I19449));
  NOT NOT1_3911(.VSS(VSS),.VDD(VDD),.Y(I19452),.A(g10560));
  NOT NOT1_3912(.VSS(VSS),.VDD(VDD),.Y(g12282),.A(I19452));
  NOT NOT1_3913(.VSS(VSS),.VDD(VDD),.Y(I19455),.A(g10606));
  NOT NOT1_3914(.VSS(VSS),.VDD(VDD),.Y(g12285),.A(I19455));
  NOT NOT1_3915(.VSS(VSS),.VDD(VDD),.Y(g12289),.A(g8469));
  NOT NOT1_3916(.VSS(VSS),.VDD(VDD),.Y(g12294),.A(g8475));
  NOT NOT1_3917(.VSS(VSS),.VDD(VDD),.Y(g12295),.A(g8478));
  NOT NOT1_3918(.VSS(VSS),.VDD(VDD),.Y(I19466),.A(g10631));
  NOT NOT1_3919(.VSS(VSS),.VDD(VDD),.Y(g12296),.A(I19466));
  NOT NOT1_3920(.VSS(VSS),.VDD(VDD),.Y(I19469),.A(g10664));
  NOT NOT1_3921(.VSS(VSS),.VDD(VDD),.Y(g12299),.A(I19469));
  NOT NOT1_3922(.VSS(VSS),.VDD(VDD),.Y(I19472),.A(g10683));
  NOT NOT1_3923(.VSS(VSS),.VDD(VDD),.Y(g12302),.A(I19472));
  NOT NOT1_3924(.VSS(VSS),.VDD(VDD),.Y(g12308),.A(g8312));
  NOT NOT1_3925(.VSS(VSS),.VDD(VDD),.Y(I19479),.A(g10549));
  NOT NOT1_3926(.VSS(VSS),.VDD(VDD),.Y(g12312),.A(I19479));
  NOT NOT1_3927(.VSS(VSS),.VDD(VDD),.Y(I19482),.A(g10500));
  NOT NOT1_3928(.VSS(VSS),.VDD(VDD),.Y(g12315),.A(I19482));
  NOT NOT1_3929(.VSS(VSS),.VDD(VDD),.Y(I19485),.A(g10617));
  NOT NOT1_3930(.VSS(VSS),.VDD(VDD),.Y(g12318),.A(I19485));
  NOT NOT1_3931(.VSS(VSS),.VDD(VDD),.Y(I19488),.A(g10653));
  NOT NOT1_3932(.VSS(VSS),.VDD(VDD),.Y(g12321),.A(I19488));
  NOT NOT1_3933(.VSS(VSS),.VDD(VDD),.Y(g12325),.A(g8494));
  NOT NOT1_3934(.VSS(VSS),.VDD(VDD),.Y(g12332),.A(g10829));
  NOT NOT1_3935(.VSS(VSS),.VDD(VDD),.Y(I19500),.A(g10424));
  NOT NOT1_3936(.VSS(VSS),.VDD(VDD),.Y(g12333),.A(I19500));
  NOT NOT1_3937(.VSS(VSS),.VDD(VDD),.Y(I19503),.A(g10486));
  NOT NOT1_3938(.VSS(VSS),.VDD(VDD),.Y(g12336),.A(I19503));
  NOT NOT1_3939(.VSS(VSS),.VDD(VDD),.Y(I19507),.A(g10606));
  NOT NOT1_3940(.VSS(VSS),.VDD(VDD),.Y(g12340),.A(I19507));
  NOT NOT1_3941(.VSS(VSS),.VDD(VDD),.Y(I19510),.A(g10574));
  NOT NOT1_3942(.VSS(VSS),.VDD(VDD),.Y(g12343),.A(I19510));
  NOT NOT1_3943(.VSS(VSS),.VDD(VDD),.Y(I19513),.A(g10664));
  NOT NOT1_3944(.VSS(VSS),.VDD(VDD),.Y(g12346),.A(I19513));
  NOT NOT1_3945(.VSS(VSS),.VDD(VDD),.Y(I19516),.A(g10683));
  NOT NOT1_3946(.VSS(VSS),.VDD(VDD),.Y(g12349),.A(I19516));
  NOT NOT1_3947(.VSS(VSS),.VDD(VDD),.Y(g12354),.A(g8381));
  NOT NOT1_3948(.VSS(VSS),.VDD(VDD),.Y(g12362),.A(g10866));
  NOT NOT1_3949(.VSS(VSS),.VDD(VDD),.Y(I19523),.A(g10500));
  NOT NOT1_3950(.VSS(VSS),.VDD(VDD),.Y(g12363),.A(I19523));
  NOT NOT1_3951(.VSS(VSS),.VDD(VDD),.Y(I19526),.A(g10560));
  NOT NOT1_3952(.VSS(VSS),.VDD(VDD),.Y(g12366),.A(I19526));
  NOT NOT1_3953(.VSS(VSS),.VDD(VDD),.Y(I19530),.A(g10653));
  NOT NOT1_3954(.VSS(VSS),.VDD(VDD),.Y(g12370),.A(I19530));
  NOT NOT1_3955(.VSS(VSS),.VDD(VDD),.Y(I19533),.A(g10631));
  NOT NOT1_3956(.VSS(VSS),.VDD(VDD),.Y(g12373),.A(I19533));
  NOT NOT1_3957(.VSS(VSS),.VDD(VDD),.Y(g12378),.A(g10847));
  NOT NOT1_3958(.VSS(VSS),.VDD(VDD),.Y(I19539),.A(g10549));
  NOT NOT1_3959(.VSS(VSS),.VDD(VDD),.Y(g12379),.A(I19539));
  NOT NOT1_3960(.VSS(VSS),.VDD(VDD),.Y(I19542),.A(g10574));
  NOT NOT1_3961(.VSS(VSS),.VDD(VDD),.Y(g12382),.A(I19542));
  NOT NOT1_3962(.VSS(VSS),.VDD(VDD),.Y(I19545),.A(g10617));
  NOT NOT1_3963(.VSS(VSS),.VDD(VDD),.Y(g12385),.A(I19545));
  NOT NOT1_3964(.VSS(VSS),.VDD(VDD),.Y(I19549),.A(g10683));
  NOT NOT1_3965(.VSS(VSS),.VDD(VDD),.Y(g12389),.A(I19549));
  NOT NOT1_3966(.VSS(VSS),.VDD(VDD),.Y(I19552),.A(g8430));
  NOT NOT1_3967(.VSS(VSS),.VDD(VDD),.Y(g12392),.A(I19552));
  NOT NOT1_3968(.VSS(VSS),.VDD(VDD),.Y(g12408),.A(g11020));
  NOT NOT1_3969(.VSS(VSS),.VDD(VDD),.Y(I19557),.A(g10606));
  NOT NOT1_3970(.VSS(VSS),.VDD(VDD),.Y(g12409),.A(I19557));
  NOT NOT1_3971(.VSS(VSS),.VDD(VDD),.Y(I19560),.A(g10631));
  NOT NOT1_3972(.VSS(VSS),.VDD(VDD),.Y(g12412),.A(I19560));
  NOT NOT1_3973(.VSS(VSS),.VDD(VDD),.Y(I19563),.A(g10664));
  NOT NOT1_3974(.VSS(VSS),.VDD(VDD),.Y(g12415),.A(I19563));
  NOT NOT1_3975(.VSS(VSS),.VDD(VDD),.Y(g12420),.A(g10986));
  NOT NOT1_3976(.VSS(VSS),.VDD(VDD),.Y(I19569),.A(g10653));
  NOT NOT1_3977(.VSS(VSS),.VDD(VDD),.Y(g12421),.A(I19569));
  NOT NOT1_3978(.VSS(VSS),.VDD(VDD),.Y(g12424),.A(g10962));
  NOT NOT1_3979(.VSS(VSS),.VDD(VDD),.Y(I19573),.A(g8835));
  NOT NOT1_3980(.VSS(VSS),.VDD(VDD),.Y(g12425),.A(I19573));
  NOT NOT1_3981(.VSS(VSS),.VDD(VDD),.Y(I19576),.A(g10683));
  NOT NOT1_3982(.VSS(VSS),.VDD(VDD),.Y(g12426),.A(I19576));
  NOT NOT1_3983(.VSS(VSS),.VDD(VDD),.Y(g12430),.A(g10905));
  NOT NOT1_3984(.VSS(VSS),.VDD(VDD),.Y(I19582),.A(g8862));
  NOT NOT1_3985(.VSS(VSS),.VDD(VDD),.Y(g12432),.A(I19582));
  NOT NOT1_3986(.VSS(VSS),.VDD(VDD),.Y(g12434),.A(g10929));
  NOT NOT1_3987(.VSS(VSS),.VDD(VDD),.Y(I19587),.A(g9173));
  NOT NOT1_3988(.VSS(VSS),.VDD(VDD),.Y(g12435),.A(I19587));
  NOT NOT1_3989(.VSS(VSS),.VDD(VDD),.Y(I19591),.A(g8900));
  NOT NOT1_3990(.VSS(VSS),.VDD(VDD),.Y(g12437),.A(I19591));
  NOT NOT1_3991(.VSS(VSS),.VDD(VDD),.Y(g12438),.A(g10846));
  NOT NOT1_3992(.VSS(VSS),.VDD(VDD),.Y(I19595),.A(g10810));
  NOT NOT1_3993(.VSS(VSS),.VDD(VDD),.Y(g12439),.A(I19595));
  NOT NOT1_3994(.VSS(VSS),.VDD(VDD),.Y(I19598),.A(g9215));
  NOT NOT1_3995(.VSS(VSS),.VDD(VDD),.Y(g12440),.A(I19598));
  NOT NOT1_3996(.VSS(VSS),.VDD(VDD),.Y(I19602),.A(g8940));
  NOT NOT1_3997(.VSS(VSS),.VDD(VDD),.Y(g12442),.A(I19602));
  NOT NOT1_3998(.VSS(VSS),.VDD(VDD),.Y(I19605),.A(g10797));
  NOT NOT1_3999(.VSS(VSS),.VDD(VDD),.Y(g12443),.A(I19605));
  NOT NOT1_4000(.VSS(VSS),.VDD(VDD),.Y(I19608),.A(g10831));
  NOT NOT1_4001(.VSS(VSS),.VDD(VDD),.Y(g12444),.A(I19608));
  NOT NOT1_4002(.VSS(VSS),.VDD(VDD),.Y(I19611),.A(g9276));
  NOT NOT1_4003(.VSS(VSS),.VDD(VDD),.Y(g12445),.A(I19611));
  NOT NOT1_4004(.VSS(VSS),.VDD(VDD),.Y(I19615),.A(g10789));
  NOT NOT1_4005(.VSS(VSS),.VDD(VDD),.Y(g12447),.A(I19615));
  NOT NOT1_4006(.VSS(VSS),.VDD(VDD),.Y(I19618),.A(g10814));
  NOT NOT1_4007(.VSS(VSS),.VDD(VDD),.Y(g12448),.A(I19618));
  NOT NOT1_4008(.VSS(VSS),.VDD(VDD),.Y(I19621),.A(g10851));
  NOT NOT1_4009(.VSS(VSS),.VDD(VDD),.Y(g12449),.A(I19621));
  NOT NOT1_4010(.VSS(VSS),.VDD(VDD),.Y(I19624),.A(g9354));
  NOT NOT1_4011(.VSS(VSS),.VDD(VDD),.Y(g12450),.A(I19624));
  NOT NOT1_4012(.VSS(VSS),.VDD(VDD),.Y(I19628),.A(g10784));
  NOT NOT1_4013(.VSS(VSS),.VDD(VDD),.Y(g12452),.A(I19628));
  NOT NOT1_4014(.VSS(VSS),.VDD(VDD),.Y(I19631),.A(g10801));
  NOT NOT1_4015(.VSS(VSS),.VDD(VDD),.Y(g12453),.A(I19631));
  NOT NOT1_4016(.VSS(VSS),.VDD(VDD),.Y(I19634),.A(g10835));
  NOT NOT1_4017(.VSS(VSS),.VDD(VDD),.Y(g12454),.A(I19634));
  NOT NOT1_4018(.VSS(VSS),.VDD(VDD),.Y(I19637),.A(g10872));
  NOT NOT1_4019(.VSS(VSS),.VDD(VDD),.Y(g12455),.A(I19637));
  NOT NOT1_4020(.VSS(VSS),.VDD(VDD),.Y(g12456),.A(g8602));
  NOT NOT1_4021(.VSS(VSS),.VDD(VDD),.Y(I19642),.A(g10793));
  NOT NOT1_4022(.VSS(VSS),.VDD(VDD),.Y(g12460),.A(I19642));
  NOT NOT1_4023(.VSS(VSS),.VDD(VDD),.Y(I19645),.A(g10818));
  NOT NOT1_4024(.VSS(VSS),.VDD(VDD),.Y(g12461),.A(I19645));
  NOT NOT1_4025(.VSS(VSS),.VDD(VDD),.Y(I19648),.A(g10855));
  NOT NOT1_4026(.VSS(VSS),.VDD(VDD),.Y(g12462),.A(I19648));
  NOT NOT1_4027(.VSS(VSS),.VDD(VDD),.Y(g12463),.A(g10730));
  NOT NOT1_4028(.VSS(VSS),.VDD(VDD),.Y(g12466),.A(g8614));
  NOT NOT1_4029(.VSS(VSS),.VDD(VDD),.Y(I19654),.A(g10805));
  NOT NOT1_4030(.VSS(VSS),.VDD(VDD),.Y(g12470),.A(I19654));
  NOT NOT1_4031(.VSS(VSS),.VDD(VDD),.Y(I19657),.A(g10839));
  NOT NOT1_4032(.VSS(VSS),.VDD(VDD),.Y(g12471),.A(I19657));
  NOT NOT1_4033(.VSS(VSS),.VDD(VDD),.Y(g12472),.A(g8617));
  NOT NOT1_4034(.VSS(VSS),.VDD(VDD),.Y(g12473),.A(g8580));
  NOT NOT1_4035(.VSS(VSS),.VDD(VDD),.Y(g12476),.A(g8622));
  NOT NOT1_4036(.VSS(VSS),.VDD(VDD),.Y(g12478),.A(g10749));
  NOT NOT1_4037(.VSS(VSS),.VDD(VDD),.Y(g12481),.A(g8627));
  NOT NOT1_4038(.VSS(VSS),.VDD(VDD),.Y(I19667),.A(g10822));
  NOT NOT1_4039(.VSS(VSS),.VDD(VDD),.Y(g12485),.A(I19667));
  NOT NOT1_4040(.VSS(VSS),.VDD(VDD),.Y(g12490),.A(g8587));
  NOT NOT1_4041(.VSS(VSS),.VDD(VDD),.Y(g12493),.A(g8632));
  NOT NOT1_4042(.VSS(VSS),.VDD(VDD),.Y(g12495),.A(g10767));
  NOT NOT1_4043(.VSS(VSS),.VDD(VDD),.Y(g12498),.A(g8637));
  NOT NOT1_4044(.VSS(VSS),.VDD(VDD),.Y(g12502),.A(g8640));
  NOT NOT1_4045(.VSS(VSS),.VDD(VDD),.Y(g12504),.A(g8643));
  NOT NOT1_4046(.VSS(VSS),.VDD(VDD),.Y(g12505),.A(g8646));
  NOT NOT1_4047(.VSS(VSS),.VDD(VDD),.Y(g12510),.A(g8594));
  NOT NOT1_4048(.VSS(VSS),.VDD(VDD),.Y(g12513),.A(g8651));
  NOT NOT1_4049(.VSS(VSS),.VDD(VDD),.Y(g12515),.A(g10773));
  NOT NOT1_4050(.VSS(VSS),.VDD(VDD),.Y(g12518),.A(g8655));
  NOT NOT1_4051(.VSS(VSS),.VDD(VDD),.Y(I19689),.A(g10016));
  NOT NOT1_4052(.VSS(VSS),.VDD(VDD),.Y(g12519),.A(I19689));
  NOT NOT1_4053(.VSS(VSS),.VDD(VDD),.Y(g12521),.A(g8659));
  NOT NOT1_4054(.VSS(VSS),.VDD(VDD),.Y(g12522),.A(g8662));
  NOT NOT1_4055(.VSS(VSS),.VDD(VDD),.Y(g12527),.A(g8605));
  NOT NOT1_4056(.VSS(VSS),.VDD(VDD),.Y(g12530),.A(g8667));
  NOT NOT1_4057(.VSS(VSS),.VDD(VDD),.Y(g12532),.A(g8670));
  NOT NOT1_4058(.VSS(VSS),.VDD(VDD),.Y(g12533),.A(g8673));
  NOT NOT1_4059(.VSS(VSS),.VDD(VDD),.Y(I19702),.A(g10125));
  NOT NOT1_4060(.VSS(VSS),.VDD(VDD),.Y(g12534),.A(I19702));
  NOT NOT1_4061(.VSS(VSS),.VDD(VDD),.Y(g12536),.A(g8678));
  NOT NOT1_4062(.VSS(VSS),.VDD(VDD),.Y(g12537),.A(g8681));
  NOT NOT1_4063(.VSS(VSS),.VDD(VDD),.Y(g12542),.A(g8684));
  NOT NOT1_4064(.VSS(VSS),.VDD(VDD),.Y(I19711),.A(g10230));
  NOT NOT1_4065(.VSS(VSS),.VDD(VDD),.Y(g12543),.A(I19711));
  NOT NOT1_4066(.VSS(VSS),.VDD(VDD),.Y(g12545),.A(g8690));
  NOT NOT1_4067(.VSS(VSS),.VDD(VDD),.Y(g12546),.A(g8693));
  NOT NOT1_4068(.VSS(VSS),.VDD(VDD),.Y(g12547),.A(g8696));
  NOT NOT1_4069(.VSS(VSS),.VDD(VDD),.Y(I19718),.A(g8726));
  NOT NOT1_4070(.VSS(VSS),.VDD(VDD),.Y(g12548),.A(I19718));
  NOT NOT1_4071(.VSS(VSS),.VDD(VDD),.Y(g12551),.A(g8700));
  NOT NOT1_4072(.VSS(VSS),.VDD(VDD),.Y(I19722),.A(g10332));
  NOT NOT1_4073(.VSS(VSS),.VDD(VDD),.Y(g12552),.A(I19722));
  NOT NOT1_4074(.VSS(VSS),.VDD(VDD),.Y(g12553),.A(g8708));
  NOT NOT1_4075(.VSS(VSS),.VDD(VDD),.Y(g12554),.A(g8711));
  NOT NOT1_4076(.VSS(VSS),.VDD(VDD),.Y(I19727),.A(g8726));
  NOT NOT1_4077(.VSS(VSS),.VDD(VDD),.Y(g12555),.A(I19727));
  NOT NOT1_4078(.VSS(VSS),.VDD(VDD),.Y(g12558),.A(g8714));
  NOT NOT1_4079(.VSS(VSS),.VDD(VDD),.Y(g12559),.A(g8719));
  NOT NOT1_4080(.VSS(VSS),.VDD(VDD),.Y(g12560),.A(g8745));
  NOT NOT1_4081(.VSS(VSS),.VDD(VDD),.Y(I19733),.A(g8726));
  NOT NOT1_4082(.VSS(VSS),.VDD(VDD),.Y(g12561),.A(I19733));
  NOT NOT1_4083(.VSS(VSS),.VDD(VDD),.Y(I19736),.A(g9184));
  NOT NOT1_4084(.VSS(VSS),.VDD(VDD),.Y(g12564),.A(I19736));
  NOT NOT1_4085(.VSS(VSS),.VDD(VDD),.Y(I19739),.A(g10694));
  NOT NOT1_4086(.VSS(VSS),.VDD(VDD),.Y(g12565),.A(I19739));
  NOT NOT1_4087(.VSS(VSS),.VDD(VDD),.Y(g12596),.A(g8748));
  NOT NOT1_4088(.VSS(VSS),.VDD(VDD),.Y(g12597),.A(g8752));
  NOT NOT1_4089(.VSS(VSS),.VDD(VDD),.Y(g12598),.A(g8757));
  NOT NOT1_4090(.VSS(VSS),.VDD(VDD),.Y(g12599),.A(g8763));
  NOT NOT1_4091(.VSS(VSS),.VDD(VDD),.Y(g12600),.A(g8766));
  NOT NOT1_4092(.VSS(VSS),.VDD(VDD),.Y(I19747),.A(g8726));
  NOT NOT1_4093(.VSS(VSS),.VDD(VDD),.Y(g12601),.A(I19747));
  NOT NOT1_4094(.VSS(VSS),.VDD(VDD),.Y(I19750),.A(g8726));
  NOT NOT1_4095(.VSS(VSS),.VDD(VDD),.Y(g12604),.A(I19750));
  NOT NOT1_4096(.VSS(VSS),.VDD(VDD),.Y(I19753),.A(g9229));
  NOT NOT1_4097(.VSS(VSS),.VDD(VDD),.Y(g12607),.A(I19753));
  NOT NOT1_4098(.VSS(VSS),.VDD(VDD),.Y(I19756),.A(g10424));
  NOT NOT1_4099(.VSS(VSS),.VDD(VDD),.Y(g12608),.A(I19756));
  NOT NOT1_4100(.VSS(VSS),.VDD(VDD),.Y(I19759),.A(g10714));
  NOT NOT1_4101(.VSS(VSS),.VDD(VDD),.Y(g12611),.A(I19759));
  NOT NOT1_4102(.VSS(VSS),.VDD(VDD),.Y(g12642),.A(g8771));
  NOT NOT1_4103(.VSS(VSS),.VDD(VDD),.Y(g12643),.A(g8775));
  NOT NOT1_4104(.VSS(VSS),.VDD(VDD),.Y(g12644),.A(g8780));
  NOT NOT1_4105(.VSS(VSS),.VDD(VDD),.Y(g12645),.A(g8785));
  NOT NOT1_4106(.VSS(VSS),.VDD(VDD),.Y(g12646),.A(g8788));
  NOT NOT1_4107(.VSS(VSS),.VDD(VDD),.Y(I19767),.A(g8726));
  NOT NOT1_4108(.VSS(VSS),.VDD(VDD),.Y(g12647),.A(I19767));
  NOT NOT1_4109(.VSS(VSS),.VDD(VDD),.Y(I19771),.A(g10038));
  NOT NOT1_4110(.VSS(VSS),.VDD(VDD),.Y(g12651),.A(I19771));
  NOT NOT1_4111(.VSS(VSS),.VDD(VDD),.Y(I19774),.A(g10500));
  NOT NOT1_4112(.VSS(VSS),.VDD(VDD),.Y(g12654),.A(I19774));
  NOT NOT1_4113(.VSS(VSS),.VDD(VDD),.Y(I19777),.A(g10735));
  NOT NOT1_4114(.VSS(VSS),.VDD(VDD),.Y(g12657),.A(I19777));
  NOT NOT1_4115(.VSS(VSS),.VDD(VDD),.Y(g12688),.A(g8794));
  NOT NOT1_4116(.VSS(VSS),.VDD(VDD),.Y(g12689),.A(g8798));
  NOT NOT1_4117(.VSS(VSS),.VDD(VDD),.Y(g12690),.A(g8802));
  NOT NOT1_4118(.VSS(VSS),.VDD(VDD),.Y(g12691),.A(g8805));
  NOT NOT1_4119(.VSS(VSS),.VDD(VDD),.Y(I19784),.A(g8726));
  NOT NOT1_4120(.VSS(VSS),.VDD(VDD),.Y(g12692),.A(I19784));
  NOT NOT1_4121(.VSS(VSS),.VDD(VDD),.Y(I19787),.A(g8726));
  NOT NOT1_4122(.VSS(VSS),.VDD(VDD),.Y(g12695),.A(I19787));
  NOT NOT1_4123(.VSS(VSS),.VDD(VDD),.Y(I19791),.A(g10486));
  NOT NOT1_4124(.VSS(VSS),.VDD(VDD),.Y(g12699),.A(I19791));
  NOT NOT1_4125(.VSS(VSS),.VDD(VDD),.Y(I19794),.A(g10676));
  NOT NOT1_4126(.VSS(VSS),.VDD(VDD),.Y(g12702),.A(I19794));
  NOT NOT1_4127(.VSS(VSS),.VDD(VDD),.Y(I19797),.A(g10147));
  NOT NOT1_4128(.VSS(VSS),.VDD(VDD),.Y(g12705),.A(I19797));
  NOT NOT1_4129(.VSS(VSS),.VDD(VDD),.Y(I19800),.A(g10574));
  NOT NOT1_4130(.VSS(VSS),.VDD(VDD),.Y(g12708),.A(I19800));
  NOT NOT1_4131(.VSS(VSS),.VDD(VDD),.Y(I19803),.A(g10754));
  NOT NOT1_4132(.VSS(VSS),.VDD(VDD),.Y(g12711),.A(I19803));
  NOT NOT1_4133(.VSS(VSS),.VDD(VDD),.Y(g12742),.A(g8813));
  NOT NOT1_4134(.VSS(VSS),.VDD(VDD),.Y(g12743),.A(g8817));
  NOT NOT1_4135(.VSS(VSS),.VDD(VDD),.Y(I19808),.A(g8726));
  NOT NOT1_4136(.VSS(VSS),.VDD(VDD),.Y(g12744),.A(I19808));
  NOT NOT1_4137(.VSS(VSS),.VDD(VDD),.Y(g12748),.A(g8823));
  NOT NOT1_4138(.VSS(VSS),.VDD(VDD),.Y(I19813),.A(g10649));
  NOT NOT1_4139(.VSS(VSS),.VDD(VDD),.Y(g12749),.A(I19813));
  NOT NOT1_4140(.VSS(VSS),.VDD(VDD),.Y(I19816),.A(g10703));
  NOT NOT1_4141(.VSS(VSS),.VDD(VDD),.Y(g12752),.A(I19816));
  NOT NOT1_4142(.VSS(VSS),.VDD(VDD),.Y(I19820),.A(g10560));
  NOT NOT1_4143(.VSS(VSS),.VDD(VDD),.Y(g12756),.A(I19820));
  NOT NOT1_4144(.VSS(VSS),.VDD(VDD),.Y(I19823),.A(g10705));
  NOT NOT1_4145(.VSS(VSS),.VDD(VDD),.Y(g12759),.A(I19823));
  NOT NOT1_4146(.VSS(VSS),.VDD(VDD),.Y(I19826),.A(g10252));
  NOT NOT1_4147(.VSS(VSS),.VDD(VDD),.Y(g12762),.A(I19826));
  NOT NOT1_4148(.VSS(VSS),.VDD(VDD),.Y(I19829),.A(g10631));
  NOT NOT1_4149(.VSS(VSS),.VDD(VDD),.Y(g12765),.A(I19829));
  NOT NOT1_4150(.VSS(VSS),.VDD(VDD),.Y(g12768),.A(g8829));
  NOT NOT1_4151(.VSS(VSS),.VDD(VDD),.Y(I19833),.A(g8726));
  NOT NOT1_4152(.VSS(VSS),.VDD(VDD),.Y(g12769),.A(I19833));
  NOT NOT1_4153(.VSS(VSS),.VDD(VDD),.Y(I19836),.A(g8726));
  NOT NOT1_4154(.VSS(VSS),.VDD(VDD),.Y(g12772),.A(I19836));
  NOT NOT1_4155(.VSS(VSS),.VDD(VDD),.Y(g12775),.A(g8832));
  NOT NOT1_4156(.VSS(VSS),.VDD(VDD),.Y(g12776),.A(g10766));
  NOT NOT1_4157(.VSS(VSS),.VDD(VDD),.Y(g12782),.A(g8836));
  NOT NOT1_4158(.VSS(VSS),.VDD(VDD),.Y(I19844),.A(g8533));
  NOT NOT1_4159(.VSS(VSS),.VDD(VDD),.Y(g12783),.A(I19844));
  NOT NOT1_4160(.VSS(VSS),.VDD(VDD),.Y(I19847),.A(g10677));
  NOT NOT1_4161(.VSS(VSS),.VDD(VDD),.Y(g12786),.A(I19847));
  NOT NOT1_4162(.VSS(VSS),.VDD(VDD),.Y(g12790),.A(g8847));
  NOT NOT1_4163(.VSS(VSS),.VDD(VDD),.Y(I19852),.A(g10679));
  NOT NOT1_4164(.VSS(VSS),.VDD(VDD),.Y(g12791),.A(I19852));
  NOT NOT1_4165(.VSS(VSS),.VDD(VDD),.Y(I19855),.A(g10723));
  NOT NOT1_4166(.VSS(VSS),.VDD(VDD),.Y(g12794),.A(I19855));
  NOT NOT1_4167(.VSS(VSS),.VDD(VDD),.Y(I19859),.A(g10617));
  NOT NOT1_4168(.VSS(VSS),.VDD(VDD),.Y(g12798),.A(I19859));
  NOT NOT1_4169(.VSS(VSS),.VDD(VDD),.Y(I19862),.A(g10725));
  NOT NOT1_4170(.VSS(VSS),.VDD(VDD),.Y(g12801),.A(I19862));
  NOT NOT1_4171(.VSS(VSS),.VDD(VDD),.Y(I19865),.A(g10354));
  NOT NOT1_4172(.VSS(VSS),.VDD(VDD),.Y(g12804),.A(I19865));
  NOT NOT1_4173(.VSS(VSS),.VDD(VDD),.Y(g12807),.A(g8853));
  NOT NOT1_4174(.VSS(VSS),.VDD(VDD),.Y(I19869),.A(g8726));
  NOT NOT1_4175(.VSS(VSS),.VDD(VDD),.Y(g12808),.A(I19869));
  NOT NOT1_4176(.VSS(VSS),.VDD(VDD),.Y(I19872),.A(g8317));
  NOT NOT1_4177(.VSS(VSS),.VDD(VDD),.Y(g12811),.A(I19872));
  NOT NOT1_4178(.VSS(VSS),.VDD(VDD),.Y(g12815),.A(g8856));
  NOT NOT1_4179(.VSS(VSS),.VDD(VDD),.Y(I19877),.A(g8547));
  NOT NOT1_4180(.VSS(VSS),.VDD(VDD),.Y(g12816),.A(I19877));
  NOT NOT1_4181(.VSS(VSS),.VDD(VDD),.Y(g12821),.A(g8863));
  NOT NOT1_4182(.VSS(VSS),.VDD(VDD),.Y(I19883),.A(g8550));
  NOT NOT1_4183(.VSS(VSS),.VDD(VDD),.Y(g12822),.A(I19883));
  NOT NOT1_4184(.VSS(VSS),.VDD(VDD),.Y(I19886),.A(g10706));
  NOT NOT1_4185(.VSS(VSS),.VDD(VDD),.Y(g12825),.A(I19886));
  NOT NOT1_4186(.VSS(VSS),.VDD(VDD),.Y(g12829),.A(g8874));
  NOT NOT1_4187(.VSS(VSS),.VDD(VDD),.Y(I19891),.A(g10708));
  NOT NOT1_4188(.VSS(VSS),.VDD(VDD),.Y(g12830),.A(I19891));
  NOT NOT1_4189(.VSS(VSS),.VDD(VDD),.Y(I19894),.A(g10744));
  NOT NOT1_4190(.VSS(VSS),.VDD(VDD),.Y(g12833),.A(I19894));
  NOT NOT1_4191(.VSS(VSS),.VDD(VDD),.Y(I19898),.A(g10664));
  NOT NOT1_4192(.VSS(VSS),.VDD(VDD),.Y(g12837),.A(I19898));
  NOT NOT1_4193(.VSS(VSS),.VDD(VDD),.Y(I19901),.A(g10746));
  NOT NOT1_4194(.VSS(VSS),.VDD(VDD),.Y(g12840),.A(I19901));
  NOT NOT1_4195(.VSS(VSS),.VDD(VDD),.Y(g12843),.A(g8879));
  NOT NOT1_4196(.VSS(VSS),.VDD(VDD),.Y(I19905),.A(g8726));
  NOT NOT1_4197(.VSS(VSS),.VDD(VDD),.Y(g12844),.A(I19905));
  NOT NOT1_4198(.VSS(VSS),.VDD(VDD),.Y(g12847),.A(g8882));
  NOT NOT1_4199(.VSS(VSS),.VDD(VDD),.Y(g12848),.A(g11059));
  NOT NOT1_4200(.VSS(VSS),.VDD(VDD),.Y(g12850),.A(g8885));
  NOT NOT1_4201(.VSS(VSS),.VDD(VDD),.Y(g12851),.A(g8888));
  NOT NOT1_4202(.VSS(VSS),.VDD(VDD),.Y(g12853),.A(g8894));
  NOT NOT1_4203(.VSS(VSS),.VDD(VDD),.Y(I19915),.A(g8560));
  NOT NOT1_4204(.VSS(VSS),.VDD(VDD),.Y(g12854),.A(I19915));
  NOT NOT1_4205(.VSS(VSS),.VDD(VDD),.Y(g12859),.A(g8901));
  NOT NOT1_4206(.VSS(VSS),.VDD(VDD),.Y(I19921),.A(g8563));
  NOT NOT1_4207(.VSS(VSS),.VDD(VDD),.Y(g12860),.A(I19921));
  NOT NOT1_4208(.VSS(VSS),.VDD(VDD),.Y(I19924),.A(g10726));
  NOT NOT1_4209(.VSS(VSS),.VDD(VDD),.Y(g12863),.A(I19924));
  NOT NOT1_4210(.VSS(VSS),.VDD(VDD),.Y(g12867),.A(g8912));
  NOT NOT1_4211(.VSS(VSS),.VDD(VDD),.Y(I19929),.A(g10728));
  NOT NOT1_4212(.VSS(VSS),.VDD(VDD),.Y(g12868),.A(I19929));
  NOT NOT1_4213(.VSS(VSS),.VDD(VDD),.Y(I19932),.A(g10763));
  NOT NOT1_4214(.VSS(VSS),.VDD(VDD),.Y(g12871),.A(I19932));
  NOT NOT1_4215(.VSS(VSS),.VDD(VDD),.Y(g12874),.A(g8915));
  NOT NOT1_4216(.VSS(VSS),.VDD(VDD),.Y(g12875),.A(g10779));
  NOT NOT1_4217(.VSS(VSS),.VDD(VDD),.Y(g12881),.A(g8918));
  NOT NOT1_4218(.VSS(VSS),.VDD(VDD),.Y(g12882),.A(g8921));
  NOT NOT1_4219(.VSS(VSS),.VDD(VDD),.Y(g12891),.A(g8925));
  NOT NOT1_4220(.VSS(VSS),.VDD(VDD),.Y(g12892),.A(g8928));
  NOT NOT1_4221(.VSS(VSS),.VDD(VDD),.Y(g12894),.A(g8934));
  NOT NOT1_4222(.VSS(VSS),.VDD(VDD),.Y(I19952),.A(g8571));
  NOT NOT1_4223(.VSS(VSS),.VDD(VDD),.Y(g12895),.A(I19952));
  NOT NOT1_4224(.VSS(VSS),.VDD(VDD),.Y(g12900),.A(g8941));
  NOT NOT1_4225(.VSS(VSS),.VDD(VDD),.Y(I19958),.A(g8574));
  NOT NOT1_4226(.VSS(VSS),.VDD(VDD),.Y(g12901),.A(I19958));
  NOT NOT1_4227(.VSS(VSS),.VDD(VDD),.Y(I19961),.A(g10747));
  NOT NOT1_4228(.VSS(VSS),.VDD(VDD),.Y(g12904),.A(I19961));
  NOT NOT1_4229(.VSS(VSS),.VDD(VDD),.Y(g12907),.A(g8949));
  NOT NOT1_4230(.VSS(VSS),.VDD(VDD),.Y(g12909),.A(g10904));
  NOT NOT1_4231(.VSS(VSS),.VDD(VDD),.Y(g12914),.A(g8952));
  NOT NOT1_4232(.VSS(VSS),.VDD(VDD),.Y(g12915),.A(g8955));
  NOT NOT1_4233(.VSS(VSS),.VDD(VDD),.Y(g12921),.A(g8958));
  NOT NOT1_4234(.VSS(VSS),.VDD(VDD),.Y(g12922),.A(g8961));
  NOT NOT1_4235(.VSS(VSS),.VDD(VDD),.Y(g12931),.A(g8965));
  NOT NOT1_4236(.VSS(VSS),.VDD(VDD),.Y(g12932),.A(g8968));
  NOT NOT1_4237(.VSS(VSS),.VDD(VDD),.Y(g12934),.A(g8974));
  NOT NOT1_4238(.VSS(VSS),.VDD(VDD),.Y(I19986),.A(g8577));
  NOT NOT1_4239(.VSS(VSS),.VDD(VDD),.Y(g12935),.A(I19986));
  NOT NOT1_4240(.VSS(VSS),.VDD(VDD),.Y(g12940),.A(g8980));
  NOT NOT1_4241(.VSS(VSS),.VDD(VDD),.Y(g12943),.A(g8984));
  NOT NOT1_4242(.VSS(VSS),.VDD(VDD),.Y(g12944),.A(g8987));
  NOT NOT1_4243(.VSS(VSS),.VDD(VDD),.Y(g12950),.A(g8990));
  NOT NOT1_4244(.VSS(VSS),.VDD(VDD),.Y(g12951),.A(g8993));
  NOT NOT1_4245(.VSS(VSS),.VDD(VDD),.Y(g12960),.A(g8997));
  NOT NOT1_4246(.VSS(VSS),.VDD(VDD),.Y(g12961),.A(g9000));
  NOT NOT1_4247(.VSS(VSS),.VDD(VDD),.Y(I20009),.A(g8313));
  NOT NOT1_4248(.VSS(VSS),.VDD(VDD),.Y(g12962),.A(I20009));
  NOT NOT1_4249(.VSS(VSS),.VDD(VDD),.Y(g12965),.A(g9006));
  NOT NOT1_4250(.VSS(VSS),.VDD(VDD),.Y(g12969),.A(g9010));
  NOT NOT1_4251(.VSS(VSS),.VDD(VDD),.Y(g12972),.A(g9013));
  NOT NOT1_4252(.VSS(VSS),.VDD(VDD),.Y(g12973),.A(g9016));
  NOT NOT1_4253(.VSS(VSS),.VDD(VDD),.Y(g12979),.A(g9019));
  NOT NOT1_4254(.VSS(VSS),.VDD(VDD),.Y(g12980),.A(g9022));
  NOT NOT1_4255(.VSS(VSS),.VDD(VDD),.Y(g12993),.A(g9035));
  NOT NOT1_4256(.VSS(VSS),.VDD(VDD),.Y(g12996),.A(g9038));
  NOT NOT1_4257(.VSS(VSS),.VDD(VDD),.Y(g12997),.A(g9041));
  NOT NOT1_4258(.VSS(VSS),.VDD(VDD),.Y(g12998),.A(g9044));
  NOT NOT1_4259(.VSS(VSS),.VDD(VDD),.Y(g13003),.A(g9058));
  NOT NOT1_4260(.VSS(VSS),.VDD(VDD),.Y(I20062),.A(g10480));
  NOT NOT1_4261(.VSS(VSS),.VDD(VDD),.Y(g13011),.A(I20062));
  NOT NOT1_4262(.VSS(VSS),.VDD(VDD),.Y(g13025),.A(g10810));
  NOT NOT1_4263(.VSS(VSS),.VDD(VDD),.Y(g13033),.A(g10797));
  NOT NOT1_4264(.VSS(VSS),.VDD(VDD),.Y(g13036),.A(g10831));
  NOT NOT1_4265(.VSS(VSS),.VDD(VDD),.Y(g13043),.A(g10789));
  NOT NOT1_4266(.VSS(VSS),.VDD(VDD),.Y(g13046),.A(g10814));
  NOT NOT1_4267(.VSS(VSS),.VDD(VDD),.Y(g13049),.A(g10851));
  NOT NOT1_4268(.VSS(VSS),.VDD(VDD),.Y(g13057),.A(g10784));
  NOT NOT1_4269(.VSS(VSS),.VDD(VDD),.Y(g13060),.A(g10801));
  NOT NOT1_4270(.VSS(VSS),.VDD(VDD),.Y(g13063),.A(g10835));
  NOT NOT1_4271(.VSS(VSS),.VDD(VDD),.Y(g13066),.A(g10872));
  NOT NOT1_4272(.VSS(VSS),.VDD(VDD),.Y(I20117),.A(g10876));
  NOT NOT1_4273(.VSS(VSS),.VDD(VDD),.Y(g13070),.A(I20117));
  NOT NOT1_4274(.VSS(VSS),.VDD(VDD),.Y(g13073),.A(g10793));
  NOT NOT1_4275(.VSS(VSS),.VDD(VDD),.Y(g13076),.A(g10818));
  NOT NOT1_4276(.VSS(VSS),.VDD(VDD),.Y(g13079),.A(g10855));
  NOT NOT1_4277(.VSS(VSS),.VDD(VDD),.Y(g13092),.A(g10805));
  NOT NOT1_4278(.VSS(VSS),.VDD(VDD),.Y(g13095),.A(g10839));
  NOT NOT1_4279(.VSS(VSS),.VDD(VDD),.Y(g13101),.A(g9128));
  NOT NOT1_4280(.VSS(VSS),.VDD(VDD),.Y(g13107),.A(g10822));
  NOT NOT1_4281(.VSS(VSS),.VDD(VDD),.Y(g13117),.A(g9134));
  NOT NOT1_4282(.VSS(VSS),.VDD(VDD),.Y(g13130),.A(g9140));
  NOT NOT1_4283(.VSS(VSS),.VDD(VDD),.Y(g13141),.A(g9146));
  NOT NOT1_4284(.VSS(VSS),.VDD(VDD),.Y(g13148),.A(g9170));
  NOT NOT1_4285(.VSS(VSS),.VDD(VDD),.Y(g13151),.A(g9184));
  NOT NOT1_4286(.VSS(VSS),.VDD(VDD),.Y(g13152),.A(g9196));
  NOT NOT1_4287(.VSS(VSS),.VDD(VDD),.Y(g13153),.A(g9199));
  NOT NOT1_4288(.VSS(VSS),.VDD(VDD),.Y(g13154),.A(g9212));
  NOT NOT1_4289(.VSS(VSS),.VDD(VDD),.Y(g13157),.A(g9229));
  NOT NOT1_4290(.VSS(VSS),.VDD(VDD),.Y(g13158),.A(g9242));
  NOT NOT1_4291(.VSS(VSS),.VDD(VDD),.Y(g13159),.A(g9245));
  NOT NOT1_4292(.VSS(VSS),.VDD(VDD),.Y(g13161),.A(g9257));
  NOT NOT1_4293(.VSS(VSS),.VDD(VDD),.Y(g13162),.A(g9260));
  NOT NOT1_4294(.VSS(VSS),.VDD(VDD),.Y(g13163),.A(g9273));
  NOT NOT1_4295(.VSS(VSS),.VDD(VDD),.Y(g13166),.A(g9290));
  NOT NOT1_4296(.VSS(VSS),.VDD(VDD),.Y(g13167),.A(g9303));
  NOT NOT1_4297(.VSS(VSS),.VDD(VDD),.Y(g13168),.A(g9306));
  NOT NOT1_4298(.VSS(VSS),.VDD(VDD),.Y(g13169),.A(g9320));
  NOT NOT1_4299(.VSS(VSS),.VDD(VDD),.Y(g13170),.A(g9323));
  NOT NOT1_4300(.VSS(VSS),.VDD(VDD),.Y(g13172),.A(g9335));
  NOT NOT1_4301(.VSS(VSS),.VDD(VDD),.Y(g13173),.A(g9338));
  NOT NOT1_4302(.VSS(VSS),.VDD(VDD),.Y(g13174),.A(g9351));
  NOT NOT1_4303(.VSS(VSS),.VDD(VDD),.Y(g13176),.A(g9368));
  NOT NOT1_4304(.VSS(VSS),.VDD(VDD),.Y(g13177),.A(g9371));
  NOT NOT1_4305(.VSS(VSS),.VDD(VDD),.Y(g13178),.A(g9384));
  NOT NOT1_4306(.VSS(VSS),.VDD(VDD),.Y(g13179),.A(g9387));
  NOT NOT1_4307(.VSS(VSS),.VDD(VDD),.Y(g13180),.A(g9401));
  NOT NOT1_4308(.VSS(VSS),.VDD(VDD),.Y(g13181),.A(g9404));
  NOT NOT1_4309(.VSS(VSS),.VDD(VDD),.Y(g13183),.A(g9416));
  NOT NOT1_4310(.VSS(VSS),.VDD(VDD),.Y(g13184),.A(g9419));
  NOT NOT1_4311(.VSS(VSS),.VDD(VDD),.Y(g13185),.A(g9443));
  NOT NOT1_4312(.VSS(VSS),.VDD(VDD),.Y(g13186),.A(g9446));
  NOT NOT1_4313(.VSS(VSS),.VDD(VDD),.Y(g13187),.A(g9450));
  NOT NOT1_4314(.VSS(VSS),.VDD(VDD),.Y(g13188),.A(g9465));
  NOT NOT1_4315(.VSS(VSS),.VDD(VDD),.Y(g13189),.A(g9468));
  NOT NOT1_4316(.VSS(VSS),.VDD(VDD),.Y(g13190),.A(g9481));
  NOT NOT1_4317(.VSS(VSS),.VDD(VDD),.Y(g13191),.A(g9484));
  NOT NOT1_4318(.VSS(VSS),.VDD(VDD),.Y(g13192),.A(g9498));
  NOT NOT1_4319(.VSS(VSS),.VDD(VDD),.Y(g13193),.A(g9501));
  NOT NOT1_4320(.VSS(VSS),.VDD(VDD),.Y(g13195),.A(g9524));
  NOT NOT1_4321(.VSS(VSS),.VDD(VDD),.Y(g13196),.A(g9528));
  NOT NOT1_4322(.VSS(VSS),.VDD(VDD),.Y(g13197),.A(g9531));
  NOT NOT1_4323(.VSS(VSS),.VDD(VDD),.Y(g13198),.A(g9585));
  NOT NOT1_4324(.VSS(VSS),.VDD(VDD),.Y(g13199),.A(g9588));
  NOT NOT1_4325(.VSS(VSS),.VDD(VDD),.Y(g13200),.A(g9592));
  NOT NOT1_4326(.VSS(VSS),.VDD(VDD),.Y(g13201),.A(g9607));
  NOT NOT1_4327(.VSS(VSS),.VDD(VDD),.Y(g13202),.A(g9610));
  NOT NOT1_4328(.VSS(VSS),.VDD(VDD),.Y(g13203),.A(g9623));
  NOT NOT1_4329(.VSS(VSS),.VDD(VDD),.Y(g13204),.A(g9626));
  NOT NOT1_4330(.VSS(VSS),.VDD(VDD),.Y(g13205),.A(g9641));
  NOT NOT1_4331(.VSS(VSS),.VDD(VDD),.Y(g13206),.A(g9644));
  NOT NOT1_4332(.VSS(VSS),.VDD(VDD),.Y(g13207),.A(g9666));
  NOT NOT1_4333(.VSS(VSS),.VDD(VDD),.Y(g13208),.A(g9670));
  NOT NOT1_4334(.VSS(VSS),.VDD(VDD),.Y(g13209),.A(g9673));
  NOT NOT1_4335(.VSS(VSS),.VDD(VDD),.Y(g13210),.A(g9727));
  NOT NOT1_4336(.VSS(VSS),.VDD(VDD),.Y(g13211),.A(g9730));
  NOT NOT1_4337(.VSS(VSS),.VDD(VDD),.Y(g13212),.A(g9734));
  NOT NOT1_4338(.VSS(VSS),.VDD(VDD),.Y(g13213),.A(g9749));
  NOT NOT1_4339(.VSS(VSS),.VDD(VDD),.Y(g13214),.A(g9752));
  NOT NOT1_4340(.VSS(VSS),.VDD(VDD),.Y(I20264),.A(g9027));
  NOT NOT1_4341(.VSS(VSS),.VDD(VDD),.Y(g13215),.A(I20264));
  NOT NOT1_4342(.VSS(VSS),.VDD(VDD),.Y(g13218),.A(g9767));
  NOT NOT1_4343(.VSS(VSS),.VDD(VDD),.Y(g13219),.A(g9770));
  NOT NOT1_4344(.VSS(VSS),.VDD(VDD),.Y(g13220),.A(g9787));
  NOT NOT1_4345(.VSS(VSS),.VDD(VDD),.Y(g13221),.A(g9790));
  NOT NOT1_4346(.VSS(VSS),.VDD(VDD),.Y(g13222),.A(g9812));
  NOT NOT1_4347(.VSS(VSS),.VDD(VDD),.Y(g13223),.A(g9816));
  NOT NOT1_4348(.VSS(VSS),.VDD(VDD),.Y(g13224),.A(g9819));
  NOT NOT1_4349(.VSS(VSS),.VDD(VDD),.Y(g13225),.A(g9873));
  NOT NOT1_4350(.VSS(VSS),.VDD(VDD),.Y(g13226),.A(g9876));
  NOT NOT1_4351(.VSS(VSS),.VDD(VDD),.Y(g13227),.A(g9880));
  NOT NOT1_4352(.VSS(VSS),.VDD(VDD),.Y(I20278),.A(g9027));
  NOT NOT1_4353(.VSS(VSS),.VDD(VDD),.Y(g13229),.A(I20278));
  NOT NOT1_4354(.VSS(VSS),.VDD(VDD),.Y(g13232),.A(g9895));
  NOT NOT1_4355(.VSS(VSS),.VDD(VDD),.Y(g13233),.A(g9898));
  NOT NOT1_4356(.VSS(VSS),.VDD(VDD),.Y(I20283),.A(g9050));
  NOT NOT1_4357(.VSS(VSS),.VDD(VDD),.Y(g13234),.A(I20283));
  NOT NOT1_4358(.VSS(VSS),.VDD(VDD),.Y(g13237),.A(g9913));
  NOT NOT1_4359(.VSS(VSS),.VDD(VDD),.Y(g13238),.A(g9916));
  NOT NOT1_4360(.VSS(VSS),.VDD(VDD),.Y(g13239),.A(g9933));
  NOT NOT1_4361(.VSS(VSS),.VDD(VDD),.Y(g13240),.A(g9936));
  NOT NOT1_4362(.VSS(VSS),.VDD(VDD),.Y(g13241),.A(g9958));
  NOT NOT1_4363(.VSS(VSS),.VDD(VDD),.Y(g13242),.A(g9962));
  NOT NOT1_4364(.VSS(VSS),.VDD(VDD),.Y(g13243),.A(g9965));
  NOT NOT1_4365(.VSS(VSS),.VDD(VDD),.Y(g13244),.A(g10004));
  NOT NOT1_4366(.VSS(VSS),.VDD(VDD),.Y(I20295),.A(g10015));
  NOT NOT1_4367(.VSS(VSS),.VDD(VDD),.Y(g13246),.A(I20295));
  NOT NOT1_4368(.VSS(VSS),.VDD(VDD),.Y(I20299),.A(g10800));
  NOT NOT1_4369(.VSS(VSS),.VDD(VDD),.Y(g13248),.A(I20299));
  NOT NOT1_4370(.VSS(VSS),.VDD(VDD),.Y(g13249),.A(g10018));
  NOT NOT1_4371(.VSS(VSS),.VDD(VDD),.Y(g13250),.A(g10021));
  NOT NOT1_4372(.VSS(VSS),.VDD(VDD),.Y(I20305),.A(g9050));
  NOT NOT1_4373(.VSS(VSS),.VDD(VDD),.Y(g13252),.A(I20305));
  NOT NOT1_4374(.VSS(VSS),.VDD(VDD),.Y(g13255),.A(g10049));
  NOT NOT1_4375(.VSS(VSS),.VDD(VDD),.Y(g13256),.A(g10052));
  NOT NOT1_4376(.VSS(VSS),.VDD(VDD),.Y(I20310),.A(g9067));
  NOT NOT1_4377(.VSS(VSS),.VDD(VDD),.Y(g13257),.A(I20310));
  NOT NOT1_4378(.VSS(VSS),.VDD(VDD),.Y(g13260),.A(g10067));
  NOT NOT1_4379(.VSS(VSS),.VDD(VDD),.Y(g13261),.A(g10070));
  NOT NOT1_4380(.VSS(VSS),.VDD(VDD),.Y(g13262),.A(g10087));
  NOT NOT1_4381(.VSS(VSS),.VDD(VDD),.Y(g13263),.A(g10090));
  NOT NOT1_4382(.VSS(VSS),.VDD(VDD),.Y(g13264),.A(g10096));
  NOT NOT1_4383(.VSS(VSS),.VDD(VDD),.Y(g13265),.A(g8568));
  NOT NOT1_4384(.VSS(VSS),.VDD(VDD),.Y(I20320),.A(g10792));
  NOT NOT1_4385(.VSS(VSS),.VDD(VDD),.Y(g13267),.A(I20320));
  NOT NOT1_4386(.VSS(VSS),.VDD(VDD),.Y(g13268),.A(g10109));
  NOT NOT1_4387(.VSS(VSS),.VDD(VDD),.Y(I20324),.A(g10124));
  NOT NOT1_4388(.VSS(VSS),.VDD(VDD),.Y(g13269),.A(I20324));
  NOT NOT1_4389(.VSS(VSS),.VDD(VDD),.Y(I20328),.A(g10817));
  NOT NOT1_4390(.VSS(VSS),.VDD(VDD),.Y(g13271),.A(I20328));
  NOT NOT1_4391(.VSS(VSS),.VDD(VDD),.Y(g13272),.A(g10127));
  NOT NOT1_4392(.VSS(VSS),.VDD(VDD),.Y(g13273),.A(g10130));
  NOT NOT1_4393(.VSS(VSS),.VDD(VDD),.Y(I20334),.A(g9067));
  NOT NOT1_4394(.VSS(VSS),.VDD(VDD),.Y(g13275),.A(I20334));
  NOT NOT1_4395(.VSS(VSS),.VDD(VDD),.Y(g13278),.A(g10158));
  NOT NOT1_4396(.VSS(VSS),.VDD(VDD),.Y(g13279),.A(g10161));
  NOT NOT1_4397(.VSS(VSS),.VDD(VDD),.Y(I20339),.A(g9084));
  NOT NOT1_4398(.VSS(VSS),.VDD(VDD),.Y(g13280),.A(I20339));
  NOT NOT1_4399(.VSS(VSS),.VDD(VDD),.Y(g13283),.A(g10176));
  NOT NOT1_4400(.VSS(VSS),.VDD(VDD),.Y(g13284),.A(g10179));
  NOT NOT1_4401(.VSS(VSS),.VDD(VDD),.Y(g13285),.A(g10189));
  NOT NOT1_4402(.VSS(VSS),.VDD(VDD),.Y(I20347),.A(g10787));
  NOT NOT1_4403(.VSS(VSS),.VDD(VDD),.Y(g13290),.A(I20347));
  NOT NOT1_4404(.VSS(VSS),.VDD(VDD),.Y(I20351),.A(g10804));
  NOT NOT1_4405(.VSS(VSS),.VDD(VDD),.Y(g13292),.A(I20351));
  NOT NOT1_4406(.VSS(VSS),.VDD(VDD),.Y(g13293),.A(g10214));
  NOT NOT1_4407(.VSS(VSS),.VDD(VDD),.Y(I20355),.A(g10229));
  NOT NOT1_4408(.VSS(VSS),.VDD(VDD),.Y(g13294),.A(I20355));
  NOT NOT1_4409(.VSS(VSS),.VDD(VDD),.Y(I20359),.A(g10838));
  NOT NOT1_4410(.VSS(VSS),.VDD(VDD),.Y(g13296),.A(I20359));
  NOT NOT1_4411(.VSS(VSS),.VDD(VDD),.Y(g13297),.A(g10232));
  NOT NOT1_4412(.VSS(VSS),.VDD(VDD),.Y(g13298),.A(g10235));
  NOT NOT1_4413(.VSS(VSS),.VDD(VDD),.Y(I20365),.A(g9084));
  NOT NOT1_4414(.VSS(VSS),.VDD(VDD),.Y(g13300),.A(I20365));
  NOT NOT1_4415(.VSS(VSS),.VDD(VDD),.Y(g13303),.A(g10263));
  NOT NOT1_4416(.VSS(VSS),.VDD(VDD),.Y(g13304),.A(g10266));
  NOT NOT1_4417(.VSS(VSS),.VDD(VDD),.Y(g13308),.A(g10273));
  NOT NOT1_4418(.VSS(VSS),.VDD(VDD),.Y(g13309),.A(g10276));
  NOT NOT1_4419(.VSS(VSS),.VDD(VDD),.Y(I20376),.A(g8569));
  NOT NOT1_4420(.VSS(VSS),.VDD(VDD),.Y(g13317),.A(I20376));
  NOT NOT1_4421(.VSS(VSS),.VDD(VDD),.Y(I20379),.A(g11213));
  NOT NOT1_4422(.VSS(VSS),.VDD(VDD),.Y(g13318),.A(I20379));
  NOT NOT1_4423(.VSS(VSS),.VDD(VDD),.Y(I20382),.A(g10907));
  NOT NOT1_4424(.VSS(VSS),.VDD(VDD),.Y(g13319),.A(I20382));
  NOT NOT1_4425(.VSS(VSS),.VDD(VDD),.Y(I20386),.A(g10796));
  NOT NOT1_4426(.VSS(VSS),.VDD(VDD),.Y(g13321),.A(I20386));
  NOT NOT1_4427(.VSS(VSS),.VDD(VDD),.Y(I20390),.A(g10821));
  NOT NOT1_4428(.VSS(VSS),.VDD(VDD),.Y(g13323),.A(I20390));
  NOT NOT1_4429(.VSS(VSS),.VDD(VDD),.Y(g13324),.A(g10316));
  NOT NOT1_4430(.VSS(VSS),.VDD(VDD),.Y(I20394),.A(g10331));
  NOT NOT1_4431(.VSS(VSS),.VDD(VDD),.Y(g13325),.A(I20394));
  NOT NOT1_4432(.VSS(VSS),.VDD(VDD),.Y(I20398),.A(g10858));
  NOT NOT1_4433(.VSS(VSS),.VDD(VDD),.Y(g13327),.A(I20398));
  NOT NOT1_4434(.VSS(VSS),.VDD(VDD),.Y(g13328),.A(g10334));
  NOT NOT1_4435(.VSS(VSS),.VDD(VDD),.Y(g13329),.A(g10337));
  NOT NOT1_4436(.VSS(VSS),.VDD(VDD),.Y(g13330),.A(g10357));
  NOT NOT1_4437(.VSS(VSS),.VDD(VDD),.Y(I20407),.A(g9027));
  NOT NOT1_4438(.VSS(VSS),.VDD(VDD),.Y(g13336),.A(I20407));
  NOT NOT1_4439(.VSS(VSS),.VDD(VDD),.Y(I20410),.A(g10887));
  NOT NOT1_4440(.VSS(VSS),.VDD(VDD),.Y(g13339),.A(I20410));
  NOT NOT1_4441(.VSS(VSS),.VDD(VDD),.Y(I20414),.A(g8575));
  NOT NOT1_4442(.VSS(VSS),.VDD(VDD),.Y(g13341),.A(I20414));
  NOT NOT1_4443(.VSS(VSS),.VDD(VDD),.Y(I20417),.A(g10933));
  NOT NOT1_4444(.VSS(VSS),.VDD(VDD),.Y(g13342),.A(I20417));
  NOT NOT1_4445(.VSS(VSS),.VDD(VDD),.Y(I20421),.A(g10808));
  NOT NOT1_4446(.VSS(VSS),.VDD(VDD),.Y(g13344),.A(I20421));
  NOT NOT1_4447(.VSS(VSS),.VDD(VDD),.Y(I20425),.A(g10842));
  NOT NOT1_4448(.VSS(VSS),.VDD(VDD),.Y(g13346),.A(I20425));
  NOT NOT1_4449(.VSS(VSS),.VDD(VDD),.Y(g13347),.A(g10409));
  NOT NOT1_4450(.VSS(VSS),.VDD(VDD),.Y(g13351),.A(g10416));
  NOT NOT1_4451(.VSS(VSS),.VDD(VDD),.Y(g13352),.A(g10419));
  NOT NOT1_4452(.VSS(VSS),.VDD(VDD),.Y(I20441),.A(g9027));
  NOT NOT1_4453(.VSS(VSS),.VDD(VDD),.Y(g13356),.A(I20441));
  NOT NOT1_4454(.VSS(VSS),.VDD(VDD),.Y(I20444),.A(g10869));
  NOT NOT1_4455(.VSS(VSS),.VDD(VDD),.Y(g13359),.A(I20444));
  NOT NOT1_4456(.VSS(VSS),.VDD(VDD),.Y(I20448),.A(g9050));
  NOT NOT1_4457(.VSS(VSS),.VDD(VDD),.Y(g13361),.A(I20448));
  NOT NOT1_4458(.VSS(VSS),.VDD(VDD),.Y(I20451),.A(g10908));
  NOT NOT1_4459(.VSS(VSS),.VDD(VDD),.Y(g13364),.A(I20451));
  NOT NOT1_4460(.VSS(VSS),.VDD(VDD),.Y(I20455),.A(g8578));
  NOT NOT1_4461(.VSS(VSS),.VDD(VDD),.Y(g13366),.A(I20455));
  NOT NOT1_4462(.VSS(VSS),.VDD(VDD),.Y(I20458),.A(g10972));
  NOT NOT1_4463(.VSS(VSS),.VDD(VDD),.Y(g13367),.A(I20458));
  NOT NOT1_4464(.VSS(VSS),.VDD(VDD),.Y(I20462),.A(g10825));
  NOT NOT1_4465(.VSS(VSS),.VDD(VDD),.Y(g13369),.A(I20462));
  NOT NOT1_4466(.VSS(VSS),.VDD(VDD),.Y(g13373),.A(g10482));
  NOT NOT1_4467(.VSS(VSS),.VDD(VDD),.Y(I20476),.A(g9027));
  NOT NOT1_4468(.VSS(VSS),.VDD(VDD),.Y(g13381),.A(I20476));
  NOT NOT1_4469(.VSS(VSS),.VDD(VDD),.Y(I20479),.A(g10849));
  NOT NOT1_4470(.VSS(VSS),.VDD(VDD),.Y(g13384),.A(I20479));
  NOT NOT1_4471(.VSS(VSS),.VDD(VDD),.Y(I20483),.A(g9050));
  NOT NOT1_4472(.VSS(VSS),.VDD(VDD),.Y(g13386),.A(I20483));
  NOT NOT1_4473(.VSS(VSS),.VDD(VDD),.Y(I20486),.A(g10889));
  NOT NOT1_4474(.VSS(VSS),.VDD(VDD),.Y(g13389),.A(I20486));
  NOT NOT1_4475(.VSS(VSS),.VDD(VDD),.Y(I20490),.A(g9067));
  NOT NOT1_4476(.VSS(VSS),.VDD(VDD),.Y(g13391),.A(I20490));
  NOT NOT1_4477(.VSS(VSS),.VDD(VDD),.Y(I20493),.A(g10934));
  NOT NOT1_4478(.VSS(VSS),.VDD(VDD),.Y(g13394),.A(I20493));
  NOT NOT1_4479(.VSS(VSS),.VDD(VDD),.Y(I20497),.A(g8579));
  NOT NOT1_4480(.VSS(VSS),.VDD(VDD),.Y(g13396),.A(I20497));
  NOT NOT1_4481(.VSS(VSS),.VDD(VDD),.Y(I20500),.A(g11007));
  NOT NOT1_4482(.VSS(VSS),.VDD(VDD),.Y(g13397),.A(I20500));
  NOT NOT1_4483(.VSS(VSS),.VDD(VDD),.Y(g13398),.A(g10542));
  NOT NOT1_4484(.VSS(VSS),.VDD(VDD),.Y(g13400),.A(g10545));
  NOT NOT1_4485(.VSS(VSS),.VDD(VDD),.Y(I20514),.A(g11769));
  NOT NOT1_4486(.VSS(VSS),.VDD(VDD),.Y(g13405),.A(I20514));
  NOT NOT1_4487(.VSS(VSS),.VDD(VDD),.Y(I20517),.A(g12425));
  NOT NOT1_4488(.VSS(VSS),.VDD(VDD),.Y(g13406),.A(I20517));
  NOT NOT1_4489(.VSS(VSS),.VDD(VDD),.Y(I20520),.A(g13246));
  NOT NOT1_4490(.VSS(VSS),.VDD(VDD),.Y(g13407),.A(I20520));
  NOT NOT1_4491(.VSS(VSS),.VDD(VDD),.Y(I20523),.A(g13317));
  NOT NOT1_4492(.VSS(VSS),.VDD(VDD),.Y(g13408),.A(I20523));
  NOT NOT1_4493(.VSS(VSS),.VDD(VDD),.Y(I20526),.A(g12519));
  NOT NOT1_4494(.VSS(VSS),.VDD(VDD),.Y(g13409),.A(I20526));
  NOT NOT1_4495(.VSS(VSS),.VDD(VDD),.Y(I20529),.A(g13319));
  NOT NOT1_4496(.VSS(VSS),.VDD(VDD),.Y(g13410),.A(I20529));
  NOT NOT1_4497(.VSS(VSS),.VDD(VDD),.Y(I20532),.A(g13339));
  NOT NOT1_4498(.VSS(VSS),.VDD(VDD),.Y(g13411),.A(I20532));
  NOT NOT1_4499(.VSS(VSS),.VDD(VDD),.Y(I20535),.A(g13359));
  NOT NOT1_4500(.VSS(VSS),.VDD(VDD),.Y(g13412),.A(I20535));
  NOT NOT1_4501(.VSS(VSS),.VDD(VDD),.Y(I20538),.A(g13384));
  NOT NOT1_4502(.VSS(VSS),.VDD(VDD),.Y(g13413),.A(I20538));
  NOT NOT1_4503(.VSS(VSS),.VDD(VDD),.Y(I20541),.A(g11599));
  NOT NOT1_4504(.VSS(VSS),.VDD(VDD),.Y(g13414),.A(I20541));
  NOT NOT1_4505(.VSS(VSS),.VDD(VDD),.Y(I20544),.A(g11628));
  NOT NOT1_4506(.VSS(VSS),.VDD(VDD),.Y(g13415),.A(I20544));
  NOT NOT1_4507(.VSS(VSS),.VDD(VDD),.Y(I20547),.A(g13248));
  NOT NOT1_4508(.VSS(VSS),.VDD(VDD),.Y(g13416),.A(I20547));
  NOT NOT1_4509(.VSS(VSS),.VDD(VDD),.Y(I20550),.A(g13267));
  NOT NOT1_4510(.VSS(VSS),.VDD(VDD),.Y(g13417),.A(I20550));
  NOT NOT1_4511(.VSS(VSS),.VDD(VDD),.Y(I20553),.A(g13290));
  NOT NOT1_4512(.VSS(VSS),.VDD(VDD),.Y(g13418),.A(I20553));
  NOT NOT1_4513(.VSS(VSS),.VDD(VDD),.Y(I20556),.A(g12435));
  NOT NOT1_4514(.VSS(VSS),.VDD(VDD),.Y(g13419),.A(I20556));
  NOT NOT1_4515(.VSS(VSS),.VDD(VDD),.Y(I20559),.A(g11937));
  NOT NOT1_4516(.VSS(VSS),.VDD(VDD),.Y(g13420),.A(I20559));
  NOT NOT1_4517(.VSS(VSS),.VDD(VDD),.Y(I20562),.A(g11786));
  NOT NOT1_4518(.VSS(VSS),.VDD(VDD),.Y(g13421),.A(I20562));
  NOT NOT1_4519(.VSS(VSS),.VDD(VDD),.Y(I20565),.A(g12432));
  NOT NOT1_4520(.VSS(VSS),.VDD(VDD),.Y(g13422),.A(I20565));
  NOT NOT1_4521(.VSS(VSS),.VDD(VDD),.Y(I20568),.A(g13269));
  NOT NOT1_4522(.VSS(VSS),.VDD(VDD),.Y(g13423),.A(I20568));
  NOT NOT1_4523(.VSS(VSS),.VDD(VDD),.Y(I20571),.A(g13341));
  NOT NOT1_4524(.VSS(VSS),.VDD(VDD),.Y(g13424),.A(I20571));
  NOT NOT1_4525(.VSS(VSS),.VDD(VDD),.Y(I20574),.A(g12534));
  NOT NOT1_4526(.VSS(VSS),.VDD(VDD),.Y(g13425),.A(I20574));
  NOT NOT1_4527(.VSS(VSS),.VDD(VDD),.Y(I20577),.A(g13342));
  NOT NOT1_4528(.VSS(VSS),.VDD(VDD),.Y(g13426),.A(I20577));
  NOT NOT1_4529(.VSS(VSS),.VDD(VDD),.Y(I20580),.A(g13364));
  NOT NOT1_4530(.VSS(VSS),.VDD(VDD),.Y(g13427),.A(I20580));
  NOT NOT1_4531(.VSS(VSS),.VDD(VDD),.Y(I20583),.A(g13389));
  NOT NOT1_4532(.VSS(VSS),.VDD(VDD),.Y(g13428),.A(I20583));
  NOT NOT1_4533(.VSS(VSS),.VDD(VDD),.Y(I20586),.A(g11606));
  NOT NOT1_4534(.VSS(VSS),.VDD(VDD),.Y(g13429),.A(I20586));
  NOT NOT1_4535(.VSS(VSS),.VDD(VDD),.Y(I20589),.A(g11629));
  NOT NOT1_4536(.VSS(VSS),.VDD(VDD),.Y(g13430),.A(I20589));
  NOT NOT1_4537(.VSS(VSS),.VDD(VDD),.Y(I20592),.A(g11651));
  NOT NOT1_4538(.VSS(VSS),.VDD(VDD),.Y(g13431),.A(I20592));
  NOT NOT1_4539(.VSS(VSS),.VDD(VDD),.Y(I20595),.A(g13271));
  NOT NOT1_4540(.VSS(VSS),.VDD(VDD),.Y(g13432),.A(I20595));
  NOT NOT1_4541(.VSS(VSS),.VDD(VDD),.Y(I20598),.A(g13292));
  NOT NOT1_4542(.VSS(VSS),.VDD(VDD),.Y(g13433),.A(I20598));
  NOT NOT1_4543(.VSS(VSS),.VDD(VDD),.Y(I20601),.A(g13321));
  NOT NOT1_4544(.VSS(VSS),.VDD(VDD),.Y(g13434),.A(I20601));
  NOT NOT1_4545(.VSS(VSS),.VDD(VDD),.Y(I20604),.A(g12440));
  NOT NOT1_4546(.VSS(VSS),.VDD(VDD),.Y(g13435),.A(I20604));
  NOT NOT1_4547(.VSS(VSS),.VDD(VDD),.Y(I20607),.A(g11990));
  NOT NOT1_4548(.VSS(VSS),.VDD(VDD),.Y(g13436),.A(I20607));
  NOT NOT1_4549(.VSS(VSS),.VDD(VDD),.Y(I20610),.A(g11812));
  NOT NOT1_4550(.VSS(VSS),.VDD(VDD),.Y(g13437),.A(I20610));
  NOT NOT1_4551(.VSS(VSS),.VDD(VDD),.Y(I20613),.A(g12437));
  NOT NOT1_4552(.VSS(VSS),.VDD(VDD),.Y(g13438),.A(I20613));
  NOT NOT1_4553(.VSS(VSS),.VDD(VDD),.Y(I20616),.A(g13294));
  NOT NOT1_4554(.VSS(VSS),.VDD(VDD),.Y(g13439),.A(I20616));
  NOT NOT1_4555(.VSS(VSS),.VDD(VDD),.Y(I20619),.A(g13366));
  NOT NOT1_4556(.VSS(VSS),.VDD(VDD),.Y(g13440),.A(I20619));
  NOT NOT1_4557(.VSS(VSS),.VDD(VDD),.Y(I20622),.A(g12543));
  NOT NOT1_4558(.VSS(VSS),.VDD(VDD),.Y(g13441),.A(I20622));
  NOT NOT1_4559(.VSS(VSS),.VDD(VDD),.Y(I20625),.A(g13367));
  NOT NOT1_4560(.VSS(VSS),.VDD(VDD),.Y(g13442),.A(I20625));
  NOT NOT1_4561(.VSS(VSS),.VDD(VDD),.Y(I20628),.A(g13394));
  NOT NOT1_4562(.VSS(VSS),.VDD(VDD),.Y(g13443),.A(I20628));
  NOT NOT1_4563(.VSS(VSS),.VDD(VDD),.Y(I20631),.A(g11611));
  NOT NOT1_4564(.VSS(VSS),.VDD(VDD),.Y(g13444),.A(I20631));
  NOT NOT1_4565(.VSS(VSS),.VDD(VDD),.Y(I20634),.A(g11636));
  NOT NOT1_4566(.VSS(VSS),.VDD(VDD),.Y(g13445),.A(I20634));
  NOT NOT1_4567(.VSS(VSS),.VDD(VDD),.Y(I20637),.A(g11652));
  NOT NOT1_4568(.VSS(VSS),.VDD(VDD),.Y(g13446),.A(I20637));
  NOT NOT1_4569(.VSS(VSS),.VDD(VDD),.Y(I20640),.A(g11670));
  NOT NOT1_4570(.VSS(VSS),.VDD(VDD),.Y(g13447),.A(I20640));
  NOT NOT1_4571(.VSS(VSS),.VDD(VDD),.Y(I20643),.A(g13296));
  NOT NOT1_4572(.VSS(VSS),.VDD(VDD),.Y(g13448),.A(I20643));
  NOT NOT1_4573(.VSS(VSS),.VDD(VDD),.Y(I20646),.A(g13323));
  NOT NOT1_4574(.VSS(VSS),.VDD(VDD),.Y(g13449),.A(I20646));
  NOT NOT1_4575(.VSS(VSS),.VDD(VDD),.Y(I20649),.A(g13344));
  NOT NOT1_4576(.VSS(VSS),.VDD(VDD),.Y(g13450),.A(I20649));
  NOT NOT1_4577(.VSS(VSS),.VDD(VDD),.Y(I20652),.A(g12445));
  NOT NOT1_4578(.VSS(VSS),.VDD(VDD),.Y(g13451),.A(I20652));
  NOT NOT1_4579(.VSS(VSS),.VDD(VDD),.Y(I20655),.A(g12059));
  NOT NOT1_4580(.VSS(VSS),.VDD(VDD),.Y(g13452),.A(I20655));
  NOT NOT1_4581(.VSS(VSS),.VDD(VDD),.Y(I20658),.A(g11845));
  NOT NOT1_4582(.VSS(VSS),.VDD(VDD),.Y(g13453),.A(I20658));
  NOT NOT1_4583(.VSS(VSS),.VDD(VDD),.Y(I20661),.A(g12442));
  NOT NOT1_4584(.VSS(VSS),.VDD(VDD),.Y(g13454),.A(I20661));
  NOT NOT1_4585(.VSS(VSS),.VDD(VDD),.Y(I20664),.A(g13325));
  NOT NOT1_4586(.VSS(VSS),.VDD(VDD),.Y(g13455),.A(I20664));
  NOT NOT1_4587(.VSS(VSS),.VDD(VDD),.Y(I20667),.A(g13396));
  NOT NOT1_4588(.VSS(VSS),.VDD(VDD),.Y(g13456),.A(I20667));
  NOT NOT1_4589(.VSS(VSS),.VDD(VDD),.Y(I20670),.A(g12552));
  NOT NOT1_4590(.VSS(VSS),.VDD(VDD),.Y(g13457),.A(I20670));
  NOT NOT1_4591(.VSS(VSS),.VDD(VDD),.Y(I20673),.A(g13397));
  NOT NOT1_4592(.VSS(VSS),.VDD(VDD),.Y(g13458),.A(I20673));
  NOT NOT1_4593(.VSS(VSS),.VDD(VDD),.Y(I20676),.A(g11616));
  NOT NOT1_4594(.VSS(VSS),.VDD(VDD),.Y(g13459),.A(I20676));
  NOT NOT1_4595(.VSS(VSS),.VDD(VDD),.Y(I20679),.A(g11641));
  NOT NOT1_4596(.VSS(VSS),.VDD(VDD),.Y(g13460),.A(I20679));
  NOT NOT1_4597(.VSS(VSS),.VDD(VDD),.Y(I20682),.A(g11659));
  NOT NOT1_4598(.VSS(VSS),.VDD(VDD),.Y(g13461),.A(I20682));
  NOT NOT1_4599(.VSS(VSS),.VDD(VDD),.Y(I20685),.A(g11671));
  NOT NOT1_4600(.VSS(VSS),.VDD(VDD),.Y(g13462),.A(I20685));
  NOT NOT1_4601(.VSS(VSS),.VDD(VDD),.Y(I20688),.A(g11682));
  NOT NOT1_4602(.VSS(VSS),.VDD(VDD),.Y(g13463),.A(I20688));
  NOT NOT1_4603(.VSS(VSS),.VDD(VDD),.Y(I20691),.A(g13327));
  NOT NOT1_4604(.VSS(VSS),.VDD(VDD),.Y(g13464),.A(I20691));
  NOT NOT1_4605(.VSS(VSS),.VDD(VDD),.Y(I20694),.A(g13346));
  NOT NOT1_4606(.VSS(VSS),.VDD(VDD),.Y(g13465),.A(I20694));
  NOT NOT1_4607(.VSS(VSS),.VDD(VDD),.Y(I20697),.A(g13369));
  NOT NOT1_4608(.VSS(VSS),.VDD(VDD),.Y(g13466),.A(I20697));
  NOT NOT1_4609(.VSS(VSS),.VDD(VDD),.Y(I20700),.A(g12450));
  NOT NOT1_4610(.VSS(VSS),.VDD(VDD),.Y(g13467),.A(I20700));
  NOT NOT1_4611(.VSS(VSS),.VDD(VDD),.Y(I20703),.A(g12123));
  NOT NOT1_4612(.VSS(VSS),.VDD(VDD),.Y(g13468),.A(I20703));
  NOT NOT1_4613(.VSS(VSS),.VDD(VDD),.Y(I20706),.A(g11490));
  NOT NOT1_4614(.VSS(VSS),.VDD(VDD),.Y(g13469),.A(I20706));
  NOT NOT1_4615(.VSS(VSS),.VDD(VDD),.Y(I20709),.A(g13070));
  NOT NOT1_4616(.VSS(VSS),.VDD(VDD),.Y(g13475),.A(I20709));
  NOT NOT1_4617(.VSS(VSS),.VDD(VDD),.Y(g13519),.A(g13228));
  NOT NOT1_4618(.VSS(VSS),.VDD(VDD),.Y(g13530),.A(g13251));
  NOT NOT1_4619(.VSS(VSS),.VDD(VDD),.Y(g13541),.A(g13274));
  NOT NOT1_4620(.VSS(VSS),.VDD(VDD),.Y(g13552),.A(g13299));
  NOT NOT1_4621(.VSS(VSS),.VDD(VDD),.Y(g13565),.A(g12192));
  NOT NOT1_4622(.VSS(VSS),.VDD(VDD),.Y(g13568),.A(g11627));
  NOT NOT1_4623(.VSS(VSS),.VDD(VDD),.Y(I20791),.A(g13149));
  NOT NOT1_4624(.VSS(VSS),.VDD(VDD),.Y(g13571),.A(I20791));
  NOT NOT1_4625(.VSS(VSS),.VDD(VDD),.Y(I20794),.A(g13111));
  NOT NOT1_4626(.VSS(VSS),.VDD(VDD),.Y(g13572),.A(I20794));
  NOT NOT1_4627(.VSS(VSS),.VDD(VDD),.Y(g13573),.A(g12247));
  NOT NOT1_4628(.VSS(VSS),.VDD(VDD),.Y(g13576),.A(g11650));
  NOT NOT1_4629(.VSS(VSS),.VDD(VDD),.Y(I20799),.A(g13155));
  NOT NOT1_4630(.VSS(VSS),.VDD(VDD),.Y(g13579),.A(I20799));
  NOT NOT1_4631(.VSS(VSS),.VDD(VDD),.Y(I20802),.A(g13160));
  NOT NOT1_4632(.VSS(VSS),.VDD(VDD),.Y(g13580),.A(I20802));
  NOT NOT1_4633(.VSS(VSS),.VDD(VDD),.Y(I20805),.A(g13124));
  NOT NOT1_4634(.VSS(VSS),.VDD(VDD),.Y(g13581),.A(I20805));
  NOT NOT1_4635(.VSS(VSS),.VDD(VDD),.Y(g13582),.A(g12290));
  NOT NOT1_4636(.VSS(VSS),.VDD(VDD),.Y(g13585),.A(g11669));
  NOT NOT1_4637(.VSS(VSS),.VDD(VDD),.Y(I20810),.A(g13164));
  NOT NOT1_4638(.VSS(VSS),.VDD(VDD),.Y(g13588),.A(I20810));
  NOT NOT1_4639(.VSS(VSS),.VDD(VDD),.Y(I20813),.A(g13265));
  NOT NOT1_4640(.VSS(VSS),.VDD(VDD),.Y(g13589),.A(I20813));
  NOT NOT1_4641(.VSS(VSS),.VDD(VDD),.Y(I20816),.A(g12487));
  NOT NOT1_4642(.VSS(VSS),.VDD(VDD),.Y(g13598),.A(I20816));
  NOT NOT1_4643(.VSS(VSS),.VDD(VDD),.Y(I20820),.A(g13171));
  NOT NOT1_4644(.VSS(VSS),.VDD(VDD),.Y(g13600),.A(I20820));
  NOT NOT1_4645(.VSS(VSS),.VDD(VDD),.Y(I20823),.A(g13135));
  NOT NOT1_4646(.VSS(VSS),.VDD(VDD),.Y(g13601),.A(I20823));
  NOT NOT1_4647(.VSS(VSS),.VDD(VDD),.Y(g13602),.A(g12326));
  NOT NOT1_4648(.VSS(VSS),.VDD(VDD),.Y(g13605),.A(g11681));
  NOT NOT1_4649(.VSS(VSS),.VDD(VDD),.Y(I20828),.A(g13175));
  NOT NOT1_4650(.VSS(VSS),.VDD(VDD),.Y(g13608),.A(I20828));
  NOT NOT1_4651(.VSS(VSS),.VDD(VDD),.Y(I20832),.A(g12507));
  NOT NOT1_4652(.VSS(VSS),.VDD(VDD),.Y(g13610),.A(I20832));
  NOT NOT1_4653(.VSS(VSS),.VDD(VDD),.Y(I20836),.A(g13182));
  NOT NOT1_4654(.VSS(VSS),.VDD(VDD),.Y(g13612),.A(I20836));
  NOT NOT1_4655(.VSS(VSS),.VDD(VDD),.Y(I20839),.A(g13143));
  NOT NOT1_4656(.VSS(VSS),.VDD(VDD),.Y(g13613),.A(I20839));
  NOT NOT1_4657(.VSS(VSS),.VDD(VDD),.Y(g13614),.A(g11690));
  NOT NOT1_4658(.VSS(VSS),.VDD(VDD),.Y(I20844),.A(g12524));
  NOT NOT1_4659(.VSS(VSS),.VDD(VDD),.Y(g13620),.A(I20844));
  NOT NOT1_4660(.VSS(VSS),.VDD(VDD),.Y(I20848),.A(g13194));
  NOT NOT1_4661(.VSS(VSS),.VDD(VDD),.Y(g13622),.A(I20848));
  NOT NOT1_4662(.VSS(VSS),.VDD(VDD),.Y(I20852),.A(g12457));
  NOT NOT1_4663(.VSS(VSS),.VDD(VDD),.Y(g13624),.A(I20852));
  NOT NOT1_4664(.VSS(VSS),.VDD(VDD),.Y(g13626),.A(g11697));
  NOT NOT1_4665(.VSS(VSS),.VDD(VDD),.Y(I20858),.A(g12539));
  NOT NOT1_4666(.VSS(VSS),.VDD(VDD),.Y(g13632),.A(I20858));
  NOT NOT1_4667(.VSS(VSS),.VDD(VDD),.Y(I20863),.A(g12467));
  NOT NOT1_4668(.VSS(VSS),.VDD(VDD),.Y(g13635),.A(I20863));
  NOT NOT1_4669(.VSS(VSS),.VDD(VDD),.Y(g13637),.A(g11703));
  NOT NOT1_4670(.VSS(VSS),.VDD(VDD),.Y(g13644),.A(g13215));
  NOT NOT1_4671(.VSS(VSS),.VDD(VDD),.Y(I20873),.A(g12482));
  NOT NOT1_4672(.VSS(VSS),.VDD(VDD),.Y(g13647),.A(I20873));
  NOT NOT1_4673(.VSS(VSS),.VDD(VDD),.Y(g13649),.A(g11711));
  NOT NOT1_4674(.VSS(VSS),.VDD(VDD),.Y(g13657),.A(g12452));
  NOT NOT1_4675(.VSS(VSS),.VDD(VDD),.Y(g13669),.A(g13229));
  NOT NOT1_4676(.VSS(VSS),.VDD(VDD),.Y(g13670),.A(g13234));
  NOT NOT1_4677(.VSS(VSS),.VDD(VDD),.Y(I20886),.A(g12499));
  NOT NOT1_4678(.VSS(VSS),.VDD(VDD),.Y(g13673),.A(I20886));
  NOT NOT1_4679(.VSS(VSS),.VDD(VDD),.Y(g13677),.A(g12447));
  NOT NOT1_4680(.VSS(VSS),.VDD(VDD),.Y(g13687),.A(g12460));
  NOT NOT1_4681(.VSS(VSS),.VDD(VDD),.Y(g13699),.A(g13252));
  NOT NOT1_4682(.VSS(VSS),.VDD(VDD),.Y(g13700),.A(g13257));
  NOT NOT1_4683(.VSS(VSS),.VDD(VDD),.Y(g13706),.A(g12443));
  NOT NOT1_4684(.VSS(VSS),.VDD(VDD),.Y(g13714),.A(g12453));
  NOT NOT1_4685(.VSS(VSS),.VDD(VDD),.Y(g13724),.A(g12470));
  NOT NOT1_4686(.VSS(VSS),.VDD(VDD),.Y(g13736),.A(g13275));
  NOT NOT1_4687(.VSS(VSS),.VDD(VDD),.Y(g13737),.A(g13280));
  NOT NOT1_4688(.VSS(VSS),.VDD(VDD),.Y(I20909),.A(g13055));
  NOT NOT1_4689(.VSS(VSS),.VDD(VDD),.Y(g13741),.A(I20909));
  NOT NOT1_4690(.VSS(VSS),.VDD(VDD),.Y(g13750),.A(g12439));
  NOT NOT1_4691(.VSS(VSS),.VDD(VDD),.Y(g13756),.A(g12448));
  NOT NOT1_4692(.VSS(VSS),.VDD(VDD),.Y(g13764),.A(g12461));
  NOT NOT1_4693(.VSS(VSS),.VDD(VDD),.Y(g13774),.A(g12485));
  NOT NOT1_4694(.VSS(VSS),.VDD(VDD),.Y(g13786),.A(g13300));
  NOT NOT1_4695(.VSS(VSS),.VDD(VDD),.Y(g13791),.A(g12444));
  NOT NOT1_4696(.VSS(VSS),.VDD(VDD),.Y(g13797),.A(g12454));
  NOT NOT1_4697(.VSS(VSS),.VDD(VDD),.Y(g13805),.A(g12471));
  NOT NOT1_4698(.VSS(VSS),.VDD(VDD),.Y(g13817),.A(g13336));
  NOT NOT1_4699(.VSS(VSS),.VDD(VDD),.Y(g13819),.A(g12449));
  NOT NOT1_4700(.VSS(VSS),.VDD(VDD),.Y(g13825),.A(g12462));
  NOT NOT1_4701(.VSS(VSS),.VDD(VDD),.Y(g13836),.A(g13356));
  NOT NOT1_4702(.VSS(VSS),.VDD(VDD),.Y(g13838),.A(g13361));
  NOT NOT1_4703(.VSS(VSS),.VDD(VDD),.Y(g13840),.A(g12455));
  NOT NOT1_4704(.VSS(VSS),.VDD(VDD),.Y(g13848),.A(g11744));
  NOT NOT1_4705(.VSS(VSS),.VDD(VDD),.Y(g13849),.A(g13381));
  NOT NOT1_4706(.VSS(VSS),.VDD(VDD),.Y(g13850),.A(g13386));
  NOT NOT1_4707(.VSS(VSS),.VDD(VDD),.Y(g13852),.A(g13391));
  NOT NOT1_4708(.VSS(VSS),.VDD(VDD),.Y(g13856),.A(g11759));
  NOT NOT1_4709(.VSS(VSS),.VDD(VDD),.Y(g13857),.A(g11760));
  NOT NOT1_4710(.VSS(VSS),.VDD(VDD),.Y(g13858),.A(g11603));
  NOT NOT1_4711(.VSS(VSS),.VDD(VDD),.Y(g13859),.A(g11608));
  NOT NOT1_4712(.VSS(VSS),.VDD(VDD),.Y(g13861),.A(g11613));
  NOT NOT1_4713(.VSS(VSS),.VDD(VDD),.Y(I20959),.A(g11713));
  NOT NOT1_4714(.VSS(VSS),.VDD(VDD),.Y(g13863),.A(I20959));
  NOT NOT1_4715(.VSS(VSS),.VDD(VDD),.Y(g13864),.A(g11767));
  NOT NOT1_4716(.VSS(VSS),.VDD(VDD),.Y(g13866),.A(g11772));
  NOT NOT1_4717(.VSS(VSS),.VDD(VDD),.Y(g13867),.A(g11773));
  NOT NOT1_4718(.VSS(VSS),.VDD(VDD),.Y(g13868),.A(g11633));
  NOT NOT1_4719(.VSS(VSS),.VDD(VDD),.Y(g13869),.A(g11638));
  NOT NOT1_4720(.VSS(VSS),.VDD(VDD),.Y(g13872),.A(g11780));
  NOT NOT1_4721(.VSS(VSS),.VDD(VDD),.Y(g13873),.A(g12698));
  NOT NOT1_4722(.VSS(VSS),.VDD(VDD),.Y(g13879),.A(g11784));
  NOT NOT1_4723(.VSS(VSS),.VDD(VDD),.Y(g13881),.A(g11789));
  NOT NOT1_4724(.VSS(VSS),.VDD(VDD),.Y(g13882),.A(g11790));
  NOT NOT1_4725(.VSS(VSS),.VDD(VDD),.Y(g13883),.A(g11656));
  NOT NOT1_4726(.VSS(VSS),.VDD(VDD),.Y(g13885),.A(g11799));
  NOT NOT1_4727(.VSS(VSS),.VDD(VDD),.Y(g13886),.A(g12747));
  NOT NOT1_4728(.VSS(VSS),.VDD(VDD),.Y(g13894),.A(g11806));
  NOT NOT1_4729(.VSS(VSS),.VDD(VDD),.Y(g13895),.A(g12755));
  NOT NOT1_4730(.VSS(VSS),.VDD(VDD),.Y(g13901),.A(g11810));
  NOT NOT1_4731(.VSS(VSS),.VDD(VDD),.Y(g13903),.A(g11815));
  NOT NOT1_4732(.VSS(VSS),.VDD(VDD),.Y(g13906),.A(g11822));
  NOT NOT1_4733(.VSS(VSS),.VDD(VDD),.Y(g13907),.A(g12781));
  NOT NOT1_4734(.VSS(VSS),.VDD(VDD),.Y(g13918),.A(g11830));
  NOT NOT1_4735(.VSS(VSS),.VDD(VDD),.Y(g13922),.A(g11831));
  NOT NOT1_4736(.VSS(VSS),.VDD(VDD),.Y(g13926),.A(g11832));
  NOT NOT1_4737(.VSS(VSS),.VDD(VDD),.Y(g13927),.A(g12789));
  NOT NOT1_4738(.VSS(VSS),.VDD(VDD),.Y(g13935),.A(g11839));
  NOT NOT1_4739(.VSS(VSS),.VDD(VDD),.Y(g13936),.A(g12797));
  NOT NOT1_4740(.VSS(VSS),.VDD(VDD),.Y(g13942),.A(g11843));
  NOT NOT1_4741(.VSS(VSS),.VDD(VDD),.Y(g13945),.A(g11855));
  NOT NOT1_4742(.VSS(VSS),.VDD(VDD),.Y(g13946),.A(g12814));
  NOT NOT1_4743(.VSS(VSS),.VDD(VDD),.Y(I21012),.A(g12503));
  NOT NOT1_4744(.VSS(VSS),.VDD(VDD),.Y(g13954),.A(I21012));
  NOT NOT1_4745(.VSS(VSS),.VDD(VDD),.Y(g13958),.A(g11863));
  NOT NOT1_4746(.VSS(VSS),.VDD(VDD),.Y(g13962),.A(g11864));
  NOT NOT1_4747(.VSS(VSS),.VDD(VDD),.Y(g13963),.A(g12820));
  NOT NOT1_4748(.VSS(VSS),.VDD(VDD),.Y(g13974),.A(g11872));
  NOT NOT1_4749(.VSS(VSS),.VDD(VDD),.Y(g13978),.A(g11873));
  NOT NOT1_4750(.VSS(VSS),.VDD(VDD),.Y(g13982),.A(g11874));
  NOT NOT1_4751(.VSS(VSS),.VDD(VDD),.Y(g13983),.A(g12828));
  NOT NOT1_4752(.VSS(VSS),.VDD(VDD),.Y(g13991),.A(g11881));
  NOT NOT1_4753(.VSS(VSS),.VDD(VDD),.Y(g13992),.A(g12836));
  NOT NOT1_4754(.VSS(VSS),.VDD(VDD),.Y(g13999),.A(g11889));
  NOT NOT1_4755(.VSS(VSS),.VDD(VDD),.Y(g14000),.A(g11890));
  NOT NOT1_4756(.VSS(VSS),.VDD(VDD),.Y(g14001),.A(g12849));
  NOT NOT1_4757(.VSS(VSS),.VDD(VDD),.Y(I21037),.A(g12486));
  NOT NOT1_4758(.VSS(VSS),.VDD(VDD),.Y(g14008),.A(I21037));
  NOT NOT1_4759(.VSS(VSS),.VDD(VDD),.Y(g14011),.A(g11896));
  NOT NOT1_4760(.VSS(VSS),.VDD(VDD),.Y(g14015),.A(g11897));
  NOT NOT1_4761(.VSS(VSS),.VDD(VDD),.Y(g14016),.A(g12852));
  NOT NOT1_4762(.VSS(VSS),.VDD(VDD),.Y(I21045),.A(g12520));
  NOT NOT1_4763(.VSS(VSS),.VDD(VDD),.Y(g14024),.A(I21045));
  NOT NOT1_4764(.VSS(VSS),.VDD(VDD),.Y(g14028),.A(g11905));
  NOT NOT1_4765(.VSS(VSS),.VDD(VDD),.Y(g14032),.A(g11906));
  NOT NOT1_4766(.VSS(VSS),.VDD(VDD),.Y(g14033),.A(g12858));
  NOT NOT1_4767(.VSS(VSS),.VDD(VDD),.Y(g14044),.A(g11914));
  NOT NOT1_4768(.VSS(VSS),.VDD(VDD),.Y(g14048),.A(g11915));
  NOT NOT1_4769(.VSS(VSS),.VDD(VDD),.Y(g14052),.A(g11916));
  NOT NOT1_4770(.VSS(VSS),.VDD(VDD),.Y(g14053),.A(g12866));
  NOT NOT1_4771(.VSS(VSS),.VDD(VDD),.Y(g14061),.A(g11928));
  NOT NOT1_4772(.VSS(VSS),.VDD(VDD),.Y(g14062),.A(g12880));
  NOT NOT1_4773(.VSS(VSS),.VDD(VDD),.Y(I21064),.A(g13147));
  NOT NOT1_4774(.VSS(VSS),.VDD(VDD),.Y(g14068),.A(I21064));
  NOT NOT1_4775(.VSS(VSS),.VDD(VDD),.Y(g14071),.A(g11934));
  NOT NOT1_4776(.VSS(VSS),.VDD(VDD),.Y(g14079),.A(g11935));
  NOT NOT1_4777(.VSS(VSS),.VDD(VDD),.Y(g14086),.A(g11938));
  NOT NOT1_4778(.VSS(VSS),.VDD(VDD),.Y(g14090),.A(g11939));
  NOT NOT1_4779(.VSS(VSS),.VDD(VDD),.Y(g14091),.A(g11940));
  NOT NOT1_4780(.VSS(VSS),.VDD(VDD),.Y(g14092),.A(g12890));
  NOT NOT1_4781(.VSS(VSS),.VDD(VDD),.Y(I21075),.A(g12506));
  NOT NOT1_4782(.VSS(VSS),.VDD(VDD),.Y(g14099),.A(I21075));
  NOT NOT1_4783(.VSS(VSS),.VDD(VDD),.Y(g14102),.A(g11946));
  NOT NOT1_4784(.VSS(VSS),.VDD(VDD),.Y(g14106),.A(g11947));
  NOT NOT1_4785(.VSS(VSS),.VDD(VDD),.Y(g14107),.A(g12893));
  NOT NOT1_4786(.VSS(VSS),.VDD(VDD),.Y(I21083),.A(g12535));
  NOT NOT1_4787(.VSS(VSS),.VDD(VDD),.Y(g14115),.A(I21083));
  NOT NOT1_4788(.VSS(VSS),.VDD(VDD),.Y(g14119),.A(g11955));
  NOT NOT1_4789(.VSS(VSS),.VDD(VDD),.Y(g14123),.A(g11956));
  NOT NOT1_4790(.VSS(VSS),.VDD(VDD),.Y(g14124),.A(g12899));
  NOT NOT1_4791(.VSS(VSS),.VDD(VDD),.Y(g14135),.A(g11964));
  NOT NOT1_4792(.VSS(VSS),.VDD(VDD),.Y(g14139),.A(g11965));
  NOT NOT1_4793(.VSS(VSS),.VDD(VDD),.Y(I21096),.A(g11749));
  NOT NOT1_4794(.VSS(VSS),.VDD(VDD),.Y(g14144),.A(I21096));
  NOT NOT1_4795(.VSS(VSS),.VDD(VDD),.Y(g14148),.A(g12912));
  NOT NOT1_4796(.VSS(VSS),.VDD(VDD),.Y(g14153),.A(g12913));
  NOT NOT1_4797(.VSS(VSS),.VDD(VDD),.Y(g14158),.A(g11974));
  NOT NOT1_4798(.VSS(VSS),.VDD(VDD),.Y(g14165),.A(g11975));
  NOT NOT1_4799(.VSS(VSS),.VDD(VDD),.Y(g14171),.A(g11979));
  NOT NOT1_4800(.VSS(VSS),.VDD(VDD),.Y(g14175),.A(g11980));
  NOT NOT1_4801(.VSS(VSS),.VDD(VDD),.Y(g14176),.A(g11981));
  NOT NOT1_4802(.VSS(VSS),.VDD(VDD),.Y(g14177),.A(g12920));
  NOT NOT1_4803(.VSS(VSS),.VDD(VDD),.Y(I21108),.A(g13150));
  NOT NOT1_4804(.VSS(VSS),.VDD(VDD),.Y(g14183),.A(I21108));
  NOT NOT1_4805(.VSS(VSS),.VDD(VDD),.Y(g14186),.A(g11987));
  NOT NOT1_4806(.VSS(VSS),.VDD(VDD),.Y(g14194),.A(g11988));
  NOT NOT1_4807(.VSS(VSS),.VDD(VDD),.Y(g14201),.A(g11991));
  NOT NOT1_4808(.VSS(VSS),.VDD(VDD),.Y(g14205),.A(g11992));
  NOT NOT1_4809(.VSS(VSS),.VDD(VDD),.Y(g14206),.A(g11993));
  NOT NOT1_4810(.VSS(VSS),.VDD(VDD),.Y(g14207),.A(g12930));
  NOT NOT1_4811(.VSS(VSS),.VDD(VDD),.Y(I21119),.A(g12523));
  NOT NOT1_4812(.VSS(VSS),.VDD(VDD),.Y(g14214),.A(I21119));
  NOT NOT1_4813(.VSS(VSS),.VDD(VDD),.Y(g14217),.A(g11999));
  NOT NOT1_4814(.VSS(VSS),.VDD(VDD),.Y(g14221),.A(g12000));
  NOT NOT1_4815(.VSS(VSS),.VDD(VDD),.Y(g14222),.A(g12933));
  NOT NOT1_4816(.VSS(VSS),.VDD(VDD),.Y(I21127),.A(g12544));
  NOT NOT1_4817(.VSS(VSS),.VDD(VDD),.Y(g14230),.A(I21127));
  NOT NOT1_4818(.VSS(VSS),.VDD(VDD),.Y(g14234),.A(g12008));
  NOT NOT1_4819(.VSS(VSS),.VDD(VDD),.Y(g14238),.A(g12939));
  NOT NOT1_4820(.VSS(VSS),.VDD(VDD),.Y(g14244),.A(g12026));
  NOT NOT1_4821(.VSS(VSS),.VDD(VDD),.Y(g14249),.A(g12034));
  NOT NOT1_4822(.VSS(VSS),.VDD(VDD),.Y(g14252),.A(g12035));
  NOT NOT1_4823(.VSS(VSS),.VDD(VDD),.Y(g14256),.A(g12036));
  NOT NOT1_4824(.VSS(VSS),.VDD(VDD),.Y(I21137),.A(g11749));
  NOT NOT1_4825(.VSS(VSS),.VDD(VDD),.Y(g14259),.A(I21137));
  NOT NOT1_4826(.VSS(VSS),.VDD(VDD),.Y(g14263),.A(g12941));
  NOT NOT1_4827(.VSS(VSS),.VDD(VDD),.Y(g14268),.A(g12942));
  NOT NOT1_4828(.VSS(VSS),.VDD(VDD),.Y(g14273),.A(g12043));
  NOT NOT1_4829(.VSS(VSS),.VDD(VDD),.Y(g14280),.A(g12044));
  NOT NOT1_4830(.VSS(VSS),.VDD(VDD),.Y(g14286),.A(g12048));
  NOT NOT1_4831(.VSS(VSS),.VDD(VDD),.Y(g14290),.A(g12049));
  NOT NOT1_4832(.VSS(VSS),.VDD(VDD),.Y(g14291),.A(g12050));
  NOT NOT1_4833(.VSS(VSS),.VDD(VDD),.Y(g14292),.A(g12949));
  NOT NOT1_4834(.VSS(VSS),.VDD(VDD),.Y(I21149),.A(g13156));
  NOT NOT1_4835(.VSS(VSS),.VDD(VDD),.Y(g14298),.A(I21149));
  NOT NOT1_4836(.VSS(VSS),.VDD(VDD),.Y(g14301),.A(g12056));
  NOT NOT1_4837(.VSS(VSS),.VDD(VDD),.Y(g14309),.A(g12057));
  NOT NOT1_4838(.VSS(VSS),.VDD(VDD),.Y(g14316),.A(g12060));
  NOT NOT1_4839(.VSS(VSS),.VDD(VDD),.Y(g14320),.A(g12061));
  NOT NOT1_4840(.VSS(VSS),.VDD(VDD),.Y(g14321),.A(g12062));
  NOT NOT1_4841(.VSS(VSS),.VDD(VDD),.Y(g14322),.A(g12959));
  NOT NOT1_4842(.VSS(VSS),.VDD(VDD),.Y(I21160),.A(g12538));
  NOT NOT1_4843(.VSS(VSS),.VDD(VDD),.Y(g14329),.A(I21160));
  NOT NOT1_4844(.VSS(VSS),.VDD(VDD),.Y(g14332),.A(g12068));
  NOT NOT1_4845(.VSS(VSS),.VDD(VDD),.Y(I21165),.A(g13110));
  NOT NOT1_4846(.VSS(VSS),.VDD(VDD),.Y(g14337),.A(I21165));
  NOT NOT1_4847(.VSS(VSS),.VDD(VDD),.Y(g14342),.A(g12967));
  NOT NOT1_4848(.VSS(VSS),.VDD(VDD),.Y(g14347),.A(g12079));
  NOT NOT1_4849(.VSS(VSS),.VDD(VDD),.Y(g14352),.A(g12081));
  NOT NOT1_4850(.VSS(VSS),.VDD(VDD),.Y(g14355),.A(g12082));
  NOT NOT1_4851(.VSS(VSS),.VDD(VDD),.Y(g14359),.A(g12083));
  NOT NOT1_4852(.VSS(VSS),.VDD(VDD),.Y(g14360),.A(g12968));
  NOT NOT1_4853(.VSS(VSS),.VDD(VDD),.Y(g14366),.A(g12090));
  NOT NOT1_4854(.VSS(VSS),.VDD(VDD),.Y(g14371),.A(g12098));
  NOT NOT1_4855(.VSS(VSS),.VDD(VDD),.Y(g14374),.A(g12099));
  NOT NOT1_4856(.VSS(VSS),.VDD(VDD),.Y(g14378),.A(g12100));
  NOT NOT1_4857(.VSS(VSS),.VDD(VDD),.Y(I21178),.A(g11749));
  NOT NOT1_4858(.VSS(VSS),.VDD(VDD),.Y(g14381),.A(I21178));
  NOT NOT1_4859(.VSS(VSS),.VDD(VDD),.Y(g14385),.A(g12970));
  NOT NOT1_4860(.VSS(VSS),.VDD(VDD),.Y(g14390),.A(g12971));
  NOT NOT1_4861(.VSS(VSS),.VDD(VDD),.Y(g14395),.A(g12107));
  NOT NOT1_4862(.VSS(VSS),.VDD(VDD),.Y(g14402),.A(g12108));
  NOT NOT1_4863(.VSS(VSS),.VDD(VDD),.Y(g14408),.A(g12112));
  NOT NOT1_4864(.VSS(VSS),.VDD(VDD),.Y(g14412),.A(g12113));
  NOT NOT1_4865(.VSS(VSS),.VDD(VDD),.Y(g14413),.A(g12114));
  NOT NOT1_4866(.VSS(VSS),.VDD(VDD),.Y(g14414),.A(g12978));
  NOT NOT1_4867(.VSS(VSS),.VDD(VDD),.Y(I21190),.A(g13165));
  NOT NOT1_4868(.VSS(VSS),.VDD(VDD),.Y(g14420),.A(I21190));
  NOT NOT1_4869(.VSS(VSS),.VDD(VDD),.Y(g14423),.A(g12120));
  NOT NOT1_4870(.VSS(VSS),.VDD(VDD),.Y(g14431),.A(g12121));
  NOT NOT1_4871(.VSS(VSS),.VDD(VDD),.Y(g14438),.A(g12124));
  NOT NOT1_4872(.VSS(VSS),.VDD(VDD),.Y(g14442),.A(g11768));
  NOT NOT1_4873(.VSS(VSS),.VDD(VDD),.Y(g14450),.A(g12146));
  NOT NOT1_4874(.VSS(VSS),.VDD(VDD),.Y(g14454),.A(g12991));
  NOT NOT1_4875(.VSS(VSS),.VDD(VDD),.Y(g14459),.A(g12151));
  NOT NOT1_4876(.VSS(VSS),.VDD(VDD),.Y(g14464),.A(g12153));
  NOT NOT1_4877(.VSS(VSS),.VDD(VDD),.Y(g14467),.A(g12154));
  NOT NOT1_4878(.VSS(VSS),.VDD(VDD),.Y(g14471),.A(g12155));
  NOT NOT1_4879(.VSS(VSS),.VDD(VDD),.Y(g14472),.A(g12992));
  NOT NOT1_4880(.VSS(VSS),.VDD(VDD),.Y(g14478),.A(g12162));
  NOT NOT1_4881(.VSS(VSS),.VDD(VDD),.Y(g14483),.A(g12170));
  NOT NOT1_4882(.VSS(VSS),.VDD(VDD),.Y(g14486),.A(g12171));
  NOT NOT1_4883(.VSS(VSS),.VDD(VDD),.Y(g14490),.A(g12172));
  NOT NOT1_4884(.VSS(VSS),.VDD(VDD),.Y(I21208),.A(g11749));
  NOT NOT1_4885(.VSS(VSS),.VDD(VDD),.Y(g14493),.A(I21208));
  NOT NOT1_4886(.VSS(VSS),.VDD(VDD),.Y(g14497),.A(g12994));
  NOT NOT1_4887(.VSS(VSS),.VDD(VDD),.Y(g14502),.A(g12995));
  NOT NOT1_4888(.VSS(VSS),.VDD(VDD),.Y(g14507),.A(g12179));
  NOT NOT1_4889(.VSS(VSS),.VDD(VDD),.Y(g14514),.A(g12180));
  NOT NOT1_4890(.VSS(VSS),.VDD(VDD),.Y(g14520),.A(g12184));
  NOT NOT1_4891(.VSS(VSS),.VDD(VDD),.Y(g14524),.A(g12185));
  NOT NOT1_4892(.VSS(VSS),.VDD(VDD),.Y(g14525),.A(g12195));
  NOT NOT1_4893(.VSS(VSS),.VDD(VDD),.Y(g14529),.A(g11785));
  NOT NOT1_4894(.VSS(VSS),.VDD(VDD),.Y(g14537),.A(g12208));
  NOT NOT1_4895(.VSS(VSS),.VDD(VDD),.Y(g14541),.A(g13001));
  NOT NOT1_4896(.VSS(VSS),.VDD(VDD),.Y(g14546),.A(g12213));
  NOT NOT1_4897(.VSS(VSS),.VDD(VDD),.Y(g14551),.A(g12215));
  NOT NOT1_4898(.VSS(VSS),.VDD(VDD),.Y(g14554),.A(g12216));
  NOT NOT1_4899(.VSS(VSS),.VDD(VDD),.Y(g14558),.A(g12217));
  NOT NOT1_4900(.VSS(VSS),.VDD(VDD),.Y(g14559),.A(g13002));
  NOT NOT1_4901(.VSS(VSS),.VDD(VDD),.Y(g14565),.A(g12224));
  NOT NOT1_4902(.VSS(VSS),.VDD(VDD),.Y(g14570),.A(g12232));
  NOT NOT1_4903(.VSS(VSS),.VDD(VDD),.Y(g14573),.A(g12233));
  NOT NOT1_4904(.VSS(VSS),.VDD(VDD),.Y(g14577),.A(g12234));
  NOT NOT1_4905(.VSS(VSS),.VDD(VDD),.Y(g14580),.A(g12250));
  NOT NOT1_4906(.VSS(VSS),.VDD(VDD),.Y(g14584),.A(g11811));
  NOT NOT1_4907(.VSS(VSS),.VDD(VDD),.Y(g14592),.A(g12263));
  NOT NOT1_4908(.VSS(VSS),.VDD(VDD),.Y(g14596),.A(g13022));
  NOT NOT1_4909(.VSS(VSS),.VDD(VDD),.Y(g14601),.A(g12268));
  NOT NOT1_4910(.VSS(VSS),.VDD(VDD),.Y(g14606),.A(g12270));
  NOT NOT1_4911(.VSS(VSS),.VDD(VDD),.Y(g14609),.A(g12271));
  NOT NOT1_4912(.VSS(VSS),.VDD(VDD),.Y(g14613),.A(g12272));
  NOT NOT1_4913(.VSS(VSS),.VDD(VDD),.Y(g14614),.A(g12293));
  NOT NOT1_4914(.VSS(VSS),.VDD(VDD),.Y(g14618),.A(g11844));
  NOT NOT1_4915(.VSS(VSS),.VDD(VDD),.Y(g14626),.A(g12306));
  NOT NOT1_4916(.VSS(VSS),.VDD(VDD),.Y(I21241),.A(g13378));
  NOT NOT1_4917(.VSS(VSS),.VDD(VDD),.Y(g14630),.A(I21241));
  NOT NOT1_4918(.VSS(VSS),.VDD(VDD),.Y(g14637),.A(g12329));
  NOT NOT1_4919(.VSS(VSS),.VDD(VDD),.Y(g14641),.A(g11823));
  NOT NOT1_4920(.VSS(VSS),.VDD(VDD),.Y(I21246),.A(g11624));
  NOT NOT1_4921(.VSS(VSS),.VDD(VDD),.Y(g14642),.A(I21246));
  NOT NOT1_4922(.VSS(VSS),.VDD(VDD),.Y(I21249),.A(g11600));
  NOT NOT1_4923(.VSS(VSS),.VDD(VDD),.Y(g14650),.A(I21249));
  NOT NOT1_4924(.VSS(VSS),.VDD(VDD),.Y(I21252),.A(g11644));
  NOT NOT1_4925(.VSS(VSS),.VDD(VDD),.Y(g14657),.A(I21252));
  NOT NOT1_4926(.VSS(VSS),.VDD(VDD),.Y(g14668),.A(g11865));
  NOT NOT1_4927(.VSS(VSS),.VDD(VDD),.Y(I21256),.A(g11647));
  NOT NOT1_4928(.VSS(VSS),.VDD(VDD),.Y(g14669),.A(I21256));
  NOT NOT1_4929(.VSS(VSS),.VDD(VDD),.Y(I21259),.A(g11630));
  NOT NOT1_4930(.VSS(VSS),.VDD(VDD),.Y(g14677),.A(I21259));
  NOT NOT1_4931(.VSS(VSS),.VDD(VDD),.Y(I21262),.A(g11713));
  NOT NOT1_4932(.VSS(VSS),.VDD(VDD),.Y(g14684),.A(I21262));
  NOT NOT1_4933(.VSS(VSS),.VDD(VDD),.Y(g14685),.A(g12245));
  NOT NOT1_4934(.VSS(VSS),.VDD(VDD),.Y(I21267),.A(g11663));
  NOT NOT1_4935(.VSS(VSS),.VDD(VDD),.Y(g14691),.A(I21267));
  NOT NOT1_4936(.VSS(VSS),.VDD(VDD),.Y(g14702),.A(g11907));
  NOT NOT1_4937(.VSS(VSS),.VDD(VDD),.Y(I21271),.A(g11666));
  NOT NOT1_4938(.VSS(VSS),.VDD(VDD),.Y(g14703),.A(I21271));
  NOT NOT1_4939(.VSS(VSS),.VDD(VDD),.Y(I21274),.A(g11653));
  NOT NOT1_4940(.VSS(VSS),.VDD(VDD),.Y(g14711),.A(I21274));
  NOT NOT1_4941(.VSS(VSS),.VDD(VDD),.Y(I21277),.A(g12430));
  NOT NOT1_4942(.VSS(VSS),.VDD(VDD),.Y(g14718),.A(I21277));
  NOT NOT1_4943(.VSS(VSS),.VDD(VDD),.Y(g14719),.A(g12288));
  NOT NOT1_4944(.VSS(VSS),.VDD(VDD),.Y(I21282),.A(g11675));
  NOT NOT1_4945(.VSS(VSS),.VDD(VDD),.Y(g14725),.A(I21282));
  NOT NOT1_4946(.VSS(VSS),.VDD(VDD),.Y(g14736),.A(g11957));
  NOT NOT1_4947(.VSS(VSS),.VDD(VDD),.Y(I21286),.A(g11678));
  NOT NOT1_4948(.VSS(VSS),.VDD(VDD),.Y(g14737),.A(I21286));
  NOT NOT1_4949(.VSS(VSS),.VDD(VDD),.Y(I21289),.A(g12434));
  NOT NOT1_4950(.VSS(VSS),.VDD(VDD),.Y(g14745),.A(I21289));
  NOT NOT1_4951(.VSS(VSS),.VDD(VDD),.Y(I21292),.A(g11888));
  NOT NOT1_4952(.VSS(VSS),.VDD(VDD),.Y(g14746),.A(I21292));
  NOT NOT1_4953(.VSS(VSS),.VDD(VDD),.Y(g14747),.A(g12324));
  NOT NOT1_4954(.VSS(VSS),.VDD(VDD),.Y(I21297),.A(g11687));
  NOT NOT1_4955(.VSS(VSS),.VDD(VDD),.Y(g14753),.A(I21297));
  NOT NOT1_4956(.VSS(VSS),.VDD(VDD),.Y(g14764),.A(g11791));
  NOT NOT1_4957(.VSS(VSS),.VDD(VDD),.Y(I21301),.A(g12438));
  NOT NOT1_4958(.VSS(VSS),.VDD(VDD),.Y(g14765),.A(I21301));
  NOT NOT1_4959(.VSS(VSS),.VDD(VDD),.Y(I21304),.A(g11927));
  NOT NOT1_4960(.VSS(VSS),.VDD(VDD),.Y(g14766),.A(I21304));
  NOT NOT1_4961(.VSS(VSS),.VDD(VDD),.Y(g14768),.A(g12352));
  NOT NOT1_4962(.VSS(VSS),.VDD(VDD),.Y(I21310),.A(g12332));
  NOT NOT1_4963(.VSS(VSS),.VDD(VDD),.Y(g14774),.A(I21310));
  NOT NOT1_4964(.VSS(VSS),.VDD(VDD),.Y(I21313),.A(g11743));
  NOT NOT1_4965(.VSS(VSS),.VDD(VDD),.Y(g14775),.A(I21313));
  NOT NOT1_4966(.VSS(VSS),.VDD(VDD),.Y(g14776),.A(g12033));
  NOT NOT1_4967(.VSS(VSS),.VDD(VDD),.Y(g14794),.A(g11848));
  NOT NOT1_4968(.VSS(VSS),.VDD(VDD),.Y(I21318),.A(g12362));
  NOT NOT1_4969(.VSS(VSS),.VDD(VDD),.Y(g14795),.A(I21318));
  NOT NOT1_4970(.VSS(VSS),.VDD(VDD),.Y(I21321),.A(g11758));
  NOT NOT1_4971(.VSS(VSS),.VDD(VDD),.Y(g14796),.A(I21321));
  NOT NOT1_4972(.VSS(VSS),.VDD(VDD),.Y(g14797),.A(g12080));
  NOT NOT1_4973(.VSS(VSS),.VDD(VDD),.Y(g14811),.A(g12097));
  NOT NOT1_4974(.VSS(VSS),.VDD(VDD),.Y(I21326),.A(g12378));
  NOT NOT1_4975(.VSS(VSS),.VDD(VDD),.Y(g14829),.A(I21326));
  NOT NOT1_4976(.VSS(VSS),.VDD(VDD),.Y(I21329),.A(g11766));
  NOT NOT1_4977(.VSS(VSS),.VDD(VDD),.Y(g14830),.A(I21329));
  NOT NOT1_4978(.VSS(VSS),.VDD(VDD),.Y(g14831),.A(g11828));
  NOT NOT1_4979(.VSS(VSS),.VDD(VDD),.Y(g14837),.A(g12145));
  NOT NOT1_4980(.VSS(VSS),.VDD(VDD),.Y(g14849),.A(g12152));
  NOT NOT1_4981(.VSS(VSS),.VDD(VDD),.Y(g14863),.A(g12169));
  NOT NOT1_4982(.VSS(VSS),.VDD(VDD),.Y(g14881),.A(g11923));
  NOT NOT1_4983(.VSS(VSS),.VDD(VDD),.Y(I21337),.A(g12408));
  NOT NOT1_4984(.VSS(VSS),.VDD(VDD),.Y(g14882),.A(I21337));
  NOT NOT1_4985(.VSS(VSS),.VDD(VDD),.Y(I21340),.A(g11779));
  NOT NOT1_4986(.VSS(VSS),.VDD(VDD),.Y(g14883),.A(I21340));
  NOT NOT1_4987(.VSS(VSS),.VDD(VDD),.Y(g14885),.A(g11860));
  NOT NOT1_4988(.VSS(VSS),.VDD(VDD),.Y(g14895),.A(g12193));
  NOT NOT1_4989(.VSS(VSS),.VDD(VDD),.Y(g14904),.A(g11870));
  NOT NOT1_4990(.VSS(VSS),.VDD(VDD),.Y(g14910),.A(g12207));
  NOT NOT1_4991(.VSS(VSS),.VDD(VDD),.Y(g14922),.A(g12214));
  NOT NOT1_4992(.VSS(VSS),.VDD(VDD),.Y(g14936),.A(g12231));
  NOT NOT1_4993(.VSS(VSS),.VDD(VDD),.Y(I21351),.A(g12420));
  NOT NOT1_4994(.VSS(VSS),.VDD(VDD),.Y(g14954),.A(I21351));
  NOT NOT1_4995(.VSS(VSS),.VDD(VDD),.Y(I21354),.A(g11798));
  NOT NOT1_4996(.VSS(VSS),.VDD(VDD),.Y(g14955),.A(I21354));
  NOT NOT1_4997(.VSS(VSS),.VDD(VDD),.Y(g14959),.A(g11976));
  NOT NOT1_4998(.VSS(VSS),.VDD(VDD),.Y(I21361),.A(g13026));
  NOT NOT1_4999(.VSS(VSS),.VDD(VDD),.Y(g14960),.A(I21361));
  NOT NOT1_5000(.VSS(VSS),.VDD(VDD),.Y(I21364),.A(g13028));
  NOT NOT1_5001(.VSS(VSS),.VDD(VDD),.Y(g14963),.A(I21364));
  NOT NOT1_5002(.VSS(VSS),.VDD(VDD),.Y(g14966),.A(g11902));
  NOT NOT1_5003(.VSS(VSS),.VDD(VDD),.Y(g14976),.A(g12248));
  NOT NOT1_5004(.VSS(VSS),.VDD(VDD),.Y(g14985),.A(g11912));
  NOT NOT1_5005(.VSS(VSS),.VDD(VDD),.Y(g14991),.A(g12262));
  NOT NOT1_5006(.VSS(VSS),.VDD(VDD),.Y(g15003),.A(g12269));
  NOT NOT1_5007(.VSS(VSS),.VDD(VDD),.Y(g15017),.A(g12009));
  NOT NOT1_5008(.VSS(VSS),.VDD(VDD),.Y(I21374),.A(g12424));
  NOT NOT1_5009(.VSS(VSS),.VDD(VDD),.Y(g15018),.A(I21374));
  NOT NOT1_5010(.VSS(VSS),.VDD(VDD),.Y(I21377),.A(g11821));
  NOT NOT1_5011(.VSS(VSS),.VDD(VDD),.Y(g15019),.A(I21377));
  NOT NOT1_5012(.VSS(VSS),.VDD(VDD),.Y(I21381),.A(g13157));
  NOT NOT1_5013(.VSS(VSS),.VDD(VDD),.Y(g15021),.A(I21381));
  NOT NOT1_5014(.VSS(VSS),.VDD(VDD),.Y(g15022),.A(g11781));
  NOT NOT1_5015(.VSS(VSS),.VDD(VDD),.Y(g15032),.A(g12027));
  NOT NOT1_5016(.VSS(VSS),.VDD(VDD),.Y(g15033),.A(g12030));
  NOT NOT1_5017(.VSS(VSS),.VDD(VDD),.Y(I21389),.A(g12883));
  NOT NOT1_5018(.VSS(VSS),.VDD(VDD),.Y(g15034),.A(I21389));
  NOT NOT1_5019(.VSS(VSS),.VDD(VDD),.Y(I21392),.A(g13020));
  NOT NOT1_5020(.VSS(VSS),.VDD(VDD),.Y(g15037),.A(I21392));
  NOT NOT1_5021(.VSS(VSS),.VDD(VDD),.Y(I21395),.A(g13034));
  NOT NOT1_5022(.VSS(VSS),.VDD(VDD),.Y(g15040),.A(I21395));
  NOT NOT1_5023(.VSS(VSS),.VDD(VDD),.Y(I21398),.A(g13021));
  NOT NOT1_5024(.VSS(VSS),.VDD(VDD),.Y(g15043),.A(I21398));
  NOT NOT1_5025(.VSS(VSS),.VDD(VDD),.Y(g15048),.A(g12045));
  NOT NOT1_5026(.VSS(VSS),.VDD(VDD),.Y(I21404),.A(g13037));
  NOT NOT1_5027(.VSS(VSS),.VDD(VDD),.Y(g15049),.A(I21404));
  NOT NOT1_5028(.VSS(VSS),.VDD(VDD),.Y(I21407),.A(g13039));
  NOT NOT1_5029(.VSS(VSS),.VDD(VDD),.Y(g15052),.A(I21407));
  NOT NOT1_5030(.VSS(VSS),.VDD(VDD),.Y(g15055),.A(g11952));
  NOT NOT1_5031(.VSS(VSS),.VDD(VDD),.Y(g15065),.A(g12291));
  NOT NOT1_5032(.VSS(VSS),.VDD(VDD),.Y(g15074),.A(g11962));
  NOT NOT1_5033(.VSS(VSS),.VDD(VDD),.Y(g15080),.A(g12305));
  NOT NOT1_5034(.VSS(VSS),.VDD(VDD),.Y(I21415),.A(g11854));
  NOT NOT1_5035(.VSS(VSS),.VDD(VDD),.Y(g15092),.A(I21415));
  NOT NOT1_5036(.VSS(VSS),.VDD(VDD),.Y(I21420),.A(g13166));
  NOT NOT1_5037(.VSS(VSS),.VDD(VDD),.Y(g15095),.A(I21420));
  NOT NOT1_5038(.VSS(VSS),.VDD(VDD),.Y(g15096),.A(g11800));
  NOT NOT1_5039(.VSS(VSS),.VDD(VDD),.Y(I21426),.A(g11661));
  NOT NOT1_5040(.VSS(VSS),.VDD(VDD),.Y(g15106),.A(I21426));
  NOT NOT1_5041(.VSS(VSS),.VDD(VDD),.Y(I21429),.A(g13027));
  NOT NOT1_5042(.VSS(VSS),.VDD(VDD),.Y(g15109),.A(I21429));
  NOT NOT1_5043(.VSS(VSS),.VDD(VDD),.Y(I21432),.A(g13044));
  NOT NOT1_5044(.VSS(VSS),.VDD(VDD),.Y(g15112),.A(I21432));
  NOT NOT1_5045(.VSS(VSS),.VDD(VDD),.Y(I21435),.A(g11662));
  NOT NOT1_5046(.VSS(VSS),.VDD(VDD),.Y(g15115),.A(I21435));
  NOT NOT1_5047(.VSS(VSS),.VDD(VDD),.Y(g15118),.A(g11807));
  NOT NOT1_5048(.VSS(VSS),.VDD(VDD),.Y(g15128),.A(g12091));
  NOT NOT1_5049(.VSS(VSS),.VDD(VDD),.Y(g15129),.A(g12094));
  NOT NOT1_5050(.VSS(VSS),.VDD(VDD),.Y(I21443),.A(g12923));
  NOT NOT1_5051(.VSS(VSS),.VDD(VDD),.Y(g15130),.A(I21443));
  NOT NOT1_5052(.VSS(VSS),.VDD(VDD),.Y(I21446),.A(g13029));
  NOT NOT1_5053(.VSS(VSS),.VDD(VDD),.Y(g15133),.A(I21446));
  NOT NOT1_5054(.VSS(VSS),.VDD(VDD),.Y(I21449),.A(g13047));
  NOT NOT1_5055(.VSS(VSS),.VDD(VDD),.Y(g15136),.A(I21449));
  NOT NOT1_5056(.VSS(VSS),.VDD(VDD),.Y(I21452),.A(g13030));
  NOT NOT1_5057(.VSS(VSS),.VDD(VDD),.Y(g15139),.A(I21452));
  NOT NOT1_5058(.VSS(VSS),.VDD(VDD),.Y(g15144),.A(g12109));
  NOT NOT1_5059(.VSS(VSS),.VDD(VDD),.Y(I21458),.A(g13050));
  NOT NOT1_5060(.VSS(VSS),.VDD(VDD),.Y(g15145),.A(I21458));
  NOT NOT1_5061(.VSS(VSS),.VDD(VDD),.Y(I21461),.A(g13052));
  NOT NOT1_5062(.VSS(VSS),.VDD(VDD),.Y(g15148),.A(I21461));
  NOT NOT1_5063(.VSS(VSS),.VDD(VDD),.Y(g15151),.A(g12005));
  NOT NOT1_5064(.VSS(VSS),.VDD(VDD),.Y(g15161),.A(g12327));
  NOT NOT1_5065(.VSS(VSS),.VDD(VDD),.Y(g15170),.A(g12125));
  NOT NOT1_5066(.VSS(VSS),.VDD(VDD),.Y(g15174),.A(g12136));
  NOT NOT1_5067(.VSS(VSS),.VDD(VDD),.Y(g15175),.A(g12139));
  NOT NOT1_5068(.VSS(VSS),.VDD(VDD),.Y(g15176),.A(g12142));
  NOT NOT1_5069(.VSS(VSS),.VDD(VDD),.Y(g15177),.A(g12339));
  NOT NOT1_5070(.VSS(VSS),.VDD(VDD),.Y(I21476),.A(g11672));
  NOT NOT1_5071(.VSS(VSS),.VDD(VDD),.Y(g15179),.A(I21476));
  NOT NOT1_5072(.VSS(VSS),.VDD(VDD),.Y(I21479),.A(g13035));
  NOT NOT1_5073(.VSS(VSS),.VDD(VDD),.Y(g15182),.A(I21479));
  NOT NOT1_5074(.VSS(VSS),.VDD(VDD),.Y(I21482),.A(g13058));
  NOT NOT1_5075(.VSS(VSS),.VDD(VDD),.Y(g15185),.A(I21482));
  NOT NOT1_5076(.VSS(VSS),.VDD(VDD),.Y(g15188),.A(g11833));
  NOT NOT1_5077(.VSS(VSS),.VDD(VDD),.Y(I21488),.A(g11673));
  NOT NOT1_5078(.VSS(VSS),.VDD(VDD),.Y(g15198),.A(I21488));
  NOT NOT1_5079(.VSS(VSS),.VDD(VDD),.Y(I21491),.A(g13038));
  NOT NOT1_5080(.VSS(VSS),.VDD(VDD),.Y(g15201),.A(I21491));
  NOT NOT1_5081(.VSS(VSS),.VDD(VDD),.Y(I21494),.A(g13061));
  NOT NOT1_5082(.VSS(VSS),.VDD(VDD),.Y(g15204),.A(I21494));
  NOT NOT1_5083(.VSS(VSS),.VDD(VDD),.Y(I21497),.A(g11674));
  NOT NOT1_5084(.VSS(VSS),.VDD(VDD),.Y(g15207),.A(I21497));
  NOT NOT1_5085(.VSS(VSS),.VDD(VDD),.Y(g15210),.A(g11840));
  NOT NOT1_5086(.VSS(VSS),.VDD(VDD),.Y(g15220),.A(g12163));
  NOT NOT1_5087(.VSS(VSS),.VDD(VDD),.Y(g15221),.A(g12166));
  NOT NOT1_5088(.VSS(VSS),.VDD(VDD),.Y(I21505),.A(g12952));
  NOT NOT1_5089(.VSS(VSS),.VDD(VDD),.Y(g15222),.A(I21505));
  NOT NOT1_5090(.VSS(VSS),.VDD(VDD),.Y(I21508),.A(g13040));
  NOT NOT1_5091(.VSS(VSS),.VDD(VDD),.Y(g15225),.A(I21508));
  NOT NOT1_5092(.VSS(VSS),.VDD(VDD),.Y(I21511),.A(g13064));
  NOT NOT1_5093(.VSS(VSS),.VDD(VDD),.Y(g15228),.A(I21511));
  NOT NOT1_5094(.VSS(VSS),.VDD(VDD),.Y(I21514),.A(g13041));
  NOT NOT1_5095(.VSS(VSS),.VDD(VDD),.Y(g15231),.A(I21514));
  NOT NOT1_5096(.VSS(VSS),.VDD(VDD),.Y(g15236),.A(g12181));
  NOT NOT1_5097(.VSS(VSS),.VDD(VDD),.Y(I21520),.A(g13067));
  NOT NOT1_5098(.VSS(VSS),.VDD(VDD),.Y(g15237),.A(I21520));
  NOT NOT1_5099(.VSS(VSS),.VDD(VDD),.Y(I21523),.A(g13069));
  NOT NOT1_5100(.VSS(VSS),.VDD(VDD),.Y(g15240),.A(I21523));
  NOT NOT1_5101(.VSS(VSS),.VDD(VDD),.Y(I21531),.A(g11683));
  NOT NOT1_5102(.VSS(VSS),.VDD(VDD),.Y(g15248),.A(I21531));
  NOT NOT1_5103(.VSS(VSS),.VDD(VDD),.Y(I21534),.A(g13045));
  NOT NOT1_5104(.VSS(VSS),.VDD(VDD),.Y(g15251),.A(I21534));
  NOT NOT1_5105(.VSS(VSS),.VDD(VDD),.Y(I21537),.A(g13071));
  NOT NOT1_5106(.VSS(VSS),.VDD(VDD),.Y(g15254),.A(I21537));
  NOT NOT1_5107(.VSS(VSS),.VDD(VDD),.Y(g15260),.A(g12198));
  NOT NOT1_5108(.VSS(VSS),.VDD(VDD),.Y(g15261),.A(g12201));
  NOT NOT1_5109(.VSS(VSS),.VDD(VDD),.Y(g15262),.A(g12204));
  NOT NOT1_5110(.VSS(VSS),.VDD(VDD),.Y(g15263),.A(g12369));
  NOT NOT1_5111(.VSS(VSS),.VDD(VDD),.Y(I21548),.A(g11684));
  NOT NOT1_5112(.VSS(VSS),.VDD(VDD),.Y(g15265),.A(I21548));
  NOT NOT1_5113(.VSS(VSS),.VDD(VDD),.Y(I21551),.A(g13048));
  NOT NOT1_5114(.VSS(VSS),.VDD(VDD),.Y(g15268),.A(I21551));
  NOT NOT1_5115(.VSS(VSS),.VDD(VDD),.Y(I21554),.A(g13074));
  NOT NOT1_5116(.VSS(VSS),.VDD(VDD),.Y(g15271),.A(I21554));
  NOT NOT1_5117(.VSS(VSS),.VDD(VDD),.Y(g15274),.A(g11875));
  NOT NOT1_5118(.VSS(VSS),.VDD(VDD),.Y(I21560),.A(g11685));
  NOT NOT1_5119(.VSS(VSS),.VDD(VDD),.Y(g15284),.A(I21560));
  NOT NOT1_5120(.VSS(VSS),.VDD(VDD),.Y(I21563),.A(g13051));
  NOT NOT1_5121(.VSS(VSS),.VDD(VDD),.Y(g15287),.A(I21563));
  NOT NOT1_5122(.VSS(VSS),.VDD(VDD),.Y(I21566),.A(g13077));
  NOT NOT1_5123(.VSS(VSS),.VDD(VDD),.Y(g15290),.A(I21566));
  NOT NOT1_5124(.VSS(VSS),.VDD(VDD),.Y(I21569),.A(g11686));
  NOT NOT1_5125(.VSS(VSS),.VDD(VDD),.Y(g15293),.A(I21569));
  NOT NOT1_5126(.VSS(VSS),.VDD(VDD),.Y(g15296),.A(g11882));
  NOT NOT1_5127(.VSS(VSS),.VDD(VDD),.Y(g15306),.A(g12225));
  NOT NOT1_5128(.VSS(VSS),.VDD(VDD),.Y(g15307),.A(g12228));
  NOT NOT1_5129(.VSS(VSS),.VDD(VDD),.Y(I21577),.A(g12981));
  NOT NOT1_5130(.VSS(VSS),.VDD(VDD),.Y(g15308),.A(I21577));
  NOT NOT1_5131(.VSS(VSS),.VDD(VDD),.Y(I21580),.A(g13053));
  NOT NOT1_5132(.VSS(VSS),.VDD(VDD),.Y(g15311),.A(I21580));
  NOT NOT1_5133(.VSS(VSS),.VDD(VDD),.Y(I21583),.A(g13080));
  NOT NOT1_5134(.VSS(VSS),.VDD(VDD),.Y(g15314),.A(I21583));
  NOT NOT1_5135(.VSS(VSS),.VDD(VDD),.Y(I21586),.A(g13054));
  NOT NOT1_5136(.VSS(VSS),.VDD(VDD),.Y(g15317),.A(I21586));
  NOT NOT1_5137(.VSS(VSS),.VDD(VDD),.Y(g15322),.A(g12239));
  NOT NOT1_5138(.VSS(VSS),.VDD(VDD),.Y(g15323),.A(g12242));
  NOT NOT1_5139(.VSS(VSS),.VDD(VDD),.Y(I21595),.A(g11691));
  NOT NOT1_5140(.VSS(VSS),.VDD(VDD),.Y(g15326),.A(I21595));
  NOT NOT1_5141(.VSS(VSS),.VDD(VDD),.Y(I21598),.A(g13059));
  NOT NOT1_5142(.VSS(VSS),.VDD(VDD),.Y(g15329),.A(I21598));
  NOT NOT1_5143(.VSS(VSS),.VDD(VDD),.Y(I21601),.A(g13087));
  NOT NOT1_5144(.VSS(VSS),.VDD(VDD),.Y(g15332),.A(I21601));
  NOT NOT1_5145(.VSS(VSS),.VDD(VDD),.Y(I21609),.A(g11692));
  NOT NOT1_5146(.VSS(VSS),.VDD(VDD),.Y(g15340),.A(I21609));
  NOT NOT1_5147(.VSS(VSS),.VDD(VDD),.Y(I21612),.A(g13062));
  NOT NOT1_5148(.VSS(VSS),.VDD(VDD),.Y(g15343),.A(I21612));
  NOT NOT1_5149(.VSS(VSS),.VDD(VDD),.Y(I21615),.A(g13090));
  NOT NOT1_5150(.VSS(VSS),.VDD(VDD),.Y(g15346),.A(I21615));
  NOT NOT1_5151(.VSS(VSS),.VDD(VDD),.Y(g15352),.A(g12253));
  NOT NOT1_5152(.VSS(VSS),.VDD(VDD),.Y(g15353),.A(g12256));
  NOT NOT1_5153(.VSS(VSS),.VDD(VDD),.Y(g15354),.A(g12259));
  NOT NOT1_5154(.VSS(VSS),.VDD(VDD),.Y(g15355),.A(g12388));
  NOT NOT1_5155(.VSS(VSS),.VDD(VDD),.Y(I21626),.A(g11693));
  NOT NOT1_5156(.VSS(VSS),.VDD(VDD),.Y(g15357),.A(I21626));
  NOT NOT1_5157(.VSS(VSS),.VDD(VDD),.Y(I21629),.A(g13065));
  NOT NOT1_5158(.VSS(VSS),.VDD(VDD),.Y(g15360),.A(I21629));
  NOT NOT1_5159(.VSS(VSS),.VDD(VDD),.Y(I21632),.A(g13093));
  NOT NOT1_5160(.VSS(VSS),.VDD(VDD),.Y(g15363),.A(I21632));
  NOT NOT1_5161(.VSS(VSS),.VDD(VDD),.Y(g15366),.A(g11917));
  NOT NOT1_5162(.VSS(VSS),.VDD(VDD),.Y(I21638),.A(g11694));
  NOT NOT1_5163(.VSS(VSS),.VDD(VDD),.Y(g15376),.A(I21638));
  NOT NOT1_5164(.VSS(VSS),.VDD(VDD),.Y(I21641),.A(g13068));
  NOT NOT1_5165(.VSS(VSS),.VDD(VDD),.Y(g15379),.A(I21641));
  NOT NOT1_5166(.VSS(VSS),.VDD(VDD),.Y(I21644),.A(g13096));
  NOT NOT1_5167(.VSS(VSS),.VDD(VDD),.Y(g15382),.A(I21644));
  NOT NOT1_5168(.VSS(VSS),.VDD(VDD),.Y(I21647),.A(g11695));
  NOT NOT1_5169(.VSS(VSS),.VDD(VDD),.Y(g15385),.A(I21647));
  NOT NOT1_5170(.VSS(VSS),.VDD(VDD),.Y(g15390),.A(g12279));
  NOT NOT1_5171(.VSS(VSS),.VDD(VDD),.Y(I21655),.A(g11696));
  NOT NOT1_5172(.VSS(VSS),.VDD(VDD),.Y(g15393),.A(I21655));
  NOT NOT1_5173(.VSS(VSS),.VDD(VDD),.Y(I21658),.A(g13072));
  NOT NOT1_5174(.VSS(VSS),.VDD(VDD),.Y(g15396),.A(I21658));
  NOT NOT1_5175(.VSS(VSS),.VDD(VDD),.Y(I21661),.A(g13098));
  NOT NOT1_5176(.VSS(VSS),.VDD(VDD),.Y(g15399),.A(I21661));
  NOT NOT1_5177(.VSS(VSS),.VDD(VDD),.Y(I21666),.A(g13100));
  NOT NOT1_5178(.VSS(VSS),.VDD(VDD),.Y(g15404),.A(I21666));
  NOT NOT1_5179(.VSS(VSS),.VDD(VDD),.Y(g15408),.A(g12282));
  NOT NOT1_5180(.VSS(VSS),.VDD(VDD),.Y(g15409),.A(g12285));
  NOT NOT1_5181(.VSS(VSS),.VDD(VDD),.Y(I21674),.A(g11698));
  NOT NOT1_5182(.VSS(VSS),.VDD(VDD),.Y(g15412),.A(I21674));
  NOT NOT1_5183(.VSS(VSS),.VDD(VDD),.Y(I21677),.A(g13075));
  NOT NOT1_5184(.VSS(VSS),.VDD(VDD),.Y(g15415),.A(I21677));
  NOT NOT1_5185(.VSS(VSS),.VDD(VDD),.Y(I21680),.A(g13102));
  NOT NOT1_5186(.VSS(VSS),.VDD(VDD),.Y(g15418),.A(I21680));
  NOT NOT1_5187(.VSS(VSS),.VDD(VDD),.Y(I21688),.A(g11699));
  NOT NOT1_5188(.VSS(VSS),.VDD(VDD),.Y(g15426),.A(I21688));
  NOT NOT1_5189(.VSS(VSS),.VDD(VDD),.Y(I21691),.A(g13078));
  NOT NOT1_5190(.VSS(VSS),.VDD(VDD),.Y(g15429),.A(I21691));
  NOT NOT1_5191(.VSS(VSS),.VDD(VDD),.Y(I21694),.A(g13105));
  NOT NOT1_5192(.VSS(VSS),.VDD(VDD),.Y(g15432),.A(I21694));
  NOT NOT1_5193(.VSS(VSS),.VDD(VDD),.Y(g15438),.A(g12296));
  NOT NOT1_5194(.VSS(VSS),.VDD(VDD),.Y(g15439),.A(g12299));
  NOT NOT1_5195(.VSS(VSS),.VDD(VDD),.Y(g15440),.A(g12302));
  NOT NOT1_5196(.VSS(VSS),.VDD(VDD),.Y(g15441),.A(g12418));
  NOT NOT1_5197(.VSS(VSS),.VDD(VDD),.Y(I21705),.A(g11700));
  NOT NOT1_5198(.VSS(VSS),.VDD(VDD),.Y(g15443),.A(I21705));
  NOT NOT1_5199(.VSS(VSS),.VDD(VDD),.Y(I21708),.A(g13081));
  NOT NOT1_5200(.VSS(VSS),.VDD(VDD),.Y(g15446),.A(I21708));
  NOT NOT1_5201(.VSS(VSS),.VDD(VDD),.Y(I21711),.A(g13108));
  NOT NOT1_5202(.VSS(VSS),.VDD(VDD),.Y(g15449),.A(I21711));
  NOT NOT1_5203(.VSS(VSS),.VDD(VDD),.Y(g15458),.A(g12312));
  NOT NOT1_5204(.VSS(VSS),.VDD(VDD),.Y(I21720),.A(g11701));
  NOT NOT1_5205(.VSS(VSS),.VDD(VDD),.Y(g15461),.A(I21720));
  NOT NOT1_5206(.VSS(VSS),.VDD(VDD),.Y(I21723),.A(g13088));
  NOT NOT1_5207(.VSS(VSS),.VDD(VDD),.Y(g15464),.A(I21723));
  NOT NOT1_5208(.VSS(VSS),.VDD(VDD),.Y(I21726),.A(g13112));
  NOT NOT1_5209(.VSS(VSS),.VDD(VDD),.Y(g15467),.A(I21726));
  NOT NOT1_5210(.VSS(VSS),.VDD(VDD),.Y(I21730),.A(g13089));
  NOT NOT1_5211(.VSS(VSS),.VDD(VDD),.Y(g15471),.A(I21730));
  NOT NOT1_5212(.VSS(VSS),.VDD(VDD),.Y(g15474),.A(g12315));
  NOT NOT1_5213(.VSS(VSS),.VDD(VDD),.Y(I21736),.A(g11702));
  NOT NOT1_5214(.VSS(VSS),.VDD(VDD),.Y(g15477),.A(I21736));
  NOT NOT1_5215(.VSS(VSS),.VDD(VDD),.Y(I21739),.A(g13091));
  NOT NOT1_5216(.VSS(VSS),.VDD(VDD),.Y(g15480),.A(I21739));
  NOT NOT1_5217(.VSS(VSS),.VDD(VDD),.Y(I21742),.A(g13114));
  NOT NOT1_5218(.VSS(VSS),.VDD(VDD),.Y(g15483),.A(I21742));
  NOT NOT1_5219(.VSS(VSS),.VDD(VDD),.Y(I21747),.A(g13116));
  NOT NOT1_5220(.VSS(VSS),.VDD(VDD),.Y(g15488),.A(I21747));
  NOT NOT1_5221(.VSS(VSS),.VDD(VDD),.Y(g15492),.A(g12318));
  NOT NOT1_5222(.VSS(VSS),.VDD(VDD),.Y(g15493),.A(g12321));
  NOT NOT1_5223(.VSS(VSS),.VDD(VDD),.Y(I21755),.A(g11704));
  NOT NOT1_5224(.VSS(VSS),.VDD(VDD),.Y(g15496),.A(I21755));
  NOT NOT1_5225(.VSS(VSS),.VDD(VDD),.Y(I21758),.A(g13094));
  NOT NOT1_5226(.VSS(VSS),.VDD(VDD),.Y(g15499),.A(I21758));
  NOT NOT1_5227(.VSS(VSS),.VDD(VDD),.Y(I21761),.A(g13118));
  NOT NOT1_5228(.VSS(VSS),.VDD(VDD),.Y(g15502),.A(I21761));
  NOT NOT1_5229(.VSS(VSS),.VDD(VDD),.Y(I21769),.A(g11705));
  NOT NOT1_5230(.VSS(VSS),.VDD(VDD),.Y(g15510),.A(I21769));
  NOT NOT1_5231(.VSS(VSS),.VDD(VDD),.Y(I21772),.A(g13097));
  NOT NOT1_5232(.VSS(VSS),.VDD(VDD),.Y(g15513),.A(I21772));
  NOT NOT1_5233(.VSS(VSS),.VDD(VDD),.Y(I21775),.A(g13121));
  NOT NOT1_5234(.VSS(VSS),.VDD(VDD),.Y(g15516),.A(I21775));
  NOT NOT1_5235(.VSS(VSS),.VDD(VDD),.Y(I21780),.A(g13305));
  NOT NOT1_5236(.VSS(VSS),.VDD(VDD),.Y(g15521),.A(I21780));
  NOT NOT1_5237(.VSS(VSS),.VDD(VDD),.Y(g15524),.A(g12333));
  NOT NOT1_5238(.VSS(VSS),.VDD(VDD),.Y(g15525),.A(g12336));
  NOT NOT1_5239(.VSS(VSS),.VDD(VDD),.Y(I21787),.A(g11707));
  NOT NOT1_5240(.VSS(VSS),.VDD(VDD),.Y(g15528),.A(I21787));
  NOT NOT1_5241(.VSS(VSS),.VDD(VDD),.Y(I21790),.A(g13099));
  NOT NOT1_5242(.VSS(VSS),.VDD(VDD),.Y(g15531),.A(I21790));
  NOT NOT1_5243(.VSS(VSS),.VDD(VDD),.Y(I21793),.A(g13123));
  NOT NOT1_5244(.VSS(VSS),.VDD(VDD),.Y(g15534),.A(I21793));
  NOT NOT1_5245(.VSS(VSS),.VDD(VDD),.Y(I21796),.A(g11708));
  NOT NOT1_5246(.VSS(VSS),.VDD(VDD),.Y(g15537),.A(I21796));
  NOT NOT1_5247(.VSS(VSS),.VDD(VDD),.Y(g15544),.A(g12340));
  NOT NOT1_5248(.VSS(VSS),.VDD(VDD),.Y(I21803),.A(g11709));
  NOT NOT1_5249(.VSS(VSS),.VDD(VDD),.Y(g15547),.A(I21803));
  NOT NOT1_5250(.VSS(VSS),.VDD(VDD),.Y(I21806),.A(g13103));
  NOT NOT1_5251(.VSS(VSS),.VDD(VDD),.Y(g15550),.A(I21806));
  NOT NOT1_5252(.VSS(VSS),.VDD(VDD),.Y(I21809),.A(g13125));
  NOT NOT1_5253(.VSS(VSS),.VDD(VDD),.Y(g15553),.A(I21809));
  NOT NOT1_5254(.VSS(VSS),.VDD(VDD),.Y(I21813),.A(g13104));
  NOT NOT1_5255(.VSS(VSS),.VDD(VDD),.Y(g15557),.A(I21813));
  NOT NOT1_5256(.VSS(VSS),.VDD(VDD),.Y(g15560),.A(g12343));
  NOT NOT1_5257(.VSS(VSS),.VDD(VDD),.Y(I21819),.A(g11710));
  NOT NOT1_5258(.VSS(VSS),.VDD(VDD),.Y(g15563),.A(I21819));
  NOT NOT1_5259(.VSS(VSS),.VDD(VDD),.Y(I21822),.A(g13106));
  NOT NOT1_5260(.VSS(VSS),.VDD(VDD),.Y(g15566),.A(I21822));
  NOT NOT1_5261(.VSS(VSS),.VDD(VDD),.Y(I21825),.A(g13127));
  NOT NOT1_5262(.VSS(VSS),.VDD(VDD),.Y(g15569),.A(I21825));
  NOT NOT1_5263(.VSS(VSS),.VDD(VDD),.Y(I21830),.A(g13129));
  NOT NOT1_5264(.VSS(VSS),.VDD(VDD),.Y(g15574),.A(I21830));
  NOT NOT1_5265(.VSS(VSS),.VDD(VDD),.Y(g15578),.A(g12346));
  NOT NOT1_5266(.VSS(VSS),.VDD(VDD),.Y(g15579),.A(g12349));
  NOT NOT1_5267(.VSS(VSS),.VDD(VDD),.Y(I21838),.A(g11712));
  NOT NOT1_5268(.VSS(VSS),.VDD(VDD),.Y(g15582),.A(I21838));
  NOT NOT1_5269(.VSS(VSS),.VDD(VDD),.Y(I21841),.A(g13109));
  NOT NOT1_5270(.VSS(VSS),.VDD(VDD),.Y(g15585),.A(I21841));
  NOT NOT1_5271(.VSS(VSS),.VDD(VDD),.Y(I21844),.A(g13131));
  NOT NOT1_5272(.VSS(VSS),.VDD(VDD),.Y(g15588),.A(I21844));
  NOT NOT1_5273(.VSS(VSS),.VDD(VDD),.Y(I21852),.A(g11716));
  NOT NOT1_5274(.VSS(VSS),.VDD(VDD),.Y(g15596),.A(I21852));
  NOT NOT1_5275(.VSS(VSS),.VDD(VDD),.Y(I21855),.A(g13113));
  NOT NOT1_5276(.VSS(VSS),.VDD(VDD),.Y(g15599),.A(I21855));
  NOT NOT1_5277(.VSS(VSS),.VDD(VDD),.Y(g15602),.A(g12363));
  NOT NOT1_5278(.VSS(VSS),.VDD(VDD),.Y(g15603),.A(g12366));
  NOT NOT1_5279(.VSS(VSS),.VDD(VDD),.Y(I21862),.A(g11717));
  NOT NOT1_5280(.VSS(VSS),.VDD(VDD),.Y(g15606),.A(I21862));
  NOT NOT1_5281(.VSS(VSS),.VDD(VDD),.Y(I21865),.A(g13115));
  NOT NOT1_5282(.VSS(VSS),.VDD(VDD),.Y(g15609),.A(I21865));
  NOT NOT1_5283(.VSS(VSS),.VDD(VDD),.Y(I21868),.A(g13134));
  NOT NOT1_5284(.VSS(VSS),.VDD(VDD),.Y(g15612),.A(I21868));
  NOT NOT1_5285(.VSS(VSS),.VDD(VDD),.Y(I21871),.A(g11718));
  NOT NOT1_5286(.VSS(VSS),.VDD(VDD),.Y(g15615),.A(I21871));
  NOT NOT1_5287(.VSS(VSS),.VDD(VDD),.Y(g15622),.A(g12370));
  NOT NOT1_5288(.VSS(VSS),.VDD(VDD),.Y(I21878),.A(g11719));
  NOT NOT1_5289(.VSS(VSS),.VDD(VDD),.Y(g15625),.A(I21878));
  NOT NOT1_5290(.VSS(VSS),.VDD(VDD),.Y(I21881),.A(g13119));
  NOT NOT1_5291(.VSS(VSS),.VDD(VDD),.Y(g15628),.A(I21881));
  NOT NOT1_5292(.VSS(VSS),.VDD(VDD),.Y(I21884),.A(g13136));
  NOT NOT1_5293(.VSS(VSS),.VDD(VDD),.Y(g15631),.A(I21884));
  NOT NOT1_5294(.VSS(VSS),.VDD(VDD),.Y(I21888),.A(g13120));
  NOT NOT1_5295(.VSS(VSS),.VDD(VDD),.Y(g15635),.A(I21888));
  NOT NOT1_5296(.VSS(VSS),.VDD(VDD),.Y(g15638),.A(g12373));
  NOT NOT1_5297(.VSS(VSS),.VDD(VDD),.Y(I21894),.A(g11720));
  NOT NOT1_5298(.VSS(VSS),.VDD(VDD),.Y(g15641),.A(I21894));
  NOT NOT1_5299(.VSS(VSS),.VDD(VDD),.Y(I21897),.A(g13122));
  NOT NOT1_5300(.VSS(VSS),.VDD(VDD),.Y(g15644),.A(I21897));
  NOT NOT1_5301(.VSS(VSS),.VDD(VDD),.Y(I21900),.A(g13138));
  NOT NOT1_5302(.VSS(VSS),.VDD(VDD),.Y(g15647),.A(I21900));
  NOT NOT1_5303(.VSS(VSS),.VDD(VDD),.Y(I21905),.A(g13140));
  NOT NOT1_5304(.VSS(VSS),.VDD(VDD),.Y(g15652),.A(I21905));
  NOT NOT1_5305(.VSS(VSS),.VDD(VDD),.Y(I21908),.A(g13082));
  NOT NOT1_5306(.VSS(VSS),.VDD(VDD),.Y(g15655),.A(I21908));
  NOT NOT1_5307(.VSS(VSS),.VDD(VDD),.Y(g15659),.A(g11706));
  NOT NOT1_5308(.VSS(VSS),.VDD(VDD),.Y(g15665),.A(g12379));
  NOT NOT1_5309(.VSS(VSS),.VDD(VDD),.Y(I21918),.A(g11721));
  NOT NOT1_5310(.VSS(VSS),.VDD(VDD),.Y(g15667),.A(I21918));
  NOT NOT1_5311(.VSS(VSS),.VDD(VDD),.Y(I21923),.A(g11722));
  NOT NOT1_5312(.VSS(VSS),.VDD(VDD),.Y(g15672),.A(I21923));
  NOT NOT1_5313(.VSS(VSS),.VDD(VDD),.Y(I21926),.A(g13126));
  NOT NOT1_5314(.VSS(VSS),.VDD(VDD),.Y(g15675),.A(I21926));
  NOT NOT1_5315(.VSS(VSS),.VDD(VDD),.Y(g15678),.A(g12382));
  NOT NOT1_5316(.VSS(VSS),.VDD(VDD),.Y(g15679),.A(g12385));
  NOT NOT1_5317(.VSS(VSS),.VDD(VDD),.Y(I21933),.A(g11723));
  NOT NOT1_5318(.VSS(VSS),.VDD(VDD),.Y(g15682),.A(I21933));
  NOT NOT1_5319(.VSS(VSS),.VDD(VDD),.Y(I21936),.A(g13128));
  NOT NOT1_5320(.VSS(VSS),.VDD(VDD),.Y(g15685),.A(I21936));
  NOT NOT1_5321(.VSS(VSS),.VDD(VDD),.Y(I21939),.A(g13142));
  NOT NOT1_5322(.VSS(VSS),.VDD(VDD),.Y(g15688),.A(I21939));
  NOT NOT1_5323(.VSS(VSS),.VDD(VDD),.Y(I21942),.A(g11724));
  NOT NOT1_5324(.VSS(VSS),.VDD(VDD),.Y(g15691),.A(I21942));
  NOT NOT1_5325(.VSS(VSS),.VDD(VDD),.Y(g15698),.A(g12389));
  NOT NOT1_5326(.VSS(VSS),.VDD(VDD),.Y(I21949),.A(g11725));
  NOT NOT1_5327(.VSS(VSS),.VDD(VDD),.Y(g15701),.A(I21949));
  NOT NOT1_5328(.VSS(VSS),.VDD(VDD),.Y(I21952),.A(g13132));
  NOT NOT1_5329(.VSS(VSS),.VDD(VDD),.Y(g15704),.A(I21952));
  NOT NOT1_5330(.VSS(VSS),.VDD(VDD),.Y(I21955),.A(g13144));
  NOT NOT1_5331(.VSS(VSS),.VDD(VDD),.Y(g15707),.A(I21955));
  NOT NOT1_5332(.VSS(VSS),.VDD(VDD),.Y(I21959),.A(g13133));
  NOT NOT1_5333(.VSS(VSS),.VDD(VDD),.Y(g15711),.A(I21959));
  NOT NOT1_5334(.VSS(VSS),.VDD(VDD),.Y(I21962),.A(g13004));
  NOT NOT1_5335(.VSS(VSS),.VDD(VDD),.Y(g15714),.A(I21962));
  NOT NOT1_5336(.VSS(VSS),.VDD(VDD),.Y(g15722),.A(g13011));
  NOT NOT1_5337(.VSS(VSS),.VDD(VDD),.Y(g15724),.A(g12409));
  NOT NOT1_5338(.VSS(VSS),.VDD(VDD),.Y(I21974),.A(g11726));
  NOT NOT1_5339(.VSS(VSS),.VDD(VDD),.Y(g15726),.A(I21974));
  NOT NOT1_5340(.VSS(VSS),.VDD(VDD),.Y(I21979),.A(g11727));
  NOT NOT1_5341(.VSS(VSS),.VDD(VDD),.Y(g15731),.A(I21979));
  NOT NOT1_5342(.VSS(VSS),.VDD(VDD),.Y(I21982),.A(g13137));
  NOT NOT1_5343(.VSS(VSS),.VDD(VDD),.Y(g15734),.A(I21982));
  NOT NOT1_5344(.VSS(VSS),.VDD(VDD),.Y(g15737),.A(g12412));
  NOT NOT1_5345(.VSS(VSS),.VDD(VDD),.Y(g15738),.A(g12415));
  NOT NOT1_5346(.VSS(VSS),.VDD(VDD),.Y(I21989),.A(g11728));
  NOT NOT1_5347(.VSS(VSS),.VDD(VDD),.Y(g15741),.A(I21989));
  NOT NOT1_5348(.VSS(VSS),.VDD(VDD),.Y(I21992),.A(g13139));
  NOT NOT1_5349(.VSS(VSS),.VDD(VDD),.Y(g15744),.A(I21992));
  NOT NOT1_5350(.VSS(VSS),.VDD(VDD),.Y(I21995),.A(g13146));
  NOT NOT1_5351(.VSS(VSS),.VDD(VDD),.Y(g15747),.A(I21995));
  NOT NOT1_5352(.VSS(VSS),.VDD(VDD),.Y(I21998),.A(g11729));
  NOT NOT1_5353(.VSS(VSS),.VDD(VDD),.Y(g15750),.A(I21998));
  NOT NOT1_5354(.VSS(VSS),.VDD(VDD),.Y(g15762),.A(g13011));
  NOT NOT1_5355(.VSS(VSS),.VDD(VDD),.Y(g15764),.A(g12421));
  NOT NOT1_5356(.VSS(VSS),.VDD(VDD),.Y(I22014),.A(g11730));
  NOT NOT1_5357(.VSS(VSS),.VDD(VDD),.Y(g15766),.A(I22014));
  NOT NOT1_5358(.VSS(VSS),.VDD(VDD),.Y(I22019),.A(g11731));
  NOT NOT1_5359(.VSS(VSS),.VDD(VDD),.Y(g15771),.A(I22019));
  NOT NOT1_5360(.VSS(VSS),.VDD(VDD),.Y(I22022),.A(g13145));
  NOT NOT1_5361(.VSS(VSS),.VDD(VDD),.Y(g15774),.A(I22022));
  NOT NOT1_5362(.VSS(VSS),.VDD(VDD),.Y(I22025),.A(g11617));
  NOT NOT1_5363(.VSS(VSS),.VDD(VDD),.Y(g15777),.A(I22025));
  NOT NOT1_5364(.VSS(VSS),.VDD(VDD),.Y(g15790),.A(g13011));
  NOT NOT1_5365(.VSS(VSS),.VDD(VDD),.Y(g15792),.A(g12426));
  NOT NOT1_5366(.VSS(VSS),.VDD(VDD),.Y(I22044),.A(g11733));
  NOT NOT1_5367(.VSS(VSS),.VDD(VDD),.Y(g15794),.A(I22044));
  NOT NOT1_5368(.VSS(VSS),.VDD(VDD),.Y(g15800),.A(g12909));
  NOT NOT1_5369(.VSS(VSS),.VDD(VDD),.Y(g15813),.A(g13011));
  NOT NOT1_5370(.VSS(VSS),.VDD(VDD),.Y(g15859),.A(g13378));
  NOT NOT1_5371(.VSS(VSS),.VDD(VDD),.Y(I22120),.A(g12909));
  NOT NOT1_5372(.VSS(VSS),.VDD(VDD),.Y(g15876),.A(I22120));
  NOT NOT1_5373(.VSS(VSS),.VDD(VDD),.Y(g15880),.A(g11624));
  NOT NOT1_5374(.VSS(VSS),.VDD(VDD),.Y(g15890),.A(g11600));
  NOT NOT1_5375(.VSS(VSS),.VDD(VDD),.Y(g15904),.A(g11644));
  NOT NOT1_5376(.VSS(VSS),.VDD(VDD),.Y(g15913),.A(g11647));
  NOT NOT1_5377(.VSS(VSS),.VDD(VDD),.Y(g15923),.A(g11630));
  NOT NOT1_5378(.VSS(VSS),.VDD(VDD),.Y(g15933),.A(g11663));
  NOT NOT1_5379(.VSS(VSS),.VDD(VDD),.Y(g15942),.A(g11666));
  NOT NOT1_5380(.VSS(VSS),.VDD(VDD),.Y(g15952),.A(g11653));
  NOT NOT1_5381(.VSS(VSS),.VDD(VDD),.Y(g15962),.A(g11675));
  NOT NOT1_5382(.VSS(VSS),.VDD(VDD),.Y(g15971),.A(g11678));
  NOT NOT1_5383(.VSS(VSS),.VDD(VDD),.Y(g15981),.A(g11687));
  NOT NOT1_5384(.VSS(VSS),.VDD(VDD),.Y(I22163),.A(g12433));
  NOT NOT1_5385(.VSS(VSS),.VDD(VDD),.Y(g15989),.A(I22163));
  NOT NOT1_5386(.VSS(VSS),.VDD(VDD),.Y(g15991),.A(g12548));
  NOT NOT1_5387(.VSS(VSS),.VDD(VDD),.Y(g15994),.A(g12555));
  NOT NOT1_5388(.VSS(VSS),.VDD(VDD),.Y(g15997),.A(g12561));
  NOT NOT1_5389(.VSS(VSS),.VDD(VDD),.Y(g16001),.A(g12601));
  NOT NOT1_5390(.VSS(VSS),.VDD(VDD),.Y(g16002),.A(g12604));
  NOT NOT1_5391(.VSS(VSS),.VDD(VDD),.Y(g16005),.A(g12608));
  NOT NOT1_5392(.VSS(VSS),.VDD(VDD),.Y(g16007),.A(g12647));
  NOT NOT1_5393(.VSS(VSS),.VDD(VDD),.Y(g16011),.A(g12651));
  NOT NOT1_5394(.VSS(VSS),.VDD(VDD),.Y(g16012),.A(g12654));
  NOT NOT1_5395(.VSS(VSS),.VDD(VDD),.Y(g16013),.A(g12692));
  NOT NOT1_5396(.VSS(VSS),.VDD(VDD),.Y(g16014),.A(g12695));
  NOT NOT1_5397(.VSS(VSS),.VDD(VDD),.Y(g16023),.A(g12699));
  NOT NOT1_5398(.VSS(VSS),.VDD(VDD),.Y(g16024),.A(g12702));
  NOT NOT1_5399(.VSS(VSS),.VDD(VDD),.Y(g16025),.A(g12705));
  NOT NOT1_5400(.VSS(VSS),.VDD(VDD),.Y(g16026),.A(g12708));
  NOT NOT1_5401(.VSS(VSS),.VDD(VDD),.Y(g16027),.A(g12744));
  NOT NOT1_5402(.VSS(VSS),.VDD(VDD),.Y(g16034),.A(g12749));
  NOT NOT1_5403(.VSS(VSS),.VDD(VDD),.Y(g16035),.A(g12752));
  NOT NOT1_5404(.VSS(VSS),.VDD(VDD),.Y(g16039),.A(g12756));
  NOT NOT1_5405(.VSS(VSS),.VDD(VDD),.Y(g16040),.A(g12759));
  NOT NOT1_5406(.VSS(VSS),.VDD(VDD),.Y(g16041),.A(g12762));
  NOT NOT1_5407(.VSS(VSS),.VDD(VDD),.Y(g16042),.A(g12765));
  NOT NOT1_5408(.VSS(VSS),.VDD(VDD),.Y(g16043),.A(g12769));
  NOT NOT1_5409(.VSS(VSS),.VDD(VDD),.Y(g16044),.A(g12772));
  NOT NOT1_5410(.VSS(VSS),.VDD(VDD),.Y(g16054),.A(g12783));
  NOT NOT1_5411(.VSS(VSS),.VDD(VDD),.Y(g16055),.A(g12786));
  NOT NOT1_5412(.VSS(VSS),.VDD(VDD),.Y(g16056),.A(g12791));
  NOT NOT1_5413(.VSS(VSS),.VDD(VDD),.Y(g16057),.A(g12794));
  NOT NOT1_5414(.VSS(VSS),.VDD(VDD),.Y(g16061),.A(g12798));
  NOT NOT1_5415(.VSS(VSS),.VDD(VDD),.Y(g16062),.A(g12801));
  NOT NOT1_5416(.VSS(VSS),.VDD(VDD),.Y(g16063),.A(g12804));
  NOT NOT1_5417(.VSS(VSS),.VDD(VDD),.Y(g16064),.A(g12808));
  NOT NOT1_5418(.VSS(VSS),.VDD(VDD),.Y(g16065),.A(g12811));
  NOT NOT1_5419(.VSS(VSS),.VDD(VDD),.Y(g16075),.A(g11861));
  NOT NOT1_5420(.VSS(VSS),.VDD(VDD),.Y(g16088),.A(g12816));
  NOT NOT1_5421(.VSS(VSS),.VDD(VDD),.Y(g16090),.A(g12822));
  NOT NOT1_5422(.VSS(VSS),.VDD(VDD),.Y(g16091),.A(g12825));
  NOT NOT1_5423(.VSS(VSS),.VDD(VDD),.Y(g16092),.A(g12830));
  NOT NOT1_5424(.VSS(VSS),.VDD(VDD),.Y(g16093),.A(g12833));
  NOT NOT1_5425(.VSS(VSS),.VDD(VDD),.Y(g16097),.A(g12837));
  NOT NOT1_5426(.VSS(VSS),.VDD(VDD),.Y(g16098),.A(g12840));
  NOT NOT1_5427(.VSS(VSS),.VDD(VDD),.Y(g16099),.A(g12844));
  NOT NOT1_5428(.VSS(VSS),.VDD(VDD),.Y(g16113),.A(g11903));
  NOT NOT1_5429(.VSS(VSS),.VDD(VDD),.Y(g16126),.A(g12854));
  NOT NOT1_5430(.VSS(VSS),.VDD(VDD),.Y(g16128),.A(g12860));
  NOT NOT1_5431(.VSS(VSS),.VDD(VDD),.Y(g16129),.A(g12863));
  NOT NOT1_5432(.VSS(VSS),.VDD(VDD),.Y(g16130),.A(g12868));
  NOT NOT1_5433(.VSS(VSS),.VDD(VDD),.Y(g16131),.A(g12871));
  NOT NOT1_5434(.VSS(VSS),.VDD(VDD),.Y(g16142),.A(g13057));
  NOT NOT1_5435(.VSS(VSS),.VDD(VDD),.Y(g16154),.A(g12194));
  NOT NOT1_5436(.VSS(VSS),.VDD(VDD),.Y(g16164),.A(g11953));
  NOT NOT1_5437(.VSS(VSS),.VDD(VDD),.Y(g16177),.A(g12895));
  NOT NOT1_5438(.VSS(VSS),.VDD(VDD),.Y(g16179),.A(g12901));
  NOT NOT1_5439(.VSS(VSS),.VDD(VDD),.Y(g16180),.A(g12904));
  NOT NOT1_5440(.VSS(VSS),.VDD(VDD),.Y(g16189),.A(g13043));
  NOT NOT1_5441(.VSS(VSS),.VDD(VDD),.Y(g16201),.A(g13073));
  NOT NOT1_5442(.VSS(VSS),.VDD(VDD),.Y(g16213),.A(g12249));
  NOT NOT1_5443(.VSS(VSS),.VDD(VDD),.Y(g16223),.A(g12006));
  NOT NOT1_5444(.VSS(VSS),.VDD(VDD),.Y(g16236),.A(g12935));
  NOT NOT1_5445(.VSS(VSS),.VDD(VDD),.Y(g16243),.A(g13033));
  NOT NOT1_5446(.VSS(VSS),.VDD(VDD),.Y(g16254),.A(g13060));
  NOT NOT1_5447(.VSS(VSS),.VDD(VDD),.Y(g16266),.A(g13092));
  NOT NOT1_5448(.VSS(VSS),.VDD(VDD),.Y(g16278),.A(g12292));
  NOT NOT1_5449(.VSS(VSS),.VDD(VDD),.Y(g16287),.A(g12962));
  NOT NOT1_5450(.VSS(VSS),.VDD(VDD),.Y(g16293),.A(g13025));
  NOT NOT1_5451(.VSS(VSS),.VDD(VDD),.Y(I22382),.A(g520));
  NOT NOT1_5452(.VSS(VSS),.VDD(VDD),.Y(g16297),.A(I22382));
  NOT NOT1_5453(.VSS(VSS),.VDD(VDD),.Y(g16302),.A(g13046));
  NOT NOT1_5454(.VSS(VSS),.VDD(VDD),.Y(g16313),.A(g13076));
  NOT NOT1_5455(.VSS(VSS),.VDD(VDD),.Y(g16325),.A(g13107));
  NOT NOT1_5456(.VSS(VSS),.VDD(VDD),.Y(g16337),.A(g12328));
  NOT NOT1_5457(.VSS(VSS),.VDD(VDD),.Y(g16351),.A(g13036));
  NOT NOT1_5458(.VSS(VSS),.VDD(VDD),.Y(I22414),.A(g1206));
  NOT NOT1_5459(.VSS(VSS),.VDD(VDD),.Y(g16355),.A(I22414));
  NOT NOT1_5460(.VSS(VSS),.VDD(VDD),.Y(g16360),.A(g13063));
  NOT NOT1_5461(.VSS(VSS),.VDD(VDD),.Y(g16371),.A(g13095));
  NOT NOT1_5462(.VSS(VSS),.VDD(VDD),.Y(g16395),.A(g13049));
  NOT NOT1_5463(.VSS(VSS),.VDD(VDD),.Y(I22444),.A(g1900));
  NOT NOT1_5464(.VSS(VSS),.VDD(VDD),.Y(g16399),.A(I22444));
  NOT NOT1_5465(.VSS(VSS),.VDD(VDD),.Y(g16404),.A(g13079));
  NOT NOT1_5466(.VSS(VSS),.VDD(VDD),.Y(g16433),.A(g13066));
  NOT NOT1_5467(.VSS(VSS),.VDD(VDD),.Y(I22475),.A(g2594));
  NOT NOT1_5468(.VSS(VSS),.VDD(VDD),.Y(g16437),.A(I22475));
  NOT NOT1_5469(.VSS(VSS),.VDD(VDD),.Y(g16466),.A(g12017));
  NOT NOT1_5470(.VSS(VSS),.VDD(VDD),.Y(I22503),.A(g13598));
  NOT NOT1_5471(.VSS(VSS),.VDD(VDD),.Y(g16467),.A(I22503));
  NOT NOT1_5472(.VSS(VSS),.VDD(VDD),.Y(I22506),.A(g13624));
  NOT NOT1_5473(.VSS(VSS),.VDD(VDD),.Y(g16468),.A(I22506));
  NOT NOT1_5474(.VSS(VSS),.VDD(VDD),.Y(I22509),.A(g13610));
  NOT NOT1_5475(.VSS(VSS),.VDD(VDD),.Y(g16469),.A(I22509));
  NOT NOT1_5476(.VSS(VSS),.VDD(VDD),.Y(I22512),.A(g13635));
  NOT NOT1_5477(.VSS(VSS),.VDD(VDD),.Y(g16470),.A(I22512));
  NOT NOT1_5478(.VSS(VSS),.VDD(VDD),.Y(I22515),.A(g13620));
  NOT NOT1_5479(.VSS(VSS),.VDD(VDD),.Y(g16471),.A(I22515));
  NOT NOT1_5480(.VSS(VSS),.VDD(VDD),.Y(I22518),.A(g13647));
  NOT NOT1_5481(.VSS(VSS),.VDD(VDD),.Y(g16472),.A(I22518));
  NOT NOT1_5482(.VSS(VSS),.VDD(VDD),.Y(I22521),.A(g13632));
  NOT NOT1_5483(.VSS(VSS),.VDD(VDD),.Y(g16473),.A(I22521));
  NOT NOT1_5484(.VSS(VSS),.VDD(VDD),.Y(I22524),.A(g13673));
  NOT NOT1_5485(.VSS(VSS),.VDD(VDD),.Y(g16474),.A(I22524));
  NOT NOT1_5486(.VSS(VSS),.VDD(VDD),.Y(I22527),.A(g13469));
  NOT NOT1_5487(.VSS(VSS),.VDD(VDD),.Y(g16475),.A(I22527));
  NOT NOT1_5488(.VSS(VSS),.VDD(VDD),.Y(I22530),.A(g14774));
  NOT NOT1_5489(.VSS(VSS),.VDD(VDD),.Y(g16476),.A(I22530));
  NOT NOT1_5490(.VSS(VSS),.VDD(VDD),.Y(I22533),.A(g14795));
  NOT NOT1_5491(.VSS(VSS),.VDD(VDD),.Y(g16477),.A(I22533));
  NOT NOT1_5492(.VSS(VSS),.VDD(VDD),.Y(I22536),.A(g14829));
  NOT NOT1_5493(.VSS(VSS),.VDD(VDD),.Y(g16478),.A(I22536));
  NOT NOT1_5494(.VSS(VSS),.VDD(VDD),.Y(I22539),.A(g14882));
  NOT NOT1_5495(.VSS(VSS),.VDD(VDD),.Y(g16479),.A(I22539));
  NOT NOT1_5496(.VSS(VSS),.VDD(VDD),.Y(I22542),.A(g14954));
  NOT NOT1_5497(.VSS(VSS),.VDD(VDD),.Y(g16480),.A(I22542));
  NOT NOT1_5498(.VSS(VSS),.VDD(VDD),.Y(I22545),.A(g15018));
  NOT NOT1_5499(.VSS(VSS),.VDD(VDD),.Y(g16481),.A(I22545));
  NOT NOT1_5500(.VSS(VSS),.VDD(VDD),.Y(I22548),.A(g14718));
  NOT NOT1_5501(.VSS(VSS),.VDD(VDD),.Y(g16482),.A(I22548));
  NOT NOT1_5502(.VSS(VSS),.VDD(VDD),.Y(I22551),.A(g14745));
  NOT NOT1_5503(.VSS(VSS),.VDD(VDD),.Y(g16483),.A(I22551));
  NOT NOT1_5504(.VSS(VSS),.VDD(VDD),.Y(I22554),.A(g14765));
  NOT NOT1_5505(.VSS(VSS),.VDD(VDD),.Y(g16484),.A(I22554));
  NOT NOT1_5506(.VSS(VSS),.VDD(VDD),.Y(I22557),.A(g14775));
  NOT NOT1_5507(.VSS(VSS),.VDD(VDD),.Y(g16485),.A(I22557));
  NOT NOT1_5508(.VSS(VSS),.VDD(VDD),.Y(I22560),.A(g14796));
  NOT NOT1_5509(.VSS(VSS),.VDD(VDD),.Y(g16486),.A(I22560));
  NOT NOT1_5510(.VSS(VSS),.VDD(VDD),.Y(I22563),.A(g14830));
  NOT NOT1_5511(.VSS(VSS),.VDD(VDD),.Y(g16487),.A(I22563));
  NOT NOT1_5512(.VSS(VSS),.VDD(VDD),.Y(I22566),.A(g14883));
  NOT NOT1_5513(.VSS(VSS),.VDD(VDD),.Y(g16488),.A(I22566));
  NOT NOT1_5514(.VSS(VSS),.VDD(VDD),.Y(I22569),.A(g14955));
  NOT NOT1_5515(.VSS(VSS),.VDD(VDD),.Y(g16489),.A(I22569));
  NOT NOT1_5516(.VSS(VSS),.VDD(VDD),.Y(I22572),.A(g15019));
  NOT NOT1_5517(.VSS(VSS),.VDD(VDD),.Y(g16490),.A(I22572));
  NOT NOT1_5518(.VSS(VSS),.VDD(VDD),.Y(I22575),.A(g15092));
  NOT NOT1_5519(.VSS(VSS),.VDD(VDD),.Y(g16491),.A(I22575));
  NOT NOT1_5520(.VSS(VSS),.VDD(VDD),.Y(I22578),.A(g14746));
  NOT NOT1_5521(.VSS(VSS),.VDD(VDD),.Y(g16492),.A(I22578));
  NOT NOT1_5522(.VSS(VSS),.VDD(VDD),.Y(I22581),.A(g14766));
  NOT NOT1_5523(.VSS(VSS),.VDD(VDD),.Y(g16493),.A(I22581));
  NOT NOT1_5524(.VSS(VSS),.VDD(VDD),.Y(I22584),.A(g15989));
  NOT NOT1_5525(.VSS(VSS),.VDD(VDD),.Y(g16494),.A(I22584));
  NOT NOT1_5526(.VSS(VSS),.VDD(VDD),.Y(I22587),.A(g14684));
  NOT NOT1_5527(.VSS(VSS),.VDD(VDD),.Y(g16495),.A(I22587));
  NOT NOT1_5528(.VSS(VSS),.VDD(VDD),.Y(I22590),.A(g13863));
  NOT NOT1_5529(.VSS(VSS),.VDD(VDD),.Y(g16496),.A(I22590));
  NOT NOT1_5530(.VSS(VSS),.VDD(VDD),.Y(I22593),.A(g15876));
  NOT NOT1_5531(.VSS(VSS),.VDD(VDD),.Y(g16497),.A(I22593));
  NOT NOT1_5532(.VSS(VSS),.VDD(VDD),.Y(g16501),.A(g14158));
  NOT NOT1_5533(.VSS(VSS),.VDD(VDD),.Y(I22599),.A(g14966));
  NOT NOT1_5534(.VSS(VSS),.VDD(VDD),.Y(g16506),.A(I22599));
  NOT NOT1_5535(.VSS(VSS),.VDD(VDD),.Y(g16507),.A(g14186));
  NOT NOT1_5536(.VSS(VSS),.VDD(VDD),.Y(I22604),.A(g15080));
  NOT NOT1_5537(.VSS(VSS),.VDD(VDD),.Y(g16514),.A(I22604));
  NOT NOT1_5538(.VSS(VSS),.VDD(VDD),.Y(g16515),.A(g14244));
  NOT NOT1_5539(.VSS(VSS),.VDD(VDD),.Y(g16523),.A(g14273));
  NOT NOT1_5540(.VSS(VSS),.VDD(VDD),.Y(I22611),.A(g15055));
  NOT NOT1_5541(.VSS(VSS),.VDD(VDD),.Y(g16528),.A(I22611));
  NOT NOT1_5542(.VSS(VSS),.VDD(VDD),.Y(g16529),.A(g14301));
  NOT NOT1_5543(.VSS(VSS),.VDD(VDD),.Y(I22618),.A(g14630));
  NOT NOT1_5544(.VSS(VSS),.VDD(VDD),.Y(g16540),.A(I22618));
  NOT NOT1_5545(.VSS(VSS),.VDD(VDD),.Y(g16543),.A(g14347));
  NOT NOT1_5546(.VSS(VSS),.VDD(VDD),.Y(g16546),.A(g14366));
  NOT NOT1_5547(.VSS(VSS),.VDD(VDD),.Y(g16554),.A(g14395));
  NOT NOT1_5548(.VSS(VSS),.VDD(VDD),.Y(I22626),.A(g15151));
  NOT NOT1_5549(.VSS(VSS),.VDD(VDD),.Y(g16559),.A(I22626));
  NOT NOT1_5550(.VSS(VSS),.VDD(VDD),.Y(g16560),.A(g14423));
  NOT NOT1_5551(.VSS(VSS),.VDD(VDD),.Y(I22640),.A(g14650));
  NOT NOT1_5552(.VSS(VSS),.VDD(VDD),.Y(g16572),.A(I22640));
  NOT NOT1_5553(.VSS(VSS),.VDD(VDD),.Y(g16575),.A(g14459));
  NOT NOT1_5554(.VSS(VSS),.VDD(VDD),.Y(g16578),.A(g14478));
  NOT NOT1_5555(.VSS(VSS),.VDD(VDD),.Y(g16586),.A(g14507));
  NOT NOT1_5556(.VSS(VSS),.VDD(VDD),.Y(I22651),.A(g14677));
  NOT NOT1_5557(.VSS(VSS),.VDD(VDD),.Y(g16596),.A(I22651));
  NOT NOT1_5558(.VSS(VSS),.VDD(VDD),.Y(g16599),.A(g14546));
  NOT NOT1_5559(.VSS(VSS),.VDD(VDD),.Y(g16602),.A(g14565));
  NOT NOT1_5560(.VSS(VSS),.VDD(VDD),.Y(I22657),.A(g14657));
  NOT NOT1_5561(.VSS(VSS),.VDD(VDD),.Y(g16608),.A(I22657));
  NOT NOT1_5562(.VSS(VSS),.VDD(VDD),.Y(I22663),.A(g14711));
  NOT NOT1_5563(.VSS(VSS),.VDD(VDD),.Y(g16616),.A(I22663));
  NOT NOT1_5564(.VSS(VSS),.VDD(VDD),.Y(g16619),.A(g14601));
  NOT NOT1_5565(.VSS(VSS),.VDD(VDD),.Y(I22667),.A(g14642));
  NOT NOT1_5566(.VSS(VSS),.VDD(VDD),.Y(g16622),.A(I22667));
  NOT NOT1_5567(.VSS(VSS),.VDD(VDD),.Y(I22671),.A(g14691));
  NOT NOT1_5568(.VSS(VSS),.VDD(VDD),.Y(g16626),.A(I22671));
  NOT NOT1_5569(.VSS(VSS),.VDD(VDD),.Y(I22676),.A(g14630));
  NOT NOT1_5570(.VSS(VSS),.VDD(VDD),.Y(g16633),.A(I22676));
  NOT NOT1_5571(.VSS(VSS),.VDD(VDD),.Y(I22679),.A(g14669));
  NOT NOT1_5572(.VSS(VSS),.VDD(VDD),.Y(g16636),.A(I22679));
  NOT NOT1_5573(.VSS(VSS),.VDD(VDD),.Y(I22683),.A(g14725));
  NOT NOT1_5574(.VSS(VSS),.VDD(VDD),.Y(g16640),.A(I22683));
  NOT NOT1_5575(.VSS(VSS),.VDD(VDD),.Y(I22687),.A(g14650));
  NOT NOT1_5576(.VSS(VSS),.VDD(VDD),.Y(g16644),.A(I22687));
  NOT NOT1_5577(.VSS(VSS),.VDD(VDD),.Y(I22690),.A(g14703));
  NOT NOT1_5578(.VSS(VSS),.VDD(VDD),.Y(g16647),.A(I22690));
  NOT NOT1_5579(.VSS(VSS),.VDD(VDD),.Y(I22694),.A(g14753));
  NOT NOT1_5580(.VSS(VSS),.VDD(VDD),.Y(g16651),.A(I22694));
  NOT NOT1_5581(.VSS(VSS),.VDD(VDD),.Y(I22699),.A(g14677));
  NOT NOT1_5582(.VSS(VSS),.VDD(VDD),.Y(g16656),.A(I22699));
  NOT NOT1_5583(.VSS(VSS),.VDD(VDD),.Y(I22702),.A(g14737));
  NOT NOT1_5584(.VSS(VSS),.VDD(VDD),.Y(g16659),.A(I22702));
  NOT NOT1_5585(.VSS(VSS),.VDD(VDD),.Y(g16665),.A(g14776));
  NOT NOT1_5586(.VSS(VSS),.VDD(VDD),.Y(I22715),.A(g14711));
  NOT NOT1_5587(.VSS(VSS),.VDD(VDD),.Y(g16673),.A(I22715));
  NOT NOT1_5588(.VSS(VSS),.VDD(VDD),.Y(I22718),.A(g14657));
  NOT NOT1_5589(.VSS(VSS),.VDD(VDD),.Y(g16676),.A(I22718));
  NOT NOT1_5590(.VSS(VSS),.VDD(VDD),.Y(g16682),.A(g14797));
  NOT NOT1_5591(.VSS(VSS),.VDD(VDD),.Y(g16686),.A(g14811));
  NOT NOT1_5592(.VSS(VSS),.VDD(VDD),.Y(I22726),.A(g14642));
  NOT NOT1_5593(.VSS(VSS),.VDD(VDD),.Y(g16694),.A(I22726));
  NOT NOT1_5594(.VSS(VSS),.VDD(VDD),.Y(g16697),.A(g14837));
  NOT NOT1_5595(.VSS(VSS),.VDD(VDD),.Y(I22730),.A(g14691));
  NOT NOT1_5596(.VSS(VSS),.VDD(VDD),.Y(g16702),.A(I22730));
  NOT NOT1_5597(.VSS(VSS),.VDD(VDD),.Y(g16708),.A(g14849));
  NOT NOT1_5598(.VSS(VSS),.VDD(VDD),.Y(g16712),.A(g14863));
  NOT NOT1_5599(.VSS(VSS),.VDD(VDD),.Y(I22737),.A(g14630));
  NOT NOT1_5600(.VSS(VSS),.VDD(VDD),.Y(g16719),.A(I22737));
  NOT NOT1_5601(.VSS(VSS),.VDD(VDD),.Y(g16722),.A(g14895));
  NOT NOT1_5602(.VSS(VSS),.VDD(VDD),.Y(I22741),.A(g14669));
  NOT NOT1_5603(.VSS(VSS),.VDD(VDD),.Y(g16725),.A(I22741));
  NOT NOT1_5604(.VSS(VSS),.VDD(VDD),.Y(g16728),.A(g14910));
  NOT NOT1_5605(.VSS(VSS),.VDD(VDD),.Y(I22745),.A(g14725));
  NOT NOT1_5606(.VSS(VSS),.VDD(VDD),.Y(g16733),.A(I22745));
  NOT NOT1_5607(.VSS(VSS),.VDD(VDD),.Y(g16739),.A(g14922));
  NOT NOT1_5608(.VSS(VSS),.VDD(VDD),.Y(g16743),.A(g14936));
  NOT NOT1_5609(.VSS(VSS),.VDD(VDD),.Y(g16749),.A(g15782));
  NOT NOT1_5610(.VSS(VSS),.VDD(VDD),.Y(I22752),.A(g14657));
  NOT NOT1_5611(.VSS(VSS),.VDD(VDD),.Y(g16758),.A(I22752));
  NOT NOT1_5612(.VSS(VSS),.VDD(VDD),.Y(I22755),.A(g14650));
  NOT NOT1_5613(.VSS(VSS),.VDD(VDD),.Y(g16761),.A(I22755));
  NOT NOT1_5614(.VSS(VSS),.VDD(VDD),.Y(g16764),.A(g14976));
  NOT NOT1_5615(.VSS(VSS),.VDD(VDD),.Y(I22759),.A(g14703));
  NOT NOT1_5616(.VSS(VSS),.VDD(VDD),.Y(g16767),.A(I22759));
  NOT NOT1_5617(.VSS(VSS),.VDD(VDD),.Y(g16770),.A(g14991));
  NOT NOT1_5618(.VSS(VSS),.VDD(VDD),.Y(I22763),.A(g14753));
  NOT NOT1_5619(.VSS(VSS),.VDD(VDD),.Y(g16775),.A(I22763));
  NOT NOT1_5620(.VSS(VSS),.VDD(VDD),.Y(g16781),.A(g15003));
  NOT NOT1_5621(.VSS(VSS),.VDD(VDD),.Y(I22768),.A(g14691));
  NOT NOT1_5622(.VSS(VSS),.VDD(VDD),.Y(g16785),.A(I22768));
  NOT NOT1_5623(.VSS(VSS),.VDD(VDD),.Y(I22771),.A(g14677));
  NOT NOT1_5624(.VSS(VSS),.VDD(VDD),.Y(g16788),.A(I22771));
  NOT NOT1_5625(.VSS(VSS),.VDD(VDD),.Y(g16791),.A(g15065));
  NOT NOT1_5626(.VSS(VSS),.VDD(VDD),.Y(I22775),.A(g14737));
  NOT NOT1_5627(.VSS(VSS),.VDD(VDD),.Y(g16794),.A(I22775));
  NOT NOT1_5628(.VSS(VSS),.VDD(VDD),.Y(g16797),.A(g15080));
  NOT NOT1_5629(.VSS(VSS),.VDD(VDD),.Y(g16804),.A(g15803));
  NOT NOT1_5630(.VSS(VSS),.VDD(VDD),.Y(g16809),.A(g15842));
  NOT NOT1_5631(.VSS(VSS),.VDD(VDD),.Y(I22783),.A(g13572));
  NOT NOT1_5632(.VSS(VSS),.VDD(VDD),.Y(g16813),.A(I22783));
  NOT NOT1_5633(.VSS(VSS),.VDD(VDD),.Y(I22786),.A(g14725));
  NOT NOT1_5634(.VSS(VSS),.VDD(VDD),.Y(g16814),.A(I22786));
  NOT NOT1_5635(.VSS(VSS),.VDD(VDD),.Y(I22789),.A(g14711));
  NOT NOT1_5636(.VSS(VSS),.VDD(VDD),.Y(g16817),.A(I22789));
  NOT NOT1_5637(.VSS(VSS),.VDD(VDD),.Y(g16820),.A(g15161));
  NOT NOT1_5638(.VSS(VSS),.VDD(VDD),.Y(g16825),.A(g15855));
  NOT NOT1_5639(.VSS(VSS),.VDD(VDD),.Y(I22797),.A(g14165));
  NOT NOT1_5640(.VSS(VSS),.VDD(VDD),.Y(g16830),.A(I22797));
  NOT NOT1_5641(.VSS(VSS),.VDD(VDD),.Y(I22800),.A(g13581));
  NOT NOT1_5642(.VSS(VSS),.VDD(VDD),.Y(g16831),.A(I22800));
  NOT NOT1_5643(.VSS(VSS),.VDD(VDD),.Y(I22803),.A(g14753));
  NOT NOT1_5644(.VSS(VSS),.VDD(VDD),.Y(g16832),.A(I22803));
  NOT NOT1_5645(.VSS(VSS),.VDD(VDD),.Y(g16836),.A(g15818));
  NOT NOT1_5646(.VSS(VSS),.VDD(VDD),.Y(g16840),.A(g15878));
  NOT NOT1_5647(.VSS(VSS),.VDD(VDD),.Y(I22810),.A(g14280));
  NOT NOT1_5648(.VSS(VSS),.VDD(VDD),.Y(g16842),.A(I22810));
  NOT NOT1_5649(.VSS(VSS),.VDD(VDD),.Y(I22813),.A(g13601));
  NOT NOT1_5650(.VSS(VSS),.VDD(VDD),.Y(g16843),.A(I22813));
  NOT NOT1_5651(.VSS(VSS),.VDD(VDD),.Y(g16846),.A(g15903));
  NOT NOT1_5652(.VSS(VSS),.VDD(VDD),.Y(I22820),.A(g14402));
  NOT NOT1_5653(.VSS(VSS),.VDD(VDD),.Y(g16848),.A(I22820));
  NOT NOT1_5654(.VSS(VSS),.VDD(VDD),.Y(I22823),.A(g13613));
  NOT NOT1_5655(.VSS(VSS),.VDD(VDD),.Y(g16849),.A(I22823));
  NOT NOT1_5656(.VSS(VSS),.VDD(VDD),.Y(I22828),.A(g14514));
  NOT NOT1_5657(.VSS(VSS),.VDD(VDD),.Y(g16852),.A(I22828));
  NOT NOT1_5658(.VSS(VSS),.VDD(VDD),.Y(I22836),.A(g13571));
  NOT NOT1_5659(.VSS(VSS),.VDD(VDD),.Y(g16858),.A(I22836));
  NOT NOT1_5660(.VSS(VSS),.VDD(VDD),.Y(I22842),.A(g13580));
  NOT NOT1_5661(.VSS(VSS),.VDD(VDD),.Y(g16862),.A(I22842));
  NOT NOT1_5662(.VSS(VSS),.VDD(VDD),.Y(I22845),.A(g13579));
  NOT NOT1_5663(.VSS(VSS),.VDD(VDD),.Y(g16863),.A(I22845));
  NOT NOT1_5664(.VSS(VSS),.VDD(VDD),.Y(g16867),.A(g13589));
  NOT NOT1_5665(.VSS(VSS),.VDD(VDD),.Y(I22852),.A(g13600));
  NOT NOT1_5666(.VSS(VSS),.VDD(VDD),.Y(g16877),.A(I22852));
  NOT NOT1_5667(.VSS(VSS),.VDD(VDD),.Y(I22855),.A(g13588));
  NOT NOT1_5668(.VSS(VSS),.VDD(VDD),.Y(g16878),.A(I22855));
  NOT NOT1_5669(.VSS(VSS),.VDD(VDD),.Y(I22860),.A(g14885));
  NOT NOT1_5670(.VSS(VSS),.VDD(VDD),.Y(g16881),.A(I22860));
  NOT NOT1_5671(.VSS(VSS),.VDD(VDD),.Y(g16884),.A(g13589));
  NOT NOT1_5672(.VSS(VSS),.VDD(VDD),.Y(g16895),.A(g13589));
  NOT NOT1_5673(.VSS(VSS),.VDD(VDD),.Y(I22866),.A(g13612));
  NOT NOT1_5674(.VSS(VSS),.VDD(VDD),.Y(g16905),.A(I22866));
  NOT NOT1_5675(.VSS(VSS),.VDD(VDD),.Y(I22869),.A(g13608));
  NOT NOT1_5676(.VSS(VSS),.VDD(VDD),.Y(g16906),.A(I22869));
  NOT NOT1_5677(.VSS(VSS),.VDD(VDD),.Y(I22875),.A(g14966));
  NOT NOT1_5678(.VSS(VSS),.VDD(VDD),.Y(g16910),.A(I22875));
  NOT NOT1_5679(.VSS(VSS),.VDD(VDD),.Y(g16913),.A(g13589));
  NOT NOT1_5680(.VSS(VSS),.VDD(VDD),.Y(g16924),.A(g13589));
  NOT NOT1_5681(.VSS(VSS),.VDD(VDD),.Y(I22881),.A(g13622));
  NOT NOT1_5682(.VSS(VSS),.VDD(VDD),.Y(g16934),.A(I22881));
  NOT NOT1_5683(.VSS(VSS),.VDD(VDD),.Y(I22893),.A(g15055));
  NOT NOT1_5684(.VSS(VSS),.VDD(VDD),.Y(g16940),.A(I22893));
  NOT NOT1_5685(.VSS(VSS),.VDD(VDD),.Y(g16943),.A(g13589));
  NOT NOT1_5686(.VSS(VSS),.VDD(VDD),.Y(g16954),.A(g13589));
  NOT NOT1_5687(.VSS(VSS),.VDD(VDD),.Y(I22912),.A(g15151));
  NOT NOT1_5688(.VSS(VSS),.VDD(VDD),.Y(g16971),.A(I22912));
  NOT NOT1_5689(.VSS(VSS),.VDD(VDD),.Y(g16974),.A(g13589));
  NOT NOT1_5690(.VSS(VSS),.VDD(VDD),.Y(g17029),.A(g14685));
  NOT NOT1_5691(.VSS(VSS),.VDD(VDD),.Y(g17057),.A(g13519));
  NOT NOT1_5692(.VSS(VSS),.VDD(VDD),.Y(g17063),.A(g14719));
  NOT NOT1_5693(.VSS(VSS),.VDD(VDD),.Y(g17092),.A(g13530));
  NOT NOT1_5694(.VSS(VSS),.VDD(VDD),.Y(g17098),.A(g14747));
  NOT NOT1_5695(.VSS(VSS),.VDD(VDD),.Y(g17130),.A(g13541));
  NOT NOT1_5696(.VSS(VSS),.VDD(VDD),.Y(g17136),.A(g14768));
  NOT NOT1_5697(.VSS(VSS),.VDD(VDD),.Y(g17157),.A(g13552));
  NOT NOT1_5698(.VSS(VSS),.VDD(VDD),.Y(I23253),.A(g13741));
  NOT NOT1_5699(.VSS(VSS),.VDD(VDD),.Y(g17189),.A(I23253));
  NOT NOT1_5700(.VSS(VSS),.VDD(VDD),.Y(I23274),.A(g13741));
  NOT NOT1_5701(.VSS(VSS),.VDD(VDD),.Y(g17200),.A(I23274));
  NOT NOT1_5702(.VSS(VSS),.VDD(VDD),.Y(g17203),.A(g13568));
  NOT NOT1_5703(.VSS(VSS),.VDD(VDD),.Y(I23287),.A(g13741));
  NOT NOT1_5704(.VSS(VSS),.VDD(VDD),.Y(g17207),.A(I23287));
  NOT NOT1_5705(.VSS(VSS),.VDD(VDD),.Y(g17208),.A(g13576));
  NOT NOT1_5706(.VSS(VSS),.VDD(VDD),.Y(I23292),.A(g13741));
  NOT NOT1_5707(.VSS(VSS),.VDD(VDD),.Y(g17212),.A(I23292));
  NOT NOT1_5708(.VSS(VSS),.VDD(VDD),.Y(g17214),.A(g13585));
  NOT NOT1_5709(.VSS(VSS),.VDD(VDD),.Y(g17217),.A(g13605));
  NOT NOT1_5710(.VSS(VSS),.VDD(VDD),.Y(I23309),.A(g16132));
  NOT NOT1_5711(.VSS(VSS),.VDD(VDD),.Y(g17227),.A(I23309));
  NOT NOT1_5712(.VSS(VSS),.VDD(VDD),.Y(I23314),.A(g15720));
  NOT NOT1_5713(.VSS(VSS),.VDD(VDD),.Y(g17230),.A(I23314));
  NOT NOT1_5714(.VSS(VSS),.VDD(VDD),.Y(I23317),.A(g16181));
  NOT NOT1_5715(.VSS(VSS),.VDD(VDD),.Y(g17233),.A(I23317));
  NOT NOT1_5716(.VSS(VSS),.VDD(VDD),.Y(I23323),.A(g15664));
  NOT NOT1_5717(.VSS(VSS),.VDD(VDD),.Y(g17237),.A(I23323));
  NOT NOT1_5718(.VSS(VSS),.VDD(VDD),.Y(I23326),.A(g15758));
  NOT NOT1_5719(.VSS(VSS),.VDD(VDD),.Y(g17240),.A(I23326));
  NOT NOT1_5720(.VSS(VSS),.VDD(VDD),.Y(I23329),.A(g15760));
  NOT NOT1_5721(.VSS(VSS),.VDD(VDD),.Y(g17243),.A(I23329));
  NOT NOT1_5722(.VSS(VSS),.VDD(VDD),.Y(I23335),.A(g16412));
  NOT NOT1_5723(.VSS(VSS),.VDD(VDD),.Y(g17249),.A(I23335));
  NOT NOT1_5724(.VSS(VSS),.VDD(VDD),.Y(I23338),.A(g15721));
  NOT NOT1_5725(.VSS(VSS),.VDD(VDD),.Y(g17252),.A(I23338));
  NOT NOT1_5726(.VSS(VSS),.VDD(VDD),.Y(I23341),.A(g15784));
  NOT NOT1_5727(.VSS(VSS),.VDD(VDD),.Y(g17255),.A(I23341));
  NOT NOT1_5728(.VSS(VSS),.VDD(VDD),.Y(g17258),.A(g16053));
  NOT NOT1_5729(.VSS(VSS),.VDD(VDD),.Y(I23345),.A(g15723));
  NOT NOT1_5730(.VSS(VSS),.VDD(VDD),.Y(g17259),.A(I23345));
  NOT NOT1_5731(.VSS(VSS),.VDD(VDD),.Y(I23348),.A(g15786));
  NOT NOT1_5732(.VSS(VSS),.VDD(VDD),.Y(g17262),.A(I23348));
  NOT NOT1_5733(.VSS(VSS),.VDD(VDD),.Y(I23351),.A(g15788));
  NOT NOT1_5734(.VSS(VSS),.VDD(VDD),.Y(g17265),.A(I23351));
  NOT NOT1_5735(.VSS(VSS),.VDD(VDD),.Y(I23358),.A(g16442));
  NOT NOT1_5736(.VSS(VSS),.VDD(VDD),.Y(g17272),.A(I23358));
  NOT NOT1_5737(.VSS(VSS),.VDD(VDD),.Y(I23361),.A(g15759));
  NOT NOT1_5738(.VSS(VSS),.VDD(VDD),.Y(g17275),.A(I23361));
  NOT NOT1_5739(.VSS(VSS),.VDD(VDD),.Y(I23364),.A(g15805));
  NOT NOT1_5740(.VSS(VSS),.VDD(VDD),.Y(g17278),.A(I23364));
  NOT NOT1_5741(.VSS(VSS),.VDD(VDD),.Y(g17281),.A(g16081));
  NOT NOT1_5742(.VSS(VSS),.VDD(VDD),.Y(I23368),.A(g16446));
  NOT NOT1_5743(.VSS(VSS),.VDD(VDD),.Y(g17282),.A(I23368));
  NOT NOT1_5744(.VSS(VSS),.VDD(VDD),.Y(I23371),.A(g15761));
  NOT NOT1_5745(.VSS(VSS),.VDD(VDD),.Y(g17285),.A(I23371));
  NOT NOT1_5746(.VSS(VSS),.VDD(VDD),.Y(I23374),.A(g15807));
  NOT NOT1_5747(.VSS(VSS),.VDD(VDD),.Y(g17288),.A(I23374));
  NOT NOT1_5748(.VSS(VSS),.VDD(VDD),.Y(I23377),.A(g15763));
  NOT NOT1_5749(.VSS(VSS),.VDD(VDD),.Y(g17291),.A(I23377));
  NOT NOT1_5750(.VSS(VSS),.VDD(VDD),.Y(I23380),.A(g15809));
  NOT NOT1_5751(.VSS(VSS),.VDD(VDD),.Y(g17294),.A(I23380));
  NOT NOT1_5752(.VSS(VSS),.VDD(VDD),.Y(I23383),.A(g15811));
  NOT NOT1_5753(.VSS(VSS),.VDD(VDD),.Y(g17297),.A(I23383));
  NOT NOT1_5754(.VSS(VSS),.VDD(VDD),.Y(I23386),.A(g13469));
  NOT NOT1_5755(.VSS(VSS),.VDD(VDD),.Y(g17300),.A(I23386));
  NOT NOT1_5756(.VSS(VSS),.VDD(VDD),.Y(I23392),.A(g13476));
  NOT NOT1_5757(.VSS(VSS),.VDD(VDD),.Y(g17304),.A(I23392));
  NOT NOT1_5758(.VSS(VSS),.VDD(VDD),.Y(I23395),.A(g15785));
  NOT NOT1_5759(.VSS(VSS),.VDD(VDD),.Y(g17307),.A(I23395));
  NOT NOT1_5760(.VSS(VSS),.VDD(VDD),.Y(I23398),.A(g15820));
  NOT NOT1_5761(.VSS(VSS),.VDD(VDD),.Y(g17310),.A(I23398));
  NOT NOT1_5762(.VSS(VSS),.VDD(VDD),.Y(g17313),.A(g16109));
  NOT NOT1_5763(.VSS(VSS),.VDD(VDD),.Y(g17314),.A(g16110));
  NOT NOT1_5764(.VSS(VSS),.VDD(VDD),.Y(I23403),.A(g13478));
  NOT NOT1_5765(.VSS(VSS),.VDD(VDD),.Y(g17315),.A(I23403));
  NOT NOT1_5766(.VSS(VSS),.VDD(VDD),.Y(I23406),.A(g15787));
  NOT NOT1_5767(.VSS(VSS),.VDD(VDD),.Y(g17318),.A(I23406));
  NOT NOT1_5768(.VSS(VSS),.VDD(VDD),.Y(I23409),.A(g15822));
  NOT NOT1_5769(.VSS(VSS),.VDD(VDD),.Y(g17321),.A(I23409));
  NOT NOT1_5770(.VSS(VSS),.VDD(VDD),.Y(I23412),.A(g13482));
  NOT NOT1_5771(.VSS(VSS),.VDD(VDD),.Y(g17324),.A(I23412));
  NOT NOT1_5772(.VSS(VSS),.VDD(VDD),.Y(I23415),.A(g15789));
  NOT NOT1_5773(.VSS(VSS),.VDD(VDD),.Y(g17327),.A(I23415));
  NOT NOT1_5774(.VSS(VSS),.VDD(VDD),.Y(I23418),.A(g15824));
  NOT NOT1_5775(.VSS(VSS),.VDD(VDD),.Y(g17330),.A(I23418));
  NOT NOT1_5776(.VSS(VSS),.VDD(VDD),.Y(I23421),.A(g15791));
  NOT NOT1_5777(.VSS(VSS),.VDD(VDD),.Y(g17333),.A(I23421));
  NOT NOT1_5778(.VSS(VSS),.VDD(VDD),.Y(I23424),.A(g15826));
  NOT NOT1_5779(.VSS(VSS),.VDD(VDD),.Y(g17336),.A(I23424));
  NOT NOT1_5780(.VSS(VSS),.VDD(VDD),.Y(I23430),.A(g13494));
  NOT NOT1_5781(.VSS(VSS),.VDD(VDD),.Y(g17342),.A(I23430));
  NOT NOT1_5782(.VSS(VSS),.VDD(VDD),.Y(I23433),.A(g15806));
  NOT NOT1_5783(.VSS(VSS),.VDD(VDD),.Y(g17345),.A(I23433));
  NOT NOT1_5784(.VSS(VSS),.VDD(VDD),.Y(I23436),.A(g15832));
  NOT NOT1_5785(.VSS(VSS),.VDD(VDD),.Y(g17348),.A(I23436));
  NOT NOT1_5786(.VSS(VSS),.VDD(VDD),.Y(g17351),.A(g16152));
  NOT NOT1_5787(.VSS(VSS),.VDD(VDD),.Y(I23442),.A(g13495));
  NOT NOT1_5788(.VSS(VSS),.VDD(VDD),.Y(g17354),.A(I23442));
  NOT NOT1_5789(.VSS(VSS),.VDD(VDD),.Y(I23445),.A(g15808));
  NOT NOT1_5790(.VSS(VSS),.VDD(VDD),.Y(g17357),.A(I23445));
  NOT NOT1_5791(.VSS(VSS),.VDD(VDD),.Y(I23448),.A(g15834));
  NOT NOT1_5792(.VSS(VSS),.VDD(VDD),.Y(g17360),.A(I23448));
  NOT NOT1_5793(.VSS(VSS),.VDD(VDD),.Y(I23451),.A(g13497));
  NOT NOT1_5794(.VSS(VSS),.VDD(VDD),.Y(g17363),.A(I23451));
  NOT NOT1_5795(.VSS(VSS),.VDD(VDD),.Y(I23454),.A(g15810));
  NOT NOT1_5796(.VSS(VSS),.VDD(VDD),.Y(g17366),.A(I23454));
  NOT NOT1_5797(.VSS(VSS),.VDD(VDD),.Y(I23457),.A(g15836));
  NOT NOT1_5798(.VSS(VSS),.VDD(VDD),.Y(g17369),.A(I23457));
  NOT NOT1_5799(.VSS(VSS),.VDD(VDD),.Y(I23460),.A(g13501));
  NOT NOT1_5800(.VSS(VSS),.VDD(VDD),.Y(g17372),.A(I23460));
  NOT NOT1_5801(.VSS(VSS),.VDD(VDD),.Y(I23463),.A(g15812));
  NOT NOT1_5802(.VSS(VSS),.VDD(VDD),.Y(g17375),.A(I23463));
  NOT NOT1_5803(.VSS(VSS),.VDD(VDD),.Y(I23466),.A(g15838));
  NOT NOT1_5804(.VSS(VSS),.VDD(VDD),.Y(g17378),.A(I23466));
  NOT NOT1_5805(.VSS(VSS),.VDD(VDD),.Y(I23472),.A(g13510));
  NOT NOT1_5806(.VSS(VSS),.VDD(VDD),.Y(g17384),.A(I23472));
  NOT NOT1_5807(.VSS(VSS),.VDD(VDD),.Y(I23475),.A(g15821));
  NOT NOT1_5808(.VSS(VSS),.VDD(VDD),.Y(g17387),.A(I23475));
  NOT NOT1_5809(.VSS(VSS),.VDD(VDD),.Y(I23478),.A(g15844));
  NOT NOT1_5810(.VSS(VSS),.VDD(VDD),.Y(g17390),.A(I23478));
  NOT NOT1_5811(.VSS(VSS),.VDD(VDD),.Y(g17394),.A(g16197));
  NOT NOT1_5812(.VSS(VSS),.VDD(VDD),.Y(I23487),.A(g13511));
  NOT NOT1_5813(.VSS(VSS),.VDD(VDD),.Y(g17399),.A(I23487));
  NOT NOT1_5814(.VSS(VSS),.VDD(VDD),.Y(I23490),.A(g15823));
  NOT NOT1_5815(.VSS(VSS),.VDD(VDD),.Y(g17402),.A(I23490));
  NOT NOT1_5816(.VSS(VSS),.VDD(VDD),.Y(I23493),.A(g15846));
  NOT NOT1_5817(.VSS(VSS),.VDD(VDD),.Y(g17405),.A(I23493));
  NOT NOT1_5818(.VSS(VSS),.VDD(VDD),.Y(I23498),.A(g13512));
  NOT NOT1_5819(.VSS(VSS),.VDD(VDD),.Y(g17410),.A(I23498));
  NOT NOT1_5820(.VSS(VSS),.VDD(VDD),.Y(I23501),.A(g15825));
  NOT NOT1_5821(.VSS(VSS),.VDD(VDD),.Y(g17413),.A(I23501));
  NOT NOT1_5822(.VSS(VSS),.VDD(VDD),.Y(I23504),.A(g15848));
  NOT NOT1_5823(.VSS(VSS),.VDD(VDD),.Y(g17416),.A(I23504));
  NOT NOT1_5824(.VSS(VSS),.VDD(VDD),.Y(I23507),.A(g13514));
  NOT NOT1_5825(.VSS(VSS),.VDD(VDD),.Y(g17419),.A(I23507));
  NOT NOT1_5826(.VSS(VSS),.VDD(VDD),.Y(I23510),.A(g15827));
  NOT NOT1_5827(.VSS(VSS),.VDD(VDD),.Y(g17422),.A(I23510));
  NOT NOT1_5828(.VSS(VSS),.VDD(VDD),.Y(I23513),.A(g15850));
  NOT NOT1_5829(.VSS(VSS),.VDD(VDD),.Y(g17425),.A(I23513));
  NOT NOT1_5830(.VSS(VSS),.VDD(VDD),.Y(I23518),.A(g15856));
  NOT NOT1_5831(.VSS(VSS),.VDD(VDD),.Y(g17430),.A(I23518));
  NOT NOT1_5832(.VSS(VSS),.VDD(VDD),.Y(I23521),.A(g13518));
  NOT NOT1_5833(.VSS(VSS),.VDD(VDD),.Y(g17433),.A(I23521));
  NOT NOT1_5834(.VSS(VSS),.VDD(VDD),.Y(I23524),.A(g15833));
  NOT NOT1_5835(.VSS(VSS),.VDD(VDD),.Y(g17436),.A(I23524));
  NOT NOT1_5836(.VSS(VSS),.VDD(VDD),.Y(I23527),.A(g15858));
  NOT NOT1_5837(.VSS(VSS),.VDD(VDD),.Y(g17439),.A(I23527));
  NOT NOT1_5838(.VSS(VSS),.VDD(VDD),.Y(I23530),.A(g14885));
  NOT NOT1_5839(.VSS(VSS),.VDD(VDD),.Y(g17442),.A(I23530));
  NOT NOT1_5840(.VSS(VSS),.VDD(VDD),.Y(g17445),.A(g16250));
  NOT NOT1_5841(.VSS(VSS),.VDD(VDD),.Y(I23539),.A(g13524));
  NOT NOT1_5842(.VSS(VSS),.VDD(VDD),.Y(g17451),.A(I23539));
  NOT NOT1_5843(.VSS(VSS),.VDD(VDD),.Y(I23542),.A(g15835));
  NOT NOT1_5844(.VSS(VSS),.VDD(VDD),.Y(g17454),.A(I23542));
  NOT NOT1_5845(.VSS(VSS),.VDD(VDD),.Y(I23545),.A(g15867));
  NOT NOT1_5846(.VSS(VSS),.VDD(VDD),.Y(g17457),.A(I23545));
  NOT NOT1_5847(.VSS(VSS),.VDD(VDD),.Y(I23553),.A(g13525));
  NOT NOT1_5848(.VSS(VSS),.VDD(VDD),.Y(g17465),.A(I23553));
  NOT NOT1_5849(.VSS(VSS),.VDD(VDD),.Y(I23556),.A(g15837));
  NOT NOT1_5850(.VSS(VSS),.VDD(VDD),.Y(g17468),.A(I23556));
  NOT NOT1_5851(.VSS(VSS),.VDD(VDD),.Y(I23559),.A(g15869));
  NOT NOT1_5852(.VSS(VSS),.VDD(VDD),.Y(g17471),.A(I23559));
  NOT NOT1_5853(.VSS(VSS),.VDD(VDD),.Y(I23564),.A(g13526));
  NOT NOT1_5854(.VSS(VSS),.VDD(VDD),.Y(g17476),.A(I23564));
  NOT NOT1_5855(.VSS(VSS),.VDD(VDD),.Y(I23567),.A(g15839));
  NOT NOT1_5856(.VSS(VSS),.VDD(VDD),.Y(g17479),.A(I23567));
  NOT NOT1_5857(.VSS(VSS),.VDD(VDD),.Y(I23570),.A(g15871));
  NOT NOT1_5858(.VSS(VSS),.VDD(VDD),.Y(g17482),.A(I23570));
  NOT NOT1_5859(.VSS(VSS),.VDD(VDD),.Y(I23575),.A(g15843));
  NOT NOT1_5860(.VSS(VSS),.VDD(VDD),.Y(g17487),.A(I23575));
  NOT NOT1_5861(.VSS(VSS),.VDD(VDD),.Y(I23578),.A(g15879));
  NOT NOT1_5862(.VSS(VSS),.VDD(VDD),.Y(g17490),.A(I23578));
  NOT NOT1_5863(.VSS(VSS),.VDD(VDD),.Y(I23581),.A(g13528));
  NOT NOT1_5864(.VSS(VSS),.VDD(VDD),.Y(g17493),.A(I23581));
  NOT NOT1_5865(.VSS(VSS),.VDD(VDD),.Y(I23584),.A(g15845));
  NOT NOT1_5866(.VSS(VSS),.VDD(VDD),.Y(g17496),.A(I23584));
  NOT NOT1_5867(.VSS(VSS),.VDD(VDD),.Y(g17499),.A(g16292));
  NOT NOT1_5868(.VSS(VSS),.VDD(VDD),.Y(I23588),.A(g14885));
  NOT NOT1_5869(.VSS(VSS),.VDD(VDD),.Y(g17500),.A(I23588));
  NOT NOT1_5870(.VSS(VSS),.VDD(VDD),.Y(I23591),.A(g14885));
  NOT NOT1_5871(.VSS(VSS),.VDD(VDD),.Y(g17503),.A(I23591));
  NOT NOT1_5872(.VSS(VSS),.VDD(VDD),.Y(I23599),.A(g15887));
  NOT NOT1_5873(.VSS(VSS),.VDD(VDD),.Y(g17511),.A(I23599));
  NOT NOT1_5874(.VSS(VSS),.VDD(VDD),.Y(I23602),.A(g13529));
  NOT NOT1_5875(.VSS(VSS),.VDD(VDD),.Y(g17514),.A(I23602));
  NOT NOT1_5876(.VSS(VSS),.VDD(VDD),.Y(I23605),.A(g15847));
  NOT NOT1_5877(.VSS(VSS),.VDD(VDD),.Y(g17517),.A(I23605));
  NOT NOT1_5878(.VSS(VSS),.VDD(VDD),.Y(I23608),.A(g15889));
  NOT NOT1_5879(.VSS(VSS),.VDD(VDD),.Y(g17520),.A(I23608));
  NOT NOT1_5880(.VSS(VSS),.VDD(VDD),.Y(I23611),.A(g14966));
  NOT NOT1_5881(.VSS(VSS),.VDD(VDD),.Y(g17523),.A(I23611));
  NOT NOT1_5882(.VSS(VSS),.VDD(VDD),.Y(I23619),.A(g13535));
  NOT NOT1_5883(.VSS(VSS),.VDD(VDD),.Y(g17531),.A(I23619));
  NOT NOT1_5884(.VSS(VSS),.VDD(VDD),.Y(I23622),.A(g15849));
  NOT NOT1_5885(.VSS(VSS),.VDD(VDD),.Y(g17534),.A(I23622));
  NOT NOT1_5886(.VSS(VSS),.VDD(VDD),.Y(I23625),.A(g15898));
  NOT NOT1_5887(.VSS(VSS),.VDD(VDD),.Y(g17537),.A(I23625));
  NOT NOT1_5888(.VSS(VSS),.VDD(VDD),.Y(I23633),.A(g13536));
  NOT NOT1_5889(.VSS(VSS),.VDD(VDD),.Y(g17545),.A(I23633));
  NOT NOT1_5890(.VSS(VSS),.VDD(VDD),.Y(I23636),.A(g15851));
  NOT NOT1_5891(.VSS(VSS),.VDD(VDD),.Y(g17548),.A(I23636));
  NOT NOT1_5892(.VSS(VSS),.VDD(VDD),.Y(I23639),.A(g15900));
  NOT NOT1_5893(.VSS(VSS),.VDD(VDD),.Y(g17551),.A(I23639));
  NOT NOT1_5894(.VSS(VSS),.VDD(VDD),.Y(I23645),.A(g13537));
  NOT NOT1_5895(.VSS(VSS),.VDD(VDD),.Y(g17557),.A(I23645));
  NOT NOT1_5896(.VSS(VSS),.VDD(VDD),.Y(I23648),.A(g15857));
  NOT NOT1_5897(.VSS(VSS),.VDD(VDD),.Y(g17560),.A(I23648));
  NOT NOT1_5898(.VSS(VSS),.VDD(VDD),.Y(I23651),.A(g13538));
  NOT NOT1_5899(.VSS(VSS),.VDD(VDD),.Y(g17563),.A(I23651));
  NOT NOT1_5900(.VSS(VSS),.VDD(VDD),.Y(g17566),.A(g16346));
  NOT NOT1_5901(.VSS(VSS),.VDD(VDD),.Y(I23655),.A(g14831));
  NOT NOT1_5902(.VSS(VSS),.VDD(VDD),.Y(g17567),.A(I23655));
  NOT NOT1_5903(.VSS(VSS),.VDD(VDD),.Y(I23658),.A(g14885));
  NOT NOT1_5904(.VSS(VSS),.VDD(VDD),.Y(g17570),.A(I23658));
  NOT NOT1_5905(.VSS(VSS),.VDD(VDD),.Y(I23661),.A(g16085));
  NOT NOT1_5906(.VSS(VSS),.VDD(VDD),.Y(g17573),.A(I23661));
  NOT NOT1_5907(.VSS(VSS),.VDD(VDD),.Y(I23667),.A(g15866));
  NOT NOT1_5908(.VSS(VSS),.VDD(VDD),.Y(g17579),.A(I23667));
  NOT NOT1_5909(.VSS(VSS),.VDD(VDD),.Y(I23670),.A(g15912));
  NOT NOT1_5910(.VSS(VSS),.VDD(VDD),.Y(g17582),.A(I23670));
  NOT NOT1_5911(.VSS(VSS),.VDD(VDD),.Y(I23673),.A(g13539));
  NOT NOT1_5912(.VSS(VSS),.VDD(VDD),.Y(g17585),.A(I23673));
  NOT NOT1_5913(.VSS(VSS),.VDD(VDD),.Y(I23676),.A(g15868));
  NOT NOT1_5914(.VSS(VSS),.VDD(VDD),.Y(g17588),.A(I23676));
  NOT NOT1_5915(.VSS(VSS),.VDD(VDD),.Y(I23679),.A(g14966));
  NOT NOT1_5916(.VSS(VSS),.VDD(VDD),.Y(g17591),.A(I23679));
  NOT NOT1_5917(.VSS(VSS),.VDD(VDD),.Y(I23682),.A(g14966));
  NOT NOT1_5918(.VSS(VSS),.VDD(VDD),.Y(g17594),.A(I23682));
  NOT NOT1_5919(.VSS(VSS),.VDD(VDD),.Y(I23689),.A(g15920));
  NOT NOT1_5920(.VSS(VSS),.VDD(VDD),.Y(g17601),.A(I23689));
  NOT NOT1_5921(.VSS(VSS),.VDD(VDD),.Y(I23692),.A(g13540));
  NOT NOT1_5922(.VSS(VSS),.VDD(VDD),.Y(g17604),.A(I23692));
  NOT NOT1_5923(.VSS(VSS),.VDD(VDD),.Y(I23695),.A(g15870));
  NOT NOT1_5924(.VSS(VSS),.VDD(VDD),.Y(g17607),.A(I23695));
  NOT NOT1_5925(.VSS(VSS),.VDD(VDD),.Y(I23698),.A(g15922));
  NOT NOT1_5926(.VSS(VSS),.VDD(VDD),.Y(g17610),.A(I23698));
  NOT NOT1_5927(.VSS(VSS),.VDD(VDD),.Y(I23701),.A(g15055));
  NOT NOT1_5928(.VSS(VSS),.VDD(VDD),.Y(g17613),.A(I23701));
  NOT NOT1_5929(.VSS(VSS),.VDD(VDD),.Y(I23709),.A(g13546));
  NOT NOT1_5930(.VSS(VSS),.VDD(VDD),.Y(g17621),.A(I23709));
  NOT NOT1_5931(.VSS(VSS),.VDD(VDD),.Y(I23712),.A(g15872));
  NOT NOT1_5932(.VSS(VSS),.VDD(VDD),.Y(g17624),.A(I23712));
  NOT NOT1_5933(.VSS(VSS),.VDD(VDD),.Y(I23715),.A(g15931));
  NOT NOT1_5934(.VSS(VSS),.VDD(VDD),.Y(g17627),.A(I23715));
  NOT NOT1_5935(.VSS(VSS),.VDD(VDD),.Y(I23725),.A(g13547));
  NOT NOT1_5936(.VSS(VSS),.VDD(VDD),.Y(g17637),.A(I23725));
  NOT NOT1_5937(.VSS(VSS),.VDD(VDD),.Y(g17640),.A(g13873));
  NOT NOT1_5938(.VSS(VSS),.VDD(VDD),.Y(I23729),.A(g14337));
  NOT NOT1_5939(.VSS(VSS),.VDD(VDD),.Y(g17645),.A(I23729));
  NOT NOT1_5940(.VSS(VSS),.VDD(VDD),.Y(g17648),.A(g16384));
  NOT NOT1_5941(.VSS(VSS),.VDD(VDD),.Y(I23733),.A(g14831));
  NOT NOT1_5942(.VSS(VSS),.VDD(VDD),.Y(g17649),.A(I23733));
  NOT NOT1_5943(.VSS(VSS),.VDD(VDD),.Y(I23739),.A(g13548));
  NOT NOT1_5944(.VSS(VSS),.VDD(VDD),.Y(g17655),.A(I23739));
  NOT NOT1_5945(.VSS(VSS),.VDD(VDD),.Y(I23742),.A(g15888));
  NOT NOT1_5946(.VSS(VSS),.VDD(VDD),.Y(g17658),.A(I23742));
  NOT NOT1_5947(.VSS(VSS),.VDD(VDD),.Y(I23745),.A(g13549));
  NOT NOT1_5948(.VSS(VSS),.VDD(VDD),.Y(g17661),.A(I23745));
  NOT NOT1_5949(.VSS(VSS),.VDD(VDD),.Y(I23748),.A(g14904));
  NOT NOT1_5950(.VSS(VSS),.VDD(VDD),.Y(g17664),.A(I23748));
  NOT NOT1_5951(.VSS(VSS),.VDD(VDD),.Y(I23751),.A(g14966));
  NOT NOT1_5952(.VSS(VSS),.VDD(VDD),.Y(g17667),.A(I23751));
  NOT NOT1_5953(.VSS(VSS),.VDD(VDD),.Y(I23754),.A(g16123));
  NOT NOT1_5954(.VSS(VSS),.VDD(VDD),.Y(g17670),.A(I23754));
  NOT NOT1_5955(.VSS(VSS),.VDD(VDD),.Y(I23760),.A(g15897));
  NOT NOT1_5956(.VSS(VSS),.VDD(VDD),.Y(g17676),.A(I23760));
  NOT NOT1_5957(.VSS(VSS),.VDD(VDD),.Y(I23763),.A(g15941));
  NOT NOT1_5958(.VSS(VSS),.VDD(VDD),.Y(g17679),.A(I23763));
  NOT NOT1_5959(.VSS(VSS),.VDD(VDD),.Y(I23766),.A(g13550));
  NOT NOT1_5960(.VSS(VSS),.VDD(VDD),.Y(g17682),.A(I23766));
  NOT NOT1_5961(.VSS(VSS),.VDD(VDD),.Y(I23769),.A(g15899));
  NOT NOT1_5962(.VSS(VSS),.VDD(VDD),.Y(g17685),.A(I23769));
  NOT NOT1_5963(.VSS(VSS),.VDD(VDD),.Y(I23772),.A(g15055));
  NOT NOT1_5964(.VSS(VSS),.VDD(VDD),.Y(g17688),.A(I23772));
  NOT NOT1_5965(.VSS(VSS),.VDD(VDD),.Y(I23775),.A(g15055));
  NOT NOT1_5966(.VSS(VSS),.VDD(VDD),.Y(g17691),.A(I23775));
  NOT NOT1_5967(.VSS(VSS),.VDD(VDD),.Y(I23782),.A(g15949));
  NOT NOT1_5968(.VSS(VSS),.VDD(VDD),.Y(g17698),.A(I23782));
  NOT NOT1_5969(.VSS(VSS),.VDD(VDD),.Y(I23785),.A(g13551));
  NOT NOT1_5970(.VSS(VSS),.VDD(VDD),.Y(g17701),.A(I23785));
  NOT NOT1_5971(.VSS(VSS),.VDD(VDD),.Y(I23788),.A(g15901));
  NOT NOT1_5972(.VSS(VSS),.VDD(VDD),.Y(g17704),.A(I23788));
  NOT NOT1_5973(.VSS(VSS),.VDD(VDD),.Y(I23791),.A(g15951));
  NOT NOT1_5974(.VSS(VSS),.VDD(VDD),.Y(g17707),.A(I23791));
  NOT NOT1_5975(.VSS(VSS),.VDD(VDD),.Y(I23794),.A(g15151));
  NOT NOT1_5976(.VSS(VSS),.VDD(VDD),.Y(g17710),.A(I23794));
  NOT NOT1_5977(.VSS(VSS),.VDD(VDD),.Y(g17720),.A(g15853));
  NOT NOT1_5978(.VSS(VSS),.VDD(VDD),.Y(g17724),.A(g13886));
  NOT NOT1_5979(.VSS(VSS),.VDD(VDD),.Y(I23817),.A(g13557));
  NOT NOT1_5980(.VSS(VSS),.VDD(VDD),.Y(g17738),.A(I23817));
  NOT NOT1_5981(.VSS(VSS),.VDD(VDD),.Y(g17741),.A(g13895));
  NOT NOT1_5982(.VSS(VSS),.VDD(VDD),.Y(I23821),.A(g14337));
  NOT NOT1_5983(.VSS(VSS),.VDD(VDD),.Y(g17746),.A(I23821));
  NOT NOT1_5984(.VSS(VSS),.VDD(VDD),.Y(I23824),.A(g14904));
  NOT NOT1_5985(.VSS(VSS),.VDD(VDD),.Y(g17749),.A(I23824));
  NOT NOT1_5986(.VSS(VSS),.VDD(VDD),.Y(I23830),.A(g13558));
  NOT NOT1_5987(.VSS(VSS),.VDD(VDD),.Y(g17755),.A(I23830));
  NOT NOT1_5988(.VSS(VSS),.VDD(VDD),.Y(I23833),.A(g15921));
  NOT NOT1_5989(.VSS(VSS),.VDD(VDD),.Y(g17758),.A(I23833));
  NOT NOT1_5990(.VSS(VSS),.VDD(VDD),.Y(I23836),.A(g13559));
  NOT NOT1_5991(.VSS(VSS),.VDD(VDD),.Y(g17761),.A(I23836));
  NOT NOT1_5992(.VSS(VSS),.VDD(VDD),.Y(I23839),.A(g14985));
  NOT NOT1_5993(.VSS(VSS),.VDD(VDD),.Y(g17764),.A(I23839));
  NOT NOT1_5994(.VSS(VSS),.VDD(VDD),.Y(I23842),.A(g15055));
  NOT NOT1_5995(.VSS(VSS),.VDD(VDD),.Y(g17767),.A(I23842));
  NOT NOT1_5996(.VSS(VSS),.VDD(VDD),.Y(I23845),.A(g16174));
  NOT NOT1_5997(.VSS(VSS),.VDD(VDD),.Y(g17770),.A(I23845));
  NOT NOT1_5998(.VSS(VSS),.VDD(VDD),.Y(I23851),.A(g15930));
  NOT NOT1_5999(.VSS(VSS),.VDD(VDD),.Y(g17776),.A(I23851));
  NOT NOT1_6000(.VSS(VSS),.VDD(VDD),.Y(I23854),.A(g15970));
  NOT NOT1_6001(.VSS(VSS),.VDD(VDD),.Y(g17779),.A(I23854));
  NOT NOT1_6002(.VSS(VSS),.VDD(VDD),.Y(I23857),.A(g13560));
  NOT NOT1_6003(.VSS(VSS),.VDD(VDD),.Y(g17782),.A(I23857));
  NOT NOT1_6004(.VSS(VSS),.VDD(VDD),.Y(I23860),.A(g15932));
  NOT NOT1_6005(.VSS(VSS),.VDD(VDD),.Y(g17785),.A(I23860));
  NOT NOT1_6006(.VSS(VSS),.VDD(VDD),.Y(I23863),.A(g15151));
  NOT NOT1_6007(.VSS(VSS),.VDD(VDD),.Y(g17788),.A(I23863));
  NOT NOT1_6008(.VSS(VSS),.VDD(VDD),.Y(I23866),.A(g15151));
  NOT NOT1_6009(.VSS(VSS),.VDD(VDD),.Y(g17791),.A(I23866));
  NOT NOT1_6010(.VSS(VSS),.VDD(VDD),.Y(I23874),.A(g15797));
  NOT NOT1_6011(.VSS(VSS),.VDD(VDD),.Y(g17799),.A(I23874));
  NOT NOT1_6012(.VSS(VSS),.VDD(VDD),.Y(g17802),.A(g13907));
  NOT NOT1_6013(.VSS(VSS),.VDD(VDD),.Y(I23888),.A(g14685));
  NOT NOT1_6014(.VSS(VSS),.VDD(VDD),.Y(g17815),.A(I23888));
  NOT NOT1_6015(.VSS(VSS),.VDD(VDD),.Y(g17825),.A(g13927));
  NOT NOT1_6016(.VSS(VSS),.VDD(VDD),.Y(I23904),.A(g13561));
  NOT NOT1_6017(.VSS(VSS),.VDD(VDD),.Y(g17839),.A(I23904));
  NOT NOT1_6018(.VSS(VSS),.VDD(VDD),.Y(g17842),.A(g13936));
  NOT NOT1_6019(.VSS(VSS),.VDD(VDD),.Y(I23908),.A(g14337));
  NOT NOT1_6020(.VSS(VSS),.VDD(VDD),.Y(g17847),.A(I23908));
  NOT NOT1_6021(.VSS(VSS),.VDD(VDD),.Y(I23911),.A(g14985));
  NOT NOT1_6022(.VSS(VSS),.VDD(VDD),.Y(g17850),.A(I23911));
  NOT NOT1_6023(.VSS(VSS),.VDD(VDD),.Y(I23917),.A(g13562));
  NOT NOT1_6024(.VSS(VSS),.VDD(VDD),.Y(g17856),.A(I23917));
  NOT NOT1_6025(.VSS(VSS),.VDD(VDD),.Y(I23920),.A(g15950));
  NOT NOT1_6026(.VSS(VSS),.VDD(VDD),.Y(g17859),.A(I23920));
  NOT NOT1_6027(.VSS(VSS),.VDD(VDD),.Y(I23923),.A(g13563));
  NOT NOT1_6028(.VSS(VSS),.VDD(VDD),.Y(g17862),.A(I23923));
  NOT NOT1_6029(.VSS(VSS),.VDD(VDD),.Y(I23926),.A(g15074));
  NOT NOT1_6030(.VSS(VSS),.VDD(VDD),.Y(g17865),.A(I23926));
  NOT NOT1_6031(.VSS(VSS),.VDD(VDD),.Y(I23929),.A(g15151));
  NOT NOT1_6032(.VSS(VSS),.VDD(VDD),.Y(g17868),.A(I23929));
  NOT NOT1_6033(.VSS(VSS),.VDD(VDD),.Y(I23932),.A(g16233));
  NOT NOT1_6034(.VSS(VSS),.VDD(VDD),.Y(g17871),.A(I23932));
  NOT NOT1_6035(.VSS(VSS),.VDD(VDD),.Y(g17878),.A(g15830));
  NOT NOT1_6036(.VSS(VSS),.VDD(VDD),.Y(g17882),.A(g13946));
  NOT NOT1_6037(.VSS(VSS),.VDD(VDD),.Y(g17892),.A(g13954));
  NOT NOT1_6038(.VSS(VSS),.VDD(VDD),.Y(g17893),.A(g14165));
  NOT NOT1_6039(.VSS(VSS),.VDD(VDD),.Y(I23954),.A(g16154));
  NOT NOT1_6040(.VSS(VSS),.VDD(VDD),.Y(g17903),.A(I23954));
  NOT NOT1_6041(.VSS(VSS),.VDD(VDD),.Y(g17914),.A(g13963));
  NOT NOT1_6042(.VSS(VSS),.VDD(VDD),.Y(I23976),.A(g14719));
  NOT NOT1_6043(.VSS(VSS),.VDD(VDD),.Y(g17927),.A(I23976));
  NOT NOT1_6044(.VSS(VSS),.VDD(VDD),.Y(g17937),.A(g13983));
  NOT NOT1_6045(.VSS(VSS),.VDD(VDD),.Y(I23992),.A(g13564));
  NOT NOT1_6046(.VSS(VSS),.VDD(VDD),.Y(g17951),.A(I23992));
  NOT NOT1_6047(.VSS(VSS),.VDD(VDD),.Y(g17954),.A(g13992));
  NOT NOT1_6048(.VSS(VSS),.VDD(VDD),.Y(I23996),.A(g14337));
  NOT NOT1_6049(.VSS(VSS),.VDD(VDD),.Y(g17959),.A(I23996));
  NOT NOT1_6050(.VSS(VSS),.VDD(VDD),.Y(I23999),.A(g15074));
  NOT NOT1_6051(.VSS(VSS),.VDD(VDD),.Y(g17962),.A(I23999));
  NOT NOT1_6052(.VSS(VSS),.VDD(VDD),.Y(g17969),.A(g15841));
  NOT NOT1_6053(.VSS(VSS),.VDD(VDD),.Y(g17974),.A(g14001));
  NOT NOT1_6054(.VSS(VSS),.VDD(VDD),.Y(g17984),.A(g14008));
  NOT NOT1_6055(.VSS(VSS),.VDD(VDD),.Y(g17988),.A(g14685));
  NOT NOT1_6056(.VSS(VSS),.VDD(VDD),.Y(g17991),.A(g14450));
  NOT NOT1_6057(.VSS(VSS),.VDD(VDD),.Y(g17993),.A(g14016));
  NOT NOT1_6058(.VSS(VSS),.VDD(VDD),.Y(g18003),.A(g14024));
  NOT NOT1_6059(.VSS(VSS),.VDD(VDD),.Y(g18004),.A(g14280));
  NOT NOT1_6060(.VSS(VSS),.VDD(VDD),.Y(I24049),.A(g16213));
  NOT NOT1_6061(.VSS(VSS),.VDD(VDD),.Y(g18014),.A(I24049));
  NOT NOT1_6062(.VSS(VSS),.VDD(VDD),.Y(g18025),.A(g14033));
  NOT NOT1_6063(.VSS(VSS),.VDD(VDD),.Y(I24071),.A(g14747));
  NOT NOT1_6064(.VSS(VSS),.VDD(VDD),.Y(g18038),.A(I24071));
  NOT NOT1_6065(.VSS(VSS),.VDD(VDD),.Y(g18048),.A(g14053));
  NOT NOT1_6066(.VSS(VSS),.VDD(VDD),.Y(g18063),.A(g15660));
  NOT NOT1_6067(.VSS(VSS),.VDD(VDD),.Y(g18070),.A(g15854));
  NOT NOT1_6068(.VSS(VSS),.VDD(VDD),.Y(g18074),.A(g14062));
  NOT NOT1_6069(.VSS(VSS),.VDD(VDD),.Y(g18084),.A(g14068));
  NOT NOT1_6070(.VSS(VSS),.VDD(VDD),.Y(g18089),.A(g14355));
  NOT NOT1_6071(.VSS(VSS),.VDD(VDD),.Y(g18091),.A(g14092));
  NOT NOT1_6072(.VSS(VSS),.VDD(VDD),.Y(g18101),.A(g14099));
  NOT NOT1_6073(.VSS(VSS),.VDD(VDD),.Y(g18105),.A(g14719));
  NOT NOT1_6074(.VSS(VSS),.VDD(VDD),.Y(g18108),.A(g14537));
  NOT NOT1_6075(.VSS(VSS),.VDD(VDD),.Y(g18110),.A(g14107));
  NOT NOT1_6076(.VSS(VSS),.VDD(VDD),.Y(g18120),.A(g14115));
  NOT NOT1_6077(.VSS(VSS),.VDD(VDD),.Y(g18121),.A(g14402));
  NOT NOT1_6078(.VSS(VSS),.VDD(VDD),.Y(I24144),.A(g16278));
  NOT NOT1_6079(.VSS(VSS),.VDD(VDD),.Y(g18131),.A(I24144));
  NOT NOT1_6080(.VSS(VSS),.VDD(VDD),.Y(g18142),.A(g14124));
  NOT NOT1_6081(.VSS(VSS),.VDD(VDD),.Y(I24166),.A(g14768));
  NOT NOT1_6082(.VSS(VSS),.VDD(VDD),.Y(g18155),.A(I24166));
  NOT NOT1_6083(.VSS(VSS),.VDD(VDD),.Y(I24171),.A(g16439));
  NOT NOT1_6084(.VSS(VSS),.VDD(VDD),.Y(g18166),.A(I24171));
  NOT NOT1_6085(.VSS(VSS),.VDD(VDD),.Y(g18170),.A(g15877));
  NOT NOT1_6086(.VSS(VSS),.VDD(VDD),.Y(g18174),.A(g14148));
  NOT NOT1_6087(.VSS(VSS),.VDD(VDD),.Y(g18179),.A(g14153));
  NOT NOT1_6088(.VSS(VSS),.VDD(VDD),.Y(g18188),.A(g14252));
  NOT NOT1_6089(.VSS(VSS),.VDD(VDD),.Y(g18190),.A(g14177));
  NOT NOT1_6090(.VSS(VSS),.VDD(VDD),.Y(g18200),.A(g14183));
  NOT NOT1_6091(.VSS(VSS),.VDD(VDD),.Y(g18205),.A(g14467));
  NOT NOT1_6092(.VSS(VSS),.VDD(VDD),.Y(g18207),.A(g14207));
  NOT NOT1_6093(.VSS(VSS),.VDD(VDD),.Y(g18217),.A(g14214));
  NOT NOT1_6094(.VSS(VSS),.VDD(VDD),.Y(g18221),.A(g14747));
  NOT NOT1_6095(.VSS(VSS),.VDD(VDD),.Y(g18224),.A(g14592));
  NOT NOT1_6096(.VSS(VSS),.VDD(VDD),.Y(g18226),.A(g14222));
  NOT NOT1_6097(.VSS(VSS),.VDD(VDD),.Y(g18236),.A(g14230));
  NOT NOT1_6098(.VSS(VSS),.VDD(VDD),.Y(g18237),.A(g14514));
  NOT NOT1_6099(.VSS(VSS),.VDD(VDD),.Y(I24247),.A(g16337));
  NOT NOT1_6100(.VSS(VSS),.VDD(VDD),.Y(g18247),.A(I24247));
  NOT NOT1_6101(.VSS(VSS),.VDD(VDD),.Y(I24258),.A(g16463));
  NOT NOT1_6102(.VSS(VSS),.VDD(VDD),.Y(g18258),.A(I24258));
  NOT NOT1_6103(.VSS(VSS),.VDD(VDD),.Y(g18261),.A(g15719));
  NOT NOT1_6104(.VSS(VSS),.VDD(VDD),.Y(g18265),.A(g14238));
  NOT NOT1_6105(.VSS(VSS),.VDD(VDD),.Y(g18275),.A(g14171));
  NOT NOT1_6106(.VSS(VSS),.VDD(VDD),.Y(I24285),.A(g15992));
  NOT NOT1_6107(.VSS(VSS),.VDD(VDD),.Y(g18278),.A(I24285));
  NOT NOT1_6108(.VSS(VSS),.VDD(VDD),.Y(g18281),.A(g14263));
  NOT NOT1_6109(.VSS(VSS),.VDD(VDD),.Y(g18286),.A(g14268));
  NOT NOT1_6110(.VSS(VSS),.VDD(VDD),.Y(g18295),.A(g14374));
  NOT NOT1_6111(.VSS(VSS),.VDD(VDD),.Y(g18297),.A(g14292));
  NOT NOT1_6112(.VSS(VSS),.VDD(VDD),.Y(g18307),.A(g14298));
  NOT NOT1_6113(.VSS(VSS),.VDD(VDD),.Y(g18312),.A(g14554));
  NOT NOT1_6114(.VSS(VSS),.VDD(VDD),.Y(g18314),.A(g14322));
  NOT NOT1_6115(.VSS(VSS),.VDD(VDD),.Y(g18324),.A(g14329));
  NOT NOT1_6116(.VSS(VSS),.VDD(VDD),.Y(g18328),.A(g14768));
  NOT NOT1_6117(.VSS(VSS),.VDD(VDD),.Y(g18331),.A(g14626));
  NOT NOT1_6118(.VSS(VSS),.VDD(VDD),.Y(I24346),.A(g15873));
  NOT NOT1_6119(.VSS(VSS),.VDD(VDD),.Y(g18334),.A(I24346));
  NOT NOT1_6120(.VSS(VSS),.VDD(VDD),.Y(g18337),.A(g15757));
  NOT NOT1_6121(.VSS(VSS),.VDD(VDD),.Y(g18341),.A(g14342));
  NOT NOT1_6122(.VSS(VSS),.VDD(VDD),.Y(g18351),.A(g13741));
  NOT NOT1_6123(.VSS(VSS),.VDD(VDD),.Y(g18353),.A(g13918));
  NOT NOT1_6124(.VSS(VSS),.VDD(VDD),.Y(I24368),.A(g15990));
  NOT NOT1_6125(.VSS(VSS),.VDD(VDD),.Y(g18355),.A(I24368));
  NOT NOT1_6126(.VSS(VSS),.VDD(VDD),.Y(g18358),.A(g14360));
  NOT NOT1_6127(.VSS(VSS),.VDD(VDD),.Y(g18368),.A(g14286));
  NOT NOT1_6128(.VSS(VSS),.VDD(VDD),.Y(I24394),.A(g15995));
  NOT NOT1_6129(.VSS(VSS),.VDD(VDD),.Y(g18371),.A(I24394));
  NOT NOT1_6130(.VSS(VSS),.VDD(VDD),.Y(g18374),.A(g14385));
  NOT NOT1_6131(.VSS(VSS),.VDD(VDD),.Y(g18379),.A(g14390));
  NOT NOT1_6132(.VSS(VSS),.VDD(VDD),.Y(g18388),.A(g14486));
  NOT NOT1_6133(.VSS(VSS),.VDD(VDD),.Y(g18390),.A(g14414));
  NOT NOT1_6134(.VSS(VSS),.VDD(VDD),.Y(g18400),.A(g14420));
  NOT NOT1_6135(.VSS(VSS),.VDD(VDD),.Y(g18405),.A(g14609));
  NOT NOT1_6136(.VSS(VSS),.VDD(VDD),.Y(g18407),.A(g15959));
  NOT NOT1_6137(.VSS(VSS),.VDD(VDD),.Y(g18414),.A(g15718));
  NOT NOT1_6138(.VSS(VSS),.VDD(VDD),.Y(g18415),.A(g15783));
  NOT NOT1_6139(.VSS(VSS),.VDD(VDD),.Y(g18429),.A(g14831));
  NOT NOT1_6140(.VSS(VSS),.VDD(VDD),.Y(I24459),.A(g13599));
  NOT NOT1_6141(.VSS(VSS),.VDD(VDD),.Y(g18432),.A(I24459));
  NOT NOT1_6142(.VSS(VSS),.VDD(VDD),.Y(g18435),.A(g14359));
  NOT NOT1_6143(.VSS(VSS),.VDD(VDD),.Y(g18436),.A(g14454));
  NOT NOT1_6144(.VSS(VSS),.VDD(VDD),.Y(g18446),.A(g13741));
  NOT NOT1_6145(.VSS(VSS),.VDD(VDD),.Y(g18448),.A(g13974));
  NOT NOT1_6146(.VSS(VSS),.VDD(VDD),.Y(I24481),.A(g15993));
  NOT NOT1_6147(.VSS(VSS),.VDD(VDD),.Y(g18450),.A(I24481));
  NOT NOT1_6148(.VSS(VSS),.VDD(VDD),.Y(g18453),.A(g14472));
  NOT NOT1_6149(.VSS(VSS),.VDD(VDD),.Y(g18463),.A(g14408));
  NOT NOT1_6150(.VSS(VSS),.VDD(VDD),.Y(I24507),.A(g15999));
  NOT NOT1_6151(.VSS(VSS),.VDD(VDD),.Y(g18466),.A(I24507));
  NOT NOT1_6152(.VSS(VSS),.VDD(VDD),.Y(g18469),.A(g14497));
  NOT NOT1_6153(.VSS(VSS),.VDD(VDD),.Y(g18474),.A(g14502));
  NOT NOT1_6154(.VSS(VSS),.VDD(VDD),.Y(g18483),.A(g14573));
  NOT NOT1_6155(.VSS(VSS),.VDD(VDD),.Y(g18485),.A(g15756));
  NOT NOT1_6156(.VSS(VSS),.VDD(VDD),.Y(g18486),.A(g15804));
  NOT NOT1_6157(.VSS(VSS),.VDD(VDD),.Y(g18490),.A(g13565));
  NOT NOT1_6158(.VSS(VSS),.VDD(VDD),.Y(g18502),.A(g14904));
  NOT NOT1_6159(.VSS(VSS),.VDD(VDD),.Y(I24560),.A(g13611));
  NOT NOT1_6160(.VSS(VSS),.VDD(VDD),.Y(g18505),.A(I24560));
  NOT NOT1_6161(.VSS(VSS),.VDD(VDD),.Y(g18508),.A(g14471));
  NOT NOT1_6162(.VSS(VSS),.VDD(VDD),.Y(g18509),.A(g14541));
  NOT NOT1_6163(.VSS(VSS),.VDD(VDD),.Y(g18519),.A(g13741));
  NOT NOT1_6164(.VSS(VSS),.VDD(VDD),.Y(g18521),.A(g14044));
  NOT NOT1_6165(.VSS(VSS),.VDD(VDD),.Y(I24582),.A(g15996));
  NOT NOT1_6166(.VSS(VSS),.VDD(VDD),.Y(g18523),.A(I24582));
  NOT NOT1_6167(.VSS(VSS),.VDD(VDD),.Y(g18526),.A(g14559));
  NOT NOT1_6168(.VSS(VSS),.VDD(VDD),.Y(g18536),.A(g14520));
  NOT NOT1_6169(.VSS(VSS),.VDD(VDD),.Y(I24608),.A(g16006));
  NOT NOT1_6170(.VSS(VSS),.VDD(VDD),.Y(g18539),.A(I24608));
  NOT NOT1_6171(.VSS(VSS),.VDD(VDD),.Y(g18543),.A(g15819));
  NOT NOT1_6172(.VSS(VSS),.VDD(VDD),.Y(g18552),.A(g16154));
  NOT NOT1_6173(.VSS(VSS),.VDD(VDD),.Y(g18554),.A(g13573));
  NOT NOT1_6174(.VSS(VSS),.VDD(VDD),.Y(g18566),.A(g14985));
  NOT NOT1_6175(.VSS(VSS),.VDD(VDD),.Y(I24662),.A(g13621));
  NOT NOT1_6176(.VSS(VSS),.VDD(VDD),.Y(g18569),.A(I24662));
  NOT NOT1_6177(.VSS(VSS),.VDD(VDD),.Y(g18572),.A(g14558));
  NOT NOT1_6178(.VSS(VSS),.VDD(VDD),.Y(g18573),.A(g14596));
  NOT NOT1_6179(.VSS(VSS),.VDD(VDD),.Y(g18583),.A(g13741));
  NOT NOT1_6180(.VSS(VSS),.VDD(VDD),.Y(g18585),.A(g14135));
  NOT NOT1_6181(.VSS(VSS),.VDD(VDD),.Y(I24684),.A(g16000));
  NOT NOT1_6182(.VSS(VSS),.VDD(VDD),.Y(g18587),.A(I24684));
  NOT NOT1_6183(.VSS(VSS),.VDD(VDD),.Y(g18593),.A(g15831));
  NOT NOT1_6184(.VSS(VSS),.VDD(VDD),.Y(g18602),.A(g16213));
  NOT NOT1_6185(.VSS(VSS),.VDD(VDD),.Y(g18604),.A(g13582));
  NOT NOT1_6186(.VSS(VSS),.VDD(VDD),.Y(g18616),.A(g15074));
  NOT NOT1_6187(.VSS(VSS),.VDD(VDD),.Y(I24732),.A(g13633));
  NOT NOT1_6188(.VSS(VSS),.VDD(VDD),.Y(g18619),.A(I24732));
  NOT NOT1_6189(.VSS(VSS),.VDD(VDD),.Y(g18622),.A(g14613));
  NOT NOT1_6190(.VSS(VSS),.VDD(VDD),.Y(g18634),.A(g16278));
  NOT NOT1_6191(.VSS(VSS),.VDD(VDD),.Y(g18636),.A(g13602));
  NOT NOT1_6192(.VSS(VSS),.VDD(VDD),.Y(g18643),.A(g16337));
  NOT NOT1_6193(.VSS(VSS),.VDD(VDD),.Y(g18646),.A(g16341));
  NOT NOT1_6194(.VSS(VSS),.VDD(VDD),.Y(g18656),.A(g14776));
  NOT NOT1_6195(.VSS(VSS),.VDD(VDD),.Y(g18670),.A(g14797));
  NOT NOT1_6196(.VSS(VSS),.VDD(VDD),.Y(g18679),.A(g14811));
  NOT NOT1_6197(.VSS(VSS),.VDD(VDD),.Y(g18691),.A(g14885));
  NOT NOT1_6198(.VSS(VSS),.VDD(VDD),.Y(g18692),.A(g14837));
  NOT NOT1_6199(.VSS(VSS),.VDD(VDD),.Y(g18699),.A(g14849));
  NOT NOT1_6200(.VSS(VSS),.VDD(VDD),.Y(g18708),.A(g14863));
  NOT NOT1_6201(.VSS(VSS),.VDD(VDD),.Y(g18720),.A(g14895));
  NOT NOT1_6202(.VSS(VSS),.VDD(VDD),.Y(g18725),.A(g13865));
  NOT NOT1_6203(.VSS(VSS),.VDD(VDD),.Y(g18727),.A(g14966));
  NOT NOT1_6204(.VSS(VSS),.VDD(VDD),.Y(g18728),.A(g14910));
  NOT NOT1_6205(.VSS(VSS),.VDD(VDD),.Y(g18735),.A(g14922));
  NOT NOT1_6206(.VSS(VSS),.VDD(VDD),.Y(g18744),.A(g14936));
  NOT NOT1_6207(.VSS(VSS),.VDD(VDD),.Y(g18756),.A(g14960));
  NOT NOT1_6208(.VSS(VSS),.VDD(VDD),.Y(g18757),.A(g14963));
  NOT NOT1_6209(.VSS(VSS),.VDD(VDD),.Y(g18758),.A(g14976));
  NOT NOT1_6210(.VSS(VSS),.VDD(VDD),.Y(g18764),.A(g15055));
  NOT NOT1_6211(.VSS(VSS),.VDD(VDD),.Y(g18765),.A(g14991));
  NOT NOT1_6212(.VSS(VSS),.VDD(VDD),.Y(g18772),.A(g15003));
  NOT NOT1_6213(.VSS(VSS),.VDD(VDD),.Y(g18783),.A(g15034));
  NOT NOT1_6214(.VSS(VSS),.VDD(VDD),.Y(g18784),.A(g15037));
  NOT NOT1_6215(.VSS(VSS),.VDD(VDD),.Y(g18785),.A(g15040));
  NOT NOT1_6216(.VSS(VSS),.VDD(VDD),.Y(g18786),.A(g15043));
  NOT NOT1_6217(.VSS(VSS),.VDD(VDD),.Y(g18787),.A(g15049));
  NOT NOT1_6218(.VSS(VSS),.VDD(VDD),.Y(g18788),.A(g15052));
  NOT NOT1_6219(.VSS(VSS),.VDD(VDD),.Y(g18789),.A(g15065));
  NOT NOT1_6220(.VSS(VSS),.VDD(VDD),.Y(g18795),.A(g15151));
  NOT NOT1_6221(.VSS(VSS),.VDD(VDD),.Y(g18796),.A(g15080));
  NOT NOT1_6222(.VSS(VSS),.VDD(VDD),.Y(g18805),.A(g15106));
  NOT NOT1_6223(.VSS(VSS),.VDD(VDD),.Y(g18806),.A(g15109));
  NOT NOT1_6224(.VSS(VSS),.VDD(VDD),.Y(g18807),.A(g15112));
  NOT NOT1_6225(.VSS(VSS),.VDD(VDD),.Y(g18808),.A(g15115));
  NOT NOT1_6226(.VSS(VSS),.VDD(VDD),.Y(g18809),.A(g15130));
  NOT NOT1_6227(.VSS(VSS),.VDD(VDD),.Y(g18810),.A(g15133));
  NOT NOT1_6228(.VSS(VSS),.VDD(VDD),.Y(g18811),.A(g15136));
  NOT NOT1_6229(.VSS(VSS),.VDD(VDD),.Y(g18812),.A(g15139));
  NOT NOT1_6230(.VSS(VSS),.VDD(VDD),.Y(g18813),.A(g15145));
  NOT NOT1_6231(.VSS(VSS),.VDD(VDD),.Y(g18814),.A(g15148));
  NOT NOT1_6232(.VSS(VSS),.VDD(VDD),.Y(g18815),.A(g15161));
  NOT NOT1_6233(.VSS(VSS),.VDD(VDD),.Y(g18822),.A(g15179));
  NOT NOT1_6234(.VSS(VSS),.VDD(VDD),.Y(g18823),.A(g15182));
  NOT NOT1_6235(.VSS(VSS),.VDD(VDD),.Y(g18824),.A(g15185));
  NOT NOT1_6236(.VSS(VSS),.VDD(VDD),.Y(g18825),.A(g15198));
  NOT NOT1_6237(.VSS(VSS),.VDD(VDD),.Y(g18826),.A(g15201));
  NOT NOT1_6238(.VSS(VSS),.VDD(VDD),.Y(g18827),.A(g15204));
  NOT NOT1_6239(.VSS(VSS),.VDD(VDD),.Y(g18828),.A(g15207));
  NOT NOT1_6240(.VSS(VSS),.VDD(VDD),.Y(g18829),.A(g15222));
  NOT NOT1_6241(.VSS(VSS),.VDD(VDD),.Y(g18830),.A(g15225));
  NOT NOT1_6242(.VSS(VSS),.VDD(VDD),.Y(g18831),.A(g15228));
  NOT NOT1_6243(.VSS(VSS),.VDD(VDD),.Y(g18832),.A(g15231));
  NOT NOT1_6244(.VSS(VSS),.VDD(VDD),.Y(g18833),.A(g15237));
  NOT NOT1_6245(.VSS(VSS),.VDD(VDD),.Y(g18834),.A(g15240));
  NOT NOT1_6246(.VSS(VSS),.VDD(VDD),.Y(g18838),.A(g15248));
  NOT NOT1_6247(.VSS(VSS),.VDD(VDD),.Y(g18839),.A(g15251));
  NOT NOT1_6248(.VSS(VSS),.VDD(VDD),.Y(g18840),.A(g15254));
  NOT NOT1_6249(.VSS(VSS),.VDD(VDD),.Y(g18841),.A(g15265));
  NOT NOT1_6250(.VSS(VSS),.VDD(VDD),.Y(g18842),.A(g15268));
  NOT NOT1_6251(.VSS(VSS),.VDD(VDD),.Y(g18843),.A(g15271));
  NOT NOT1_6252(.VSS(VSS),.VDD(VDD),.Y(g18844),.A(g15284));
  NOT NOT1_6253(.VSS(VSS),.VDD(VDD),.Y(g18845),.A(g15287));
  NOT NOT1_6254(.VSS(VSS),.VDD(VDD),.Y(g18846),.A(g15290));
  NOT NOT1_6255(.VSS(VSS),.VDD(VDD),.Y(g18847),.A(g15293));
  NOT NOT1_6256(.VSS(VSS),.VDD(VDD),.Y(g18848),.A(g15308));
  NOT NOT1_6257(.VSS(VSS),.VDD(VDD),.Y(g18849),.A(g15311));
  NOT NOT1_6258(.VSS(VSS),.VDD(VDD),.Y(g18850),.A(g15314));
  NOT NOT1_6259(.VSS(VSS),.VDD(VDD),.Y(g18851),.A(g15317));
  NOT NOT1_6260(.VSS(VSS),.VDD(VDD),.Y(g18853),.A(g15326));
  NOT NOT1_6261(.VSS(VSS),.VDD(VDD),.Y(g18854),.A(g15329));
  NOT NOT1_6262(.VSS(VSS),.VDD(VDD),.Y(g18855),.A(g15332));
  NOT NOT1_6263(.VSS(VSS),.VDD(VDD),.Y(g18856),.A(g15340));
  NOT NOT1_6264(.VSS(VSS),.VDD(VDD),.Y(g18857),.A(g15343));
  NOT NOT1_6265(.VSS(VSS),.VDD(VDD),.Y(g18858),.A(g15346));
  NOT NOT1_6266(.VSS(VSS),.VDD(VDD),.Y(g18859),.A(g15357));
  NOT NOT1_6267(.VSS(VSS),.VDD(VDD),.Y(g18860),.A(g15360));
  NOT NOT1_6268(.VSS(VSS),.VDD(VDD),.Y(g18861),.A(g15363));
  NOT NOT1_6269(.VSS(VSS),.VDD(VDD),.Y(g18862),.A(g15376));
  NOT NOT1_6270(.VSS(VSS),.VDD(VDD),.Y(g18863),.A(g15379));
  NOT NOT1_6271(.VSS(VSS),.VDD(VDD),.Y(g18864),.A(g15382));
  NOT NOT1_6272(.VSS(VSS),.VDD(VDD),.Y(g18865),.A(g15385));
  NOT NOT1_6273(.VSS(VSS),.VDD(VDD),.Y(I24894),.A(g14797));
  NOT NOT1_6274(.VSS(VSS),.VDD(VDD),.Y(g18869),.A(I24894));
  NOT NOT1_6275(.VSS(VSS),.VDD(VDD),.Y(g18870),.A(g15393));
  NOT NOT1_6276(.VSS(VSS),.VDD(VDD),.Y(g18871),.A(g15396));
  NOT NOT1_6277(.VSS(VSS),.VDD(VDD),.Y(g18872),.A(g15399));
  NOT NOT1_6278(.VSS(VSS),.VDD(VDD),.Y(g18873),.A(g15404));
  NOT NOT1_6279(.VSS(VSS),.VDD(VDD),.Y(g18874),.A(g15412));
  NOT NOT1_6280(.VSS(VSS),.VDD(VDD),.Y(g18875),.A(g15415));
  NOT NOT1_6281(.VSS(VSS),.VDD(VDD),.Y(g18876),.A(g15418));
  NOT NOT1_6282(.VSS(VSS),.VDD(VDD),.Y(g18877),.A(g15426));
  NOT NOT1_6283(.VSS(VSS),.VDD(VDD),.Y(g18878),.A(g15429));
  NOT NOT1_6284(.VSS(VSS),.VDD(VDD),.Y(g18879),.A(g15432));
  NOT NOT1_6285(.VSS(VSS),.VDD(VDD),.Y(g18880),.A(g15443));
  NOT NOT1_6286(.VSS(VSS),.VDD(VDD),.Y(g18881),.A(g15446));
  NOT NOT1_6287(.VSS(VSS),.VDD(VDD),.Y(g18882),.A(g15449));
  NOT NOT1_6288(.VSS(VSS),.VDD(VDD),.Y(g18884),.A(g13469));
  NOT NOT1_6289(.VSS(VSS),.VDD(VDD),.Y(I24913),.A(g15800));
  NOT NOT1_6290(.VSS(VSS),.VDD(VDD),.Y(g18886),.A(I24913));
  NOT NOT1_6291(.VSS(VSS),.VDD(VDD),.Y(I24916),.A(g14776));
  NOT NOT1_6292(.VSS(VSS),.VDD(VDD),.Y(g18890),.A(I24916));
  NOT NOT1_6293(.VSS(VSS),.VDD(VDD),.Y(g18891),.A(g15461));
  NOT NOT1_6294(.VSS(VSS),.VDD(VDD),.Y(g18892),.A(g15464));
  NOT NOT1_6295(.VSS(VSS),.VDD(VDD),.Y(g18893),.A(g15467));
  NOT NOT1_6296(.VSS(VSS),.VDD(VDD),.Y(g18894),.A(g15471));
  NOT NOT1_6297(.VSS(VSS),.VDD(VDD),.Y(I24923),.A(g14849));
  NOT NOT1_6298(.VSS(VSS),.VDD(VDD),.Y(g18895),.A(I24923));
  NOT NOT1_6299(.VSS(VSS),.VDD(VDD),.Y(g18896),.A(g15477));
  NOT NOT1_6300(.VSS(VSS),.VDD(VDD),.Y(g18897),.A(g15480));
  NOT NOT1_6301(.VSS(VSS),.VDD(VDD),.Y(g18898),.A(g15483));
  NOT NOT1_6302(.VSS(VSS),.VDD(VDD),.Y(g18899),.A(g15488));
  NOT NOT1_6303(.VSS(VSS),.VDD(VDD),.Y(g18900),.A(g15496));
  NOT NOT1_6304(.VSS(VSS),.VDD(VDD),.Y(g18901),.A(g15499));
  NOT NOT1_6305(.VSS(VSS),.VDD(VDD),.Y(g18902),.A(g15502));
  NOT NOT1_6306(.VSS(VSS),.VDD(VDD),.Y(g18903),.A(g15510));
  NOT NOT1_6307(.VSS(VSS),.VDD(VDD),.Y(g18904),.A(g15513));
  NOT NOT1_6308(.VSS(VSS),.VDD(VDD),.Y(g18905),.A(g15516));
  NOT NOT1_6309(.VSS(VSS),.VDD(VDD),.Y(g18908),.A(g15521));
  NOT NOT1_6310(.VSS(VSS),.VDD(VDD),.Y(g18909),.A(g15528));
  NOT NOT1_6311(.VSS(VSS),.VDD(VDD),.Y(g18910),.A(g15531));
  NOT NOT1_6312(.VSS(VSS),.VDD(VDD),.Y(g18911),.A(g15534));
  NOT NOT1_6313(.VSS(VSS),.VDD(VDD),.Y(g18912),.A(g15537));
  NOT NOT1_6314(.VSS(VSS),.VDD(VDD),.Y(I24943),.A(g14811));
  NOT NOT1_6315(.VSS(VSS),.VDD(VDD),.Y(g18913),.A(I24943));
  NOT NOT1_6316(.VSS(VSS),.VDD(VDD),.Y(g18914),.A(g15547));
  NOT NOT1_6317(.VSS(VSS),.VDD(VDD),.Y(g18915),.A(g15550));
  NOT NOT1_6318(.VSS(VSS),.VDD(VDD),.Y(g18916),.A(g15553));
  NOT NOT1_6319(.VSS(VSS),.VDD(VDD),.Y(g18917),.A(g15557));
  NOT NOT1_6320(.VSS(VSS),.VDD(VDD),.Y(I24950),.A(g14922));
  NOT NOT1_6321(.VSS(VSS),.VDD(VDD),.Y(g18918),.A(I24950));
  NOT NOT1_6322(.VSS(VSS),.VDD(VDD),.Y(g18919),.A(g15563));
  NOT NOT1_6323(.VSS(VSS),.VDD(VDD),.Y(g18920),.A(g15566));
  NOT NOT1_6324(.VSS(VSS),.VDD(VDD),.Y(g18921),.A(g15569));
  NOT NOT1_6325(.VSS(VSS),.VDD(VDD),.Y(g18922),.A(g15574));
  NOT NOT1_6326(.VSS(VSS),.VDD(VDD),.Y(g18923),.A(g15582));
  NOT NOT1_6327(.VSS(VSS),.VDD(VDD),.Y(g18924),.A(g15585));
  NOT NOT1_6328(.VSS(VSS),.VDD(VDD),.Y(g18925),.A(g15588));
  NOT NOT1_6329(.VSS(VSS),.VDD(VDD),.Y(g18926),.A(g15596));
  NOT NOT1_6330(.VSS(VSS),.VDD(VDD),.Y(g18927),.A(g15599));
  NOT NOT1_6331(.VSS(VSS),.VDD(VDD),.Y(g18928),.A(g15606));
  NOT NOT1_6332(.VSS(VSS),.VDD(VDD),.Y(g18929),.A(g15609));
  NOT NOT1_6333(.VSS(VSS),.VDD(VDD),.Y(g18930),.A(g15612));
  NOT NOT1_6334(.VSS(VSS),.VDD(VDD),.Y(g18931),.A(g15615));
  NOT NOT1_6335(.VSS(VSS),.VDD(VDD),.Y(I24966),.A(g14863));
  NOT NOT1_6336(.VSS(VSS),.VDD(VDD),.Y(g18932),.A(I24966));
  NOT NOT1_6337(.VSS(VSS),.VDD(VDD),.Y(g18933),.A(g15625));
  NOT NOT1_6338(.VSS(VSS),.VDD(VDD),.Y(g18934),.A(g15628));
  NOT NOT1_6339(.VSS(VSS),.VDD(VDD),.Y(g18935),.A(g15631));
  NOT NOT1_6340(.VSS(VSS),.VDD(VDD),.Y(g18936),.A(g15635));
  NOT NOT1_6341(.VSS(VSS),.VDD(VDD),.Y(I24973),.A(g15003));
  NOT NOT1_6342(.VSS(VSS),.VDD(VDD),.Y(g18937),.A(I24973));
  NOT NOT1_6343(.VSS(VSS),.VDD(VDD),.Y(g18938),.A(g15641));
  NOT NOT1_6344(.VSS(VSS),.VDD(VDD),.Y(g18939),.A(g15644));
  NOT NOT1_6345(.VSS(VSS),.VDD(VDD),.Y(g18940),.A(g15647));
  NOT NOT1_6346(.VSS(VSS),.VDD(VDD),.Y(g18941),.A(g15652));
  NOT NOT1_6347(.VSS(VSS),.VDD(VDD),.Y(g18943),.A(g15655));
  NOT NOT1_6348(.VSS(VSS),.VDD(VDD),.Y(I24982),.A(g14347));
  NOT NOT1_6349(.VSS(VSS),.VDD(VDD),.Y(g18944),.A(I24982));
  NOT NOT1_6350(.VSS(VSS),.VDD(VDD),.Y(g18945),.A(g15667));
  NOT NOT1_6351(.VSS(VSS),.VDD(VDD),.Y(g18946),.A(g15672));
  NOT NOT1_6352(.VSS(VSS),.VDD(VDD),.Y(g18947),.A(g15675));
  NOT NOT1_6353(.VSS(VSS),.VDD(VDD),.Y(g18948),.A(g15682));
  NOT NOT1_6354(.VSS(VSS),.VDD(VDD),.Y(g18949),.A(g15685));
  NOT NOT1_6355(.VSS(VSS),.VDD(VDD),.Y(g18950),.A(g15688));
  NOT NOT1_6356(.VSS(VSS),.VDD(VDD),.Y(g18951),.A(g15691));
  NOT NOT1_6357(.VSS(VSS),.VDD(VDD),.Y(I24992),.A(g14936));
  NOT NOT1_6358(.VSS(VSS),.VDD(VDD),.Y(g18952),.A(I24992));
  NOT NOT1_6359(.VSS(VSS),.VDD(VDD),.Y(g18953),.A(g15701));
  NOT NOT1_6360(.VSS(VSS),.VDD(VDD),.Y(g18954),.A(g15704));
  NOT NOT1_6361(.VSS(VSS),.VDD(VDD),.Y(g18955),.A(g15707));
  NOT NOT1_6362(.VSS(VSS),.VDD(VDD),.Y(g18956),.A(g15711));
  NOT NOT1_6363(.VSS(VSS),.VDD(VDD),.Y(g18958),.A(g15714));
  NOT NOT1_6364(.VSS(VSS),.VDD(VDD),.Y(I25001),.A(g14244));
  NOT NOT1_6365(.VSS(VSS),.VDD(VDD),.Y(g18959),.A(I25001));
  NOT NOT1_6366(.VSS(VSS),.VDD(VDD),.Y(I25004),.A(g14459));
  NOT NOT1_6367(.VSS(VSS),.VDD(VDD),.Y(g18960),.A(I25004));
  NOT NOT1_6368(.VSS(VSS),.VDD(VDD),.Y(g18961),.A(g15726));
  NOT NOT1_6369(.VSS(VSS),.VDD(VDD),.Y(g18962),.A(g15731));
  NOT NOT1_6370(.VSS(VSS),.VDD(VDD),.Y(g18963),.A(g15734));
  NOT NOT1_6371(.VSS(VSS),.VDD(VDD),.Y(g18964),.A(g15741));
  NOT NOT1_6372(.VSS(VSS),.VDD(VDD),.Y(g18965),.A(g15744));
  NOT NOT1_6373(.VSS(VSS),.VDD(VDD),.Y(g18966),.A(g15747));
  NOT NOT1_6374(.VSS(VSS),.VDD(VDD),.Y(g18967),.A(g15750));
  NOT NOT1_6375(.VSS(VSS),.VDD(VDD),.Y(I25015),.A(g14158));
  NOT NOT1_6376(.VSS(VSS),.VDD(VDD),.Y(g18969),.A(I25015));
  NOT NOT1_6377(.VSS(VSS),.VDD(VDD),.Y(I25018),.A(g14366));
  NOT NOT1_6378(.VSS(VSS),.VDD(VDD),.Y(g18970),.A(I25018));
  NOT NOT1_6379(.VSS(VSS),.VDD(VDD),.Y(I25021),.A(g14546));
  NOT NOT1_6380(.VSS(VSS),.VDD(VDD),.Y(g18971),.A(I25021));
  NOT NOT1_6381(.VSS(VSS),.VDD(VDD),.Y(g18972),.A(g15766));
  NOT NOT1_6382(.VSS(VSS),.VDD(VDD),.Y(g18973),.A(g15771));
  NOT NOT1_6383(.VSS(VSS),.VDD(VDD),.Y(g18974),.A(g15774));
  NOT NOT1_6384(.VSS(VSS),.VDD(VDD),.Y(g18976),.A(g15777));
  NOT NOT1_6385(.VSS(VSS),.VDD(VDD),.Y(I25037),.A(g14071));
  NOT NOT1_6386(.VSS(VSS),.VDD(VDD),.Y(g18981),.A(I25037));
  NOT NOT1_6387(.VSS(VSS),.VDD(VDD),.Y(I25041),.A(g14895));
  NOT NOT1_6388(.VSS(VSS),.VDD(VDD),.Y(g18983),.A(I25041));
  NOT NOT1_6389(.VSS(VSS),.VDD(VDD),.Y(I25044),.A(g14273));
  NOT NOT1_6390(.VSS(VSS),.VDD(VDD),.Y(g18984),.A(I25044));
  NOT NOT1_6391(.VSS(VSS),.VDD(VDD),.Y(I25047),.A(g14478));
  NOT NOT1_6392(.VSS(VSS),.VDD(VDD),.Y(g18985),.A(I25047));
  NOT NOT1_6393(.VSS(VSS),.VDD(VDD),.Y(I25050),.A(g14601));
  NOT NOT1_6394(.VSS(VSS),.VDD(VDD),.Y(g18986),.A(I25050));
  NOT NOT1_6395(.VSS(VSS),.VDD(VDD),.Y(g18987),.A(g15794));
  NOT NOT1_6396(.VSS(VSS),.VDD(VDD),.Y(I25054),.A(g14837));
  NOT NOT1_6397(.VSS(VSS),.VDD(VDD),.Y(g18988),.A(I25054));
  NOT NOT1_6398(.VSS(VSS),.VDD(VDD),.Y(I25057),.A(g14186));
  NOT NOT1_6399(.VSS(VSS),.VDD(VDD),.Y(g18989),.A(I25057));
  NOT NOT1_6400(.VSS(VSS),.VDD(VDD),.Y(I25061),.A(g14976));
  NOT NOT1_6401(.VSS(VSS),.VDD(VDD),.Y(g18991),.A(I25061));
  NOT NOT1_6402(.VSS(VSS),.VDD(VDD),.Y(I25064),.A(g14395));
  NOT NOT1_6403(.VSS(VSS),.VDD(VDD),.Y(g18992),.A(I25064));
  NOT NOT1_6404(.VSS(VSS),.VDD(VDD),.Y(I25067),.A(g14565));
  NOT NOT1_6405(.VSS(VSS),.VDD(VDD),.Y(g18993),.A(I25067));
  NOT NOT1_6406(.VSS(VSS),.VDD(VDD),.Y(I25071),.A(g14910));
  NOT NOT1_6407(.VSS(VSS),.VDD(VDD),.Y(g18995),.A(I25071));
  NOT NOT1_6408(.VSS(VSS),.VDD(VDD),.Y(I25074),.A(g14301));
  NOT NOT1_6409(.VSS(VSS),.VDD(VDD),.Y(g18996),.A(I25074));
  NOT NOT1_6410(.VSS(VSS),.VDD(VDD),.Y(I25078),.A(g15065));
  NOT NOT1_6411(.VSS(VSS),.VDD(VDD),.Y(g18998),.A(I25078));
  NOT NOT1_6412(.VSS(VSS),.VDD(VDD),.Y(I25081),.A(g14507));
  NOT NOT1_6413(.VSS(VSS),.VDD(VDD),.Y(g18999),.A(I25081));
  NOT NOT1_6414(.VSS(VSS),.VDD(VDD),.Y(I25084),.A(g14885));
  NOT NOT1_6415(.VSS(VSS),.VDD(VDD),.Y(g19000),.A(I25084));
  NOT NOT1_6416(.VSS(VSS),.VDD(VDD),.Y(g19001),.A(g14071));
  NOT NOT1_6417(.VSS(VSS),.VDD(VDD),.Y(I25089),.A(g14991));
  NOT NOT1_6418(.VSS(VSS),.VDD(VDD),.Y(g19008),.A(I25089));
  NOT NOT1_6419(.VSS(VSS),.VDD(VDD),.Y(I25092),.A(g14423));
  NOT NOT1_6420(.VSS(VSS),.VDD(VDD),.Y(g19009),.A(I25092));
  NOT NOT1_6421(.VSS(VSS),.VDD(VDD),.Y(I25096),.A(g15161));
  NOT NOT1_6422(.VSS(VSS),.VDD(VDD),.Y(g19011),.A(I25096));
  NOT NOT1_6423(.VSS(VSS),.VDD(VDD),.Y(I25099),.A(g19000));
  NOT NOT1_6424(.VSS(VSS),.VDD(VDD),.Y(g19012),.A(I25099));
  NOT NOT1_6425(.VSS(VSS),.VDD(VDD),.Y(I25102),.A(g18944));
  NOT NOT1_6426(.VSS(VSS),.VDD(VDD),.Y(g19013),.A(I25102));
  NOT NOT1_6427(.VSS(VSS),.VDD(VDD),.Y(I25105),.A(g18959));
  NOT NOT1_6428(.VSS(VSS),.VDD(VDD),.Y(g19014),.A(I25105));
  NOT NOT1_6429(.VSS(VSS),.VDD(VDD),.Y(I25108),.A(g18969));
  NOT NOT1_6430(.VSS(VSS),.VDD(VDD),.Y(g19015),.A(I25108));
  NOT NOT1_6431(.VSS(VSS),.VDD(VDD),.Y(I25111),.A(g18981));
  NOT NOT1_6432(.VSS(VSS),.VDD(VDD),.Y(g19016),.A(I25111));
  NOT NOT1_6433(.VSS(VSS),.VDD(VDD),.Y(I25114),.A(g18983));
  NOT NOT1_6434(.VSS(VSS),.VDD(VDD),.Y(g19017),.A(I25114));
  NOT NOT1_6435(.VSS(VSS),.VDD(VDD),.Y(I25117),.A(g18988));
  NOT NOT1_6436(.VSS(VSS),.VDD(VDD),.Y(g19018),.A(I25117));
  NOT NOT1_6437(.VSS(VSS),.VDD(VDD),.Y(I25120),.A(g18869));
  NOT NOT1_6438(.VSS(VSS),.VDD(VDD),.Y(g19019),.A(I25120));
  NOT NOT1_6439(.VSS(VSS),.VDD(VDD),.Y(I25123),.A(g18890));
  NOT NOT1_6440(.VSS(VSS),.VDD(VDD),.Y(g19020),.A(I25123));
  NOT NOT1_6441(.VSS(VSS),.VDD(VDD),.Y(I25126),.A(g16858));
  NOT NOT1_6442(.VSS(VSS),.VDD(VDD),.Y(g19021),.A(I25126));
  NOT NOT1_6443(.VSS(VSS),.VDD(VDD),.Y(I25129),.A(g16813));
  NOT NOT1_6444(.VSS(VSS),.VDD(VDD),.Y(g19022),.A(I25129));
  NOT NOT1_6445(.VSS(VSS),.VDD(VDD),.Y(I25132),.A(g16862));
  NOT NOT1_6446(.VSS(VSS),.VDD(VDD),.Y(g19023),.A(I25132));
  NOT NOT1_6447(.VSS(VSS),.VDD(VDD),.Y(I25135),.A(g16506));
  NOT NOT1_6448(.VSS(VSS),.VDD(VDD),.Y(g19024),.A(I25135));
  NOT NOT1_6449(.VSS(VSS),.VDD(VDD),.Y(I25138),.A(g18960));
  NOT NOT1_6450(.VSS(VSS),.VDD(VDD),.Y(g19025),.A(I25138));
  NOT NOT1_6451(.VSS(VSS),.VDD(VDD),.Y(I25141),.A(g18970));
  NOT NOT1_6452(.VSS(VSS),.VDD(VDD),.Y(g19026),.A(I25141));
  NOT NOT1_6453(.VSS(VSS),.VDD(VDD),.Y(I25144),.A(g18984));
  NOT NOT1_6454(.VSS(VSS),.VDD(VDD),.Y(g19027),.A(I25144));
  NOT NOT1_6455(.VSS(VSS),.VDD(VDD),.Y(I25147),.A(g18989));
  NOT NOT1_6456(.VSS(VSS),.VDD(VDD),.Y(g19028),.A(I25147));
  NOT NOT1_6457(.VSS(VSS),.VDD(VDD),.Y(I25150),.A(g18991));
  NOT NOT1_6458(.VSS(VSS),.VDD(VDD),.Y(g19029),.A(I25150));
  NOT NOT1_6459(.VSS(VSS),.VDD(VDD),.Y(I25153),.A(g18995));
  NOT NOT1_6460(.VSS(VSS),.VDD(VDD),.Y(g19030),.A(I25153));
  NOT NOT1_6461(.VSS(VSS),.VDD(VDD),.Y(I25156),.A(g18895));
  NOT NOT1_6462(.VSS(VSS),.VDD(VDD),.Y(g19031),.A(I25156));
  NOT NOT1_6463(.VSS(VSS),.VDD(VDD),.Y(I25159),.A(g18913));
  NOT NOT1_6464(.VSS(VSS),.VDD(VDD),.Y(g19032),.A(I25159));
  NOT NOT1_6465(.VSS(VSS),.VDD(VDD),.Y(I25162),.A(g16863));
  NOT NOT1_6466(.VSS(VSS),.VDD(VDD),.Y(g19033),.A(I25162));
  NOT NOT1_6467(.VSS(VSS),.VDD(VDD),.Y(I25165),.A(g16831));
  NOT NOT1_6468(.VSS(VSS),.VDD(VDD),.Y(g19034),.A(I25165));
  NOT NOT1_6469(.VSS(VSS),.VDD(VDD),.Y(I25168),.A(g16877));
  NOT NOT1_6470(.VSS(VSS),.VDD(VDD),.Y(g19035),.A(I25168));
  NOT NOT1_6471(.VSS(VSS),.VDD(VDD),.Y(I25171),.A(g16528));
  NOT NOT1_6472(.VSS(VSS),.VDD(VDD),.Y(g19036),.A(I25171));
  NOT NOT1_6473(.VSS(VSS),.VDD(VDD),.Y(I25174),.A(g18971));
  NOT NOT1_6474(.VSS(VSS),.VDD(VDD),.Y(g19037),.A(I25174));
  NOT NOT1_6475(.VSS(VSS),.VDD(VDD),.Y(I25177),.A(g18985));
  NOT NOT1_6476(.VSS(VSS),.VDD(VDD),.Y(g19038),.A(I25177));
  NOT NOT1_6477(.VSS(VSS),.VDD(VDD),.Y(I25180),.A(g18992));
  NOT NOT1_6478(.VSS(VSS),.VDD(VDD),.Y(g19039),.A(I25180));
  NOT NOT1_6479(.VSS(VSS),.VDD(VDD),.Y(I25183),.A(g18996));
  NOT NOT1_6480(.VSS(VSS),.VDD(VDD),.Y(g19040),.A(I25183));
  NOT NOT1_6481(.VSS(VSS),.VDD(VDD),.Y(I25186),.A(g18998));
  NOT NOT1_6482(.VSS(VSS),.VDD(VDD),.Y(g19041),.A(I25186));
  NOT NOT1_6483(.VSS(VSS),.VDD(VDD),.Y(I25189),.A(g19008));
  NOT NOT1_6484(.VSS(VSS),.VDD(VDD),.Y(g19042),.A(I25189));
  NOT NOT1_6485(.VSS(VSS),.VDD(VDD),.Y(I25192),.A(g18918));
  NOT NOT1_6486(.VSS(VSS),.VDD(VDD),.Y(g19043),.A(I25192));
  NOT NOT1_6487(.VSS(VSS),.VDD(VDD),.Y(I25195),.A(g18932));
  NOT NOT1_6488(.VSS(VSS),.VDD(VDD),.Y(g19044),.A(I25195));
  NOT NOT1_6489(.VSS(VSS),.VDD(VDD),.Y(I25198),.A(g16878));
  NOT NOT1_6490(.VSS(VSS),.VDD(VDD),.Y(g19045),.A(I25198));
  NOT NOT1_6491(.VSS(VSS),.VDD(VDD),.Y(I25201),.A(g16843));
  NOT NOT1_6492(.VSS(VSS),.VDD(VDD),.Y(g19046),.A(I25201));
  NOT NOT1_6493(.VSS(VSS),.VDD(VDD),.Y(I25204),.A(g16905));
  NOT NOT1_6494(.VSS(VSS),.VDD(VDD),.Y(g19047),.A(I25204));
  NOT NOT1_6495(.VSS(VSS),.VDD(VDD),.Y(I25207),.A(g16559));
  NOT NOT1_6496(.VSS(VSS),.VDD(VDD),.Y(g19048),.A(I25207));
  NOT NOT1_6497(.VSS(VSS),.VDD(VDD),.Y(I25210),.A(g18986));
  NOT NOT1_6498(.VSS(VSS),.VDD(VDD),.Y(g19049),.A(I25210));
  NOT NOT1_6499(.VSS(VSS),.VDD(VDD),.Y(I25213),.A(g18993));
  NOT NOT1_6500(.VSS(VSS),.VDD(VDD),.Y(g19050),.A(I25213));
  NOT NOT1_6501(.VSS(VSS),.VDD(VDD),.Y(I25216),.A(g18999));
  NOT NOT1_6502(.VSS(VSS),.VDD(VDD),.Y(g19051),.A(I25216));
  NOT NOT1_6503(.VSS(VSS),.VDD(VDD),.Y(I25219),.A(g19009));
  NOT NOT1_6504(.VSS(VSS),.VDD(VDD),.Y(g19052),.A(I25219));
  NOT NOT1_6505(.VSS(VSS),.VDD(VDD),.Y(I25222),.A(g19011));
  NOT NOT1_6506(.VSS(VSS),.VDD(VDD),.Y(g19053),.A(I25222));
  NOT NOT1_6507(.VSS(VSS),.VDD(VDD),.Y(I25225),.A(g16514));
  NOT NOT1_6508(.VSS(VSS),.VDD(VDD),.Y(g19054),.A(I25225));
  NOT NOT1_6509(.VSS(VSS),.VDD(VDD),.Y(I25228),.A(g18937));
  NOT NOT1_6510(.VSS(VSS),.VDD(VDD),.Y(g19055),.A(I25228));
  NOT NOT1_6511(.VSS(VSS),.VDD(VDD),.Y(I25231),.A(g18952));
  NOT NOT1_6512(.VSS(VSS),.VDD(VDD),.Y(g19056),.A(I25231));
  NOT NOT1_6513(.VSS(VSS),.VDD(VDD),.Y(I25234),.A(g16906));
  NOT NOT1_6514(.VSS(VSS),.VDD(VDD),.Y(g19057),.A(I25234));
  NOT NOT1_6515(.VSS(VSS),.VDD(VDD),.Y(I25237),.A(g16849));
  NOT NOT1_6516(.VSS(VSS),.VDD(VDD),.Y(g19058),.A(I25237));
  NOT NOT1_6517(.VSS(VSS),.VDD(VDD),.Y(I25240),.A(g16934));
  NOT NOT1_6518(.VSS(VSS),.VDD(VDD),.Y(g19059),.A(I25240));
  NOT NOT1_6519(.VSS(VSS),.VDD(VDD),.Y(I25243),.A(g17227));
  NOT NOT1_6520(.VSS(VSS),.VDD(VDD),.Y(g19060),.A(I25243));
  NOT NOT1_6521(.VSS(VSS),.VDD(VDD),.Y(I25246),.A(g17233));
  NOT NOT1_6522(.VSS(VSS),.VDD(VDD),.Y(g19061),.A(I25246));
  NOT NOT1_6523(.VSS(VSS),.VDD(VDD),.Y(I25249),.A(g17300));
  NOT NOT1_6524(.VSS(VSS),.VDD(VDD),.Y(g19062),.A(I25249));
  NOT NOT1_6525(.VSS(VSS),.VDD(VDD),.Y(I25253),.A(g17124));
  NOT NOT1_6526(.VSS(VSS),.VDD(VDD),.Y(g19064),.A(I25253));
  NOT NOT1_6527(.VSS(VSS),.VDD(VDD),.Y(g19070),.A(g18583));
  NOT NOT1_6528(.VSS(VSS),.VDD(VDD),.Y(I25258),.A(g16974));
  NOT NOT1_6529(.VSS(VSS),.VDD(VDD),.Y(g19075),.A(I25258));
  NOT NOT1_6530(.VSS(VSS),.VDD(VDD),.Y(g19078),.A(g18619));
  NOT NOT1_6531(.VSS(VSS),.VDD(VDD),.Y(I25264),.A(g17151));
  NOT NOT1_6532(.VSS(VSS),.VDD(VDD),.Y(g19081),.A(I25264));
  NOT NOT1_6533(.VSS(VSS),.VDD(VDD),.Y(I25272),.A(g17051));
  NOT NOT1_6534(.VSS(VSS),.VDD(VDD),.Y(g19091),.A(I25272));
  NOT NOT1_6535(.VSS(VSS),.VDD(VDD),.Y(g19096),.A(g18980));
  NOT NOT1_6536(.VSS(VSS),.VDD(VDD),.Y(I25283),.A(g17086));
  NOT NOT1_6537(.VSS(VSS),.VDD(VDD),.Y(g19098),.A(I25283));
  NOT NOT1_6538(.VSS(VSS),.VDD(VDD),.Y(I25294),.A(g17124));
  NOT NOT1_6539(.VSS(VSS),.VDD(VDD),.Y(g19105),.A(I25294));
  NOT NOT1_6540(.VSS(VSS),.VDD(VDD),.Y(I25303),.A(g17151));
  NOT NOT1_6541(.VSS(VSS),.VDD(VDD),.Y(g19110),.A(I25303));
  NOT NOT1_6542(.VSS(VSS),.VDD(VDD),.Y(I25308),.A(g16867));
  NOT NOT1_6543(.VSS(VSS),.VDD(VDD),.Y(g19113),.A(I25308));
  NOT NOT1_6544(.VSS(VSS),.VDD(VDD),.Y(I25315),.A(g16895));
  NOT NOT1_6545(.VSS(VSS),.VDD(VDD),.Y(g19118),.A(I25315));
  NOT NOT1_6546(.VSS(VSS),.VDD(VDD),.Y(I25320),.A(g16924));
  NOT NOT1_6547(.VSS(VSS),.VDD(VDD),.Y(g19125),.A(I25320));
  NOT NOT1_6548(.VSS(VSS),.VDD(VDD),.Y(I25325),.A(g16954));
  NOT NOT1_6549(.VSS(VSS),.VDD(VDD),.Y(g19132),.A(I25325));
  NOT NOT1_6550(.VSS(VSS),.VDD(VDD),.Y(I25334),.A(g17645));
  NOT NOT1_6551(.VSS(VSS),.VDD(VDD),.Y(g19145),.A(I25334));
  NOT NOT1_6552(.VSS(VSS),.VDD(VDD),.Y(I25338),.A(g17746));
  NOT NOT1_6553(.VSS(VSS),.VDD(VDD),.Y(g19147),.A(I25338));
  NOT NOT1_6554(.VSS(VSS),.VDD(VDD),.Y(I25344),.A(g17847));
  NOT NOT1_6555(.VSS(VSS),.VDD(VDD),.Y(g19151),.A(I25344));
  NOT NOT1_6556(.VSS(VSS),.VDD(VDD),.Y(I25351),.A(g17959));
  NOT NOT1_6557(.VSS(VSS),.VDD(VDD),.Y(g19156),.A(I25351));
  NOT NOT1_6558(.VSS(VSS),.VDD(VDD),.Y(I25355),.A(g18669));
  NOT NOT1_6559(.VSS(VSS),.VDD(VDD),.Y(g19158),.A(I25355));
  NOT NOT1_6560(.VSS(VSS),.VDD(VDD),.Y(I25358),.A(g18678));
  NOT NOT1_6561(.VSS(VSS),.VDD(VDD),.Y(g19159),.A(I25358));
  NOT NOT1_6562(.VSS(VSS),.VDD(VDD),.Y(I25365),.A(g18707));
  NOT NOT1_6563(.VSS(VSS),.VDD(VDD),.Y(g19164),.A(I25365));
  NOT NOT1_6564(.VSS(VSS),.VDD(VDD),.Y(I25371),.A(g18719));
  NOT NOT1_6565(.VSS(VSS),.VDD(VDD),.Y(g19168),.A(I25371));
  NOT NOT1_6566(.VSS(VSS),.VDD(VDD),.Y(I25374),.A(g18726));
  NOT NOT1_6567(.VSS(VSS),.VDD(VDD),.Y(g19169),.A(I25374));
  NOT NOT1_6568(.VSS(VSS),.VDD(VDD),.Y(I25377),.A(g18743));
  NOT NOT1_6569(.VSS(VSS),.VDD(VDD),.Y(g19170),.A(I25377));
  NOT NOT1_6570(.VSS(VSS),.VDD(VDD),.Y(I25383),.A(g18755));
  NOT NOT1_6571(.VSS(VSS),.VDD(VDD),.Y(g19174),.A(I25383));
  NOT NOT1_6572(.VSS(VSS),.VDD(VDD),.Y(I25386),.A(g18763));
  NOT NOT1_6573(.VSS(VSS),.VDD(VDD),.Y(g19175),.A(I25386));
  NOT NOT1_6574(.VSS(VSS),.VDD(VDD),.Y(I25389),.A(g18780));
  NOT NOT1_6575(.VSS(VSS),.VDD(VDD),.Y(g19176),.A(I25389));
  NOT NOT1_6576(.VSS(VSS),.VDD(VDD),.Y(I25395),.A(g18782));
  NOT NOT1_6577(.VSS(VSS),.VDD(VDD),.Y(g19180),.A(I25395));
  NOT NOT1_6578(.VSS(VSS),.VDD(VDD),.Y(I25399),.A(g18794));
  NOT NOT1_6579(.VSS(VSS),.VDD(VDD),.Y(g19182),.A(I25399));
  NOT NOT1_6580(.VSS(VSS),.VDD(VDD),.Y(I25402),.A(g18821));
  NOT NOT1_6581(.VSS(VSS),.VDD(VDD),.Y(g19183),.A(I25402));
  NOT NOT1_6582(.VSS(VSS),.VDD(VDD),.Y(I25406),.A(g18804));
  NOT NOT1_6583(.VSS(VSS),.VDD(VDD),.Y(g19185),.A(I25406));
  NOT NOT1_6584(.VSS(VSS),.VDD(VDD),.Y(I25412),.A(g18820));
  NOT NOT1_6585(.VSS(VSS),.VDD(VDD),.Y(g19189),.A(I25412));
  NOT NOT1_6586(.VSS(VSS),.VDD(VDD),.Y(I25415),.A(g18835));
  NOT NOT1_6587(.VSS(VSS),.VDD(VDD),.Y(g19190),.A(I25415));
  NOT NOT1_6588(.VSS(VSS),.VDD(VDD),.Y(I25423),.A(g18852));
  NOT NOT1_6589(.VSS(VSS),.VDD(VDD),.Y(g19196),.A(I25423));
  NOT NOT1_6590(.VSS(VSS),.VDD(VDD),.Y(I25426),.A(g18836));
  NOT NOT1_6591(.VSS(VSS),.VDD(VDD),.Y(g19197),.A(I25426));
  NOT NOT1_6592(.VSS(VSS),.VDD(VDD),.Y(I25429),.A(g18975));
  NOT NOT1_6593(.VSS(VSS),.VDD(VDD),.Y(g19198),.A(I25429));
  NOT NOT1_6594(.VSS(VSS),.VDD(VDD),.Y(I25432),.A(g18837));
  NOT NOT1_6595(.VSS(VSS),.VDD(VDD),.Y(g19199),.A(I25432));
  NOT NOT1_6596(.VSS(VSS),.VDD(VDD),.Y(I25442),.A(g18866));
  NOT NOT1_6597(.VSS(VSS),.VDD(VDD),.Y(g19207),.A(I25442));
  NOT NOT1_6598(.VSS(VSS),.VDD(VDD),.Y(I25445),.A(g18968));
  NOT NOT1_6599(.VSS(VSS),.VDD(VDD),.Y(g19208),.A(I25445));
  NOT NOT1_6600(.VSS(VSS),.VDD(VDD),.Y(I25456),.A(g18883));
  NOT NOT1_6601(.VSS(VSS),.VDD(VDD),.Y(g19217),.A(I25456));
  NOT NOT1_6602(.VSS(VSS),.VDD(VDD),.Y(I25459),.A(g18867));
  NOT NOT1_6603(.VSS(VSS),.VDD(VDD),.Y(g19218),.A(I25459));
  NOT NOT1_6604(.VSS(VSS),.VDD(VDD),.Y(I25463),.A(g18868));
  NOT NOT1_6605(.VSS(VSS),.VDD(VDD),.Y(g19220),.A(I25463));
  NOT NOT1_6606(.VSS(VSS),.VDD(VDD),.Y(I25474),.A(g18885));
  NOT NOT1_6607(.VSS(VSS),.VDD(VDD),.Y(g19229),.A(I25474));
  NOT NOT1_6608(.VSS(VSS),.VDD(VDD),.Y(I25486),.A(g18754));
  NOT NOT1_6609(.VSS(VSS),.VDD(VDD),.Y(g19237),.A(I25486));
  NOT NOT1_6610(.VSS(VSS),.VDD(VDD),.Y(I25489),.A(g18906));
  NOT NOT1_6611(.VSS(VSS),.VDD(VDD),.Y(g19238),.A(I25489));
  NOT NOT1_6612(.VSS(VSS),.VDD(VDD),.Y(I25492),.A(g18907));
  NOT NOT1_6613(.VSS(VSS),.VDD(VDD),.Y(g19239),.A(I25492));
  NOT NOT1_6614(.VSS(VSS),.VDD(VDD),.Y(I25506),.A(g18781));
  NOT NOT1_6615(.VSS(VSS),.VDD(VDD),.Y(g19247),.A(I25506));
  NOT NOT1_6616(.VSS(VSS),.VDD(VDD),.Y(I25510),.A(g18542));
  NOT NOT1_6617(.VSS(VSS),.VDD(VDD),.Y(g19249),.A(I25510));
  NOT NOT1_6618(.VSS(VSS),.VDD(VDD),.Y(g19251),.A(g16540));
  NOT NOT1_6619(.VSS(VSS),.VDD(VDD),.Y(I25525),.A(g18803));
  NOT NOT1_6620(.VSS(VSS),.VDD(VDD),.Y(g19258),.A(I25525));
  NOT NOT1_6621(.VSS(VSS),.VDD(VDD),.Y(I25528),.A(g18942));
  NOT NOT1_6622(.VSS(VSS),.VDD(VDD),.Y(g19259),.A(I25528));
  NOT NOT1_6623(.VSS(VSS),.VDD(VDD),.Y(g19265),.A(g16572));
  NOT NOT1_6624(.VSS(VSS),.VDD(VDD),.Y(I25557),.A(g18957));
  NOT NOT1_6625(.VSS(VSS),.VDD(VDD),.Y(g19270),.A(I25557));
  NOT NOT1_6626(.VSS(VSS),.VDD(VDD),.Y(I25567),.A(g17186));
  NOT NOT1_6627(.VSS(VSS),.VDD(VDD),.Y(g19272),.A(I25567));
  NOT NOT1_6628(.VSS(VSS),.VDD(VDD),.Y(g19280),.A(g16596));
  NOT NOT1_6629(.VSS(VSS),.VDD(VDD),.Y(g19287),.A(g16608));
  NOT NOT1_6630(.VSS(VSS),.VDD(VDD),.Y(I25612),.A(g17197));
  NOT NOT1_6631(.VSS(VSS),.VDD(VDD),.Y(g19291),.A(I25612));
  NOT NOT1_6632(.VSS(VSS),.VDD(VDD),.Y(g19299),.A(g16616));
  NOT NOT1_6633(.VSS(VSS),.VDD(VDD),.Y(g19301),.A(g16622));
  NOT NOT1_6634(.VSS(VSS),.VDD(VDD),.Y(g19302),.A(g17025));
  NOT NOT1_6635(.VSS(VSS),.VDD(VDD),.Y(g19305),.A(g16626));
  NOT NOT1_6636(.VSS(VSS),.VDD(VDD),.Y(I25660),.A(g17204));
  NOT NOT1_6637(.VSS(VSS),.VDD(VDD),.Y(g19309),.A(I25660));
  NOT NOT1_6638(.VSS(VSS),.VDD(VDD),.Y(g19319),.A(g16633));
  NOT NOT1_6639(.VSS(VSS),.VDD(VDD),.Y(g19322),.A(g16636));
  NOT NOT1_6640(.VSS(VSS),.VDD(VDD),.Y(g19323),.A(g17059));
  NOT NOT1_6641(.VSS(VSS),.VDD(VDD),.Y(g19326),.A(g16640));
  NOT NOT1_6642(.VSS(VSS),.VDD(VDD),.Y(I25717),.A(g17209));
  NOT NOT1_6643(.VSS(VSS),.VDD(VDD),.Y(g19330),.A(I25717));
  NOT NOT1_6644(.VSS(VSS),.VDD(VDD),.Y(I25728),.A(g17118));
  NOT NOT1_6645(.VSS(VSS),.VDD(VDD),.Y(g19335),.A(I25728));
  NOT NOT1_6646(.VSS(VSS),.VDD(VDD),.Y(g19346),.A(g16644));
  NOT NOT1_6647(.VSS(VSS),.VDD(VDD),.Y(g19349),.A(g16647));
  NOT NOT1_6648(.VSS(VSS),.VDD(VDD),.Y(g19350),.A(g17094));
  NOT NOT1_6649(.VSS(VSS),.VDD(VDD),.Y(g19353),.A(g16651));
  NOT NOT1_6650(.VSS(VSS),.VDD(VDD),.Y(I25768),.A(g17139));
  NOT NOT1_6651(.VSS(VSS),.VDD(VDD),.Y(g19358),.A(I25768));
  NOT NOT1_6652(.VSS(VSS),.VDD(VDD),.Y(I25778),.A(g17145));
  NOT NOT1_6653(.VSS(VSS),.VDD(VDD),.Y(g19369),.A(I25778));
  NOT NOT1_6654(.VSS(VSS),.VDD(VDD),.Y(g19380),.A(g16656));
  NOT NOT1_6655(.VSS(VSS),.VDD(VDD),.Y(g19383),.A(g16659));
  NOT NOT1_6656(.VSS(VSS),.VDD(VDD),.Y(g19384),.A(g17132));
  NOT NOT1_6657(.VSS(VSS),.VDD(VDD),.Y(g19387),.A(g16567));
  NOT NOT1_6658(.VSS(VSS),.VDD(VDD),.Y(g19388),.A(g17139));
  NOT NOT1_6659(.VSS(VSS),.VDD(VDD),.Y(I25816),.A(g17162));
  NOT NOT1_6660(.VSS(VSS),.VDD(VDD),.Y(g19390),.A(I25816));
  NOT NOT1_6661(.VSS(VSS),.VDD(VDD),.Y(I25826),.A(g17168));
  NOT NOT1_6662(.VSS(VSS),.VDD(VDD),.Y(g19401),.A(I25826));
  NOT NOT1_6663(.VSS(VSS),.VDD(VDD),.Y(g19412),.A(g16673));
  NOT NOT1_6664(.VSS(VSS),.VDD(VDD),.Y(g19415),.A(g16676));
  NOT NOT1_6665(.VSS(VSS),.VDD(VDD),.Y(g19417),.A(g16591));
  NOT NOT1_6666(.VSS(VSS),.VDD(VDD),.Y(g19418),.A(g17162));
  NOT NOT1_6667(.VSS(VSS),.VDD(VDD),.Y(I25862),.A(g17177));
  NOT NOT1_6668(.VSS(VSS),.VDD(VDD),.Y(g19420),.A(I25862));
  NOT NOT1_6669(.VSS(VSS),.VDD(VDD),.Y(I25872),.A(g17183));
  NOT NOT1_6670(.VSS(VSS),.VDD(VDD),.Y(g19431),.A(I25872));
  NOT NOT1_6671(.VSS(VSS),.VDD(VDD),.Y(g19441),.A(g17213));
  NOT NOT1_6672(.VSS(VSS),.VDD(VDD),.Y(g19444),.A(g17985));
  NOT NOT1_6673(.VSS(VSS),.VDD(VDD),.Y(g19448),.A(g16694));
  NOT NOT1_6674(.VSS(VSS),.VDD(VDD),.Y(g19452),.A(g16702));
  NOT NOT1_6675(.VSS(VSS),.VDD(VDD),.Y(g19454),.A(g16611));
  NOT NOT1_6676(.VSS(VSS),.VDD(VDD),.Y(g19455),.A(g17177));
  NOT NOT1_6677(.VSS(VSS),.VDD(VDD),.Y(I25904),.A(g17194));
  NOT NOT1_6678(.VSS(VSS),.VDD(VDD),.Y(g19457),.A(I25904));
  NOT NOT1_6679(.VSS(VSS),.VDD(VDD),.Y(g19467),.A(g16719));
  NOT NOT1_6680(.VSS(VSS),.VDD(VDD),.Y(g19468),.A(g17216));
  NOT NOT1_6681(.VSS(VSS),.VDD(VDD),.Y(g19471),.A(g18102));
  NOT NOT1_6682(.VSS(VSS),.VDD(VDD),.Y(g19475),.A(g16725));
  NOT NOT1_6683(.VSS(VSS),.VDD(VDD),.Y(g19479),.A(g16733));
  NOT NOT1_6684(.VSS(VSS),.VDD(VDD),.Y(g19481),.A(g16629));
  NOT NOT1_6685(.VSS(VSS),.VDD(VDD),.Y(g19482),.A(g17194));
  NOT NOT1_6686(.VSS(VSS),.VDD(VDD),.Y(g19483),.A(g16758));
  NOT NOT1_6687(.VSS(VSS),.VDD(VDD),.Y(g19484),.A(g16867));
  NOT NOT1_6688(.VSS(VSS),.VDD(VDD),.Y(g19490),.A(g16761));
  NOT NOT1_6689(.VSS(VSS),.VDD(VDD),.Y(g19491),.A(g17219));
  NOT NOT1_6690(.VSS(VSS),.VDD(VDD),.Y(g19494),.A(g18218));
  NOT NOT1_6691(.VSS(VSS),.VDD(VDD),.Y(g19498),.A(g16767));
  NOT NOT1_6692(.VSS(VSS),.VDD(VDD),.Y(g19502),.A(g16775));
  NOT NOT1_6693(.VSS(VSS),.VDD(VDD),.Y(g19504),.A(g16785));
  NOT NOT1_6694(.VSS(VSS),.VDD(VDD),.Y(g19505),.A(g16895));
  NOT NOT1_6695(.VSS(VSS),.VDD(VDD),.Y(g19511),.A(g16788));
  NOT NOT1_6696(.VSS(VSS),.VDD(VDD),.Y(g19512),.A(g17221));
  NOT NOT1_6697(.VSS(VSS),.VDD(VDD),.Y(g19515),.A(g18325));
  NOT NOT1_6698(.VSS(VSS),.VDD(VDD),.Y(g19519),.A(g16794));
  NOT NOT1_6699(.VSS(VSS),.VDD(VDD),.Y(g19523),.A(g16814));
  NOT NOT1_6700(.VSS(VSS),.VDD(VDD),.Y(g19524),.A(g16924));
  NOT NOT1_6701(.VSS(VSS),.VDD(VDD),.Y(g19530),.A(g16817));
  NOT NOT1_6702(.VSS(VSS),.VDD(VDD),.Y(g19533),.A(g16832));
  NOT NOT1_6703(.VSS(VSS),.VDD(VDD),.Y(g19534),.A(g16954));
  NOT NOT1_6704(.VSS(VSS),.VDD(VDD),.Y(I25966),.A(g16654));
  NOT NOT1_6705(.VSS(VSS),.VDD(VDD),.Y(g19543),.A(I25966));
  NOT NOT1_6706(.VSS(VSS),.VDD(VDD),.Y(I25971),.A(g16671));
  NOT NOT1_6707(.VSS(VSS),.VDD(VDD),.Y(g19546),.A(I25971));
  NOT NOT1_6708(.VSS(VSS),.VDD(VDD),.Y(I25977),.A(g16692));
  NOT NOT1_6709(.VSS(VSS),.VDD(VDD),.Y(g19550),.A(I25977));
  NOT NOT1_6710(.VSS(VSS),.VDD(VDD),.Y(I25985),.A(g16718));
  NOT NOT1_6711(.VSS(VSS),.VDD(VDD),.Y(g19556),.A(I25985));
  NOT NOT1_6712(.VSS(VSS),.VDD(VDD),.Y(I25994),.A(g16860));
  NOT NOT1_6713(.VSS(VSS),.VDD(VDD),.Y(g19563),.A(I25994));
  NOT NOT1_6714(.VSS(VSS),.VDD(VDD),.Y(I26006),.A(g16866));
  NOT NOT1_6715(.VSS(VSS),.VDD(VDD),.Y(g19573),.A(I26006));
  NOT NOT1_6716(.VSS(VSS),.VDD(VDD),.Y(g19577),.A(g16881));
  NOT NOT1_6717(.VSS(VSS),.VDD(VDD),.Y(g19578),.A(g16884));
  NOT NOT1_6718(.VSS(VSS),.VDD(VDD),.Y(I26025),.A(g16803));
  NOT NOT1_6719(.VSS(VSS),.VDD(VDD),.Y(g19595),.A(I26025));
  NOT NOT1_6720(.VSS(VSS),.VDD(VDD),.Y(I26028),.A(g16566));
  NOT NOT1_6721(.VSS(VSS),.VDD(VDD),.Y(g19596),.A(I26028));
  NOT NOT1_6722(.VSS(VSS),.VDD(VDD),.Y(g19607),.A(g16910));
  NOT NOT1_6723(.VSS(VSS),.VDD(VDD),.Y(g19608),.A(g16913));
  NOT NOT1_6724(.VSS(VSS),.VDD(VDD),.Y(I26051),.A(g16824));
  NOT NOT1_6725(.VSS(VSS),.VDD(VDD),.Y(g19622),.A(I26051));
  NOT NOT1_6726(.VSS(VSS),.VDD(VDD),.Y(g19640),.A(g16940));
  NOT NOT1_6727(.VSS(VSS),.VDD(VDD),.Y(g19641),.A(g16943));
  NOT NOT1_6728(.VSS(VSS),.VDD(VDD),.Y(I26078),.A(g16835));
  NOT NOT1_6729(.VSS(VSS),.VDD(VDD),.Y(g19652),.A(I26078));
  NOT NOT1_6730(.VSS(VSS),.VDD(VDD),.Y(I26085),.A(g18085));
  NOT NOT1_6731(.VSS(VSS),.VDD(VDD),.Y(g19657),.A(I26085));
  NOT NOT1_6732(.VSS(VSS),.VDD(VDD),.Y(g19680),.A(g16971));
  NOT NOT1_6733(.VSS(VSS),.VDD(VDD),.Y(g19681),.A(g16974));
  NOT NOT1_6734(.VSS(VSS),.VDD(VDD),.Y(I26112),.A(g16844));
  NOT NOT1_6735(.VSS(VSS),.VDD(VDD),.Y(g19689),.A(I26112));
  NOT NOT1_6736(.VSS(VSS),.VDD(VDD),.Y(I26115),.A(g16845));
  NOT NOT1_6737(.VSS(VSS),.VDD(VDD),.Y(g19690),.A(I26115));
  NOT NOT1_6738(.VSS(VSS),.VDD(VDD),.Y(I26123),.A(g17503));
  NOT NOT1_6739(.VSS(VSS),.VDD(VDD),.Y(g19696),.A(I26123));
  NOT NOT1_6740(.VSS(VSS),.VDD(VDD),.Y(I26134),.A(g18201));
  NOT NOT1_6741(.VSS(VSS),.VDD(VDD),.Y(g19705),.A(I26134));
  NOT NOT1_6742(.VSS(VSS),.VDD(VDD),.Y(I26154),.A(g16851));
  NOT NOT1_6743(.VSS(VSS),.VDD(VDD),.Y(g19725),.A(I26154));
  NOT NOT1_6744(.VSS(VSS),.VDD(VDD),.Y(I26171),.A(g17594));
  NOT NOT1_6745(.VSS(VSS),.VDD(VDD),.Y(g19740),.A(I26171));
  NOT NOT1_6746(.VSS(VSS),.VDD(VDD),.Y(I26182),.A(g18308));
  NOT NOT1_6747(.VSS(VSS),.VDD(VDD),.Y(g19749),.A(I26182));
  NOT NOT1_6748(.VSS(VSS),.VDD(VDD),.Y(I26195),.A(g16853));
  NOT NOT1_6749(.VSS(VSS),.VDD(VDD),.Y(g19762),.A(I26195));
  NOT NOT1_6750(.VSS(VSS),.VDD(VDD),.Y(I26198),.A(g16854));
  NOT NOT1_6751(.VSS(VSS),.VDD(VDD),.Y(g19763),.A(I26198));
  NOT NOT1_6752(.VSS(VSS),.VDD(VDD),.Y(I26220),.A(g17691));
  NOT NOT1_6753(.VSS(VSS),.VDD(VDD),.Y(g19783),.A(I26220));
  NOT NOT1_6754(.VSS(VSS),.VDD(VDD),.Y(I26231),.A(g18401));
  NOT NOT1_6755(.VSS(VSS),.VDD(VDD),.Y(g19792),.A(I26231));
  NOT NOT1_6756(.VSS(VSS),.VDD(VDD),.Y(I26237),.A(g16857));
  NOT NOT1_6757(.VSS(VSS),.VDD(VDD),.Y(g19798),.A(I26237));
  NOT NOT1_6758(.VSS(VSS),.VDD(VDD),.Y(I26266),.A(g17791));
  NOT NOT1_6759(.VSS(VSS),.VDD(VDD),.Y(g19825),.A(I26266));
  NOT NOT1_6760(.VSS(VSS),.VDD(VDD),.Y(g19830),.A(g18886));
  NOT NOT1_6761(.VSS(VSS),.VDD(VDD),.Y(I26276),.A(g16861));
  NOT NOT1_6762(.VSS(VSS),.VDD(VDD),.Y(g19838),.A(I26276));
  NOT NOT1_6763(.VSS(VSS),.VDD(VDD),.Y(I26334),.A(g18977));
  NOT NOT1_6764(.VSS(VSS),.VDD(VDD),.Y(g19890),.A(I26334));
  NOT NOT1_6765(.VSS(VSS),.VDD(VDD),.Y(I26337),.A(g16880));
  NOT NOT1_6766(.VSS(VSS),.VDD(VDD),.Y(g19893),.A(I26337));
  NOT NOT1_6767(.VSS(VSS),.VDD(VDD),.Y(I26340),.A(g17025));
  NOT NOT1_6768(.VSS(VSS),.VDD(VDD),.Y(g19894),.A(I26340));
  NOT NOT1_6769(.VSS(VSS),.VDD(VDD),.Y(I26365),.A(g18626));
  NOT NOT1_6770(.VSS(VSS),.VDD(VDD),.Y(g19915),.A(I26365));
  NOT NOT1_6771(.VSS(VSS),.VDD(VDD),.Y(g19918),.A(g18646));
  NOT NOT1_6772(.VSS(VSS),.VDD(VDD),.Y(I26369),.A(g17059));
  NOT NOT1_6773(.VSS(VSS),.VDD(VDD),.Y(g19919),.A(I26369));
  NOT NOT1_6774(.VSS(VSS),.VDD(VDD),.Y(g19933),.A(g18548));
  NOT NOT1_6775(.VSS(VSS),.VDD(VDD),.Y(I26388),.A(g17094));
  NOT NOT1_6776(.VSS(VSS),.VDD(VDD),.Y(g19934),.A(I26388));
  NOT NOT1_6777(.VSS(VSS),.VDD(VDD),.Y(I26401),.A(g17012));
  NOT NOT1_6778(.VSS(VSS),.VDD(VDD),.Y(g19945),.A(I26401));
  NOT NOT1_6779(.VSS(VSS),.VDD(VDD),.Y(g19948),.A(g17896));
  NOT NOT1_6780(.VSS(VSS),.VDD(VDD),.Y(g19950),.A(g18598));
  NOT NOT1_6781(.VSS(VSS),.VDD(VDD),.Y(I26407),.A(g17132));
  NOT NOT1_6782(.VSS(VSS),.VDD(VDD),.Y(g19951),.A(I26407));
  NOT NOT1_6783(.VSS(VSS),.VDD(VDD),.Y(I26413),.A(g16643));
  NOT NOT1_6784(.VSS(VSS),.VDD(VDD),.Y(g19957),.A(I26413));
  NOT NOT1_6785(.VSS(VSS),.VDD(VDD),.Y(I26420),.A(g17042));
  NOT NOT1_6786(.VSS(VSS),.VDD(VDD),.Y(g19972),.A(I26420));
  NOT NOT1_6787(.VSS(VSS),.VDD(VDD),.Y(g19975),.A(g18007));
  NOT NOT1_6788(.VSS(VSS),.VDD(VDD),.Y(g19977),.A(g18630));
  NOT NOT1_6789(.VSS(VSS),.VDD(VDD),.Y(I26426),.A(g16536));
  NOT NOT1_6790(.VSS(VSS),.VDD(VDD),.Y(g19978),.A(I26426));
  NOT NOT1_6791(.VSS(VSS),.VDD(VDD),.Y(I26437),.A(g16655));
  NOT NOT1_6792(.VSS(VSS),.VDD(VDD),.Y(g19987),.A(I26437));
  NOT NOT1_6793(.VSS(VSS),.VDD(VDD),.Y(I26444),.A(g17076));
  NOT NOT1_6794(.VSS(VSS),.VDD(VDD),.Y(g20002),.A(I26444));
  NOT NOT1_6795(.VSS(VSS),.VDD(VDD),.Y(g20005),.A(g18124));
  NOT NOT1_6796(.VSS(VSS),.VDD(VDD),.Y(g20007),.A(g18639));
  NOT NOT1_6797(.VSS(VSS),.VDD(VDD),.Y(I26458),.A(g17985));
  NOT NOT1_6798(.VSS(VSS),.VDD(VDD),.Y(g20016),.A(I26458));
  NOT NOT1_6799(.VSS(VSS),.VDD(VDD),.Y(I26469),.A(g16672));
  NOT NOT1_6800(.VSS(VSS),.VDD(VDD),.Y(g20025),.A(I26469));
  NOT NOT1_6801(.VSS(VSS),.VDD(VDD),.Y(I26476),.A(g17111));
  NOT NOT1_6802(.VSS(VSS),.VDD(VDD),.Y(g20040),.A(I26476));
  NOT NOT1_6803(.VSS(VSS),.VDD(VDD),.Y(g20043),.A(g18240));
  NOT NOT1_6804(.VSS(VSS),.VDD(VDD),.Y(I26481),.A(g18590));
  NOT NOT1_6805(.VSS(VSS),.VDD(VDD),.Y(g20045),.A(I26481));
  NOT NOT1_6806(.VSS(VSS),.VDD(VDD),.Y(I26494),.A(g18102));
  NOT NOT1_6807(.VSS(VSS),.VDD(VDD),.Y(g20058),.A(I26494));
  NOT NOT1_6808(.VSS(VSS),.VDD(VDD),.Y(I26505),.A(g16693));
  NOT NOT1_6809(.VSS(VSS),.VDD(VDD),.Y(g20067),.A(I26505));
  NOT NOT1_6810(.VSS(VSS),.VDD(VDD),.Y(I26512),.A(g16802));
  NOT NOT1_6811(.VSS(VSS),.VDD(VDD),.Y(g20082),.A(I26512));
  NOT NOT1_6812(.VSS(VSS),.VDD(VDD),.Y(g20083),.A(g17968));
  NOT NOT1_6813(.VSS(VSS),.VDD(VDD),.Y(I26535),.A(g18218));
  NOT NOT1_6814(.VSS(VSS),.VDD(VDD),.Y(g20099),.A(I26535));
  NOT NOT1_6815(.VSS(VSS),.VDD(VDD),.Y(I26545),.A(g16823));
  NOT NOT1_6816(.VSS(VSS),.VDD(VDD),.Y(g20105),.A(I26545));
  NOT NOT1_6817(.VSS(VSS),.VDD(VDD),.Y(I26574),.A(g18325));
  NOT NOT1_6818(.VSS(VSS),.VDD(VDD),.Y(g20124),.A(I26574));
  NOT NOT1_6819(.VSS(VSS),.VDD(VDD),.Y(g20127),.A(g18623));
  NOT NOT1_6820(.VSS(VSS),.VDD(VDD),.Y(g20140),.A(g16830));
  NOT NOT1_6821(.VSS(VSS),.VDD(VDD),.Y(g20163),.A(g17973));
  NOT NOT1_6822(.VSS(VSS),.VDD(VDD),.Y(I26612),.A(g17645));
  NOT NOT1_6823(.VSS(VSS),.VDD(VDD),.Y(g20164),.A(I26612));
  NOT NOT1_6824(.VSS(VSS),.VDD(VDD),.Y(g20178),.A(g16842));
  NOT NOT1_6825(.VSS(VSS),.VDD(VDD),.Y(g20193),.A(g18691));
  NOT NOT1_6826(.VSS(VSS),.VDD(VDD),.Y(I26642),.A(g17746));
  NOT NOT1_6827(.VSS(VSS),.VDD(VDD),.Y(g20198),.A(I26642));
  NOT NOT1_6828(.VSS(VSS),.VDD(VDD),.Y(g20212),.A(g16848));
  NOT NOT1_6829(.VSS(VSS),.VDD(VDD),.Y(g20223),.A(g18727));
  NOT NOT1_6830(.VSS(VSS),.VDD(VDD),.Y(I26664),.A(g17847));
  NOT NOT1_6831(.VSS(VSS),.VDD(VDD),.Y(g20228),.A(I26664));
  NOT NOT1_6832(.VSS(VSS),.VDD(VDD),.Y(g20242),.A(g16852));
  NOT NOT1_6833(.VSS(VSS),.VDD(VDD),.Y(g20250),.A(g18764));
  NOT NOT1_6834(.VSS(VSS),.VDD(VDD),.Y(I26679),.A(g17959));
  NOT NOT1_6835(.VSS(VSS),.VDD(VDD),.Y(g20255),.A(I26679));
  NOT NOT1_6836(.VSS(VSS),.VDD(VDD),.Y(g20269),.A(g17230));
  NOT NOT1_6837(.VSS(VSS),.VDD(VDD),.Y(g20273),.A(g18795));
  NOT NOT1_6838(.VSS(VSS),.VDD(VDD),.Y(g20278),.A(g17237));
  NOT NOT1_6839(.VSS(VSS),.VDD(VDD),.Y(g20279),.A(g17240));
  NOT NOT1_6840(.VSS(VSS),.VDD(VDD),.Y(g20281),.A(g17243));
  NOT NOT1_6841(.VSS(VSS),.VDD(VDD),.Y(g20286),.A(g17249));
  NOT NOT1_6842(.VSS(VSS),.VDD(VDD),.Y(g20287),.A(g17252));
  NOT NOT1_6843(.VSS(VSS),.VDD(VDD),.Y(g20288),.A(g17255));
  NOT NOT1_6844(.VSS(VSS),.VDD(VDD),.Y(g20289),.A(g17259));
  NOT NOT1_6845(.VSS(VSS),.VDD(VDD),.Y(g20290),.A(g17262));
  NOT NOT1_6846(.VSS(VSS),.VDD(VDD),.Y(g20292),.A(g17265));
  NOT NOT1_6847(.VSS(VSS),.VDD(VDD),.Y(I26714),.A(g17720));
  NOT NOT1_6848(.VSS(VSS),.VDD(VDD),.Y(g20295),.A(I26714));
  NOT NOT1_6849(.VSS(VSS),.VDD(VDD),.Y(g20296),.A(g17272));
  NOT NOT1_6850(.VSS(VSS),.VDD(VDD),.Y(g20297),.A(g17275));
  NOT NOT1_6851(.VSS(VSS),.VDD(VDD),.Y(g20298),.A(g17278));
  NOT NOT1_6852(.VSS(VSS),.VDD(VDD),.Y(g20302),.A(g17282));
  NOT NOT1_6853(.VSS(VSS),.VDD(VDD),.Y(g20303),.A(g17285));
  NOT NOT1_6854(.VSS(VSS),.VDD(VDD),.Y(g20304),.A(g17288));
  NOT NOT1_6855(.VSS(VSS),.VDD(VDD),.Y(g20305),.A(g17291));
  NOT NOT1_6856(.VSS(VSS),.VDD(VDD),.Y(g20306),.A(g17294));
  NOT NOT1_6857(.VSS(VSS),.VDD(VDD),.Y(g20308),.A(g17297));
  NOT NOT1_6858(.VSS(VSS),.VDD(VDD),.Y(g20311),.A(g17304));
  NOT NOT1_6859(.VSS(VSS),.VDD(VDD),.Y(g20312),.A(g17307));
  NOT NOT1_6860(.VSS(VSS),.VDD(VDD),.Y(g20313),.A(g17310));
  NOT NOT1_6861(.VSS(VSS),.VDD(VDD),.Y(g20315),.A(g17315));
  NOT NOT1_6862(.VSS(VSS),.VDD(VDD),.Y(g20316),.A(g17318));
  NOT NOT1_6863(.VSS(VSS),.VDD(VDD),.Y(g20317),.A(g17321));
  NOT NOT1_6864(.VSS(VSS),.VDD(VDD),.Y(g20321),.A(g17324));
  NOT NOT1_6865(.VSS(VSS),.VDD(VDD),.Y(g20322),.A(g17327));
  NOT NOT1_6866(.VSS(VSS),.VDD(VDD),.Y(g20323),.A(g17330));
  NOT NOT1_6867(.VSS(VSS),.VDD(VDD),.Y(g20324),.A(g17333));
  NOT NOT1_6868(.VSS(VSS),.VDD(VDD),.Y(g20325),.A(g17336));
  NOT NOT1_6869(.VSS(VSS),.VDD(VDD),.Y(g20327),.A(g17342));
  NOT NOT1_6870(.VSS(VSS),.VDD(VDD),.Y(g20328),.A(g17345));
  NOT NOT1_6871(.VSS(VSS),.VDD(VDD),.Y(g20329),.A(g17348));
  NOT NOT1_6872(.VSS(VSS),.VDD(VDD),.Y(g20330),.A(g17354));
  NOT NOT1_6873(.VSS(VSS),.VDD(VDD),.Y(g20331),.A(g17357));
  NOT NOT1_6874(.VSS(VSS),.VDD(VDD),.Y(g20332),.A(g17360));
  NOT NOT1_6875(.VSS(VSS),.VDD(VDD),.Y(g20334),.A(g17363));
  NOT NOT1_6876(.VSS(VSS),.VDD(VDD),.Y(g20335),.A(g17366));
  NOT NOT1_6877(.VSS(VSS),.VDD(VDD),.Y(g20336),.A(g17369));
  NOT NOT1_6878(.VSS(VSS),.VDD(VDD),.Y(g20340),.A(g17372));
  NOT NOT1_6879(.VSS(VSS),.VDD(VDD),.Y(g20341),.A(g17375));
  NOT NOT1_6880(.VSS(VSS),.VDD(VDD),.Y(g20342),.A(g17378));
  NOT NOT1_6881(.VSS(VSS),.VDD(VDD),.Y(g20344),.A(g17384));
  NOT NOT1_6882(.VSS(VSS),.VDD(VDD),.Y(g20345),.A(g17387));
  NOT NOT1_6883(.VSS(VSS),.VDD(VDD),.Y(g20346),.A(g17390));
  NOT NOT1_6884(.VSS(VSS),.VDD(VDD),.Y(g20347),.A(g17399));
  NOT NOT1_6885(.VSS(VSS),.VDD(VDD),.Y(g20348),.A(g17402));
  NOT NOT1_6886(.VSS(VSS),.VDD(VDD),.Y(g20349),.A(g17405));
  NOT NOT1_6887(.VSS(VSS),.VDD(VDD),.Y(g20350),.A(g17410));
  NOT NOT1_6888(.VSS(VSS),.VDD(VDD),.Y(g20351),.A(g17413));
  NOT NOT1_6889(.VSS(VSS),.VDD(VDD),.Y(g20352),.A(g17416));
  NOT NOT1_6890(.VSS(VSS),.VDD(VDD),.Y(g20354),.A(g17419));
  NOT NOT1_6891(.VSS(VSS),.VDD(VDD),.Y(g20355),.A(g17422));
  NOT NOT1_6892(.VSS(VSS),.VDD(VDD),.Y(g20356),.A(g17425));
  NOT NOT1_6893(.VSS(VSS),.VDD(VDD),.Y(I26777),.A(g17222));
  NOT NOT1_6894(.VSS(VSS),.VDD(VDD),.Y(g20360),.A(I26777));
  NOT NOT1_6895(.VSS(VSS),.VDD(VDD),.Y(g20361),.A(g17430));
  NOT NOT1_6896(.VSS(VSS),.VDD(VDD),.Y(g20362),.A(g17433));
  NOT NOT1_6897(.VSS(VSS),.VDD(VDD),.Y(g20363),.A(g17436));
  NOT NOT1_6898(.VSS(VSS),.VDD(VDD),.Y(g20364),.A(g17439));
  NOT NOT1_6899(.VSS(VSS),.VDD(VDD),.Y(g20365),.A(g17442));
  NOT NOT1_6900(.VSS(VSS),.VDD(VDD),.Y(g20366),.A(g17451));
  NOT NOT1_6901(.VSS(VSS),.VDD(VDD),.Y(g20367),.A(g17454));
  NOT NOT1_6902(.VSS(VSS),.VDD(VDD),.Y(g20368),.A(g17457));
  NOT NOT1_6903(.VSS(VSS),.VDD(VDD),.Y(g20369),.A(g17465));
  NOT NOT1_6904(.VSS(VSS),.VDD(VDD),.Y(g20370),.A(g17468));
  NOT NOT1_6905(.VSS(VSS),.VDD(VDD),.Y(g20371),.A(g17471));
  NOT NOT1_6906(.VSS(VSS),.VDD(VDD),.Y(g20372),.A(g17476));
  NOT NOT1_6907(.VSS(VSS),.VDD(VDD),.Y(g20373),.A(g17479));
  NOT NOT1_6908(.VSS(VSS),.VDD(VDD),.Y(g20374),.A(g17482));
  NOT NOT1_6909(.VSS(VSS),.VDD(VDD),.Y(I26796),.A(g17224));
  NOT NOT1_6910(.VSS(VSS),.VDD(VDD),.Y(g20377),.A(I26796));
  NOT NOT1_6911(.VSS(VSS),.VDD(VDD),.Y(g20378),.A(g17487));
  NOT NOT1_6912(.VSS(VSS),.VDD(VDD),.Y(g20379),.A(g17490));
  NOT NOT1_6913(.VSS(VSS),.VDD(VDD),.Y(g20380),.A(g17493));
  NOT NOT1_6914(.VSS(VSS),.VDD(VDD),.Y(g20381),.A(g17496));
  NOT NOT1_6915(.VSS(VSS),.VDD(VDD),.Y(g20382),.A(g17500));
  NOT NOT1_6916(.VSS(VSS),.VDD(VDD),.Y(g20383),.A(g17503));
  NOT NOT1_6917(.VSS(VSS),.VDD(VDD),.Y(g20384),.A(g17511));
  NOT NOT1_6918(.VSS(VSS),.VDD(VDD),.Y(g20385),.A(g17514));
  NOT NOT1_6919(.VSS(VSS),.VDD(VDD),.Y(g20386),.A(g17517));
  NOT NOT1_6920(.VSS(VSS),.VDD(VDD),.Y(g20387),.A(g17520));
  NOT NOT1_6921(.VSS(VSS),.VDD(VDD),.Y(g20388),.A(g17523));
  NOT NOT1_6922(.VSS(VSS),.VDD(VDD),.Y(g20389),.A(g17531));
  NOT NOT1_6923(.VSS(VSS),.VDD(VDD),.Y(g20390),.A(g17534));
  NOT NOT1_6924(.VSS(VSS),.VDD(VDD),.Y(g20391),.A(g17537));
  NOT NOT1_6925(.VSS(VSS),.VDD(VDD),.Y(g20392),.A(g17545));
  NOT NOT1_6926(.VSS(VSS),.VDD(VDD),.Y(g20393),.A(g17548));
  NOT NOT1_6927(.VSS(VSS),.VDD(VDD),.Y(g20394),.A(g17551));
  NOT NOT1_6928(.VSS(VSS),.VDD(VDD),.Y(I26816),.A(g17225));
  NOT NOT1_6929(.VSS(VSS),.VDD(VDD),.Y(g20395),.A(I26816));
  NOT NOT1_6930(.VSS(VSS),.VDD(VDD),.Y(I26819),.A(g17226));
  NOT NOT1_6931(.VSS(VSS),.VDD(VDD),.Y(g20396),.A(I26819));
  NOT NOT1_6932(.VSS(VSS),.VDD(VDD),.Y(g20397),.A(g17557));
  NOT NOT1_6933(.VSS(VSS),.VDD(VDD),.Y(g20398),.A(g17560));
  NOT NOT1_6934(.VSS(VSS),.VDD(VDD),.Y(g20399),.A(g17563));
  NOT NOT1_6935(.VSS(VSS),.VDD(VDD),.Y(g20400),.A(g17567));
  NOT NOT1_6936(.VSS(VSS),.VDD(VDD),.Y(g20401),.A(g17570));
  NOT NOT1_6937(.VSS(VSS),.VDD(VDD),.Y(g20402),.A(g17573));
  NOT NOT1_6938(.VSS(VSS),.VDD(VDD),.Y(g20403),.A(g17579));
  NOT NOT1_6939(.VSS(VSS),.VDD(VDD),.Y(g20404),.A(g17582));
  NOT NOT1_6940(.VSS(VSS),.VDD(VDD),.Y(g20405),.A(g17585));
  NOT NOT1_6941(.VSS(VSS),.VDD(VDD),.Y(g20406),.A(g17588));
  NOT NOT1_6942(.VSS(VSS),.VDD(VDD),.Y(g20407),.A(g17591));
  NOT NOT1_6943(.VSS(VSS),.VDD(VDD),.Y(g20408),.A(g17594));
  NOT NOT1_6944(.VSS(VSS),.VDD(VDD),.Y(g20409),.A(g17601));
  NOT NOT1_6945(.VSS(VSS),.VDD(VDD),.Y(g20410),.A(g17604));
  NOT NOT1_6946(.VSS(VSS),.VDD(VDD),.Y(g20411),.A(g17607));
  NOT NOT1_6947(.VSS(VSS),.VDD(VDD),.Y(g20412),.A(g17610));
  NOT NOT1_6948(.VSS(VSS),.VDD(VDD),.Y(g20413),.A(g17613));
  NOT NOT1_6949(.VSS(VSS),.VDD(VDD),.Y(g20414),.A(g17621));
  NOT NOT1_6950(.VSS(VSS),.VDD(VDD),.Y(g20415),.A(g17624));
  NOT NOT1_6951(.VSS(VSS),.VDD(VDD),.Y(g20416),.A(g17627));
  NOT NOT1_6952(.VSS(VSS),.VDD(VDD),.Y(I26843),.A(g17228));
  NOT NOT1_6953(.VSS(VSS),.VDD(VDD),.Y(g20418),.A(I26843));
  NOT NOT1_6954(.VSS(VSS),.VDD(VDD),.Y(I26846),.A(g17229));
  NOT NOT1_6955(.VSS(VSS),.VDD(VDD),.Y(g20419),.A(I26846));
  NOT NOT1_6956(.VSS(VSS),.VDD(VDD),.Y(g20420),.A(g17637));
  NOT NOT1_6957(.VSS(VSS),.VDD(VDD),.Y(g20421),.A(g17649));
  NOT NOT1_6958(.VSS(VSS),.VDD(VDD),.Y(g20422),.A(g17655));
  NOT NOT1_6959(.VSS(VSS),.VDD(VDD),.Y(g20423),.A(g17658));
  NOT NOT1_6960(.VSS(VSS),.VDD(VDD),.Y(g20424),.A(g17661));
  NOT NOT1_6961(.VSS(VSS),.VDD(VDD),.Y(g20425),.A(g17664));
  NOT NOT1_6962(.VSS(VSS),.VDD(VDD),.Y(g20426),.A(g17667));
  NOT NOT1_6963(.VSS(VSS),.VDD(VDD),.Y(g20427),.A(g17670));
  NOT NOT1_6964(.VSS(VSS),.VDD(VDD),.Y(g20428),.A(g17676));
  NOT NOT1_6965(.VSS(VSS),.VDD(VDD),.Y(g20429),.A(g17679));
  NOT NOT1_6966(.VSS(VSS),.VDD(VDD),.Y(g20430),.A(g17682));
  NOT NOT1_6967(.VSS(VSS),.VDD(VDD),.Y(g20431),.A(g17685));
  NOT NOT1_6968(.VSS(VSS),.VDD(VDD),.Y(g20432),.A(g17688));
  NOT NOT1_6969(.VSS(VSS),.VDD(VDD),.Y(g20433),.A(g17691));
  NOT NOT1_6970(.VSS(VSS),.VDD(VDD),.Y(g20434),.A(g17698));
  NOT NOT1_6971(.VSS(VSS),.VDD(VDD),.Y(g20435),.A(g17701));
  NOT NOT1_6972(.VSS(VSS),.VDD(VDD),.Y(g20436),.A(g17704));
  NOT NOT1_6973(.VSS(VSS),.VDD(VDD),.Y(g20437),.A(g17707));
  NOT NOT1_6974(.VSS(VSS),.VDD(VDD),.Y(g20438),.A(g17710));
  NOT NOT1_6975(.VSS(VSS),.VDD(VDD),.Y(I26868),.A(g17234));
  NOT NOT1_6976(.VSS(VSS),.VDD(VDD),.Y(g20439),.A(I26868));
  NOT NOT1_6977(.VSS(VSS),.VDD(VDD),.Y(I26871),.A(g17235));
  NOT NOT1_6978(.VSS(VSS),.VDD(VDD),.Y(g20440),.A(I26871));
  NOT NOT1_6979(.VSS(VSS),.VDD(VDD),.Y(I26874),.A(g17236));
  NOT NOT1_6980(.VSS(VSS),.VDD(VDD),.Y(g20441),.A(I26874));
  NOT NOT1_6981(.VSS(VSS),.VDD(VDD),.Y(g20442),.A(g17738));
  NOT NOT1_6982(.VSS(VSS),.VDD(VDD),.Y(g20443),.A(g17749));
  NOT NOT1_6983(.VSS(VSS),.VDD(VDD),.Y(g20444),.A(g17755));
  NOT NOT1_6984(.VSS(VSS),.VDD(VDD),.Y(g20445),.A(g17758));
  NOT NOT1_6985(.VSS(VSS),.VDD(VDD),.Y(g20446),.A(g17761));
  NOT NOT1_6986(.VSS(VSS),.VDD(VDD),.Y(g20447),.A(g17764));
  NOT NOT1_6987(.VSS(VSS),.VDD(VDD),.Y(g20448),.A(g17767));
  NOT NOT1_6988(.VSS(VSS),.VDD(VDD),.Y(g20449),.A(g17770));
  NOT NOT1_6989(.VSS(VSS),.VDD(VDD),.Y(g20450),.A(g17776));
  NOT NOT1_6990(.VSS(VSS),.VDD(VDD),.Y(g20451),.A(g17779));
  NOT NOT1_6991(.VSS(VSS),.VDD(VDD),.Y(g20452),.A(g17782));
  NOT NOT1_6992(.VSS(VSS),.VDD(VDD),.Y(g20453),.A(g17785));
  NOT NOT1_6993(.VSS(VSS),.VDD(VDD),.Y(g20454),.A(g17788));
  NOT NOT1_6994(.VSS(VSS),.VDD(VDD),.Y(g20455),.A(g17791));
  NOT NOT1_6995(.VSS(VSS),.VDD(VDD),.Y(g20456),.A(g17799));
  NOT NOT1_6996(.VSS(VSS),.VDD(VDD),.Y(I26892),.A(g17246));
  NOT NOT1_6997(.VSS(VSS),.VDD(VDD),.Y(g20457),.A(I26892));
  NOT NOT1_6998(.VSS(VSS),.VDD(VDD),.Y(I26895),.A(g17247));
  NOT NOT1_6999(.VSS(VSS),.VDD(VDD),.Y(g20458),.A(I26895));
  NOT NOT1_7000(.VSS(VSS),.VDD(VDD),.Y(I26898),.A(g17248));
  NOT NOT1_7001(.VSS(VSS),.VDD(VDD),.Y(g20459),.A(I26898));
  NOT NOT1_7002(.VSS(VSS),.VDD(VDD),.Y(g20461),.A(g17839));
  NOT NOT1_7003(.VSS(VSS),.VDD(VDD),.Y(g20462),.A(g17850));
  NOT NOT1_7004(.VSS(VSS),.VDD(VDD),.Y(g20463),.A(g17856));
  NOT NOT1_7005(.VSS(VSS),.VDD(VDD),.Y(g20464),.A(g17859));
  NOT NOT1_7006(.VSS(VSS),.VDD(VDD),.Y(g20465),.A(g17862));
  NOT NOT1_7007(.VSS(VSS),.VDD(VDD),.Y(g20466),.A(g17865));
  NOT NOT1_7008(.VSS(VSS),.VDD(VDD),.Y(g20467),.A(g17868));
  NOT NOT1_7009(.VSS(VSS),.VDD(VDD),.Y(g20468),.A(g17871));
  NOT NOT1_7010(.VSS(VSS),.VDD(VDD),.Y(I26910),.A(g17269));
  NOT NOT1_7011(.VSS(VSS),.VDD(VDD),.Y(g20469),.A(I26910));
  NOT NOT1_7012(.VSS(VSS),.VDD(VDD),.Y(I26913),.A(g17270));
  NOT NOT1_7013(.VSS(VSS),.VDD(VDD),.Y(g20470),.A(I26913));
  NOT NOT1_7014(.VSS(VSS),.VDD(VDD),.Y(I26916),.A(g17271));
  NOT NOT1_7015(.VSS(VSS),.VDD(VDD),.Y(g20471),.A(I26916));
  NOT NOT1_7016(.VSS(VSS),.VDD(VDD),.Y(g20476),.A(g17951));
  NOT NOT1_7017(.VSS(VSS),.VDD(VDD),.Y(g20477),.A(g17962));
  NOT NOT1_7018(.VSS(VSS),.VDD(VDD),.Y(I26923),.A(g17302));
  NOT NOT1_7019(.VSS(VSS),.VDD(VDD),.Y(g20478),.A(I26923));
  NOT NOT1_7020(.VSS(VSS),.VDD(VDD),.Y(I26926),.A(g17303));
  NOT NOT1_7021(.VSS(VSS),.VDD(VDD),.Y(g20479),.A(I26926));
  NOT NOT1_7022(.VSS(VSS),.VDD(VDD),.Y(I26931),.A(g17340));
  NOT NOT1_7023(.VSS(VSS),.VDD(VDD),.Y(g20484),.A(I26931));
  NOT NOT1_7024(.VSS(VSS),.VDD(VDD),.Y(I26934),.A(g17341));
  NOT NOT1_7025(.VSS(VSS),.VDD(VDD),.Y(g20485),.A(I26934));
  NOT NOT1_7026(.VSS(VSS),.VDD(VDD),.Y(g20490),.A(g18166));
  NOT NOT1_7027(.VSS(VSS),.VDD(VDD),.Y(I26940),.A(g17383));
  NOT NOT1_7028(.VSS(VSS),.VDD(VDD),.Y(g20491),.A(I26940));
  NOT NOT1_7029(.VSS(VSS),.VDD(VDD),.Y(g20496),.A(g18258));
  NOT NOT1_7030(.VSS(VSS),.VDD(VDD),.Y(I26947),.A(g17429));
  NOT NOT1_7031(.VSS(VSS),.VDD(VDD),.Y(g20498),.A(I26947));
  NOT NOT1_7032(.VSS(VSS),.VDD(VDD),.Y(g20500),.A(g18278));
  NOT NOT1_7033(.VSS(VSS),.VDD(VDD),.Y(g20501),.A(g18334));
  NOT NOT1_7034(.VSS(VSS),.VDD(VDD),.Y(g20504),.A(g18355));
  NOT NOT1_7035(.VSS(VSS),.VDD(VDD),.Y(g20505),.A(g18371));
  NOT NOT1_7036(.VSS(VSS),.VDD(VDD),.Y(g20507),.A(g18351));
  NOT NOT1_7037(.VSS(VSS),.VDD(VDD),.Y(I26960),.A(g16884));
  NOT NOT1_7038(.VSS(VSS),.VDD(VDD),.Y(g20513),.A(I26960));
  NOT NOT1_7039(.VSS(VSS),.VDD(VDD),.Y(g20516),.A(g18432));
  NOT NOT1_7040(.VSS(VSS),.VDD(VDD),.Y(g20517),.A(g18450));
  NOT NOT1_7041(.VSS(VSS),.VDD(VDD),.Y(g20518),.A(g18466));
  NOT NOT1_7042(.VSS(VSS),.VDD(VDD),.Y(I26966),.A(g17051));
  NOT NOT1_7043(.VSS(VSS),.VDD(VDD),.Y(g20519),.A(I26966));
  NOT NOT1_7044(.VSS(VSS),.VDD(VDD),.Y(g20526),.A(g18446));
  NOT NOT1_7045(.VSS(VSS),.VDD(VDD),.Y(I26972),.A(g16913));
  NOT NOT1_7046(.VSS(VSS),.VDD(VDD),.Y(g20531),.A(I26972));
  NOT NOT1_7047(.VSS(VSS),.VDD(VDD),.Y(g20534),.A(g18505));
  NOT NOT1_7048(.VSS(VSS),.VDD(VDD),.Y(g20535),.A(g18523));
  NOT NOT1_7049(.VSS(VSS),.VDD(VDD),.Y(g20536),.A(g18539));
  NOT NOT1_7050(.VSS(VSS),.VDD(VDD),.Y(I26980),.A(g17086));
  NOT NOT1_7051(.VSS(VSS),.VDD(VDD),.Y(g20539),.A(I26980));
  NOT NOT1_7052(.VSS(VSS),.VDD(VDD),.Y(g20545),.A(g18519));
  NOT NOT1_7053(.VSS(VSS),.VDD(VDD),.Y(I26985),.A(g16943));
  NOT NOT1_7054(.VSS(VSS),.VDD(VDD),.Y(g20550),.A(I26985));
  NOT NOT1_7055(.VSS(VSS),.VDD(VDD),.Y(g20553),.A(g18569));
  NOT NOT1_7056(.VSS(VSS),.VDD(VDD),.Y(g20554),.A(g18587));
  NOT NOT1_7057(.VSS(VSS),.VDD(VDD),.Y(I26990),.A(g19145));
  NOT NOT1_7058(.VSS(VSS),.VDD(VDD),.Y(g20555),.A(I26990));
  NOT NOT1_7059(.VSS(VSS),.VDD(VDD),.Y(I26993),.A(g19159));
  NOT NOT1_7060(.VSS(VSS),.VDD(VDD),.Y(g20556),.A(I26993));
  NOT NOT1_7061(.VSS(VSS),.VDD(VDD),.Y(I26996),.A(g19169));
  NOT NOT1_7062(.VSS(VSS),.VDD(VDD),.Y(g20557),.A(I26996));
  NOT NOT1_7063(.VSS(VSS),.VDD(VDD),.Y(I26999),.A(g19543));
  NOT NOT1_7064(.VSS(VSS),.VDD(VDD),.Y(g20558),.A(I26999));
  NOT NOT1_7065(.VSS(VSS),.VDD(VDD),.Y(I27002),.A(g19147));
  NOT NOT1_7066(.VSS(VSS),.VDD(VDD),.Y(g20559),.A(I27002));
  NOT NOT1_7067(.VSS(VSS),.VDD(VDD),.Y(I27005),.A(g19164));
  NOT NOT1_7068(.VSS(VSS),.VDD(VDD),.Y(g20560),.A(I27005));
  NOT NOT1_7069(.VSS(VSS),.VDD(VDD),.Y(I27008),.A(g19175));
  NOT NOT1_7070(.VSS(VSS),.VDD(VDD),.Y(g20561),.A(I27008));
  NOT NOT1_7071(.VSS(VSS),.VDD(VDD),.Y(I27011),.A(g19546));
  NOT NOT1_7072(.VSS(VSS),.VDD(VDD),.Y(g20562),.A(I27011));
  NOT NOT1_7073(.VSS(VSS),.VDD(VDD),.Y(I27014),.A(g19151));
  NOT NOT1_7074(.VSS(VSS),.VDD(VDD),.Y(g20563),.A(I27014));
  NOT NOT1_7075(.VSS(VSS),.VDD(VDD),.Y(I27017),.A(g19170));
  NOT NOT1_7076(.VSS(VSS),.VDD(VDD),.Y(g20564),.A(I27017));
  NOT NOT1_7077(.VSS(VSS),.VDD(VDD),.Y(I27020),.A(g19182));
  NOT NOT1_7078(.VSS(VSS),.VDD(VDD),.Y(g20565),.A(I27020));
  NOT NOT1_7079(.VSS(VSS),.VDD(VDD),.Y(I27023),.A(g19550));
  NOT NOT1_7080(.VSS(VSS),.VDD(VDD),.Y(g20566),.A(I27023));
  NOT NOT1_7081(.VSS(VSS),.VDD(VDD),.Y(I27026),.A(g19156));
  NOT NOT1_7082(.VSS(VSS),.VDD(VDD),.Y(g20567),.A(I27026));
  NOT NOT1_7083(.VSS(VSS),.VDD(VDD),.Y(I27029),.A(g19176));
  NOT NOT1_7084(.VSS(VSS),.VDD(VDD),.Y(g20568),.A(I27029));
  NOT NOT1_7085(.VSS(VSS),.VDD(VDD),.Y(I27032),.A(g19189));
  NOT NOT1_7086(.VSS(VSS),.VDD(VDD),.Y(g20569),.A(I27032));
  NOT NOT1_7087(.VSS(VSS),.VDD(VDD),.Y(I27035),.A(g19556));
  NOT NOT1_7088(.VSS(VSS),.VDD(VDD),.Y(g20570),.A(I27035));
  NOT NOT1_7089(.VSS(VSS),.VDD(VDD),.Y(I27038),.A(g20082));
  NOT NOT1_7090(.VSS(VSS),.VDD(VDD),.Y(g20571),.A(I27038));
  NOT NOT1_7091(.VSS(VSS),.VDD(VDD),.Y(I27041),.A(g19237));
  NOT NOT1_7092(.VSS(VSS),.VDD(VDD),.Y(g20572),.A(I27041));
  NOT NOT1_7093(.VSS(VSS),.VDD(VDD),.Y(I27044),.A(g19247));
  NOT NOT1_7094(.VSS(VSS),.VDD(VDD),.Y(g20573),.A(I27044));
  NOT NOT1_7095(.VSS(VSS),.VDD(VDD),.Y(I27047),.A(g19258));
  NOT NOT1_7096(.VSS(VSS),.VDD(VDD),.Y(g20574),.A(I27047));
  NOT NOT1_7097(.VSS(VSS),.VDD(VDD),.Y(I27050),.A(g19183));
  NOT NOT1_7098(.VSS(VSS),.VDD(VDD),.Y(g20575),.A(I27050));
  NOT NOT1_7099(.VSS(VSS),.VDD(VDD),.Y(I27053),.A(g19190));
  NOT NOT1_7100(.VSS(VSS),.VDD(VDD),.Y(g20576),.A(I27053));
  NOT NOT1_7101(.VSS(VSS),.VDD(VDD),.Y(I27056),.A(g19196));
  NOT NOT1_7102(.VSS(VSS),.VDD(VDD),.Y(g20577),.A(I27056));
  NOT NOT1_7103(.VSS(VSS),.VDD(VDD),.Y(I27059),.A(g19207));
  NOT NOT1_7104(.VSS(VSS),.VDD(VDD),.Y(g20578),.A(I27059));
  NOT NOT1_7105(.VSS(VSS),.VDD(VDD),.Y(I27062),.A(g19217));
  NOT NOT1_7106(.VSS(VSS),.VDD(VDD),.Y(g20579),.A(I27062));
  NOT NOT1_7107(.VSS(VSS),.VDD(VDD),.Y(I27065),.A(g19270));
  NOT NOT1_7108(.VSS(VSS),.VDD(VDD),.Y(g20580),.A(I27065));
  NOT NOT1_7109(.VSS(VSS),.VDD(VDD),.Y(I27068),.A(g19197));
  NOT NOT1_7110(.VSS(VSS),.VDD(VDD),.Y(g20581),.A(I27068));
  NOT NOT1_7111(.VSS(VSS),.VDD(VDD),.Y(I27071),.A(g19218));
  NOT NOT1_7112(.VSS(VSS),.VDD(VDD),.Y(g20582),.A(I27071));
  NOT NOT1_7113(.VSS(VSS),.VDD(VDD),.Y(I27074),.A(g19238));
  NOT NOT1_7114(.VSS(VSS),.VDD(VDD),.Y(g20583),.A(I27074));
  NOT NOT1_7115(.VSS(VSS),.VDD(VDD),.Y(I27077),.A(g19259));
  NOT NOT1_7116(.VSS(VSS),.VDD(VDD),.Y(g20584),.A(I27077));
  NOT NOT1_7117(.VSS(VSS),.VDD(VDD),.Y(I27080),.A(g19198));
  NOT NOT1_7118(.VSS(VSS),.VDD(VDD),.Y(g20585),.A(I27080));
  NOT NOT1_7119(.VSS(VSS),.VDD(VDD),.Y(I27083),.A(g19208));
  NOT NOT1_7120(.VSS(VSS),.VDD(VDD),.Y(g20586),.A(I27083));
  NOT NOT1_7121(.VSS(VSS),.VDD(VDD),.Y(I27086),.A(g19229));
  NOT NOT1_7122(.VSS(VSS),.VDD(VDD),.Y(g20587),.A(I27086));
  NOT NOT1_7123(.VSS(VSS),.VDD(VDD),.Y(I27089),.A(g20105));
  NOT NOT1_7124(.VSS(VSS),.VDD(VDD),.Y(g20588),.A(I27089));
  NOT NOT1_7125(.VSS(VSS),.VDD(VDD),.Y(I27092),.A(g19174));
  NOT NOT1_7126(.VSS(VSS),.VDD(VDD),.Y(g20589),.A(I27092));
  NOT NOT1_7127(.VSS(VSS),.VDD(VDD),.Y(I27095),.A(g19185));
  NOT NOT1_7128(.VSS(VSS),.VDD(VDD),.Y(g20590),.A(I27095));
  NOT NOT1_7129(.VSS(VSS),.VDD(VDD),.Y(I27098),.A(g19199));
  NOT NOT1_7130(.VSS(VSS),.VDD(VDD),.Y(g20591),.A(I27098));
  NOT NOT1_7131(.VSS(VSS),.VDD(VDD),.Y(I27101),.A(g19220));
  NOT NOT1_7132(.VSS(VSS),.VDD(VDD),.Y(g20592),.A(I27101));
  NOT NOT1_7133(.VSS(VSS),.VDD(VDD),.Y(I27104),.A(g19239));
  NOT NOT1_7134(.VSS(VSS),.VDD(VDD),.Y(g20593),.A(I27104));
  NOT NOT1_7135(.VSS(VSS),.VDD(VDD),.Y(I27107),.A(g19249));
  NOT NOT1_7136(.VSS(VSS),.VDD(VDD),.Y(g20594),.A(I27107));
  NOT NOT1_7137(.VSS(VSS),.VDD(VDD),.Y(I27110),.A(g19622));
  NOT NOT1_7138(.VSS(VSS),.VDD(VDD),.Y(g20595),.A(I27110));
  NOT NOT1_7139(.VSS(VSS),.VDD(VDD),.Y(I27113),.A(g19689));
  NOT NOT1_7140(.VSS(VSS),.VDD(VDD),.Y(g20596),.A(I27113));
  NOT NOT1_7141(.VSS(VSS),.VDD(VDD),.Y(I27116),.A(g19762));
  NOT NOT1_7142(.VSS(VSS),.VDD(VDD),.Y(g20597),.A(I27116));
  NOT NOT1_7143(.VSS(VSS),.VDD(VDD),.Y(I27119),.A(g19563));
  NOT NOT1_7144(.VSS(VSS),.VDD(VDD),.Y(g20598),.A(I27119));
  NOT NOT1_7145(.VSS(VSS),.VDD(VDD),.Y(I27122),.A(g19595));
  NOT NOT1_7146(.VSS(VSS),.VDD(VDD),.Y(g20599),.A(I27122));
  NOT NOT1_7147(.VSS(VSS),.VDD(VDD),.Y(I27125),.A(g19652));
  NOT NOT1_7148(.VSS(VSS),.VDD(VDD),.Y(g20600),.A(I27125));
  NOT NOT1_7149(.VSS(VSS),.VDD(VDD),.Y(I27128),.A(g19725));
  NOT NOT1_7150(.VSS(VSS),.VDD(VDD),.Y(g20601),.A(I27128));
  NOT NOT1_7151(.VSS(VSS),.VDD(VDD),.Y(I27131),.A(g19798));
  NOT NOT1_7152(.VSS(VSS),.VDD(VDD),.Y(g20602),.A(I27131));
  NOT NOT1_7153(.VSS(VSS),.VDD(VDD),.Y(I27134),.A(g19573));
  NOT NOT1_7154(.VSS(VSS),.VDD(VDD),.Y(g20603),.A(I27134));
  NOT NOT1_7155(.VSS(VSS),.VDD(VDD),.Y(I27137),.A(g19596));
  NOT NOT1_7156(.VSS(VSS),.VDD(VDD),.Y(g20604),.A(I27137));
  NOT NOT1_7157(.VSS(VSS),.VDD(VDD),.Y(I27140),.A(g19690));
  NOT NOT1_7158(.VSS(VSS),.VDD(VDD),.Y(g20605),.A(I27140));
  NOT NOT1_7159(.VSS(VSS),.VDD(VDD),.Y(I27143),.A(g19763));
  NOT NOT1_7160(.VSS(VSS),.VDD(VDD),.Y(g20606),.A(I27143));
  NOT NOT1_7161(.VSS(VSS),.VDD(VDD),.Y(I27146),.A(g19838));
  NOT NOT1_7162(.VSS(VSS),.VDD(VDD),.Y(g20607),.A(I27146));
  NOT NOT1_7163(.VSS(VSS),.VDD(VDD),.Y(I27149),.A(g19893));
  NOT NOT1_7164(.VSS(VSS),.VDD(VDD),.Y(g20608),.A(I27149));
  NOT NOT1_7165(.VSS(VSS),.VDD(VDD),.Y(I27152),.A(g20360));
  NOT NOT1_7166(.VSS(VSS),.VDD(VDD),.Y(g20609),.A(I27152));
  NOT NOT1_7167(.VSS(VSS),.VDD(VDD),.Y(I27155),.A(g20395));
  NOT NOT1_7168(.VSS(VSS),.VDD(VDD),.Y(g20610),.A(I27155));
  NOT NOT1_7169(.VSS(VSS),.VDD(VDD),.Y(I27158),.A(g20439));
  NOT NOT1_7170(.VSS(VSS),.VDD(VDD),.Y(g20611),.A(I27158));
  NOT NOT1_7171(.VSS(VSS),.VDD(VDD),.Y(I27161),.A(g20377));
  NOT NOT1_7172(.VSS(VSS),.VDD(VDD),.Y(g20612),.A(I27161));
  NOT NOT1_7173(.VSS(VSS),.VDD(VDD),.Y(I27164),.A(g20418));
  NOT NOT1_7174(.VSS(VSS),.VDD(VDD),.Y(g20613),.A(I27164));
  NOT NOT1_7175(.VSS(VSS),.VDD(VDD),.Y(I27167),.A(g20457));
  NOT NOT1_7176(.VSS(VSS),.VDD(VDD),.Y(g20614),.A(I27167));
  NOT NOT1_7177(.VSS(VSS),.VDD(VDD),.Y(I27170),.A(g20396));
  NOT NOT1_7178(.VSS(VSS),.VDD(VDD),.Y(g20615),.A(I27170));
  NOT NOT1_7179(.VSS(VSS),.VDD(VDD),.Y(I27173),.A(g20440));
  NOT NOT1_7180(.VSS(VSS),.VDD(VDD),.Y(g20616),.A(I27173));
  NOT NOT1_7181(.VSS(VSS),.VDD(VDD),.Y(I27176),.A(g20469));
  NOT NOT1_7182(.VSS(VSS),.VDD(VDD),.Y(g20617),.A(I27176));
  NOT NOT1_7183(.VSS(VSS),.VDD(VDD),.Y(I27179),.A(g20419));
  NOT NOT1_7184(.VSS(VSS),.VDD(VDD),.Y(g20618),.A(I27179));
  NOT NOT1_7185(.VSS(VSS),.VDD(VDD),.Y(I27182),.A(g20458));
  NOT NOT1_7186(.VSS(VSS),.VDD(VDD),.Y(g20619),.A(I27182));
  NOT NOT1_7187(.VSS(VSS),.VDD(VDD),.Y(I27185),.A(g20478));
  NOT NOT1_7188(.VSS(VSS),.VDD(VDD),.Y(g20620),.A(I27185));
  NOT NOT1_7189(.VSS(VSS),.VDD(VDD),.Y(I27188),.A(g20441));
  NOT NOT1_7190(.VSS(VSS),.VDD(VDD),.Y(g20621),.A(I27188));
  NOT NOT1_7191(.VSS(VSS),.VDD(VDD),.Y(I27191),.A(g20470));
  NOT NOT1_7192(.VSS(VSS),.VDD(VDD),.Y(g20622),.A(I27191));
  NOT NOT1_7193(.VSS(VSS),.VDD(VDD),.Y(I27194),.A(g20484));
  NOT NOT1_7194(.VSS(VSS),.VDD(VDD),.Y(g20623),.A(I27194));
  NOT NOT1_7195(.VSS(VSS),.VDD(VDD),.Y(I27197),.A(g20459));
  NOT NOT1_7196(.VSS(VSS),.VDD(VDD),.Y(g20624),.A(I27197));
  NOT NOT1_7197(.VSS(VSS),.VDD(VDD),.Y(I27200),.A(g20479));
  NOT NOT1_7198(.VSS(VSS),.VDD(VDD),.Y(g20625),.A(I27200));
  NOT NOT1_7199(.VSS(VSS),.VDD(VDD),.Y(I27203),.A(g20491));
  NOT NOT1_7200(.VSS(VSS),.VDD(VDD),.Y(g20626),.A(I27203));
  NOT NOT1_7201(.VSS(VSS),.VDD(VDD),.Y(I27206),.A(g20471));
  NOT NOT1_7202(.VSS(VSS),.VDD(VDD),.Y(g20627),.A(I27206));
  NOT NOT1_7203(.VSS(VSS),.VDD(VDD),.Y(I27209),.A(g20485));
  NOT NOT1_7204(.VSS(VSS),.VDD(VDD),.Y(g20628),.A(I27209));
  NOT NOT1_7205(.VSS(VSS),.VDD(VDD),.Y(I27212),.A(g20498));
  NOT NOT1_7206(.VSS(VSS),.VDD(VDD),.Y(g20629),.A(I27212));
  NOT NOT1_7207(.VSS(VSS),.VDD(VDD),.Y(I27215),.A(g19158));
  NOT NOT1_7208(.VSS(VSS),.VDD(VDD),.Y(g20630),.A(I27215));
  NOT NOT1_7209(.VSS(VSS),.VDD(VDD),.Y(I27218),.A(g19168));
  NOT NOT1_7210(.VSS(VSS),.VDD(VDD),.Y(g20631),.A(I27218));
  NOT NOT1_7211(.VSS(VSS),.VDD(VDD),.Y(I27221),.A(g19180));
  NOT NOT1_7212(.VSS(VSS),.VDD(VDD),.Y(g20632),.A(I27221));
  NOT NOT1_7213(.VSS(VSS),.VDD(VDD),.Y(I27225),.A(g19358));
  NOT NOT1_7214(.VSS(VSS),.VDD(VDD),.Y(g20634),.A(I27225));
  NOT NOT1_7215(.VSS(VSS),.VDD(VDD),.Y(I27228),.A(g19390));
  NOT NOT1_7216(.VSS(VSS),.VDD(VDD),.Y(g20637),.A(I27228));
  NOT NOT1_7217(.VSS(VSS),.VDD(VDD),.Y(I27232),.A(g19401));
  NOT NOT1_7218(.VSS(VSS),.VDD(VDD),.Y(g20641),.A(I27232));
  NOT NOT1_7219(.VSS(VSS),.VDD(VDD),.Y(I27235),.A(g19420));
  NOT NOT1_7220(.VSS(VSS),.VDD(VDD),.Y(g20644),.A(I27235));
  NOT NOT1_7221(.VSS(VSS),.VDD(VDD),.Y(I27240),.A(g19335));
  NOT NOT1_7222(.VSS(VSS),.VDD(VDD),.Y(g20649),.A(I27240));
  NOT NOT1_7223(.VSS(VSS),.VDD(VDD),.Y(I27243),.A(g19335));
  NOT NOT1_7224(.VSS(VSS),.VDD(VDD),.Y(g20652),.A(I27243));
  NOT NOT1_7225(.VSS(VSS),.VDD(VDD),.Y(I27246),.A(g19335));
  NOT NOT1_7226(.VSS(VSS),.VDD(VDD),.Y(g20655),.A(I27246));
  NOT NOT1_7227(.VSS(VSS),.VDD(VDD),.Y(I27250),.A(g19390));
  NOT NOT1_7228(.VSS(VSS),.VDD(VDD),.Y(g20659),.A(I27250));
  NOT NOT1_7229(.VSS(VSS),.VDD(VDD),.Y(I27253),.A(g19420));
  NOT NOT1_7230(.VSS(VSS),.VDD(VDD),.Y(g20662),.A(I27253));
  NOT NOT1_7231(.VSS(VSS),.VDD(VDD),.Y(I27257),.A(g19431));
  NOT NOT1_7232(.VSS(VSS),.VDD(VDD),.Y(g20666),.A(I27257));
  NOT NOT1_7233(.VSS(VSS),.VDD(VDD),.Y(I27260),.A(g19457));
  NOT NOT1_7234(.VSS(VSS),.VDD(VDD),.Y(g20669),.A(I27260));
  NOT NOT1_7235(.VSS(VSS),.VDD(VDD),.Y(I27264),.A(g19358));
  NOT NOT1_7236(.VSS(VSS),.VDD(VDD),.Y(g20673),.A(I27264));
  NOT NOT1_7237(.VSS(VSS),.VDD(VDD),.Y(I27267),.A(g19358));
  NOT NOT1_7238(.VSS(VSS),.VDD(VDD),.Y(g20676),.A(I27267));
  NOT NOT1_7239(.VSS(VSS),.VDD(VDD),.Y(I27270),.A(g19335));
  NOT NOT1_7240(.VSS(VSS),.VDD(VDD),.Y(g20679),.A(I27270));
  NOT NOT1_7241(.VSS(VSS),.VDD(VDD),.Y(I27275),.A(g19369));
  NOT NOT1_7242(.VSS(VSS),.VDD(VDD),.Y(g20684),.A(I27275));
  NOT NOT1_7243(.VSS(VSS),.VDD(VDD),.Y(I27278),.A(g19369));
  NOT NOT1_7244(.VSS(VSS),.VDD(VDD),.Y(g20687),.A(I27278));
  NOT NOT1_7245(.VSS(VSS),.VDD(VDD),.Y(I27281),.A(g19369));
  NOT NOT1_7246(.VSS(VSS),.VDD(VDD),.Y(g20690),.A(I27281));
  NOT NOT1_7247(.VSS(VSS),.VDD(VDD),.Y(I27285),.A(g19420));
  NOT NOT1_7248(.VSS(VSS),.VDD(VDD),.Y(g20694),.A(I27285));
  NOT NOT1_7249(.VSS(VSS),.VDD(VDD),.Y(I27288),.A(g19457));
  NOT NOT1_7250(.VSS(VSS),.VDD(VDD),.Y(g20697),.A(I27288));
  NOT NOT1_7251(.VSS(VSS),.VDD(VDD),.Y(I27293),.A(g19335));
  NOT NOT1_7252(.VSS(VSS),.VDD(VDD),.Y(g20704),.A(I27293));
  NOT NOT1_7253(.VSS(VSS),.VDD(VDD),.Y(I27297),.A(g19390));
  NOT NOT1_7254(.VSS(VSS),.VDD(VDD),.Y(g20708),.A(I27297));
  NOT NOT1_7255(.VSS(VSS),.VDD(VDD),.Y(I27300),.A(g19390));
  NOT NOT1_7256(.VSS(VSS),.VDD(VDD),.Y(g20711),.A(I27300));
  NOT NOT1_7257(.VSS(VSS),.VDD(VDD),.Y(I27303),.A(g19369));
  NOT NOT1_7258(.VSS(VSS),.VDD(VDD),.Y(g20714),.A(I27303));
  NOT NOT1_7259(.VSS(VSS),.VDD(VDD),.Y(I27308),.A(g19401));
  NOT NOT1_7260(.VSS(VSS),.VDD(VDD),.Y(g20719),.A(I27308));
  NOT NOT1_7261(.VSS(VSS),.VDD(VDD),.Y(I27311),.A(g19401));
  NOT NOT1_7262(.VSS(VSS),.VDD(VDD),.Y(g20722),.A(I27311));
  NOT NOT1_7263(.VSS(VSS),.VDD(VDD),.Y(I27314),.A(g19401));
  NOT NOT1_7264(.VSS(VSS),.VDD(VDD),.Y(g20725),.A(I27314));
  NOT NOT1_7265(.VSS(VSS),.VDD(VDD),.Y(I27318),.A(g19457));
  NOT NOT1_7266(.VSS(VSS),.VDD(VDD),.Y(g20729),.A(I27318));
  NOT NOT1_7267(.VSS(VSS),.VDD(VDD),.Y(I27321),.A(g19335));
  NOT NOT1_7268(.VSS(VSS),.VDD(VDD),.Y(g20732),.A(I27321));
  NOT NOT1_7269(.VSS(VSS),.VDD(VDD),.Y(I27324),.A(g19358));
  NOT NOT1_7270(.VSS(VSS),.VDD(VDD),.Y(g20735),.A(I27324));
  NOT NOT1_7271(.VSS(VSS),.VDD(VDD),.Y(I27328),.A(g19369));
  NOT NOT1_7272(.VSS(VSS),.VDD(VDD),.Y(g20739),.A(I27328));
  NOT NOT1_7273(.VSS(VSS),.VDD(VDD),.Y(I27332),.A(g19420));
  NOT NOT1_7274(.VSS(VSS),.VDD(VDD),.Y(g20743),.A(I27332));
  NOT NOT1_7275(.VSS(VSS),.VDD(VDD),.Y(I27335),.A(g19420));
  NOT NOT1_7276(.VSS(VSS),.VDD(VDD),.Y(g20746),.A(I27335));
  NOT NOT1_7277(.VSS(VSS),.VDD(VDD),.Y(I27338),.A(g19401));
  NOT NOT1_7278(.VSS(VSS),.VDD(VDD),.Y(g20749),.A(I27338));
  NOT NOT1_7279(.VSS(VSS),.VDD(VDD),.Y(I27343),.A(g19431));
  NOT NOT1_7280(.VSS(VSS),.VDD(VDD),.Y(g20754),.A(I27343));
  NOT NOT1_7281(.VSS(VSS),.VDD(VDD),.Y(I27346),.A(g19431));
  NOT NOT1_7282(.VSS(VSS),.VDD(VDD),.Y(g20757),.A(I27346));
  NOT NOT1_7283(.VSS(VSS),.VDD(VDD),.Y(I27349),.A(g19431));
  NOT NOT1_7284(.VSS(VSS),.VDD(VDD),.Y(g20760),.A(I27349));
  NOT NOT1_7285(.VSS(VSS),.VDD(VDD),.Y(I27352),.A(g19358));
  NOT NOT1_7286(.VSS(VSS),.VDD(VDD),.Y(g20763),.A(I27352));
  NOT NOT1_7287(.VSS(VSS),.VDD(VDD),.Y(I27355),.A(g19335));
  NOT NOT1_7288(.VSS(VSS),.VDD(VDD),.Y(g20766),.A(I27355));
  NOT NOT1_7289(.VSS(VSS),.VDD(VDD),.Y(I27358),.A(g19369));
  NOT NOT1_7290(.VSS(VSS),.VDD(VDD),.Y(g20769),.A(I27358));
  NOT NOT1_7291(.VSS(VSS),.VDD(VDD),.Y(I27361),.A(g19390));
  NOT NOT1_7292(.VSS(VSS),.VDD(VDD),.Y(g20772),.A(I27361));
  NOT NOT1_7293(.VSS(VSS),.VDD(VDD),.Y(I27365),.A(g19401));
  NOT NOT1_7294(.VSS(VSS),.VDD(VDD),.Y(g20776),.A(I27365));
  NOT NOT1_7295(.VSS(VSS),.VDD(VDD),.Y(I27369),.A(g19457));
  NOT NOT1_7296(.VSS(VSS),.VDD(VDD),.Y(g20780),.A(I27369));
  NOT NOT1_7297(.VSS(VSS),.VDD(VDD),.Y(I27372),.A(g19457));
  NOT NOT1_7298(.VSS(VSS),.VDD(VDD),.Y(g20783),.A(I27372));
  NOT NOT1_7299(.VSS(VSS),.VDD(VDD),.Y(I27375),.A(g19431));
  NOT NOT1_7300(.VSS(VSS),.VDD(VDD),.Y(g20786),.A(I27375));
  NOT NOT1_7301(.VSS(VSS),.VDD(VDD),.Y(I27379),.A(g19358));
  NOT NOT1_7302(.VSS(VSS),.VDD(VDD),.Y(g20790),.A(I27379));
  NOT NOT1_7303(.VSS(VSS),.VDD(VDD),.Y(I27382),.A(g19390));
  NOT NOT1_7304(.VSS(VSS),.VDD(VDD),.Y(g20793),.A(I27382));
  NOT NOT1_7305(.VSS(VSS),.VDD(VDD),.Y(I27385),.A(g19369));
  NOT NOT1_7306(.VSS(VSS),.VDD(VDD),.Y(g20796),.A(I27385));
  NOT NOT1_7307(.VSS(VSS),.VDD(VDD),.Y(I27388),.A(g19401));
  NOT NOT1_7308(.VSS(VSS),.VDD(VDD),.Y(g20799),.A(I27388));
  NOT NOT1_7309(.VSS(VSS),.VDD(VDD),.Y(I27391),.A(g19420));
  NOT NOT1_7310(.VSS(VSS),.VDD(VDD),.Y(g20802),.A(I27391));
  NOT NOT1_7311(.VSS(VSS),.VDD(VDD),.Y(I27395),.A(g19431));
  NOT NOT1_7312(.VSS(VSS),.VDD(VDD),.Y(g20806),.A(I27395));
  NOT NOT1_7313(.VSS(VSS),.VDD(VDD),.Y(I27399),.A(g19390));
  NOT NOT1_7314(.VSS(VSS),.VDD(VDD),.Y(g20810),.A(I27399));
  NOT NOT1_7315(.VSS(VSS),.VDD(VDD),.Y(I27402),.A(g19420));
  NOT NOT1_7316(.VSS(VSS),.VDD(VDD),.Y(g20813),.A(I27402));
  NOT NOT1_7317(.VSS(VSS),.VDD(VDD),.Y(I27405),.A(g19401));
  NOT NOT1_7318(.VSS(VSS),.VDD(VDD),.Y(g20816),.A(I27405));
  NOT NOT1_7319(.VSS(VSS),.VDD(VDD),.Y(I27408),.A(g19431));
  NOT NOT1_7320(.VSS(VSS),.VDD(VDD),.Y(g20819),.A(I27408));
  NOT NOT1_7321(.VSS(VSS),.VDD(VDD),.Y(I27411),.A(g19457));
  NOT NOT1_7322(.VSS(VSS),.VDD(VDD),.Y(g20822),.A(I27411));
  NOT NOT1_7323(.VSS(VSS),.VDD(VDD),.Y(I27416),.A(g19420));
  NOT NOT1_7324(.VSS(VSS),.VDD(VDD),.Y(g20827),.A(I27416));
  NOT NOT1_7325(.VSS(VSS),.VDD(VDD),.Y(I27419),.A(g19457));
  NOT NOT1_7326(.VSS(VSS),.VDD(VDD),.Y(g20830),.A(I27419));
  NOT NOT1_7327(.VSS(VSS),.VDD(VDD),.Y(I27422),.A(g19431));
  NOT NOT1_7328(.VSS(VSS),.VDD(VDD),.Y(g20833),.A(I27422));
  NOT NOT1_7329(.VSS(VSS),.VDD(VDD),.Y(I27426),.A(g19457));
  NOT NOT1_7330(.VSS(VSS),.VDD(VDD),.Y(g20837),.A(I27426));
  NOT NOT1_7331(.VSS(VSS),.VDD(VDD),.Y(g20842),.A(g19441));
  NOT NOT1_7332(.VSS(VSS),.VDD(VDD),.Y(g20850),.A(g19468));
  NOT NOT1_7333(.VSS(VSS),.VDD(VDD),.Y(g20858),.A(g19491));
  NOT NOT1_7334(.VSS(VSS),.VDD(VDD),.Y(g20866),.A(g19512));
  NOT NOT1_7335(.VSS(VSS),.VDD(VDD),.Y(g20885),.A(g19865));
  NOT NOT1_7336(.VSS(VSS),.VDD(VDD),.Y(g20904),.A(g19896));
  NOT NOT1_7337(.VSS(VSS),.VDD(VDD),.Y(g20928),.A(g19921));
  NOT NOT1_7338(.VSS(VSS),.VDD(VDD),.Y(I27488),.A(g20310));
  NOT NOT1_7339(.VSS(VSS),.VDD(VDD),.Y(g20942),.A(I27488));
  NOT NOT1_7340(.VSS(VSS),.VDD(VDD),.Y(I27491),.A(g20314));
  NOT NOT1_7341(.VSS(VSS),.VDD(VDD),.Y(g20943),.A(I27491));
  NOT NOT1_7342(.VSS(VSS),.VDD(VDD),.Y(g20956),.A(g19936));
  NOT NOT1_7343(.VSS(VSS),.VDD(VDD),.Y(I27516),.A(g20333));
  NOT NOT1_7344(.VSS(VSS),.VDD(VDD),.Y(g20971),.A(I27516));
  NOT NOT1_7345(.VSS(VSS),.VDD(VDD),.Y(I27531),.A(g20343));
  NOT NOT1_7346(.VSS(VSS),.VDD(VDD),.Y(g20984),.A(I27531));
  NOT NOT1_7347(.VSS(VSS),.VDD(VDD),.Y(I27534),.A(g20083));
  NOT NOT1_7348(.VSS(VSS),.VDD(VDD),.Y(g20985),.A(I27534));
  NOT NOT1_7349(.VSS(VSS),.VDD(VDD),.Y(I27537),.A(g19957));
  NOT NOT1_7350(.VSS(VSS),.VDD(VDD),.Y(g20986),.A(I27537));
  NOT NOT1_7351(.VSS(VSS),.VDD(VDD),.Y(I27549),.A(g20353));
  NOT NOT1_7352(.VSS(VSS),.VDD(VDD),.Y(g20998),.A(I27549));
  NOT NOT1_7353(.VSS(VSS),.VDD(VDD),.Y(I27565),.A(g19987));
  NOT NOT1_7354(.VSS(VSS),.VDD(VDD),.Y(g21012),.A(I27565));
  NOT NOT1_7355(.VSS(VSS),.VDD(VDD),.Y(I27577),.A(g20375));
  NOT NOT1_7356(.VSS(VSS),.VDD(VDD),.Y(g21024),.A(I27577));
  NOT NOT1_7357(.VSS(VSS),.VDD(VDD),.Y(I27585),.A(g20376));
  NOT NOT1_7358(.VSS(VSS),.VDD(VDD),.Y(g21030),.A(I27585));
  NOT NOT1_7359(.VSS(VSS),.VDD(VDD),.Y(I27593),.A(g20025));
  NOT NOT1_7360(.VSS(VSS),.VDD(VDD),.Y(g21036),.A(I27593));
  NOT NOT1_7361(.VSS(VSS),.VDD(VDD),.Y(g21050),.A(g20513));
  NOT NOT1_7362(.VSS(VSS),.VDD(VDD),.Y(I27614),.A(g20067));
  NOT NOT1_7363(.VSS(VSS),.VDD(VDD),.Y(g21057),.A(I27614));
  NOT NOT1_7364(.VSS(VSS),.VDD(VDD),.Y(I27621),.A(g20417));
  NOT NOT1_7365(.VSS(VSS),.VDD(VDD),.Y(g21064),.A(I27621));
  NOT NOT1_7366(.VSS(VSS),.VDD(VDD),.Y(g21066),.A(g20519));
  NOT NOT1_7367(.VSS(VSS),.VDD(VDD),.Y(g21069),.A(g20531));
  NOT NOT1_7368(.VSS(VSS),.VDD(VDD),.Y(g21076),.A(g20539));
  NOT NOT1_7369(.VSS(VSS),.VDD(VDD),.Y(g21079),.A(g20550));
  NOT NOT1_7370(.VSS(VSS),.VDD(VDD),.Y(I27646),.A(g20507));
  NOT NOT1_7371(.VSS(VSS),.VDD(VDD),.Y(g21087),.A(I27646));
  NOT NOT1_7372(.VSS(VSS),.VDD(VDD),.Y(g21090),.A(g19064));
  NOT NOT1_7373(.VSS(VSS),.VDD(VDD),.Y(g21093),.A(g19075));
  NOT NOT1_7374(.VSS(VSS),.VDD(VDD),.Y(I27658),.A(g20526));
  NOT NOT1_7375(.VSS(VSS),.VDD(VDD),.Y(g21099),.A(I27658));
  NOT NOT1_7376(.VSS(VSS),.VDD(VDD),.Y(g21102),.A(g19081));
  NOT NOT1_7377(.VSS(VSS),.VDD(VDD),.Y(I27667),.A(g20507));
  NOT NOT1_7378(.VSS(VSS),.VDD(VDD),.Y(g21108),.A(I27667));
  NOT NOT1_7379(.VSS(VSS),.VDD(VDD),.Y(I27672),.A(g20545));
  NOT NOT1_7380(.VSS(VSS),.VDD(VDD),.Y(g21113),.A(I27672));
  NOT NOT1_7381(.VSS(VSS),.VDD(VDD),.Y(I27684),.A(g20526));
  NOT NOT1_7382(.VSS(VSS),.VDD(VDD),.Y(g21125),.A(I27684));
  NOT NOT1_7383(.VSS(VSS),.VDD(VDD),.Y(I27689),.A(g19070));
  NOT NOT1_7384(.VSS(VSS),.VDD(VDD),.Y(g21130),.A(I27689));
  NOT NOT1_7385(.VSS(VSS),.VDD(VDD),.Y(I27705),.A(g20545));
  NOT NOT1_7386(.VSS(VSS),.VDD(VDD),.Y(g21144),.A(I27705));
  NOT NOT1_7387(.VSS(VSS),.VDD(VDD),.Y(I27727),.A(g19070));
  NOT NOT1_7388(.VSS(VSS),.VDD(VDD),.Y(g21164),.A(I27727));
  NOT NOT1_7389(.VSS(VSS),.VDD(VDD),.Y(I27749),.A(g19954));
  NOT NOT1_7390(.VSS(VSS),.VDD(VDD),.Y(g21184),.A(I27749));
  NOT NOT1_7391(.VSS(VSS),.VDD(VDD),.Y(g21187),.A(g19113));
  NOT NOT1_7392(.VSS(VSS),.VDD(VDD),.Y(I27766),.A(g19984));
  NOT NOT1_7393(.VSS(VSS),.VDD(VDD),.Y(g21199),.A(I27766));
  NOT NOT1_7394(.VSS(VSS),.VDD(VDD),.Y(g21202),.A(g19118));
  NOT NOT1_7395(.VSS(VSS),.VDD(VDD),.Y(I27779),.A(g20022));
  NOT NOT1_7396(.VSS(VSS),.VDD(VDD),.Y(g21214),.A(I27779));
  NOT NOT1_7397(.VSS(VSS),.VDD(VDD),.Y(g21217),.A(g19125));
  NOT NOT1_7398(.VSS(VSS),.VDD(VDD),.Y(I27785),.A(g20064));
  NOT NOT1_7399(.VSS(VSS),.VDD(VDD),.Y(g21222),.A(I27785));
  NOT NOT1_7400(.VSS(VSS),.VDD(VDD),.Y(g21225),.A(g19132));
  NOT NOT1_7401(.VSS(VSS),.VDD(VDD),.Y(g21241),.A(g19945));
  NOT NOT1_7402(.VSS(VSS),.VDD(VDD),.Y(g21249),.A(g19972));
  NOT NOT1_7403(.VSS(VSS),.VDD(VDD),.Y(g21258),.A(g20002));
  NOT NOT1_7404(.VSS(VSS),.VDD(VDD),.Y(g21266),.A(g20040));
  NOT NOT1_7405(.VSS(VSS),.VDD(VDD),.Y(I27822),.A(g19865));
  NOT NOT1_7406(.VSS(VSS),.VDD(VDD),.Y(g21271),.A(I27822));
  NOT NOT1_7407(.VSS(VSS),.VDD(VDD),.Y(I27827),.A(g19896));
  NOT NOT1_7408(.VSS(VSS),.VDD(VDD),.Y(g21278),.A(I27827));
  NOT NOT1_7409(.VSS(VSS),.VDD(VDD),.Y(I27832),.A(g19921));
  NOT NOT1_7410(.VSS(VSS),.VDD(VDD),.Y(g21285),.A(I27832));
  NOT NOT1_7411(.VSS(VSS),.VDD(VDD),.Y(I27838),.A(g19936));
  NOT NOT1_7412(.VSS(VSS),.VDD(VDD),.Y(g21293),.A(I27838));
  NOT NOT1_7413(.VSS(VSS),.VDD(VDD),.Y(I27868),.A(g19144));
  NOT NOT1_7414(.VSS(VSS),.VDD(VDD),.Y(g21327),.A(I27868));
  NOT NOT1_7415(.VSS(VSS),.VDD(VDD),.Y(I27897),.A(g19149));
  NOT NOT1_7416(.VSS(VSS),.VDD(VDD),.Y(g21358),.A(I27897));
  NOT NOT1_7417(.VSS(VSS),.VDD(VDD),.Y(I27900),.A(g19096));
  NOT NOT1_7418(.VSS(VSS),.VDD(VDD),.Y(g21359),.A(I27900));
  NOT NOT1_7419(.VSS(VSS),.VDD(VDD),.Y(I27917),.A(g19153));
  NOT NOT1_7420(.VSS(VSS),.VDD(VDD),.Y(g21376),.A(I27917));
  NOT NOT1_7421(.VSS(VSS),.VDD(VDD),.Y(I27920),.A(g19154));
  NOT NOT1_7422(.VSS(VSS),.VDD(VDD),.Y(g21377),.A(I27920));
  NOT NOT1_7423(.VSS(VSS),.VDD(VDD),.Y(I27927),.A(g19957));
  NOT NOT1_7424(.VSS(VSS),.VDD(VDD),.Y(g21382),.A(I27927));
  NOT NOT1_7425(.VSS(VSS),.VDD(VDD),.Y(I27942),.A(g19157));
  NOT NOT1_7426(.VSS(VSS),.VDD(VDD),.Y(g21399),.A(I27942));
  NOT NOT1_7427(.VSS(VSS),.VDD(VDD),.Y(g21400),.A(g19918));
  NOT NOT1_7428(.VSS(VSS),.VDD(VDD),.Y(I27949),.A(g19957));
  NOT NOT1_7429(.VSS(VSS),.VDD(VDD),.Y(g21404),.A(I27949));
  NOT NOT1_7430(.VSS(VSS),.VDD(VDD),.Y(I27958),.A(g19987));
  NOT NOT1_7431(.VSS(VSS),.VDD(VDD),.Y(g21415),.A(I27958));
  NOT NOT1_7432(.VSS(VSS),.VDD(VDD),.Y(I27969),.A(g19162));
  NOT NOT1_7433(.VSS(VSS),.VDD(VDD),.Y(g21426),.A(I27969));
  NOT NOT1_7434(.VSS(VSS),.VDD(VDD),.Y(I27972),.A(g19163));
  NOT NOT1_7435(.VSS(VSS),.VDD(VDD),.Y(g21427),.A(I27972));
  NOT NOT1_7436(.VSS(VSS),.VDD(VDD),.Y(I27976),.A(g19957));
  NOT NOT1_7437(.VSS(VSS),.VDD(VDD),.Y(g21429),.A(I27976));
  NOT NOT1_7438(.VSS(VSS),.VDD(VDD),.Y(I27984),.A(g19987));
  NOT NOT1_7439(.VSS(VSS),.VDD(VDD),.Y(g21441),.A(I27984));
  NOT NOT1_7440(.VSS(VSS),.VDD(VDD),.Y(I27992),.A(g20025));
  NOT NOT1_7441(.VSS(VSS),.VDD(VDD),.Y(g21449),.A(I27992));
  NOT NOT1_7442(.VSS(VSS),.VDD(VDD),.Y(I28000),.A(g19167));
  NOT NOT1_7443(.VSS(VSS),.VDD(VDD),.Y(g21457),.A(I28000));
  NOT NOT1_7444(.VSS(VSS),.VDD(VDD),.Y(I28003),.A(g19957));
  NOT NOT1_7445(.VSS(VSS),.VDD(VDD),.Y(g21458),.A(I28003));
  NOT NOT1_7446(.VSS(VSS),.VDD(VDD),.Y(g21461),.A(g19957));
  NOT NOT1_7447(.VSS(VSS),.VDD(VDD),.Y(I28009),.A(g20473));
  NOT NOT1_7448(.VSS(VSS),.VDD(VDD),.Y(g21473),.A(I28009));
  NOT NOT1_7449(.VSS(VSS),.VDD(VDD),.Y(I28013),.A(g19987));
  NOT NOT1_7450(.VSS(VSS),.VDD(VDD),.Y(g21477),.A(I28013));
  NOT NOT1_7451(.VSS(VSS),.VDD(VDD),.Y(I28019),.A(g20025));
  NOT NOT1_7452(.VSS(VSS),.VDD(VDD),.Y(g21483),.A(I28019));
  NOT NOT1_7453(.VSS(VSS),.VDD(VDD),.Y(I28027),.A(g20067));
  NOT NOT1_7454(.VSS(VSS),.VDD(VDD),.Y(g21491),.A(I28027));
  NOT NOT1_7455(.VSS(VSS),.VDD(VDD),.Y(I28031),.A(g19172));
  NOT NOT1_7456(.VSS(VSS),.VDD(VDD),.Y(g21495),.A(I28031));
  NOT NOT1_7457(.VSS(VSS),.VDD(VDD),.Y(I28034),.A(g19173));
  NOT NOT1_7458(.VSS(VSS),.VDD(VDD),.Y(g21496),.A(I28034));
  NOT NOT1_7459(.VSS(VSS),.VDD(VDD),.Y(I28038),.A(g19957));
  NOT NOT1_7460(.VSS(VSS),.VDD(VDD),.Y(g21498),.A(I28038));
  NOT NOT1_7461(.VSS(VSS),.VDD(VDD),.Y(I28043),.A(g19987));
  NOT NOT1_7462(.VSS(VSS),.VDD(VDD),.Y(g21505),.A(I28043));
  NOT NOT1_7463(.VSS(VSS),.VDD(VDD),.Y(g21508),.A(g19987));
  NOT NOT1_7464(.VSS(VSS),.VDD(VDD),.Y(I28047),.A(g20481));
  NOT NOT1_7465(.VSS(VSS),.VDD(VDD),.Y(g21514),.A(I28047));
  NOT NOT1_7466(.VSS(VSS),.VDD(VDD),.Y(I28051),.A(g20025));
  NOT NOT1_7467(.VSS(VSS),.VDD(VDD),.Y(g21518),.A(I28051));
  NOT NOT1_7468(.VSS(VSS),.VDD(VDD),.Y(I28057),.A(g20067));
  NOT NOT1_7469(.VSS(VSS),.VDD(VDD),.Y(g21524),.A(I28057));
  NOT NOT1_7470(.VSS(VSS),.VDD(VDD),.Y(I28061),.A(g19178));
  NOT NOT1_7471(.VSS(VSS),.VDD(VDD),.Y(g21528),.A(I28061));
  NOT NOT1_7472(.VSS(VSS),.VDD(VDD),.Y(g21529),.A(g19272));
  NOT NOT1_7473(.VSS(VSS),.VDD(VDD),.Y(I28065),.A(g19957));
  NOT NOT1_7474(.VSS(VSS),.VDD(VDD),.Y(g21530),.A(I28065));
  NOT NOT1_7475(.VSS(VSS),.VDD(VDD),.Y(I28072),.A(g19987));
  NOT NOT1_7476(.VSS(VSS),.VDD(VDD),.Y(g21537),.A(I28072));
  NOT NOT1_7477(.VSS(VSS),.VDD(VDD),.Y(I28076),.A(g20025));
  NOT NOT1_7478(.VSS(VSS),.VDD(VDD),.Y(g21541),.A(I28076));
  NOT NOT1_7479(.VSS(VSS),.VDD(VDD),.Y(g21544),.A(g20025));
  NOT NOT1_7480(.VSS(VSS),.VDD(VDD),.Y(I28080),.A(g20487));
  NOT NOT1_7481(.VSS(VSS),.VDD(VDD),.Y(g21550),.A(I28080));
  NOT NOT1_7482(.VSS(VSS),.VDD(VDD),.Y(I28084),.A(g20067));
  NOT NOT1_7483(.VSS(VSS),.VDD(VDD),.Y(g21554),.A(I28084));
  NOT NOT1_7484(.VSS(VSS),.VDD(VDD),.Y(I28087),.A(g19184));
  NOT NOT1_7485(.VSS(VSS),.VDD(VDD),.Y(g21557),.A(I28087));
  NOT NOT1_7486(.VSS(VSS),.VDD(VDD),.Y(I28090),.A(g20008));
  NOT NOT1_7487(.VSS(VSS),.VDD(VDD),.Y(g21558),.A(I28090));
  NOT NOT1_7488(.VSS(VSS),.VDD(VDD),.Y(I28093),.A(g19957));
  NOT NOT1_7489(.VSS(VSS),.VDD(VDD),.Y(g21561),.A(I28093));
  NOT NOT1_7490(.VSS(VSS),.VDD(VDD),.Y(g21565),.A(g19291));
  NOT NOT1_7491(.VSS(VSS),.VDD(VDD),.Y(I28100),.A(g19987));
  NOT NOT1_7492(.VSS(VSS),.VDD(VDD),.Y(g21566),.A(I28100));
  NOT NOT1_7493(.VSS(VSS),.VDD(VDD),.Y(I28107),.A(g20025));
  NOT NOT1_7494(.VSS(VSS),.VDD(VDD),.Y(g21573),.A(I28107));
  NOT NOT1_7495(.VSS(VSS),.VDD(VDD),.Y(I28111),.A(g20067));
  NOT NOT1_7496(.VSS(VSS),.VDD(VDD),.Y(g21577),.A(I28111));
  NOT NOT1_7497(.VSS(VSS),.VDD(VDD),.Y(g21580),.A(g20067));
  NOT NOT1_7498(.VSS(VSS),.VDD(VDD),.Y(I28115),.A(g20493));
  NOT NOT1_7499(.VSS(VSS),.VDD(VDD),.Y(g21586),.A(I28115));
  NOT NOT1_7500(.VSS(VSS),.VDD(VDD),.Y(I28119),.A(g19957));
  NOT NOT1_7501(.VSS(VSS),.VDD(VDD),.Y(g21590),.A(I28119));
  NOT NOT1_7502(.VSS(VSS),.VDD(VDD),.Y(I28123),.A(g19987));
  NOT NOT1_7503(.VSS(VSS),.VDD(VDD),.Y(g21594),.A(I28123));
  NOT NOT1_7504(.VSS(VSS),.VDD(VDD),.Y(g21598),.A(g19309));
  NOT NOT1_7505(.VSS(VSS),.VDD(VDD),.Y(I28130),.A(g20025));
  NOT NOT1_7506(.VSS(VSS),.VDD(VDD),.Y(g21599),.A(I28130));
  NOT NOT1_7507(.VSS(VSS),.VDD(VDD),.Y(I28137),.A(g20067));
  NOT NOT1_7508(.VSS(VSS),.VDD(VDD),.Y(g21606),.A(I28137));
  NOT NOT1_7509(.VSS(VSS),.VDD(VDD),.Y(I28143),.A(g19957));
  NOT NOT1_7510(.VSS(VSS),.VDD(VDD),.Y(g21612),.A(I28143));
  NOT NOT1_7511(.VSS(VSS),.VDD(VDD),.Y(I28148),.A(g19987));
  NOT NOT1_7512(.VSS(VSS),.VDD(VDD),.Y(g21619),.A(I28148));
  NOT NOT1_7513(.VSS(VSS),.VDD(VDD),.Y(I28152),.A(g20025));
  NOT NOT1_7514(.VSS(VSS),.VDD(VDD),.Y(g21623),.A(I28152));
  NOT NOT1_7515(.VSS(VSS),.VDD(VDD),.Y(g21627),.A(g19330));
  NOT NOT1_7516(.VSS(VSS),.VDD(VDD),.Y(I28159),.A(g20067));
  NOT NOT1_7517(.VSS(VSS),.VDD(VDD),.Y(g21628),.A(I28159));
  NOT NOT1_7518(.VSS(VSS),.VDD(VDD),.Y(I28169),.A(g19987));
  NOT NOT1_7519(.VSS(VSS),.VDD(VDD),.Y(g21640),.A(I28169));
  NOT NOT1_7520(.VSS(VSS),.VDD(VDD),.Y(I28174),.A(g20025));
  NOT NOT1_7521(.VSS(VSS),.VDD(VDD),.Y(g21647),.A(I28174));
  NOT NOT1_7522(.VSS(VSS),.VDD(VDD),.Y(I28178),.A(g20067));
  NOT NOT1_7523(.VSS(VSS),.VDD(VDD),.Y(g21651),.A(I28178));
  NOT NOT1_7524(.VSS(VSS),.VDD(VDD),.Y(I28184),.A(g19103));
  NOT NOT1_7525(.VSS(VSS),.VDD(VDD),.Y(g21655),.A(I28184));
  NOT NOT1_7526(.VSS(VSS),.VDD(VDD),.Y(g21661),.A(g19091));
  NOT NOT1_7527(.VSS(VSS),.VDD(VDD),.Y(I28201),.A(g20025));
  NOT NOT1_7528(.VSS(VSS),.VDD(VDD),.Y(g21671),.A(I28201));
  NOT NOT1_7529(.VSS(VSS),.VDD(VDD),.Y(I28206),.A(g20067));
  NOT NOT1_7530(.VSS(VSS),.VDD(VDD),.Y(g21678),.A(I28206));
  NOT NOT1_7531(.VSS(VSS),.VDD(VDD),.Y(I28210),.A(g20537));
  NOT NOT1_7532(.VSS(VSS),.VDD(VDD),.Y(g21682),.A(I28210));
  NOT NOT1_7533(.VSS(VSS),.VDD(VDD),.Y(g21690),.A(g19098));
  NOT NOT1_7534(.VSS(VSS),.VDD(VDD),.Y(I28229),.A(g20067));
  NOT NOT1_7535(.VSS(VSS),.VDD(VDD),.Y(g21700),.A(I28229));
  NOT NOT1_7536(.VSS(VSS),.VDD(VDD),.Y(I28235),.A(g20153));
  NOT NOT1_7537(.VSS(VSS),.VDD(VDD),.Y(g21708),.A(I28235));
  NOT NOT1_7538(.VSS(VSS),.VDD(VDD),.Y(g21716),.A(g19894));
  NOT NOT1_7539(.VSS(VSS),.VDD(VDD),.Y(g21726),.A(g19105));
  NOT NOT1_7540(.VSS(VSS),.VDD(VDD),.Y(g21742),.A(g19919));
  NOT NOT1_7541(.VSS(VSS),.VDD(VDD),.Y(g21752),.A(g19110));
  NOT NOT1_7542(.VSS(VSS),.VDD(VDD),.Y(g21766),.A(g19934));
  NOT NOT1_7543(.VSS(VSS),.VDD(VDD),.Y(g21782),.A(g19951));
  NOT NOT1_7544(.VSS(VSS),.VDD(VDD),.Y(I28314),.A(g19152));
  NOT NOT1_7545(.VSS(VSS),.VDD(VDD),.Y(g21795),.A(I28314));
  NOT NOT1_7546(.VSS(VSS),.VDD(VDD),.Y(I28357),.A(g20497));
  NOT NOT1_7547(.VSS(VSS),.VDD(VDD),.Y(g21824),.A(I28357));
  NOT NOT1_7548(.VSS(VSS),.VDD(VDD),.Y(I28360),.A(g20163));
  NOT NOT1_7549(.VSS(VSS),.VDD(VDD),.Y(g21825),.A(I28360));
  NOT NOT1_7550(.VSS(VSS),.VDD(VDD),.Y(g21861),.A(g19657));
  NOT NOT1_7551(.VSS(VSS),.VDD(VDD),.Y(g21867),.A(g19705));
  NOT NOT1_7552(.VSS(VSS),.VDD(VDD),.Y(g21872),.A(g19749));
  NOT NOT1_7553(.VSS(VSS),.VDD(VDD),.Y(g21876),.A(g19792));
  NOT NOT1_7554(.VSS(VSS),.VDD(VDD),.Y(g21883),.A(g19890));
  NOT NOT1_7555(.VSS(VSS),.VDD(VDD),.Y(g21886),.A(g19915));
  NOT NOT1_7556(.VSS(VSS),.VDD(VDD),.Y(g21895),.A(g19945));
  NOT NOT1_7557(.VSS(VSS),.VDD(VDD),.Y(g21902),.A(g19978));
  NOT NOT1_7558(.VSS(VSS),.VDD(VDD),.Y(g21907),.A(g19972));
  NOT NOT1_7559(.VSS(VSS),.VDD(VDD),.Y(I28432),.A(g19335));
  NOT NOT1_7560(.VSS(VSS),.VDD(VDD),.Y(g21914),.A(I28432));
  NOT NOT1_7561(.VSS(VSS),.VDD(VDD),.Y(I28435),.A(g19358));
  NOT NOT1_7562(.VSS(VSS),.VDD(VDD),.Y(g21917),.A(I28435));
  NOT NOT1_7563(.VSS(VSS),.VDD(VDD),.Y(g21921),.A(g20002));
  NOT NOT1_7564(.VSS(VSS),.VDD(VDD),.Y(g21927),.A(g20045));
  NOT NOT1_7565(.VSS(VSS),.VDD(VDD),.Y(I28443),.A(g19358));
  NOT NOT1_7566(.VSS(VSS),.VDD(VDD),.Y(g21928),.A(I28443));
  NOT NOT1_7567(.VSS(VSS),.VDD(VDD),.Y(I28447),.A(g19369));
  NOT NOT1_7568(.VSS(VSS),.VDD(VDD),.Y(g21932),.A(I28447));
  NOT NOT1_7569(.VSS(VSS),.VDD(VDD),.Y(I28450),.A(g19390));
  NOT NOT1_7570(.VSS(VSS),.VDD(VDD),.Y(g21935),.A(I28450));
  NOT NOT1_7571(.VSS(VSS),.VDD(VDD),.Y(g21939),.A(g20040));
  NOT NOT1_7572(.VSS(VSS),.VDD(VDD),.Y(I28455),.A(g20943));
  NOT NOT1_7573(.VSS(VSS),.VDD(VDD),.Y(g21943),.A(I28455));
  NOT NOT1_7574(.VSS(VSS),.VDD(VDD),.Y(I28458),.A(g20971));
  NOT NOT1_7575(.VSS(VSS),.VDD(VDD),.Y(g21944),.A(I28458));
  NOT NOT1_7576(.VSS(VSS),.VDD(VDD),.Y(I28461),.A(g20998));
  NOT NOT1_7577(.VSS(VSS),.VDD(VDD),.Y(g21945),.A(I28461));
  NOT NOT1_7578(.VSS(VSS),.VDD(VDD),.Y(I28464),.A(g21024));
  NOT NOT1_7579(.VSS(VSS),.VDD(VDD),.Y(g21946),.A(I28464));
  NOT NOT1_7580(.VSS(VSS),.VDD(VDD),.Y(I28467),.A(g20942));
  NOT NOT1_7581(.VSS(VSS),.VDD(VDD),.Y(g21947),.A(I28467));
  NOT NOT1_7582(.VSS(VSS),.VDD(VDD),.Y(I28470),.A(g20984));
  NOT NOT1_7583(.VSS(VSS),.VDD(VDD),.Y(g21948),.A(I28470));
  NOT NOT1_7584(.VSS(VSS),.VDD(VDD),.Y(I28473),.A(g21030));
  NOT NOT1_7585(.VSS(VSS),.VDD(VDD),.Y(g21949),.A(I28473));
  NOT NOT1_7586(.VSS(VSS),.VDD(VDD),.Y(I28476),.A(g21064));
  NOT NOT1_7587(.VSS(VSS),.VDD(VDD),.Y(g21950),.A(I28476));
  NOT NOT1_7588(.VSS(VSS),.VDD(VDD),.Y(I28479),.A(g21795));
  NOT NOT1_7589(.VSS(VSS),.VDD(VDD),.Y(g21951),.A(I28479));
  NOT NOT1_7590(.VSS(VSS),.VDD(VDD),.Y(I28482),.A(g21376));
  NOT NOT1_7591(.VSS(VSS),.VDD(VDD),.Y(g21952),.A(I28482));
  NOT NOT1_7592(.VSS(VSS),.VDD(VDD),.Y(I28485),.A(g21426));
  NOT NOT1_7593(.VSS(VSS),.VDD(VDD),.Y(g21953),.A(I28485));
  NOT NOT1_7594(.VSS(VSS),.VDD(VDD),.Y(I28488),.A(g21495));
  NOT NOT1_7595(.VSS(VSS),.VDD(VDD),.Y(g21954),.A(I28488));
  NOT NOT1_7596(.VSS(VSS),.VDD(VDD),.Y(I28491),.A(g21327));
  NOT NOT1_7597(.VSS(VSS),.VDD(VDD),.Y(g21955),.A(I28491));
  NOT NOT1_7598(.VSS(VSS),.VDD(VDD),.Y(I28494),.A(g21358));
  NOT NOT1_7599(.VSS(VSS),.VDD(VDD),.Y(g21956),.A(I28494));
  NOT NOT1_7600(.VSS(VSS),.VDD(VDD),.Y(I28497),.A(g21399));
  NOT NOT1_7601(.VSS(VSS),.VDD(VDD),.Y(g21957),.A(I28497));
  NOT NOT1_7602(.VSS(VSS),.VDD(VDD),.Y(I28500),.A(g21457));
  NOT NOT1_7603(.VSS(VSS),.VDD(VDD),.Y(g21958),.A(I28500));
  NOT NOT1_7604(.VSS(VSS),.VDD(VDD),.Y(I28503),.A(g21528));
  NOT NOT1_7605(.VSS(VSS),.VDD(VDD),.Y(g21959),.A(I28503));
  NOT NOT1_7606(.VSS(VSS),.VDD(VDD),.Y(I28506),.A(g21377));
  NOT NOT1_7607(.VSS(VSS),.VDD(VDD),.Y(g21960),.A(I28506));
  NOT NOT1_7608(.VSS(VSS),.VDD(VDD),.Y(I28509),.A(g21427));
  NOT NOT1_7609(.VSS(VSS),.VDD(VDD),.Y(g21961),.A(I28509));
  NOT NOT1_7610(.VSS(VSS),.VDD(VDD),.Y(I28512),.A(g21496));
  NOT NOT1_7611(.VSS(VSS),.VDD(VDD),.Y(g21962),.A(I28512));
  NOT NOT1_7612(.VSS(VSS),.VDD(VDD),.Y(I28515),.A(g21557));
  NOT NOT1_7613(.VSS(VSS),.VDD(VDD),.Y(g21963),.A(I28515));
  NOT NOT1_7614(.VSS(VSS),.VDD(VDD),.Y(I28518),.A(g20985));
  NOT NOT1_7615(.VSS(VSS),.VDD(VDD),.Y(g21964),.A(I28518));
  NOT NOT1_7616(.VSS(VSS),.VDD(VDD),.Y(I28521),.A(g21824));
  NOT NOT1_7617(.VSS(VSS),.VDD(VDD),.Y(g21965),.A(I28521));
  NOT NOT1_7618(.VSS(VSS),.VDD(VDD),.Y(I28524),.A(g21359));
  NOT NOT1_7619(.VSS(VSS),.VDD(VDD),.Y(g21966),.A(I28524));
  NOT NOT1_7620(.VSS(VSS),.VDD(VDD),.Y(I28527),.A(g21407));
  NOT NOT1_7621(.VSS(VSS),.VDD(VDD),.Y(g21967),.A(I28527));
  NOT NOT1_7622(.VSS(VSS),.VDD(VDD),.Y(I28541),.A(g21467));
  NOT NOT1_7623(.VSS(VSS),.VDD(VDD),.Y(g21982),.A(I28541));
  NOT NOT1_7624(.VSS(VSS),.VDD(VDD),.Y(I28550),.A(g21432));
  NOT NOT1_7625(.VSS(VSS),.VDD(VDD),.Y(g21995),.A(I28550));
  NOT NOT1_7626(.VSS(VSS),.VDD(VDD),.Y(I28557),.A(g21407));
  NOT NOT1_7627(.VSS(VSS),.VDD(VDD),.Y(g22003),.A(I28557));
  NOT NOT1_7628(.VSS(VSS),.VDD(VDD),.Y(I28564),.A(g21385));
  NOT NOT1_7629(.VSS(VSS),.VDD(VDD),.Y(g22014),.A(I28564));
  NOT NOT1_7630(.VSS(VSS),.VDD(VDD),.Y(I28628),.A(g21842));
  NOT NOT1_7631(.VSS(VSS),.VDD(VDD),.Y(g22082),.A(I28628));
  NOT NOT1_7632(.VSS(VSS),.VDD(VDD),.Y(I28649),.A(g21843));
  NOT NOT1_7633(.VSS(VSS),.VDD(VDD),.Y(g22107),.A(I28649));
  NOT NOT1_7634(.VSS(VSS),.VDD(VDD),.Y(I28671),.A(g21845));
  NOT NOT1_7635(.VSS(VSS),.VDD(VDD),.Y(g22133),.A(I28671));
  NOT NOT1_7636(.VSS(VSS),.VDD(VDD),.Y(I28693),.A(g21847));
  NOT NOT1_7637(.VSS(VSS),.VDD(VDD),.Y(g22156),.A(I28693));
  NOT NOT1_7638(.VSS(VSS),.VDD(VDD),.Y(I28712),.A(g21851));
  NOT NOT1_7639(.VSS(VSS),.VDD(VDD),.Y(g22176),.A(I28712));
  NOT NOT1_7640(.VSS(VSS),.VDD(VDD),.Y(g22212),.A(g21914));
  NOT NOT1_7641(.VSS(VSS),.VDD(VDD),.Y(g22213),.A(g21917));
  NOT NOT1_7642(.VSS(VSS),.VDD(VDD),.Y(g22217),.A(g21928));
  NOT NOT1_7643(.VSS(VSS),.VDD(VDD),.Y(I28781),.A(g21331));
  NOT NOT1_7644(.VSS(VSS),.VDD(VDD),.Y(g22219),.A(I28781));
  NOT NOT1_7645(.VSS(VSS),.VDD(VDD),.Y(g22221),.A(g21932));
  NOT NOT1_7646(.VSS(VSS),.VDD(VDD),.Y(g22222),.A(g21935));
  NOT NOT1_7647(.VSS(VSS),.VDD(VDD),.Y(I28789),.A(g21878));
  NOT NOT1_7648(.VSS(VSS),.VDD(VDD),.Y(g22225),.A(I28789));
  NOT NOT1_7649(.VSS(VSS),.VDD(VDD),.Y(I28792),.A(g21880));
  NOT NOT1_7650(.VSS(VSS),.VDD(VDD),.Y(g22226),.A(I28792));
  NOT NOT1_7651(.VSS(VSS),.VDD(VDD),.Y(g22230),.A(g20634));
  NOT NOT1_7652(.VSS(VSS),.VDD(VDD),.Y(I28800),.A(g21316));
  NOT NOT1_7653(.VSS(VSS),.VDD(VDD),.Y(g22232),.A(I28800));
  NOT NOT1_7654(.VSS(VSS),.VDD(VDD),.Y(g22233),.A(g20637));
  NOT NOT1_7655(.VSS(VSS),.VDD(VDD),.Y(g22236),.A(g20641));
  NOT NOT1_7656(.VSS(VSS),.VDD(VDD),.Y(g22237),.A(g20644));
  NOT NOT1_7657(.VSS(VSS),.VDD(VDD),.Y(g22239),.A(g20649));
  NOT NOT1_7658(.VSS(VSS),.VDD(VDD),.Y(g22240),.A(g20652));
  NOT NOT1_7659(.VSS(VSS),.VDD(VDD),.Y(g22241),.A(g20655));
  NOT NOT1_7660(.VSS(VSS),.VDD(VDD),.Y(I28813),.A(g21502));
  NOT NOT1_7661(.VSS(VSS),.VDD(VDD),.Y(g22243),.A(I28813));
  NOT NOT1_7662(.VSS(VSS),.VDD(VDD),.Y(g22246),.A(g20659));
  NOT NOT1_7663(.VSS(VSS),.VDD(VDD),.Y(g22248),.A(g20662));
  NOT NOT1_7664(.VSS(VSS),.VDD(VDD),.Y(g22251),.A(g20666));
  NOT NOT1_7665(.VSS(VSS),.VDD(VDD),.Y(g22252),.A(g20669));
  NOT NOT1_7666(.VSS(VSS),.VDD(VDD),.Y(I28825),.A(g21882));
  NOT NOT1_7667(.VSS(VSS),.VDD(VDD),.Y(g22253),.A(I28825));
  NOT NOT1_7668(.VSS(VSS),.VDD(VDD),.Y(g22256),.A(g20673));
  NOT NOT1_7669(.VSS(VSS),.VDD(VDD),.Y(g22257),.A(g20676));
  NOT NOT1_7670(.VSS(VSS),.VDD(VDD),.Y(g22258),.A(g20679));
  NOT NOT1_7671(.VSS(VSS),.VDD(VDD),.Y(I28833),.A(g21470));
  NOT NOT1_7672(.VSS(VSS),.VDD(VDD),.Y(g22259),.A(I28833));
  NOT NOT1_7673(.VSS(VSS),.VDD(VDD),.Y(g22260),.A(g20684));
  NOT NOT1_7674(.VSS(VSS),.VDD(VDD),.Y(g22261),.A(g20687));
  NOT NOT1_7675(.VSS(VSS),.VDD(VDD),.Y(g22262),.A(g20690));
  NOT NOT1_7676(.VSS(VSS),.VDD(VDD),.Y(g22266),.A(g20694));
  NOT NOT1_7677(.VSS(VSS),.VDD(VDD),.Y(g22268),.A(g20697));
  NOT NOT1_7678(.VSS(VSS),.VDD(VDD),.Y(g22271),.A(g20704));
  NOT NOT1_7679(.VSS(VSS),.VDD(VDD),.Y(g22274),.A(g20708));
  NOT NOT1_7680(.VSS(VSS),.VDD(VDD),.Y(g22275),.A(g20711));
  NOT NOT1_7681(.VSS(VSS),.VDD(VDD),.Y(g22276),.A(g20714));
  NOT NOT1_7682(.VSS(VSS),.VDD(VDD),.Y(g22277),.A(g20719));
  NOT NOT1_7683(.VSS(VSS),.VDD(VDD),.Y(g22278),.A(g20722));
  NOT NOT1_7684(.VSS(VSS),.VDD(VDD),.Y(g22279),.A(g20725));
  NOT NOT1_7685(.VSS(VSS),.VDD(VDD),.Y(g22283),.A(g20729));
  NOT NOT1_7686(.VSS(VSS),.VDD(VDD),.Y(g22286),.A(g20732));
  NOT NOT1_7687(.VSS(VSS),.VDD(VDD),.Y(g22287),.A(g20735));
  NOT NOT1_7688(.VSS(VSS),.VDD(VDD),.Y(g22290),.A(g20739));
  NOT NOT1_7689(.VSS(VSS),.VDD(VDD),.Y(g22293),.A(g20743));
  NOT NOT1_7690(.VSS(VSS),.VDD(VDD),.Y(g22294),.A(g20746));
  NOT NOT1_7691(.VSS(VSS),.VDD(VDD),.Y(g22295),.A(g20749));
  NOT NOT1_7692(.VSS(VSS),.VDD(VDD),.Y(g22296),.A(g20754));
  NOT NOT1_7693(.VSS(VSS),.VDD(VDD),.Y(g22297),.A(g20757));
  NOT NOT1_7694(.VSS(VSS),.VDD(VDD),.Y(g22298),.A(g20760));
  NOT NOT1_7695(.VSS(VSS),.VDD(VDD),.Y(I28876),.A(g21238));
  NOT NOT1_7696(.VSS(VSS),.VDD(VDD),.Y(g22300),.A(I28876));
  NOT NOT1_7697(.VSS(VSS),.VDD(VDD),.Y(g22303),.A(g20763));
  NOT NOT1_7698(.VSS(VSS),.VDD(VDD),.Y(g22304),.A(g20766));
  NOT NOT1_7699(.VSS(VSS),.VDD(VDD),.Y(g22306),.A(g20769));
  NOT NOT1_7700(.VSS(VSS),.VDD(VDD),.Y(g22307),.A(g20772));
  NOT NOT1_7701(.VSS(VSS),.VDD(VDD),.Y(g22310),.A(g20776));
  NOT NOT1_7702(.VSS(VSS),.VDD(VDD),.Y(g22313),.A(g20780));
  NOT NOT1_7703(.VSS(VSS),.VDD(VDD),.Y(g22314),.A(g20783));
  NOT NOT1_7704(.VSS(VSS),.VDD(VDD),.Y(g22315),.A(g20786));
  NOT NOT1_7705(.VSS(VSS),.VDD(VDD),.Y(g22316),.A(g21149));
  NOT NOT1_7706(.VSS(VSS),.VDD(VDD),.Y(g22318),.A(g20790));
  NOT NOT1_7707(.VSS(VSS),.VDD(VDD),.Y(g22319),.A(g21228));
  NOT NOT1_7708(.VSS(VSS),.VDD(VDD),.Y(I28896),.A(g21246));
  NOT NOT1_7709(.VSS(VSS),.VDD(VDD),.Y(g22328),.A(I28896));
  NOT NOT1_7710(.VSS(VSS),.VDD(VDD),.Y(g22331),.A(g20793));
  NOT NOT1_7711(.VSS(VSS),.VDD(VDD),.Y(g22332),.A(g20796));
  NOT NOT1_7712(.VSS(VSS),.VDD(VDD),.Y(g22334),.A(g20799));
  NOT NOT1_7713(.VSS(VSS),.VDD(VDD),.Y(g22335),.A(g20802));
  NOT NOT1_7714(.VSS(VSS),.VDD(VDD),.Y(g22338),.A(g20806));
  NOT NOT1_7715(.VSS(VSS),.VDD(VDD),.Y(g22341),.A(g21169));
  NOT NOT1_7716(.VSS(VSS),.VDD(VDD),.Y(g22343),.A(g20810));
  NOT NOT1_7717(.VSS(VSS),.VDD(VDD),.Y(g22344),.A(g21233));
  NOT NOT1_7718(.VSS(VSS),.VDD(VDD),.Y(I28913),.A(g21255));
  NOT NOT1_7719(.VSS(VSS),.VDD(VDD),.Y(g22353),.A(I28913));
  NOT NOT1_7720(.VSS(VSS),.VDD(VDD),.Y(g22356),.A(g20813));
  NOT NOT1_7721(.VSS(VSS),.VDD(VDD),.Y(g22357),.A(g20816));
  NOT NOT1_7722(.VSS(VSS),.VDD(VDD),.Y(g22359),.A(g20819));
  NOT NOT1_7723(.VSS(VSS),.VDD(VDD),.Y(g22360),.A(g20822));
  NOT NOT1_7724(.VSS(VSS),.VDD(VDD),.Y(g22364),.A(g21189));
  NOT NOT1_7725(.VSS(VSS),.VDD(VDD),.Y(g22366),.A(g20827));
  NOT NOT1_7726(.VSS(VSS),.VDD(VDD),.Y(g22367),.A(g21242));
  NOT NOT1_7727(.VSS(VSS),.VDD(VDD),.Y(I28928),.A(g21263));
  NOT NOT1_7728(.VSS(VSS),.VDD(VDD),.Y(g22376),.A(I28928));
  NOT NOT1_7729(.VSS(VSS),.VDD(VDD),.Y(g22379),.A(g20830));
  NOT NOT1_7730(.VSS(VSS),.VDD(VDD),.Y(g22380),.A(g20833));
  NOT NOT1_7731(.VSS(VSS),.VDD(VDD),.Y(g22384),.A(g21204));
  NOT NOT1_7732(.VSS(VSS),.VDD(VDD),.Y(g22386),.A(g20837));
  NOT NOT1_7733(.VSS(VSS),.VDD(VDD),.Y(g22387),.A(g21250));
  NOT NOT1_7734(.VSS(VSS),.VDD(VDD),.Y(g22401),.A(g21533));
  NOT NOT1_7735(.VSS(VSS),.VDD(VDD),.Y(g22402),.A(g21569));
  NOT NOT1_7736(.VSS(VSS),.VDD(VDD),.Y(g22403),.A(g21602));
  NOT NOT1_7737(.VSS(VSS),.VDD(VDD),.Y(g22404),.A(g21631));
  NOT NOT1_7738(.VSS(VSS),.VDD(VDD),.Y(I28949),.A(g21685));
  NOT NOT1_7739(.VSS(VSS),.VDD(VDD),.Y(g22405),.A(I28949));
  NOT NOT1_7740(.VSS(VSS),.VDD(VDD),.Y(g22408),.A(g20986));
  NOT NOT1_7741(.VSS(VSS),.VDD(VDD),.Y(I28953),.A(g21659));
  NOT NOT1_7742(.VSS(VSS),.VDD(VDD),.Y(g22409),.A(I28953));
  NOT NOT1_7743(.VSS(VSS),.VDD(VDD),.Y(I28956),.A(g21714));
  NOT NOT1_7744(.VSS(VSS),.VDD(VDD),.Y(g22412),.A(I28956));
  NOT NOT1_7745(.VSS(VSS),.VDD(VDD),.Y(I28959),.A(g21636));
  NOT NOT1_7746(.VSS(VSS),.VDD(VDD),.Y(g22415),.A(I28959));
  NOT NOT1_7747(.VSS(VSS),.VDD(VDD),.Y(I28962),.A(g21721));
  NOT NOT1_7748(.VSS(VSS),.VDD(VDD),.Y(g22418),.A(I28962));
  NOT NOT1_7749(.VSS(VSS),.VDD(VDD),.Y(g22421),.A(g21012));
  NOT NOT1_7750(.VSS(VSS),.VDD(VDD),.Y(I28966),.A(g20633));
  NOT NOT1_7751(.VSS(VSS),.VDD(VDD),.Y(g22422),.A(I28966));
  NOT NOT1_7752(.VSS(VSS),.VDD(VDD),.Y(I28969),.A(g21686));
  NOT NOT1_7753(.VSS(VSS),.VDD(VDD),.Y(g22425),.A(I28969));
  NOT NOT1_7754(.VSS(VSS),.VDD(VDD),.Y(I28972),.A(g21736));
  NOT NOT1_7755(.VSS(VSS),.VDD(VDD),.Y(g22428),.A(I28972));
  NOT NOT1_7756(.VSS(VSS),.VDD(VDD),.Y(I28975),.A(g21688));
  NOT NOT1_7757(.VSS(VSS),.VDD(VDD),.Y(g22431),.A(I28975));
  NOT NOT1_7758(.VSS(VSS),.VDD(VDD),.Y(I28978),.A(g21740));
  NOT NOT1_7759(.VSS(VSS),.VDD(VDD),.Y(g22434),.A(I28978));
  NOT NOT1_7760(.VSS(VSS),.VDD(VDD),.Y(I28981),.A(g21667));
  NOT NOT1_7761(.VSS(VSS),.VDD(VDD),.Y(g22437),.A(I28981));
  NOT NOT1_7762(.VSS(VSS),.VDD(VDD),.Y(I28984),.A(g21747));
  NOT NOT1_7763(.VSS(VSS),.VDD(VDD),.Y(g22440),.A(I28984));
  NOT NOT1_7764(.VSS(VSS),.VDD(VDD),.Y(g22443),.A(g21036));
  NOT NOT1_7765(.VSS(VSS),.VDD(VDD),.Y(I28988),.A(g20874));
  NOT NOT1_7766(.VSS(VSS),.VDD(VDD),.Y(g22444),.A(I28988));
  NOT NOT1_7767(.VSS(VSS),.VDD(VDD),.Y(I28991),.A(g20648));
  NOT NOT1_7768(.VSS(VSS),.VDD(VDD),.Y(g22445),.A(I28991));
  NOT NOT1_7769(.VSS(VSS),.VDD(VDD),.Y(I28994),.A(g21715));
  NOT NOT1_7770(.VSS(VSS),.VDD(VDD),.Y(g22448),.A(I28994));
  NOT NOT1_7771(.VSS(VSS),.VDD(VDD),.Y(I28997),.A(g21759));
  NOT NOT1_7772(.VSS(VSS),.VDD(VDD),.Y(g22451),.A(I28997));
  NOT NOT1_7773(.VSS(VSS),.VDD(VDD),.Y(I29001),.A(g20658));
  NOT NOT1_7774(.VSS(VSS),.VDD(VDD),.Y(g22455),.A(I29001));
  NOT NOT1_7775(.VSS(VSS),.VDD(VDD),.Y(I29004),.A(g21722));
  NOT NOT1_7776(.VSS(VSS),.VDD(VDD),.Y(g22458),.A(I29004));
  NOT NOT1_7777(.VSS(VSS),.VDD(VDD),.Y(I29007),.A(g21760));
  NOT NOT1_7778(.VSS(VSS),.VDD(VDD),.Y(g22461),.A(I29007));
  NOT NOT1_7779(.VSS(VSS),.VDD(VDD),.Y(I29010),.A(g21724));
  NOT NOT1_7780(.VSS(VSS),.VDD(VDD),.Y(g22464),.A(I29010));
  NOT NOT1_7781(.VSS(VSS),.VDD(VDD),.Y(I29013),.A(g21764));
  NOT NOT1_7782(.VSS(VSS),.VDD(VDD),.Y(g22467),.A(I29013));
  NOT NOT1_7783(.VSS(VSS),.VDD(VDD),.Y(I29016),.A(g21696));
  NOT NOT1_7784(.VSS(VSS),.VDD(VDD),.Y(g22470),.A(I29016));
  NOT NOT1_7785(.VSS(VSS),.VDD(VDD),.Y(I29019),.A(g21771));
  NOT NOT1_7786(.VSS(VSS),.VDD(VDD),.Y(g22473),.A(I29019));
  NOT NOT1_7787(.VSS(VSS),.VDD(VDD),.Y(g22476),.A(g21057));
  NOT NOT1_7788(.VSS(VSS),.VDD(VDD),.Y(I29023),.A(g20672));
  NOT NOT1_7789(.VSS(VSS),.VDD(VDD),.Y(g22477),.A(I29023));
  NOT NOT1_7790(.VSS(VSS),.VDD(VDD),.Y(I29026),.A(g21737));
  NOT NOT1_7791(.VSS(VSS),.VDD(VDD),.Y(g22480),.A(I29026));
  NOT NOT1_7792(.VSS(VSS),.VDD(VDD),.Y(I29030),.A(g20683));
  NOT NOT1_7793(.VSS(VSS),.VDD(VDD),.Y(g22484),.A(I29030));
  NOT NOT1_7794(.VSS(VSS),.VDD(VDD),.Y(I29033),.A(g21741));
  NOT NOT1_7795(.VSS(VSS),.VDD(VDD),.Y(g22487),.A(I29033));
  NOT NOT1_7796(.VSS(VSS),.VDD(VDD),.Y(I29036),.A(g21775));
  NOT NOT1_7797(.VSS(VSS),.VDD(VDD),.Y(g22490),.A(I29036));
  NOT NOT1_7798(.VSS(VSS),.VDD(VDD),.Y(I29040),.A(g20693));
  NOT NOT1_7799(.VSS(VSS),.VDD(VDD),.Y(g22494),.A(I29040));
  NOT NOT1_7800(.VSS(VSS),.VDD(VDD),.Y(I29043),.A(g21748));
  NOT NOT1_7801(.VSS(VSS),.VDD(VDD),.Y(g22497),.A(I29043));
  NOT NOT1_7802(.VSS(VSS),.VDD(VDD),.Y(I29046),.A(g21776));
  NOT NOT1_7803(.VSS(VSS),.VDD(VDD),.Y(g22500),.A(I29046));
  NOT NOT1_7804(.VSS(VSS),.VDD(VDD),.Y(I29049),.A(g21750));
  NOT NOT1_7805(.VSS(VSS),.VDD(VDD),.Y(g22503),.A(I29049));
  NOT NOT1_7806(.VSS(VSS),.VDD(VDD),.Y(I29052),.A(g21780));
  NOT NOT1_7807(.VSS(VSS),.VDD(VDD),.Y(g22506),.A(I29052));
  NOT NOT1_7808(.VSS(VSS),.VDD(VDD),.Y(I29055),.A(g21732));
  NOT NOT1_7809(.VSS(VSS),.VDD(VDD),.Y(g22509),.A(I29055));
  NOT NOT1_7810(.VSS(VSS),.VDD(VDD),.Y(I29058),.A(g20703));
  NOT NOT1_7811(.VSS(VSS),.VDD(VDD),.Y(g22512),.A(I29058));
  NOT NOT1_7812(.VSS(VSS),.VDD(VDD),.Y(I29064),.A(g20875));
  NOT NOT1_7813(.VSS(VSS),.VDD(VDD),.Y(g22518),.A(I29064));
  NOT NOT1_7814(.VSS(VSS),.VDD(VDD),.Y(I29067),.A(g20876));
  NOT NOT1_7815(.VSS(VSS),.VDD(VDD),.Y(g22519),.A(I29067));
  NOT NOT1_7816(.VSS(VSS),.VDD(VDD),.Y(I29070),.A(g20707));
  NOT NOT1_7817(.VSS(VSS),.VDD(VDD),.Y(g22520),.A(I29070));
  NOT NOT1_7818(.VSS(VSS),.VDD(VDD),.Y(I29073),.A(g21761));
  NOT NOT1_7819(.VSS(VSS),.VDD(VDD),.Y(g22523),.A(I29073));
  NOT NOT1_7820(.VSS(VSS),.VDD(VDD),.Y(I29077),.A(g20718));
  NOT NOT1_7821(.VSS(VSS),.VDD(VDD),.Y(g22527),.A(I29077));
  NOT NOT1_7822(.VSS(VSS),.VDD(VDD),.Y(I29080),.A(g21765));
  NOT NOT1_7823(.VSS(VSS),.VDD(VDD),.Y(g22530),.A(I29080));
  NOT NOT1_7824(.VSS(VSS),.VDD(VDD),.Y(I29083),.A(g21790));
  NOT NOT1_7825(.VSS(VSS),.VDD(VDD),.Y(g22533),.A(I29083));
  NOT NOT1_7826(.VSS(VSS),.VDD(VDD),.Y(I29087),.A(g20728));
  NOT NOT1_7827(.VSS(VSS),.VDD(VDD),.Y(g22537),.A(I29087));
  NOT NOT1_7828(.VSS(VSS),.VDD(VDD),.Y(I29090),.A(g21772));
  NOT NOT1_7829(.VSS(VSS),.VDD(VDD),.Y(g22540),.A(I29090));
  NOT NOT1_7830(.VSS(VSS),.VDD(VDD),.Y(I29093),.A(g21791));
  NOT NOT1_7831(.VSS(VSS),.VDD(VDD),.Y(g22543),.A(I29093));
  NOT NOT1_7832(.VSS(VSS),.VDD(VDD),.Y(g22547),.A(g21087));
  NOT NOT1_7833(.VSS(VSS),.VDD(VDD),.Y(I29098),.A(g20879));
  NOT NOT1_7834(.VSS(VSS),.VDD(VDD),.Y(g22548),.A(I29098));
  NOT NOT1_7835(.VSS(VSS),.VDD(VDD),.Y(I29101),.A(g20880));
  NOT NOT1_7836(.VSS(VSS),.VDD(VDD),.Y(g22549),.A(I29101));
  NOT NOT1_7837(.VSS(VSS),.VDD(VDD),.Y(I29104),.A(g20881));
  NOT NOT1_7838(.VSS(VSS),.VDD(VDD),.Y(g22550),.A(I29104));
  NOT NOT1_7839(.VSS(VSS),.VDD(VDD),.Y(I29107),.A(g21435));
  NOT NOT1_7840(.VSS(VSS),.VDD(VDD),.Y(g22551),.A(I29107));
  NOT NOT1_7841(.VSS(VSS),.VDD(VDD),.Y(I29110),.A(g20738));
  NOT NOT1_7842(.VSS(VSS),.VDD(VDD),.Y(g22552),.A(I29110));
  NOT NOT1_7843(.VSS(VSS),.VDD(VDD),.Y(I29116),.A(g20882));
  NOT NOT1_7844(.VSS(VSS),.VDD(VDD),.Y(g22558),.A(I29116));
  NOT NOT1_7845(.VSS(VSS),.VDD(VDD),.Y(I29119),.A(g20883));
  NOT NOT1_7846(.VSS(VSS),.VDD(VDD),.Y(g22559),.A(I29119));
  NOT NOT1_7847(.VSS(VSS),.VDD(VDD),.Y(I29122),.A(g20742));
  NOT NOT1_7848(.VSS(VSS),.VDD(VDD),.Y(g22560),.A(I29122));
  NOT NOT1_7849(.VSS(VSS),.VDD(VDD),.Y(I29125),.A(g21777));
  NOT NOT1_7850(.VSS(VSS),.VDD(VDD),.Y(g22563),.A(I29125));
  NOT NOT1_7851(.VSS(VSS),.VDD(VDD),.Y(I29129),.A(g20753));
  NOT NOT1_7852(.VSS(VSS),.VDD(VDD),.Y(g22567),.A(I29129));
  NOT NOT1_7853(.VSS(VSS),.VDD(VDD),.Y(I29132),.A(g21781));
  NOT NOT1_7854(.VSS(VSS),.VDD(VDD),.Y(g22570),.A(I29132));
  NOT NOT1_7855(.VSS(VSS),.VDD(VDD),.Y(I29135),.A(g21804));
  NOT NOT1_7856(.VSS(VSS),.VDD(VDD),.Y(g22573),.A(I29135));
  NOT NOT1_7857(.VSS(VSS),.VDD(VDD),.Y(I29142),.A(g20682));
  NOT NOT1_7858(.VSS(VSS),.VDD(VDD),.Y(g22582),.A(I29142));
  NOT NOT1_7859(.VSS(VSS),.VDD(VDD),.Y(I29145),.A(g20891));
  NOT NOT1_7860(.VSS(VSS),.VDD(VDD),.Y(g22583),.A(I29145));
  NOT NOT1_7861(.VSS(VSS),.VDD(VDD),.Y(I29148),.A(g20892));
  NOT NOT1_7862(.VSS(VSS),.VDD(VDD),.Y(g22584),.A(I29148));
  NOT NOT1_7863(.VSS(VSS),.VDD(VDD),.Y(I29151),.A(g20893));
  NOT NOT1_7864(.VSS(VSS),.VDD(VDD),.Y(g22585),.A(I29151));
  NOT NOT1_7865(.VSS(VSS),.VDD(VDD),.Y(I29154),.A(g20894));
  NOT NOT1_7866(.VSS(VSS),.VDD(VDD),.Y(g22586),.A(I29154));
  NOT NOT1_7867(.VSS(VSS),.VDD(VDD),.Y(g22588),.A(g21099));
  NOT NOT1_7868(.VSS(VSS),.VDD(VDD),.Y(I29159),.A(g20896));
  NOT NOT1_7869(.VSS(VSS),.VDD(VDD),.Y(g22589),.A(I29159));
  NOT NOT1_7870(.VSS(VSS),.VDD(VDD),.Y(I29162),.A(g20897));
  NOT NOT1_7871(.VSS(VSS),.VDD(VDD),.Y(g22590),.A(I29162));
  NOT NOT1_7872(.VSS(VSS),.VDD(VDD),.Y(I29165),.A(g20898));
  NOT NOT1_7873(.VSS(VSS),.VDD(VDD),.Y(g22591),.A(I29165));
  NOT NOT1_7874(.VSS(VSS),.VDD(VDD),.Y(I29168),.A(g20775));
  NOT NOT1_7875(.VSS(VSS),.VDD(VDD),.Y(g22592),.A(I29168));
  NOT NOT1_7876(.VSS(VSS),.VDD(VDD),.Y(I29174),.A(g20899));
  NOT NOT1_7877(.VSS(VSS),.VDD(VDD),.Y(g22598),.A(I29174));
  NOT NOT1_7878(.VSS(VSS),.VDD(VDD),.Y(I29177),.A(g20900));
  NOT NOT1_7879(.VSS(VSS),.VDD(VDD),.Y(g22599),.A(I29177));
  NOT NOT1_7880(.VSS(VSS),.VDD(VDD),.Y(I29180),.A(g20779));
  NOT NOT1_7881(.VSS(VSS),.VDD(VDD),.Y(g22600),.A(I29180));
  NOT NOT1_7882(.VSS(VSS),.VDD(VDD),.Y(I29183),.A(g21792));
  NOT NOT1_7883(.VSS(VSS),.VDD(VDD),.Y(g22603),.A(I29183));
  NOT NOT1_7884(.VSS(VSS),.VDD(VDD),.Y(g22609),.A(g21108));
  NOT NOT1_7885(.VSS(VSS),.VDD(VDD),.Y(I29191),.A(g20901));
  NOT NOT1_7886(.VSS(VSS),.VDD(VDD),.Y(g22611),.A(I29191));
  NOT NOT1_7887(.VSS(VSS),.VDD(VDD),.Y(I29194),.A(g20902));
  NOT NOT1_7888(.VSS(VSS),.VDD(VDD),.Y(g22612),.A(I29194));
  NOT NOT1_7889(.VSS(VSS),.VDD(VDD),.Y(I29197),.A(g20903));
  NOT NOT1_7890(.VSS(VSS),.VDD(VDD),.Y(g22613),.A(I29197));
  NOT NOT1_7891(.VSS(VSS),.VDD(VDD),.Y(I29203),.A(g20717));
  NOT NOT1_7892(.VSS(VSS),.VDD(VDD),.Y(g22619),.A(I29203));
  NOT NOT1_7893(.VSS(VSS),.VDD(VDD),.Y(I29206),.A(g20910));
  NOT NOT1_7894(.VSS(VSS),.VDD(VDD),.Y(g22620),.A(I29206));
  NOT NOT1_7895(.VSS(VSS),.VDD(VDD),.Y(I29209),.A(g20911));
  NOT NOT1_7896(.VSS(VSS),.VDD(VDD),.Y(g22621),.A(I29209));
  NOT NOT1_7897(.VSS(VSS),.VDD(VDD),.Y(I29212),.A(g20912));
  NOT NOT1_7898(.VSS(VSS),.VDD(VDD),.Y(g22622),.A(I29212));
  NOT NOT1_7899(.VSS(VSS),.VDD(VDD),.Y(I29215),.A(g20913));
  NOT NOT1_7900(.VSS(VSS),.VDD(VDD),.Y(g22623),.A(I29215));
  NOT NOT1_7901(.VSS(VSS),.VDD(VDD),.Y(g22625),.A(g21113));
  NOT NOT1_7902(.VSS(VSS),.VDD(VDD),.Y(I29220),.A(g20915));
  NOT NOT1_7903(.VSS(VSS),.VDD(VDD),.Y(g22626),.A(I29220));
  NOT NOT1_7904(.VSS(VSS),.VDD(VDD),.Y(I29223),.A(g20916));
  NOT NOT1_7905(.VSS(VSS),.VDD(VDD),.Y(g22627),.A(I29223));
  NOT NOT1_7906(.VSS(VSS),.VDD(VDD),.Y(I29226),.A(g20917));
  NOT NOT1_7907(.VSS(VSS),.VDD(VDD),.Y(g22628),.A(I29226));
  NOT NOT1_7908(.VSS(VSS),.VDD(VDD),.Y(I29229),.A(g20805));
  NOT NOT1_7909(.VSS(VSS),.VDD(VDD),.Y(g22629),.A(I29229));
  NOT NOT1_7910(.VSS(VSS),.VDD(VDD),.Y(I29235),.A(g20918));
  NOT NOT1_7911(.VSS(VSS),.VDD(VDD),.Y(g22635),.A(I29235));
  NOT NOT1_7912(.VSS(VSS),.VDD(VDD),.Y(I29238),.A(g20919));
  NOT NOT1_7913(.VSS(VSS),.VDD(VDD),.Y(g22636),.A(I29238));
  NOT NOT1_7914(.VSS(VSS),.VDD(VDD),.Y(I29243),.A(g20921));
  NOT NOT1_7915(.VSS(VSS),.VDD(VDD),.Y(g22639),.A(I29243));
  NOT NOT1_7916(.VSS(VSS),.VDD(VDD),.Y(I29246),.A(g20922));
  NOT NOT1_7917(.VSS(VSS),.VDD(VDD),.Y(g22640),.A(I29246));
  NOT NOT1_7918(.VSS(VSS),.VDD(VDD),.Y(I29249),.A(g20923));
  NOT NOT1_7919(.VSS(VSS),.VDD(VDD),.Y(g22641),.A(I29249));
  NOT NOT1_7920(.VSS(VSS),.VDD(VDD),.Y(I29252),.A(g20924));
  NOT NOT1_7921(.VSS(VSS),.VDD(VDD),.Y(g22642),.A(I29252));
  NOT NOT1_7922(.VSS(VSS),.VDD(VDD),.Y(g22645),.A(g21125));
  NOT NOT1_7923(.VSS(VSS),.VDD(VDD),.Y(I29259),.A(g20925));
  NOT NOT1_7924(.VSS(VSS),.VDD(VDD),.Y(g22647),.A(I29259));
  NOT NOT1_7925(.VSS(VSS),.VDD(VDD),.Y(I29262),.A(g20926));
  NOT NOT1_7926(.VSS(VSS),.VDD(VDD),.Y(g22648),.A(I29262));
  NOT NOT1_7927(.VSS(VSS),.VDD(VDD),.Y(I29265),.A(g20927));
  NOT NOT1_7928(.VSS(VSS),.VDD(VDD),.Y(g22649),.A(I29265));
  NOT NOT1_7929(.VSS(VSS),.VDD(VDD),.Y(I29271),.A(g20752));
  NOT NOT1_7930(.VSS(VSS),.VDD(VDD),.Y(g22655),.A(I29271));
  NOT NOT1_7931(.VSS(VSS),.VDD(VDD),.Y(I29274),.A(g20934));
  NOT NOT1_7932(.VSS(VSS),.VDD(VDD),.Y(g22656),.A(I29274));
  NOT NOT1_7933(.VSS(VSS),.VDD(VDD),.Y(I29277),.A(g20935));
  NOT NOT1_7934(.VSS(VSS),.VDD(VDD),.Y(g22657),.A(I29277));
  NOT NOT1_7935(.VSS(VSS),.VDD(VDD),.Y(I29280),.A(g20936));
  NOT NOT1_7936(.VSS(VSS),.VDD(VDD),.Y(g22658),.A(I29280));
  NOT NOT1_7937(.VSS(VSS),.VDD(VDD),.Y(I29283),.A(g20937));
  NOT NOT1_7938(.VSS(VSS),.VDD(VDD),.Y(g22659),.A(I29283));
  NOT NOT1_7939(.VSS(VSS),.VDD(VDD),.Y(g22661),.A(g21130));
  NOT NOT1_7940(.VSS(VSS),.VDD(VDD),.Y(I29288),.A(g20939));
  NOT NOT1_7941(.VSS(VSS),.VDD(VDD),.Y(g22662),.A(I29288));
  NOT NOT1_7942(.VSS(VSS),.VDD(VDD),.Y(I29291),.A(g20940));
  NOT NOT1_7943(.VSS(VSS),.VDD(VDD),.Y(g22663),.A(I29291));
  NOT NOT1_7944(.VSS(VSS),.VDD(VDD),.Y(I29294),.A(g20941));
  NOT NOT1_7945(.VSS(VSS),.VDD(VDD),.Y(g22664),.A(I29294));
  NOT NOT1_7946(.VSS(VSS),.VDD(VDD),.Y(I29301),.A(g20944));
  NOT NOT1_7947(.VSS(VSS),.VDD(VDD),.Y(g22669),.A(I29301));
  NOT NOT1_7948(.VSS(VSS),.VDD(VDD),.Y(I29304),.A(g20945));
  NOT NOT1_7949(.VSS(VSS),.VDD(VDD),.Y(g22670),.A(I29304));
  NOT NOT1_7950(.VSS(VSS),.VDD(VDD),.Y(I29307),.A(g20946));
  NOT NOT1_7951(.VSS(VSS),.VDD(VDD),.Y(g22671),.A(I29307));
  NOT NOT1_7952(.VSS(VSS),.VDD(VDD),.Y(I29310),.A(g20947));
  NOT NOT1_7953(.VSS(VSS),.VDD(VDD),.Y(g22672),.A(I29310));
  NOT NOT1_7954(.VSS(VSS),.VDD(VDD),.Y(I29313),.A(g20948));
  NOT NOT1_7955(.VSS(VSS),.VDD(VDD),.Y(g22673),.A(I29313));
  NOT NOT1_7956(.VSS(VSS),.VDD(VDD),.Y(I29317),.A(g20949));
  NOT NOT1_7957(.VSS(VSS),.VDD(VDD),.Y(g22675),.A(I29317));
  NOT NOT1_7958(.VSS(VSS),.VDD(VDD),.Y(I29320),.A(g20950));
  NOT NOT1_7959(.VSS(VSS),.VDD(VDD),.Y(g22676),.A(I29320));
  NOT NOT1_7960(.VSS(VSS),.VDD(VDD),.Y(I29323),.A(g20951));
  NOT NOT1_7961(.VSS(VSS),.VDD(VDD),.Y(g22677),.A(I29323));
  NOT NOT1_7962(.VSS(VSS),.VDD(VDD),.Y(I29326),.A(g20952));
  NOT NOT1_7963(.VSS(VSS),.VDD(VDD),.Y(g22678),.A(I29326));
  NOT NOT1_7964(.VSS(VSS),.VDD(VDD),.Y(g22681),.A(g21144));
  NOT NOT1_7965(.VSS(VSS),.VDD(VDD),.Y(I29333),.A(g20953));
  NOT NOT1_7966(.VSS(VSS),.VDD(VDD),.Y(g22683),.A(I29333));
  NOT NOT1_7967(.VSS(VSS),.VDD(VDD),.Y(I29336),.A(g20954));
  NOT NOT1_7968(.VSS(VSS),.VDD(VDD),.Y(g22684),.A(I29336));
  NOT NOT1_7969(.VSS(VSS),.VDD(VDD),.Y(I29339),.A(g20955));
  NOT NOT1_7970(.VSS(VSS),.VDD(VDD),.Y(g22685),.A(I29339));
  NOT NOT1_7971(.VSS(VSS),.VDD(VDD),.Y(I29345),.A(g20789));
  NOT NOT1_7972(.VSS(VSS),.VDD(VDD),.Y(g22691),.A(I29345));
  NOT NOT1_7973(.VSS(VSS),.VDD(VDD),.Y(I29348),.A(g20962));
  NOT NOT1_7974(.VSS(VSS),.VDD(VDD),.Y(g22692),.A(I29348));
  NOT NOT1_7975(.VSS(VSS),.VDD(VDD),.Y(I29351),.A(g20963));
  NOT NOT1_7976(.VSS(VSS),.VDD(VDD),.Y(g22693),.A(I29351));
  NOT NOT1_7977(.VSS(VSS),.VDD(VDD),.Y(I29354),.A(g20964));
  NOT NOT1_7978(.VSS(VSS),.VDD(VDD),.Y(g22694),.A(I29354));
  NOT NOT1_7979(.VSS(VSS),.VDD(VDD),.Y(I29357),.A(g20965));
  NOT NOT1_7980(.VSS(VSS),.VDD(VDD),.Y(g22695),.A(I29357));
  NOT NOT1_7981(.VSS(VSS),.VDD(VDD),.Y(I29360),.A(g21796));
  NOT NOT1_7982(.VSS(VSS),.VDD(VDD),.Y(g22696),.A(I29360));
  NOT NOT1_7983(.VSS(VSS),.VDD(VDD),.Y(I29366),.A(g20966));
  NOT NOT1_7984(.VSS(VSS),.VDD(VDD),.Y(g22702),.A(I29366));
  NOT NOT1_7985(.VSS(VSS),.VDD(VDD),.Y(I29369),.A(g20967));
  NOT NOT1_7986(.VSS(VSS),.VDD(VDD),.Y(g22703),.A(I29369));
  NOT NOT1_7987(.VSS(VSS),.VDD(VDD),.Y(I29372),.A(g20968));
  NOT NOT1_7988(.VSS(VSS),.VDD(VDD),.Y(g22704),.A(I29372));
  NOT NOT1_7989(.VSS(VSS),.VDD(VDD),.Y(I29375),.A(g20969));
  NOT NOT1_7990(.VSS(VSS),.VDD(VDD),.Y(g22705),.A(I29375));
  NOT NOT1_7991(.VSS(VSS),.VDD(VDD),.Y(I29378),.A(g20970));
  NOT NOT1_7992(.VSS(VSS),.VDD(VDD),.Y(g22706),.A(I29378));
  NOT NOT1_7993(.VSS(VSS),.VDD(VDD),.Y(I29383),.A(g20972));
  NOT NOT1_7994(.VSS(VSS),.VDD(VDD),.Y(g22709),.A(I29383));
  NOT NOT1_7995(.VSS(VSS),.VDD(VDD),.Y(I29386),.A(g20973));
  NOT NOT1_7996(.VSS(VSS),.VDD(VDD),.Y(g22710),.A(I29386));
  NOT NOT1_7997(.VSS(VSS),.VDD(VDD),.Y(I29389),.A(g20974));
  NOT NOT1_7998(.VSS(VSS),.VDD(VDD),.Y(g22711),.A(I29389));
  NOT NOT1_7999(.VSS(VSS),.VDD(VDD),.Y(I29392),.A(g20975));
  NOT NOT1_8000(.VSS(VSS),.VDD(VDD),.Y(g22712),.A(I29392));
  NOT NOT1_8001(.VSS(VSS),.VDD(VDD),.Y(I29395),.A(g20976));
  NOT NOT1_8002(.VSS(VSS),.VDD(VDD),.Y(g22713),.A(I29395));
  NOT NOT1_8003(.VSS(VSS),.VDD(VDD),.Y(I29399),.A(g20977));
  NOT NOT1_8004(.VSS(VSS),.VDD(VDD),.Y(g22715),.A(I29399));
  NOT NOT1_8005(.VSS(VSS),.VDD(VDD),.Y(I29402),.A(g20978));
  NOT NOT1_8006(.VSS(VSS),.VDD(VDD),.Y(g22716),.A(I29402));
  NOT NOT1_8007(.VSS(VSS),.VDD(VDD),.Y(I29405),.A(g20979));
  NOT NOT1_8008(.VSS(VSS),.VDD(VDD),.Y(g22717),.A(I29405));
  NOT NOT1_8009(.VSS(VSS),.VDD(VDD),.Y(I29408),.A(g20980));
  NOT NOT1_8010(.VSS(VSS),.VDD(VDD),.Y(g22718),.A(I29408));
  NOT NOT1_8011(.VSS(VSS),.VDD(VDD),.Y(g22721),.A(g21164));
  NOT NOT1_8012(.VSS(VSS),.VDD(VDD),.Y(I29415),.A(g20981));
  NOT NOT1_8013(.VSS(VSS),.VDD(VDD),.Y(g22723),.A(I29415));
  NOT NOT1_8014(.VSS(VSS),.VDD(VDD),.Y(I29418),.A(g20982));
  NOT NOT1_8015(.VSS(VSS),.VDD(VDD),.Y(g22724),.A(I29418));
  NOT NOT1_8016(.VSS(VSS),.VDD(VDD),.Y(I29421),.A(g20983));
  NOT NOT1_8017(.VSS(VSS),.VDD(VDD),.Y(g22725),.A(I29421));
  NOT NOT1_8018(.VSS(VSS),.VDD(VDD),.Y(I29426),.A(g20989));
  NOT NOT1_8019(.VSS(VSS),.VDD(VDD),.Y(g22728),.A(I29426));
  NOT NOT1_8020(.VSS(VSS),.VDD(VDD),.Y(I29429),.A(g20990));
  NOT NOT1_8021(.VSS(VSS),.VDD(VDD),.Y(g22729),.A(I29429));
  NOT NOT1_8022(.VSS(VSS),.VDD(VDD),.Y(I29432),.A(g20991));
  NOT NOT1_8023(.VSS(VSS),.VDD(VDD),.Y(g22730),.A(I29432));
  NOT NOT1_8024(.VSS(VSS),.VDD(VDD),.Y(I29435),.A(g20992));
  NOT NOT1_8025(.VSS(VSS),.VDD(VDD),.Y(g22731),.A(I29435));
  NOT NOT1_8026(.VSS(VSS),.VDD(VDD),.Y(I29439),.A(g20993));
  NOT NOT1_8027(.VSS(VSS),.VDD(VDD),.Y(g22733),.A(I29439));
  NOT NOT1_8028(.VSS(VSS),.VDD(VDD),.Y(I29442),.A(g20994));
  NOT NOT1_8029(.VSS(VSS),.VDD(VDD),.Y(g22734),.A(I29442));
  NOT NOT1_8030(.VSS(VSS),.VDD(VDD),.Y(I29445),.A(g20995));
  NOT NOT1_8031(.VSS(VSS),.VDD(VDD),.Y(g22735),.A(I29445));
  NOT NOT1_8032(.VSS(VSS),.VDD(VDD),.Y(I29448),.A(g20996));
  NOT NOT1_8033(.VSS(VSS),.VDD(VDD),.Y(g22736),.A(I29448));
  NOT NOT1_8034(.VSS(VSS),.VDD(VDD),.Y(I29451),.A(g20997));
  NOT NOT1_8035(.VSS(VSS),.VDD(VDD),.Y(g22737),.A(I29451));
  NOT NOT1_8036(.VSS(VSS),.VDD(VDD),.Y(I29456),.A(g20999));
  NOT NOT1_8037(.VSS(VSS),.VDD(VDD),.Y(g22740),.A(I29456));
  NOT NOT1_8038(.VSS(VSS),.VDD(VDD),.Y(I29459),.A(g21000));
  NOT NOT1_8039(.VSS(VSS),.VDD(VDD),.Y(g22741),.A(I29459));
  NOT NOT1_8040(.VSS(VSS),.VDD(VDD),.Y(I29462),.A(g21001));
  NOT NOT1_8041(.VSS(VSS),.VDD(VDD),.Y(g22742),.A(I29462));
  NOT NOT1_8042(.VSS(VSS),.VDD(VDD),.Y(I29465),.A(g21002));
  NOT NOT1_8043(.VSS(VSS),.VDD(VDD),.Y(g22743),.A(I29465));
  NOT NOT1_8044(.VSS(VSS),.VDD(VDD),.Y(I29468),.A(g21003));
  NOT NOT1_8045(.VSS(VSS),.VDD(VDD),.Y(g22744),.A(I29468));
  NOT NOT1_8046(.VSS(VSS),.VDD(VDD),.Y(I29472),.A(g21004));
  NOT NOT1_8047(.VSS(VSS),.VDD(VDD),.Y(g22746),.A(I29472));
  NOT NOT1_8048(.VSS(VSS),.VDD(VDD),.Y(I29475),.A(g21005));
  NOT NOT1_8049(.VSS(VSS),.VDD(VDD),.Y(g22747),.A(I29475));
  NOT NOT1_8050(.VSS(VSS),.VDD(VDD),.Y(I29478),.A(g21006));
  NOT NOT1_8051(.VSS(VSS),.VDD(VDD),.Y(g22748),.A(I29478));
  NOT NOT1_8052(.VSS(VSS),.VDD(VDD),.Y(I29481),.A(g21007));
  NOT NOT1_8053(.VSS(VSS),.VDD(VDD),.Y(g22749),.A(I29481));
  NOT NOT1_8054(.VSS(VSS),.VDD(VDD),.Y(I29484),.A(g21903));
  NOT NOT1_8055(.VSS(VSS),.VDD(VDD),.Y(g22750),.A(I29484));
  NOT NOT1_8056(.VSS(VSS),.VDD(VDD),.Y(g22753),.A(g21184));
  NOT NOT1_8057(.VSS(VSS),.VDD(VDD),.Y(I29490),.A(g21009));
  NOT NOT1_8058(.VSS(VSS),.VDD(VDD),.Y(g22756),.A(I29490));
  NOT NOT1_8059(.VSS(VSS),.VDD(VDD),.Y(I29493),.A(g21010));
  NOT NOT1_8060(.VSS(VSS),.VDD(VDD),.Y(g22757),.A(I29493));
  NOT NOT1_8061(.VSS(VSS),.VDD(VDD),.Y(I29496),.A(g21011));
  NOT NOT1_8062(.VSS(VSS),.VDD(VDD),.Y(g22758),.A(I29496));
  NOT NOT1_8063(.VSS(VSS),.VDD(VDD),.Y(I29500),.A(g21015));
  NOT NOT1_8064(.VSS(VSS),.VDD(VDD),.Y(g22760),.A(I29500));
  NOT NOT1_8065(.VSS(VSS),.VDD(VDD),.Y(I29503),.A(g21016));
  NOT NOT1_8066(.VSS(VSS),.VDD(VDD),.Y(g22761),.A(I29503));
  NOT NOT1_8067(.VSS(VSS),.VDD(VDD),.Y(I29506),.A(g21017));
  NOT NOT1_8068(.VSS(VSS),.VDD(VDD),.Y(g22762),.A(I29506));
  NOT NOT1_8069(.VSS(VSS),.VDD(VDD),.Y(I29509),.A(g21018));
  NOT NOT1_8070(.VSS(VSS),.VDD(VDD),.Y(g22763),.A(I29509));
  NOT NOT1_8071(.VSS(VSS),.VDD(VDD),.Y(I29513),.A(g21019));
  NOT NOT1_8072(.VSS(VSS),.VDD(VDD),.Y(g22765),.A(I29513));
  NOT NOT1_8073(.VSS(VSS),.VDD(VDD),.Y(I29516),.A(g21020));
  NOT NOT1_8074(.VSS(VSS),.VDD(VDD),.Y(g22766),.A(I29516));
  NOT NOT1_8075(.VSS(VSS),.VDD(VDD),.Y(I29519),.A(g21021));
  NOT NOT1_8076(.VSS(VSS),.VDD(VDD),.Y(g22767),.A(I29519));
  NOT NOT1_8077(.VSS(VSS),.VDD(VDD),.Y(I29522),.A(g21022));
  NOT NOT1_8078(.VSS(VSS),.VDD(VDD),.Y(g22768),.A(I29522));
  NOT NOT1_8079(.VSS(VSS),.VDD(VDD),.Y(I29525),.A(g21023));
  NOT NOT1_8080(.VSS(VSS),.VDD(VDD),.Y(g22769),.A(I29525));
  NOT NOT1_8081(.VSS(VSS),.VDD(VDD),.Y(I29530),.A(g21025));
  NOT NOT1_8082(.VSS(VSS),.VDD(VDD),.Y(g22772),.A(I29530));
  NOT NOT1_8083(.VSS(VSS),.VDD(VDD),.Y(I29533),.A(g21026));
  NOT NOT1_8084(.VSS(VSS),.VDD(VDD),.Y(g22773),.A(I29533));
  NOT NOT1_8085(.VSS(VSS),.VDD(VDD),.Y(I29536),.A(g21027));
  NOT NOT1_8086(.VSS(VSS),.VDD(VDD),.Y(g22774),.A(I29536));
  NOT NOT1_8087(.VSS(VSS),.VDD(VDD),.Y(I29539),.A(g21028));
  NOT NOT1_8088(.VSS(VSS),.VDD(VDD),.Y(g22775),.A(I29539));
  NOT NOT1_8089(.VSS(VSS),.VDD(VDD),.Y(I29542),.A(g21029));
  NOT NOT1_8090(.VSS(VSS),.VDD(VDD),.Y(g22776),.A(I29542));
  NOT NOT1_8091(.VSS(VSS),.VDD(VDD),.Y(g22777),.A(g21796));
  NOT NOT1_8092(.VSS(VSS),.VDD(VDD),.Y(I29547),.A(g21031));
  NOT NOT1_8093(.VSS(VSS),.VDD(VDD),.Y(g22785),.A(I29547));
  NOT NOT1_8094(.VSS(VSS),.VDD(VDD),.Y(I29550),.A(g21032));
  NOT NOT1_8095(.VSS(VSS),.VDD(VDD),.Y(g22786),.A(I29550));
  NOT NOT1_8096(.VSS(VSS),.VDD(VDD),.Y(g22787),.A(g21199));
  NOT NOT1_8097(.VSS(VSS),.VDD(VDD),.Y(I29556),.A(g21033));
  NOT NOT1_8098(.VSS(VSS),.VDD(VDD),.Y(g22790),.A(I29556));
  NOT NOT1_8099(.VSS(VSS),.VDD(VDD),.Y(I29559),.A(g21034));
  NOT NOT1_8100(.VSS(VSS),.VDD(VDD),.Y(g22791),.A(I29559));
  NOT NOT1_8101(.VSS(VSS),.VDD(VDD),.Y(I29562),.A(g21035));
  NOT NOT1_8102(.VSS(VSS),.VDD(VDD),.Y(g22792),.A(I29562));
  NOT NOT1_8103(.VSS(VSS),.VDD(VDD),.Y(I29566),.A(g21039));
  NOT NOT1_8104(.VSS(VSS),.VDD(VDD),.Y(g22794),.A(I29566));
  NOT NOT1_8105(.VSS(VSS),.VDD(VDD),.Y(I29569),.A(g21040));
  NOT NOT1_8106(.VSS(VSS),.VDD(VDD),.Y(g22795),.A(I29569));
  NOT NOT1_8107(.VSS(VSS),.VDD(VDD),.Y(I29572),.A(g21041));
  NOT NOT1_8108(.VSS(VSS),.VDD(VDD),.Y(g22796),.A(I29572));
  NOT NOT1_8109(.VSS(VSS),.VDD(VDD),.Y(I29575),.A(g21042));
  NOT NOT1_8110(.VSS(VSS),.VDD(VDD),.Y(g22797),.A(I29575));
  NOT NOT1_8111(.VSS(VSS),.VDD(VDD),.Y(I29579),.A(g21043));
  NOT NOT1_8112(.VSS(VSS),.VDD(VDD),.Y(g22799),.A(I29579));
  NOT NOT1_8113(.VSS(VSS),.VDD(VDD),.Y(I29582),.A(g21044));
  NOT NOT1_8114(.VSS(VSS),.VDD(VDD),.Y(g22800),.A(I29582));
  NOT NOT1_8115(.VSS(VSS),.VDD(VDD),.Y(I29585),.A(g21045));
  NOT NOT1_8116(.VSS(VSS),.VDD(VDD),.Y(g22801),.A(I29585));
  NOT NOT1_8117(.VSS(VSS),.VDD(VDD),.Y(I29588),.A(g21046));
  NOT NOT1_8118(.VSS(VSS),.VDD(VDD),.Y(g22802),.A(I29588));
  NOT NOT1_8119(.VSS(VSS),.VDD(VDD),.Y(I29591),.A(g21047));
  NOT NOT1_8120(.VSS(VSS),.VDD(VDD),.Y(g22803),.A(I29591));
  NOT NOT1_8121(.VSS(VSS),.VDD(VDD),.Y(g22805),.A(g21894));
  NOT NOT1_8122(.VSS(VSS),.VDD(VDD),.Y(g22806),.A(g21615));
  NOT NOT1_8123(.VSS(VSS),.VDD(VDD),.Y(I29600),.A(g21720));
  NOT NOT1_8124(.VSS(VSS),.VDD(VDD),.Y(g22812),.A(I29600));
  NOT NOT1_8125(.VSS(VSS),.VDD(VDD),.Y(I29603),.A(g21051));
  NOT NOT1_8126(.VSS(VSS),.VDD(VDD),.Y(g22824),.A(I29603));
  NOT NOT1_8127(.VSS(VSS),.VDD(VDD),.Y(I29606),.A(g21364));
  NOT NOT1_8128(.VSS(VSS),.VDD(VDD),.Y(g22825),.A(I29606));
  NOT NOT1_8129(.VSS(VSS),.VDD(VDD),.Y(I29610),.A(g21052));
  NOT NOT1_8130(.VSS(VSS),.VDD(VDD),.Y(g22827),.A(I29610));
  NOT NOT1_8131(.VSS(VSS),.VDD(VDD),.Y(I29613),.A(g21053));
  NOT NOT1_8132(.VSS(VSS),.VDD(VDD),.Y(g22828),.A(I29613));
  NOT NOT1_8133(.VSS(VSS),.VDD(VDD),.Y(g22829),.A(g21214));
  NOT NOT1_8134(.VSS(VSS),.VDD(VDD),.Y(I29619),.A(g21054));
  NOT NOT1_8135(.VSS(VSS),.VDD(VDD),.Y(g22832),.A(I29619));
  NOT NOT1_8136(.VSS(VSS),.VDD(VDD),.Y(I29622),.A(g21055));
  NOT NOT1_8137(.VSS(VSS),.VDD(VDD),.Y(g22833),.A(I29622));
  NOT NOT1_8138(.VSS(VSS),.VDD(VDD),.Y(I29625),.A(g21056));
  NOT NOT1_8139(.VSS(VSS),.VDD(VDD),.Y(g22834),.A(I29625));
  NOT NOT1_8140(.VSS(VSS),.VDD(VDD),.Y(I29629),.A(g21060));
  NOT NOT1_8141(.VSS(VSS),.VDD(VDD),.Y(g22836),.A(I29629));
  NOT NOT1_8142(.VSS(VSS),.VDD(VDD),.Y(I29632),.A(g21061));
  NOT NOT1_8143(.VSS(VSS),.VDD(VDD),.Y(g22837),.A(I29632));
  NOT NOT1_8144(.VSS(VSS),.VDD(VDD),.Y(I29635),.A(g21062));
  NOT NOT1_8145(.VSS(VSS),.VDD(VDD),.Y(g22838),.A(I29635));
  NOT NOT1_8146(.VSS(VSS),.VDD(VDD),.Y(I29638),.A(g21063));
  NOT NOT1_8147(.VSS(VSS),.VDD(VDD),.Y(g22839),.A(I29638));
  NOT NOT1_8148(.VSS(VSS),.VDD(VDD),.Y(I29641),.A(g20825));
  NOT NOT1_8149(.VSS(VSS),.VDD(VDD),.Y(g22840),.A(I29641));
  NOT NOT1_8150(.VSS(VSS),.VDD(VDD),.Y(g22843),.A(g21889));
  NOT NOT1_8151(.VSS(VSS),.VDD(VDD),.Y(g22847),.A(g21643));
  NOT NOT1_8152(.VSS(VSS),.VDD(VDD),.Y(I29653),.A(g21746));
  NOT NOT1_8153(.VSS(VSS),.VDD(VDD),.Y(g22852),.A(I29653));
  NOT NOT1_8154(.VSS(VSS),.VDD(VDD),.Y(I29656),.A(g21070));
  NOT NOT1_8155(.VSS(VSS),.VDD(VDD),.Y(g22864),.A(I29656));
  NOT NOT1_8156(.VSS(VSS),.VDD(VDD),.Y(I29660),.A(g21071));
  NOT NOT1_8157(.VSS(VSS),.VDD(VDD),.Y(g22866),.A(I29660));
  NOT NOT1_8158(.VSS(VSS),.VDD(VDD),.Y(I29663),.A(g21072));
  NOT NOT1_8159(.VSS(VSS),.VDD(VDD),.Y(g22867),.A(I29663));
  NOT NOT1_8160(.VSS(VSS),.VDD(VDD),.Y(g22868),.A(g21222));
  NOT NOT1_8161(.VSS(VSS),.VDD(VDD),.Y(I29669),.A(g21073));
  NOT NOT1_8162(.VSS(VSS),.VDD(VDD),.Y(g22871),.A(I29669));
  NOT NOT1_8163(.VSS(VSS),.VDD(VDD),.Y(I29672),.A(g21074));
  NOT NOT1_8164(.VSS(VSS),.VDD(VDD),.Y(g22872),.A(I29672));
  NOT NOT1_8165(.VSS(VSS),.VDD(VDD),.Y(I29675),.A(g21075));
  NOT NOT1_8166(.VSS(VSS),.VDD(VDD),.Y(g22873),.A(I29675));
  NOT NOT1_8167(.VSS(VSS),.VDD(VDD),.Y(g22875),.A(g21884));
  NOT NOT1_8168(.VSS(VSS),.VDD(VDD),.Y(g22882),.A(g21674));
  NOT NOT1_8169(.VSS(VSS),.VDD(VDD),.Y(I29687),.A(g21770));
  NOT NOT1_8170(.VSS(VSS),.VDD(VDD),.Y(g22887),.A(I29687));
  NOT NOT1_8171(.VSS(VSS),.VDD(VDD),.Y(I29690),.A(g21080));
  NOT NOT1_8172(.VSS(VSS),.VDD(VDD),.Y(g22899),.A(I29690));
  NOT NOT1_8173(.VSS(VSS),.VDD(VDD),.Y(I29694),.A(g21081));
  NOT NOT1_8174(.VSS(VSS),.VDD(VDD),.Y(g22901),.A(I29694));
  NOT NOT1_8175(.VSS(VSS),.VDD(VDD),.Y(I29697),.A(g21082));
  NOT NOT1_8176(.VSS(VSS),.VDD(VDD),.Y(g22902),.A(I29697));
  NOT NOT1_8177(.VSS(VSS),.VDD(VDD),.Y(I29700),.A(g20700));
  NOT NOT1_8178(.VSS(VSS),.VDD(VDD),.Y(g22903),.A(I29700));
  NOT NOT1_8179(.VSS(VSS),.VDD(VDD),.Y(g22907),.A(g21711));
  NOT NOT1_8180(.VSS(VSS),.VDD(VDD),.Y(g22917),.A(g21703));
  NOT NOT1_8181(.VSS(VSS),.VDD(VDD),.Y(I29712),.A(g21786));
  NOT NOT1_8182(.VSS(VSS),.VDD(VDD),.Y(g22922),.A(I29712));
  NOT NOT1_8183(.VSS(VSS),.VDD(VDD),.Y(I29715),.A(g21094));
  NOT NOT1_8184(.VSS(VSS),.VDD(VDD),.Y(g22934),.A(I29715));
  NOT NOT1_8185(.VSS(VSS),.VDD(VDD),.Y(I29724),.A(g21851));
  NOT NOT1_8186(.VSS(VSS),.VDD(VDD),.Y(g22945),.A(I29724));
  NOT NOT1_8187(.VSS(VSS),.VDD(VDD),.Y(I29727),.A(g20877));
  NOT NOT1_8188(.VSS(VSS),.VDD(VDD),.Y(g22948),.A(I29727));
  NOT NOT1_8189(.VSS(VSS),.VDD(VDD),.Y(g22949),.A(g21665));
  NOT NOT1_8190(.VSS(VSS),.VDD(VDD),.Y(g22954),.A(g21739));
  NOT NOT1_8191(.VSS(VSS),.VDD(VDD),.Y(g22958),.A(g21694));
  NOT NOT1_8192(.VSS(VSS),.VDD(VDD),.Y(g22962),.A(g21763));
  NOT NOT1_8193(.VSS(VSS),.VDD(VDD),.Y(g22966),.A(g21730));
  NOT NOT1_8194(.VSS(VSS),.VDD(VDD),.Y(I29736),.A(g20884));
  NOT NOT1_8195(.VSS(VSS),.VDD(VDD),.Y(g22970),.A(I29736));
  NOT NOT1_8196(.VSS(VSS),.VDD(VDD),.Y(g22971),.A(g21779));
  NOT NOT1_8197(.VSS(VSS),.VDD(VDD),.Y(g22975),.A(g21756));
  NOT NOT1_8198(.VSS(VSS),.VDD(VDD),.Y(I29741),.A(g21346));
  NOT NOT1_8199(.VSS(VSS),.VDD(VDD),.Y(g22979),.A(I29741));
  NOT NOT1_8200(.VSS(VSS),.VDD(VDD),.Y(g22980),.A(g21794));
  NOT NOT1_8201(.VSS(VSS),.VDD(VDD),.Y(g22986),.A(g21382));
  NOT NOT1_8202(.VSS(VSS),.VDD(VDD),.Y(g22988),.A(g21404));
  NOT NOT1_8203(.VSS(VSS),.VDD(VDD),.Y(g22989),.A(g21415));
  NOT NOT1_8204(.VSS(VSS),.VDD(VDD),.Y(g22991),.A(g21429));
  NOT NOT1_8205(.VSS(VSS),.VDD(VDD),.Y(g22995),.A(g21441));
  NOT NOT1_8206(.VSS(VSS),.VDD(VDD),.Y(g22996),.A(g21449));
  NOT NOT1_8207(.VSS(VSS),.VDD(VDD),.Y(g22998),.A(g21458));
  NOT NOT1_8208(.VSS(VSS),.VDD(VDD),.Y(g23001),.A(g21473));
  NOT NOT1_8209(.VSS(VSS),.VDD(VDD),.Y(g23002),.A(g21477));
  NOT NOT1_8210(.VSS(VSS),.VDD(VDD),.Y(g23006),.A(g21483));
  NOT NOT1_8211(.VSS(VSS),.VDD(VDD),.Y(g23007),.A(g21491));
  NOT NOT1_8212(.VSS(VSS),.VDD(VDD),.Y(g23008),.A(g21498));
  NOT NOT1_8213(.VSS(VSS),.VDD(VDD),.Y(g23012),.A(g21505));
  NOT NOT1_8214(.VSS(VSS),.VDD(VDD),.Y(g23015),.A(g21514));
  NOT NOT1_8215(.VSS(VSS),.VDD(VDD),.Y(g23016),.A(g21518));
  NOT NOT1_8216(.VSS(VSS),.VDD(VDD),.Y(g23020),.A(g21524));
  NOT NOT1_8217(.VSS(VSS),.VDD(VDD),.Y(g23021),.A(g21530));
  NOT NOT1_8218(.VSS(VSS),.VDD(VDD),.Y(g23024),.A(g21537));
  NOT NOT1_8219(.VSS(VSS),.VDD(VDD),.Y(g23028),.A(g21541));
  NOT NOT1_8220(.VSS(VSS),.VDD(VDD),.Y(g23031),.A(g21550));
  NOT NOT1_8221(.VSS(VSS),.VDD(VDD),.Y(g23032),.A(g21554));
  NOT NOT1_8222(.VSS(VSS),.VDD(VDD),.Y(g23036),.A(g21558));
  NOT NOT1_8223(.VSS(VSS),.VDD(VDD),.Y(g23037),.A(g21561));
  NOT NOT1_8224(.VSS(VSS),.VDD(VDD),.Y(g23038),.A(g21566));
  NOT NOT1_8225(.VSS(VSS),.VDD(VDD),.Y(g23041),.A(g21573));
  NOT NOT1_8226(.VSS(VSS),.VDD(VDD),.Y(g23045),.A(g21577));
  NOT NOT1_8227(.VSS(VSS),.VDD(VDD),.Y(g23048),.A(g21586));
  NOT NOT1_8228(.VSS(VSS),.VDD(VDD),.Y(g23049),.A(g21590));
  NOT NOT1_8229(.VSS(VSS),.VDD(VDD),.Y(I29797),.A(g21432));
  NOT NOT1_8230(.VSS(VSS),.VDD(VDD),.Y(g23050),.A(I29797));
  NOT NOT1_8231(.VSS(VSS),.VDD(VDD),.Y(I29802),.A(g21435));
  NOT NOT1_8232(.VSS(VSS),.VDD(VDD),.Y(g23055),.A(I29802));
  NOT NOT1_8233(.VSS(VSS),.VDD(VDD),.Y(g23056),.A(g21594));
  NOT NOT1_8234(.VSS(VSS),.VDD(VDD),.Y(g23057),.A(g21599));
  NOT NOT1_8235(.VSS(VSS),.VDD(VDD),.Y(g23060),.A(g21606));
  NOT NOT1_8236(.VSS(VSS),.VDD(VDD),.Y(g23064),.A(g21612));
  NOT NOT1_8237(.VSS(VSS),.VDD(VDD),.Y(I29812),.A(g21467));
  NOT NOT1_8238(.VSS(VSS),.VDD(VDD),.Y(g23065),.A(I29812));
  NOT NOT1_8239(.VSS(VSS),.VDD(VDD),.Y(I29817),.A(g21470));
  NOT NOT1_8240(.VSS(VSS),.VDD(VDD),.Y(g23068),.A(I29817));
  NOT NOT1_8241(.VSS(VSS),.VDD(VDD),.Y(g23069),.A(g21619));
  NOT NOT1_8242(.VSS(VSS),.VDD(VDD),.Y(g23074),.A(g21623));
  NOT NOT1_8243(.VSS(VSS),.VDD(VDD),.Y(g23075),.A(g21628));
  NOT NOT1_8244(.VSS(VSS),.VDD(VDD),.Y(I29827),.A(g21502));
  NOT NOT1_8245(.VSS(VSS),.VDD(VDD),.Y(g23078),.A(I29827));
  NOT NOT1_8246(.VSS(VSS),.VDD(VDD),.Y(g23079),.A(g21640));
  NOT NOT1_8247(.VSS(VSS),.VDD(VDD),.Y(g23082),.A(g21647));
  NOT NOT1_8248(.VSS(VSS),.VDD(VDD),.Y(g23087),.A(g21651));
  NOT NOT1_8249(.VSS(VSS),.VDD(VDD),.Y(g23088),.A(g21655));
  NOT NOT1_8250(.VSS(VSS),.VDD(VDD),.Y(I29841),.A(g21316));
  NOT NOT1_8251(.VSS(VSS),.VDD(VDD),.Y(g23094),.A(I29841));
  NOT NOT1_8252(.VSS(VSS),.VDD(VDD),.Y(g23095),.A(g21671));
  NOT NOT1_8253(.VSS(VSS),.VDD(VDD),.Y(g23098),.A(g21678));
  NOT NOT1_8254(.VSS(VSS),.VDD(VDD),.Y(g23103),.A(g21682));
  NOT NOT1_8255(.VSS(VSS),.VDD(VDD),.Y(I29852),.A(g21331));
  NOT NOT1_8256(.VSS(VSS),.VDD(VDD),.Y(g23105),.A(I29852));
  NOT NOT1_8257(.VSS(VSS),.VDD(VDD),.Y(g23112),.A(g21700));
  NOT NOT1_8258(.VSS(VSS),.VDD(VDD),.Y(g23115),.A(g21708));
  NOT NOT1_8259(.VSS(VSS),.VDD(VDD),.Y(I29863),.A(g21346));
  NOT NOT1_8260(.VSS(VSS),.VDD(VDD),.Y(g23116),.A(I29863));
  NOT NOT1_8261(.VSS(VSS),.VDD(VDD),.Y(I29872),.A(g21364));
  NOT NOT1_8262(.VSS(VSS),.VDD(VDD),.Y(g23125),.A(I29872));
  NOT NOT1_8263(.VSS(VSS),.VDD(VDD),.Y(I29881),.A(g21385));
  NOT NOT1_8264(.VSS(VSS),.VDD(VDD),.Y(g23134),.A(I29881));
  NOT NOT1_8265(.VSS(VSS),.VDD(VDD),.Y(g23140),.A(g21825));
  NOT NOT1_8266(.VSS(VSS),.VDD(VDD),.Y(g23141),.A(g21825));
  NOT NOT1_8267(.VSS(VSS),.VDD(VDD),.Y(g23142),.A(g21825));
  NOT NOT1_8268(.VSS(VSS),.VDD(VDD),.Y(g23143),.A(g21825));
  NOT NOT1_8269(.VSS(VSS),.VDD(VDD),.Y(g23144),.A(g21825));
  NOT NOT1_8270(.VSS(VSS),.VDD(VDD),.Y(g23145),.A(g21825));
  NOT NOT1_8271(.VSS(VSS),.VDD(VDD),.Y(g23146),.A(g21825));
  NOT NOT1_8272(.VSS(VSS),.VDD(VDD),.Y(g23147),.A(g21825));
  NOT NOT1_8273(.VSS(VSS),.VDD(VDD),.Y(I29897),.A(g23116));
  NOT NOT1_8274(.VSS(VSS),.VDD(VDD),.Y(g23148),.A(I29897));
  NOT NOT1_8275(.VSS(VSS),.VDD(VDD),.Y(I29900),.A(g23125));
  NOT NOT1_8276(.VSS(VSS),.VDD(VDD),.Y(g23149),.A(I29900));
  NOT NOT1_8277(.VSS(VSS),.VDD(VDD),.Y(I29903),.A(g23134));
  NOT NOT1_8278(.VSS(VSS),.VDD(VDD),.Y(g23150),.A(I29903));
  NOT NOT1_8279(.VSS(VSS),.VDD(VDD),.Y(I29906),.A(g21967));
  NOT NOT1_8280(.VSS(VSS),.VDD(VDD),.Y(g23151),.A(I29906));
  NOT NOT1_8281(.VSS(VSS),.VDD(VDD),.Y(I29909),.A(g23050));
  NOT NOT1_8282(.VSS(VSS),.VDD(VDD),.Y(g23152),.A(I29909));
  NOT NOT1_8283(.VSS(VSS),.VDD(VDD),.Y(I29912),.A(g23065));
  NOT NOT1_8284(.VSS(VSS),.VDD(VDD),.Y(g23153),.A(I29912));
  NOT NOT1_8285(.VSS(VSS),.VDD(VDD),.Y(I29915),.A(g23055));
  NOT NOT1_8286(.VSS(VSS),.VDD(VDD),.Y(g23154),.A(I29915));
  NOT NOT1_8287(.VSS(VSS),.VDD(VDD),.Y(I29918),.A(g23068));
  NOT NOT1_8288(.VSS(VSS),.VDD(VDD),.Y(g23155),.A(I29918));
  NOT NOT1_8289(.VSS(VSS),.VDD(VDD),.Y(I29921),.A(g23078));
  NOT NOT1_8290(.VSS(VSS),.VDD(VDD),.Y(g23156),.A(I29921));
  NOT NOT1_8291(.VSS(VSS),.VDD(VDD),.Y(I29924),.A(g23094));
  NOT NOT1_8292(.VSS(VSS),.VDD(VDD),.Y(g23157),.A(I29924));
  NOT NOT1_8293(.VSS(VSS),.VDD(VDD),.Y(I29927),.A(g23105));
  NOT NOT1_8294(.VSS(VSS),.VDD(VDD),.Y(g23158),.A(I29927));
  NOT NOT1_8295(.VSS(VSS),.VDD(VDD),.Y(I29930),.A(g22176));
  NOT NOT1_8296(.VSS(VSS),.VDD(VDD),.Y(g23159),.A(I29930));
  NOT NOT1_8297(.VSS(VSS),.VDD(VDD),.Y(I29933),.A(g22082));
  NOT NOT1_8298(.VSS(VSS),.VDD(VDD),.Y(g23160),.A(I29933));
  NOT NOT1_8299(.VSS(VSS),.VDD(VDD),.Y(I29936),.A(g22582));
  NOT NOT1_8300(.VSS(VSS),.VDD(VDD),.Y(g23161),.A(I29936));
  NOT NOT1_8301(.VSS(VSS),.VDD(VDD),.Y(I29939),.A(g22518));
  NOT NOT1_8302(.VSS(VSS),.VDD(VDD),.Y(g23162),.A(I29939));
  NOT NOT1_8303(.VSS(VSS),.VDD(VDD),.Y(I29942),.A(g22548));
  NOT NOT1_8304(.VSS(VSS),.VDD(VDD),.Y(g23163),.A(I29942));
  NOT NOT1_8305(.VSS(VSS),.VDD(VDD),.Y(I29945),.A(g22583));
  NOT NOT1_8306(.VSS(VSS),.VDD(VDD),.Y(g23164),.A(I29945));
  NOT NOT1_8307(.VSS(VSS),.VDD(VDD),.Y(I29948),.A(g22549));
  NOT NOT1_8308(.VSS(VSS),.VDD(VDD),.Y(g23165),.A(I29948));
  NOT NOT1_8309(.VSS(VSS),.VDD(VDD),.Y(I29951),.A(g22584));
  NOT NOT1_8310(.VSS(VSS),.VDD(VDD),.Y(g23166),.A(I29951));
  NOT NOT1_8311(.VSS(VSS),.VDD(VDD),.Y(I29954),.A(g22611));
  NOT NOT1_8312(.VSS(VSS),.VDD(VDD),.Y(g23167),.A(I29954));
  NOT NOT1_8313(.VSS(VSS),.VDD(VDD),.Y(I29957),.A(g22585));
  NOT NOT1_8314(.VSS(VSS),.VDD(VDD),.Y(g23168),.A(I29957));
  NOT NOT1_8315(.VSS(VSS),.VDD(VDD),.Y(I29960),.A(g22612));
  NOT NOT1_8316(.VSS(VSS),.VDD(VDD),.Y(g23169),.A(I29960));
  NOT NOT1_8317(.VSS(VSS),.VDD(VDD),.Y(I29963),.A(g22639));
  NOT NOT1_8318(.VSS(VSS),.VDD(VDD),.Y(g23170),.A(I29963));
  NOT NOT1_8319(.VSS(VSS),.VDD(VDD),.Y(I29966),.A(g22613));
  NOT NOT1_8320(.VSS(VSS),.VDD(VDD),.Y(g23171),.A(I29966));
  NOT NOT1_8321(.VSS(VSS),.VDD(VDD),.Y(I29969),.A(g22640));
  NOT NOT1_8322(.VSS(VSS),.VDD(VDD),.Y(g23172),.A(I29969));
  NOT NOT1_8323(.VSS(VSS),.VDD(VDD),.Y(I29972),.A(g22669));
  NOT NOT1_8324(.VSS(VSS),.VDD(VDD),.Y(g23173),.A(I29972));
  NOT NOT1_8325(.VSS(VSS),.VDD(VDD),.Y(I29975),.A(g22641));
  NOT NOT1_8326(.VSS(VSS),.VDD(VDD),.Y(g23174),.A(I29975));
  NOT NOT1_8327(.VSS(VSS),.VDD(VDD),.Y(I29978),.A(g22670));
  NOT NOT1_8328(.VSS(VSS),.VDD(VDD),.Y(g23175),.A(I29978));
  NOT NOT1_8329(.VSS(VSS),.VDD(VDD),.Y(I29981),.A(g22702));
  NOT NOT1_8330(.VSS(VSS),.VDD(VDD),.Y(g23176),.A(I29981));
  NOT NOT1_8331(.VSS(VSS),.VDD(VDD),.Y(I29984),.A(g22671));
  NOT NOT1_8332(.VSS(VSS),.VDD(VDD),.Y(g23177),.A(I29984));
  NOT NOT1_8333(.VSS(VSS),.VDD(VDD),.Y(I29987),.A(g22703));
  NOT NOT1_8334(.VSS(VSS),.VDD(VDD),.Y(g23178),.A(I29987));
  NOT NOT1_8335(.VSS(VSS),.VDD(VDD),.Y(I29990),.A(g22728));
  NOT NOT1_8336(.VSS(VSS),.VDD(VDD),.Y(g23179),.A(I29990));
  NOT NOT1_8337(.VSS(VSS),.VDD(VDD),.Y(I29993),.A(g22704));
  NOT NOT1_8338(.VSS(VSS),.VDD(VDD),.Y(g23180),.A(I29993));
  NOT NOT1_8339(.VSS(VSS),.VDD(VDD),.Y(I29996),.A(g22729));
  NOT NOT1_8340(.VSS(VSS),.VDD(VDD),.Y(g23181),.A(I29996));
  NOT NOT1_8341(.VSS(VSS),.VDD(VDD),.Y(I29999),.A(g22756));
  NOT NOT1_8342(.VSS(VSS),.VDD(VDD),.Y(g23182),.A(I29999));
  NOT NOT1_8343(.VSS(VSS),.VDD(VDD),.Y(I30002),.A(g22730));
  NOT NOT1_8344(.VSS(VSS),.VDD(VDD),.Y(g23183),.A(I30002));
  NOT NOT1_8345(.VSS(VSS),.VDD(VDD),.Y(I30005),.A(g22757));
  NOT NOT1_8346(.VSS(VSS),.VDD(VDD),.Y(g23184),.A(I30005));
  NOT NOT1_8347(.VSS(VSS),.VDD(VDD),.Y(I30008),.A(g22785));
  NOT NOT1_8348(.VSS(VSS),.VDD(VDD),.Y(g23185),.A(I30008));
  NOT NOT1_8349(.VSS(VSS),.VDD(VDD),.Y(I30011),.A(g22758));
  NOT NOT1_8350(.VSS(VSS),.VDD(VDD),.Y(g23186),.A(I30011));
  NOT NOT1_8351(.VSS(VSS),.VDD(VDD),.Y(I30014),.A(g22786));
  NOT NOT1_8352(.VSS(VSS),.VDD(VDD),.Y(g23187),.A(I30014));
  NOT NOT1_8353(.VSS(VSS),.VDD(VDD),.Y(I30017),.A(g22824));
  NOT NOT1_8354(.VSS(VSS),.VDD(VDD),.Y(g23188),.A(I30017));
  NOT NOT1_8355(.VSS(VSS),.VDD(VDD),.Y(I30020),.A(g22519));
  NOT NOT1_8356(.VSS(VSS),.VDD(VDD),.Y(g23189),.A(I30020));
  NOT NOT1_8357(.VSS(VSS),.VDD(VDD),.Y(I30023),.A(g22550));
  NOT NOT1_8358(.VSS(VSS),.VDD(VDD),.Y(g23190),.A(I30023));
  NOT NOT1_8359(.VSS(VSS),.VDD(VDD),.Y(I30026),.A(g22586));
  NOT NOT1_8360(.VSS(VSS),.VDD(VDD),.Y(g23191),.A(I30026));
  NOT NOT1_8361(.VSS(VSS),.VDD(VDD),.Y(I30029),.A(g22642));
  NOT NOT1_8362(.VSS(VSS),.VDD(VDD),.Y(g23192),.A(I30029));
  NOT NOT1_8363(.VSS(VSS),.VDD(VDD),.Y(I30032),.A(g22672));
  NOT NOT1_8364(.VSS(VSS),.VDD(VDD),.Y(g23193),.A(I30032));
  NOT NOT1_8365(.VSS(VSS),.VDD(VDD),.Y(I30035),.A(g22705));
  NOT NOT1_8366(.VSS(VSS),.VDD(VDD),.Y(g23194),.A(I30035));
  NOT NOT1_8367(.VSS(VSS),.VDD(VDD),.Y(I30038),.A(g22673));
  NOT NOT1_8368(.VSS(VSS),.VDD(VDD),.Y(g23195),.A(I30038));
  NOT NOT1_8369(.VSS(VSS),.VDD(VDD),.Y(I30041),.A(g22706));
  NOT NOT1_8370(.VSS(VSS),.VDD(VDD),.Y(g23196),.A(I30041));
  NOT NOT1_8371(.VSS(VSS),.VDD(VDD),.Y(I30044),.A(g22731));
  NOT NOT1_8372(.VSS(VSS),.VDD(VDD),.Y(g23197),.A(I30044));
  NOT NOT1_8373(.VSS(VSS),.VDD(VDD),.Y(I30047),.A(g22107));
  NOT NOT1_8374(.VSS(VSS),.VDD(VDD),.Y(g23198),.A(I30047));
  NOT NOT1_8375(.VSS(VSS),.VDD(VDD),.Y(I30050),.A(g22619));
  NOT NOT1_8376(.VSS(VSS),.VDD(VDD),.Y(g23199),.A(I30050));
  NOT NOT1_8377(.VSS(VSS),.VDD(VDD),.Y(I30053),.A(g22558));
  NOT NOT1_8378(.VSS(VSS),.VDD(VDD),.Y(g23200),.A(I30053));
  NOT NOT1_8379(.VSS(VSS),.VDD(VDD),.Y(I30056),.A(g22589));
  NOT NOT1_8380(.VSS(VSS),.VDD(VDD),.Y(g23201),.A(I30056));
  NOT NOT1_8381(.VSS(VSS),.VDD(VDD),.Y(I30059),.A(g22620));
  NOT NOT1_8382(.VSS(VSS),.VDD(VDD),.Y(g23202),.A(I30059));
  NOT NOT1_8383(.VSS(VSS),.VDD(VDD),.Y(I30062),.A(g22590));
  NOT NOT1_8384(.VSS(VSS),.VDD(VDD),.Y(g23203),.A(I30062));
  NOT NOT1_8385(.VSS(VSS),.VDD(VDD),.Y(I30065),.A(g22621));
  NOT NOT1_8386(.VSS(VSS),.VDD(VDD),.Y(g23204),.A(I30065));
  NOT NOT1_8387(.VSS(VSS),.VDD(VDD),.Y(I30068),.A(g22647));
  NOT NOT1_8388(.VSS(VSS),.VDD(VDD),.Y(g23205),.A(I30068));
  NOT NOT1_8389(.VSS(VSS),.VDD(VDD),.Y(I30071),.A(g22622));
  NOT NOT1_8390(.VSS(VSS),.VDD(VDD),.Y(g23206),.A(I30071));
  NOT NOT1_8391(.VSS(VSS),.VDD(VDD),.Y(I30074),.A(g22648));
  NOT NOT1_8392(.VSS(VSS),.VDD(VDD),.Y(g23207),.A(I30074));
  NOT NOT1_8393(.VSS(VSS),.VDD(VDD),.Y(I30077),.A(g22675));
  NOT NOT1_8394(.VSS(VSS),.VDD(VDD),.Y(g23208),.A(I30077));
  NOT NOT1_8395(.VSS(VSS),.VDD(VDD),.Y(I30080),.A(g22649));
  NOT NOT1_8396(.VSS(VSS),.VDD(VDD),.Y(g23209),.A(I30080));
  NOT NOT1_8397(.VSS(VSS),.VDD(VDD),.Y(I30083),.A(g22676));
  NOT NOT1_8398(.VSS(VSS),.VDD(VDD),.Y(g23210),.A(I30083));
  NOT NOT1_8399(.VSS(VSS),.VDD(VDD),.Y(I30086),.A(g22709));
  NOT NOT1_8400(.VSS(VSS),.VDD(VDD),.Y(g23211),.A(I30086));
  NOT NOT1_8401(.VSS(VSS),.VDD(VDD),.Y(I30089),.A(g22677));
  NOT NOT1_8402(.VSS(VSS),.VDD(VDD),.Y(g23212),.A(I30089));
  NOT NOT1_8403(.VSS(VSS),.VDD(VDD),.Y(I30092),.A(g22710));
  NOT NOT1_8404(.VSS(VSS),.VDD(VDD),.Y(g23213),.A(I30092));
  NOT NOT1_8405(.VSS(VSS),.VDD(VDD),.Y(I30095),.A(g22733));
  NOT NOT1_8406(.VSS(VSS),.VDD(VDD),.Y(g23214),.A(I30095));
  NOT NOT1_8407(.VSS(VSS),.VDD(VDD),.Y(I30098),.A(g22711));
  NOT NOT1_8408(.VSS(VSS),.VDD(VDD),.Y(g23215),.A(I30098));
  NOT NOT1_8409(.VSS(VSS),.VDD(VDD),.Y(I30101),.A(g22734));
  NOT NOT1_8410(.VSS(VSS),.VDD(VDD),.Y(g23216),.A(I30101));
  NOT NOT1_8411(.VSS(VSS),.VDD(VDD),.Y(I30104),.A(g22760));
  NOT NOT1_8412(.VSS(VSS),.VDD(VDD),.Y(g23217),.A(I30104));
  NOT NOT1_8413(.VSS(VSS),.VDD(VDD),.Y(I30107),.A(g22735));
  NOT NOT1_8414(.VSS(VSS),.VDD(VDD),.Y(g23218),.A(I30107));
  NOT NOT1_8415(.VSS(VSS),.VDD(VDD),.Y(I30110),.A(g22761));
  NOT NOT1_8416(.VSS(VSS),.VDD(VDD),.Y(g23219),.A(I30110));
  NOT NOT1_8417(.VSS(VSS),.VDD(VDD),.Y(I30113),.A(g22790));
  NOT NOT1_8418(.VSS(VSS),.VDD(VDD),.Y(g23220),.A(I30113));
  NOT NOT1_8419(.VSS(VSS),.VDD(VDD),.Y(I30116),.A(g22762));
  NOT NOT1_8420(.VSS(VSS),.VDD(VDD),.Y(g23221),.A(I30116));
  NOT NOT1_8421(.VSS(VSS),.VDD(VDD),.Y(I30119),.A(g22791));
  NOT NOT1_8422(.VSS(VSS),.VDD(VDD),.Y(g23222),.A(I30119));
  NOT NOT1_8423(.VSS(VSS),.VDD(VDD),.Y(I30122),.A(g22827));
  NOT NOT1_8424(.VSS(VSS),.VDD(VDD),.Y(g23223),.A(I30122));
  NOT NOT1_8425(.VSS(VSS),.VDD(VDD),.Y(I30125),.A(g22792));
  NOT NOT1_8426(.VSS(VSS),.VDD(VDD),.Y(g23224),.A(I30125));
  NOT NOT1_8427(.VSS(VSS),.VDD(VDD),.Y(I30128),.A(g22828));
  NOT NOT1_8428(.VSS(VSS),.VDD(VDD),.Y(g23225),.A(I30128));
  NOT NOT1_8429(.VSS(VSS),.VDD(VDD),.Y(I30131),.A(g22864));
  NOT NOT1_8430(.VSS(VSS),.VDD(VDD),.Y(g23226),.A(I30131));
  NOT NOT1_8431(.VSS(VSS),.VDD(VDD),.Y(I30134),.A(g22559));
  NOT NOT1_8432(.VSS(VSS),.VDD(VDD),.Y(g23227),.A(I30134));
  NOT NOT1_8433(.VSS(VSS),.VDD(VDD),.Y(I30137),.A(g22591));
  NOT NOT1_8434(.VSS(VSS),.VDD(VDD),.Y(g23228),.A(I30137));
  NOT NOT1_8435(.VSS(VSS),.VDD(VDD),.Y(I30140),.A(g22623));
  NOT NOT1_8436(.VSS(VSS),.VDD(VDD),.Y(g23229),.A(I30140));
  NOT NOT1_8437(.VSS(VSS),.VDD(VDD),.Y(I30143),.A(g22678));
  NOT NOT1_8438(.VSS(VSS),.VDD(VDD),.Y(g23230),.A(I30143));
  NOT NOT1_8439(.VSS(VSS),.VDD(VDD),.Y(I30146),.A(g22712));
  NOT NOT1_8440(.VSS(VSS),.VDD(VDD),.Y(g23231),.A(I30146));
  NOT NOT1_8441(.VSS(VSS),.VDD(VDD),.Y(I30149),.A(g22736));
  NOT NOT1_8442(.VSS(VSS),.VDD(VDD),.Y(g23232),.A(I30149));
  NOT NOT1_8443(.VSS(VSS),.VDD(VDD),.Y(I30152),.A(g22713));
  NOT NOT1_8444(.VSS(VSS),.VDD(VDD),.Y(g23233),.A(I30152));
  NOT NOT1_8445(.VSS(VSS),.VDD(VDD),.Y(I30155),.A(g22737));
  NOT NOT1_8446(.VSS(VSS),.VDD(VDD),.Y(g23234),.A(I30155));
  NOT NOT1_8447(.VSS(VSS),.VDD(VDD),.Y(I30158),.A(g22763));
  NOT NOT1_8448(.VSS(VSS),.VDD(VDD),.Y(g23235),.A(I30158));
  NOT NOT1_8449(.VSS(VSS),.VDD(VDD),.Y(I30161),.A(g22133));
  NOT NOT1_8450(.VSS(VSS),.VDD(VDD),.Y(g23236),.A(I30161));
  NOT NOT1_8451(.VSS(VSS),.VDD(VDD),.Y(I30164),.A(g22655));
  NOT NOT1_8452(.VSS(VSS),.VDD(VDD),.Y(g23237),.A(I30164));
  NOT NOT1_8453(.VSS(VSS),.VDD(VDD),.Y(I30167),.A(g22598));
  NOT NOT1_8454(.VSS(VSS),.VDD(VDD),.Y(g23238),.A(I30167));
  NOT NOT1_8455(.VSS(VSS),.VDD(VDD),.Y(I30170),.A(g22626));
  NOT NOT1_8456(.VSS(VSS),.VDD(VDD),.Y(g23239),.A(I30170));
  NOT NOT1_8457(.VSS(VSS),.VDD(VDD),.Y(I30173),.A(g22656));
  NOT NOT1_8458(.VSS(VSS),.VDD(VDD),.Y(g23240),.A(I30173));
  NOT NOT1_8459(.VSS(VSS),.VDD(VDD),.Y(I30176),.A(g22627));
  NOT NOT1_8460(.VSS(VSS),.VDD(VDD),.Y(g23241),.A(I30176));
  NOT NOT1_8461(.VSS(VSS),.VDD(VDD),.Y(I30179),.A(g22657));
  NOT NOT1_8462(.VSS(VSS),.VDD(VDD),.Y(g23242),.A(I30179));
  NOT NOT1_8463(.VSS(VSS),.VDD(VDD),.Y(I30182),.A(g22683));
  NOT NOT1_8464(.VSS(VSS),.VDD(VDD),.Y(g23243),.A(I30182));
  NOT NOT1_8465(.VSS(VSS),.VDD(VDD),.Y(I30185),.A(g22658));
  NOT NOT1_8466(.VSS(VSS),.VDD(VDD),.Y(g23244),.A(I30185));
  NOT NOT1_8467(.VSS(VSS),.VDD(VDD),.Y(I30188),.A(g22684));
  NOT NOT1_8468(.VSS(VSS),.VDD(VDD),.Y(g23245),.A(I30188));
  NOT NOT1_8469(.VSS(VSS),.VDD(VDD),.Y(I30191),.A(g22715));
  NOT NOT1_8470(.VSS(VSS),.VDD(VDD),.Y(g23246),.A(I30191));
  NOT NOT1_8471(.VSS(VSS),.VDD(VDD),.Y(I30194),.A(g22685));
  NOT NOT1_8472(.VSS(VSS),.VDD(VDD),.Y(g23247),.A(I30194));
  NOT NOT1_8473(.VSS(VSS),.VDD(VDD),.Y(I30197),.A(g22716));
  NOT NOT1_8474(.VSS(VSS),.VDD(VDD),.Y(g23248),.A(I30197));
  NOT NOT1_8475(.VSS(VSS),.VDD(VDD),.Y(I30200),.A(g22740));
  NOT NOT1_8476(.VSS(VSS),.VDD(VDD),.Y(g23249),.A(I30200));
  NOT NOT1_8477(.VSS(VSS),.VDD(VDD),.Y(I30203),.A(g22717));
  NOT NOT1_8478(.VSS(VSS),.VDD(VDD),.Y(g23250),.A(I30203));
  NOT NOT1_8479(.VSS(VSS),.VDD(VDD),.Y(I30206),.A(g22741));
  NOT NOT1_8480(.VSS(VSS),.VDD(VDD),.Y(g23251),.A(I30206));
  NOT NOT1_8481(.VSS(VSS),.VDD(VDD),.Y(I30209),.A(g22765));
  NOT NOT1_8482(.VSS(VSS),.VDD(VDD),.Y(g23252),.A(I30209));
  NOT NOT1_8483(.VSS(VSS),.VDD(VDD),.Y(I30212),.A(g22742));
  NOT NOT1_8484(.VSS(VSS),.VDD(VDD),.Y(g23253),.A(I30212));
  NOT NOT1_8485(.VSS(VSS),.VDD(VDD),.Y(I30215),.A(g22766));
  NOT NOT1_8486(.VSS(VSS),.VDD(VDD),.Y(g23254),.A(I30215));
  NOT NOT1_8487(.VSS(VSS),.VDD(VDD),.Y(I30218),.A(g22794));
  NOT NOT1_8488(.VSS(VSS),.VDD(VDD),.Y(g23255),.A(I30218));
  NOT NOT1_8489(.VSS(VSS),.VDD(VDD),.Y(I30221),.A(g22767));
  NOT NOT1_8490(.VSS(VSS),.VDD(VDD),.Y(g23256),.A(I30221));
  NOT NOT1_8491(.VSS(VSS),.VDD(VDD),.Y(I30224),.A(g22795));
  NOT NOT1_8492(.VSS(VSS),.VDD(VDD),.Y(g23257),.A(I30224));
  NOT NOT1_8493(.VSS(VSS),.VDD(VDD),.Y(I30227),.A(g22832));
  NOT NOT1_8494(.VSS(VSS),.VDD(VDD),.Y(g23258),.A(I30227));
  NOT NOT1_8495(.VSS(VSS),.VDD(VDD),.Y(I30230),.A(g22796));
  NOT NOT1_8496(.VSS(VSS),.VDD(VDD),.Y(g23259),.A(I30230));
  NOT NOT1_8497(.VSS(VSS),.VDD(VDD),.Y(I30233),.A(g22833));
  NOT NOT1_8498(.VSS(VSS),.VDD(VDD),.Y(g23260),.A(I30233));
  NOT NOT1_8499(.VSS(VSS),.VDD(VDD),.Y(I30236),.A(g22866));
  NOT NOT1_8500(.VSS(VSS),.VDD(VDD),.Y(g23261),.A(I30236));
  NOT NOT1_8501(.VSS(VSS),.VDD(VDD),.Y(I30239),.A(g22834));
  NOT NOT1_8502(.VSS(VSS),.VDD(VDD),.Y(g23262),.A(I30239));
  NOT NOT1_8503(.VSS(VSS),.VDD(VDD),.Y(I30242),.A(g22867));
  NOT NOT1_8504(.VSS(VSS),.VDD(VDD),.Y(g23263),.A(I30242));
  NOT NOT1_8505(.VSS(VSS),.VDD(VDD),.Y(I30245),.A(g22899));
  NOT NOT1_8506(.VSS(VSS),.VDD(VDD),.Y(g23264),.A(I30245));
  NOT NOT1_8507(.VSS(VSS),.VDD(VDD),.Y(I30248),.A(g22599));
  NOT NOT1_8508(.VSS(VSS),.VDD(VDD),.Y(g23265),.A(I30248));
  NOT NOT1_8509(.VSS(VSS),.VDD(VDD),.Y(I30251),.A(g22628));
  NOT NOT1_8510(.VSS(VSS),.VDD(VDD),.Y(g23266),.A(I30251));
  NOT NOT1_8511(.VSS(VSS),.VDD(VDD),.Y(I30254),.A(g22659));
  NOT NOT1_8512(.VSS(VSS),.VDD(VDD),.Y(g23267),.A(I30254));
  NOT NOT1_8513(.VSS(VSS),.VDD(VDD),.Y(I30257),.A(g22718));
  NOT NOT1_8514(.VSS(VSS),.VDD(VDD),.Y(g23268),.A(I30257));
  NOT NOT1_8515(.VSS(VSS),.VDD(VDD),.Y(I30260),.A(g22743));
  NOT NOT1_8516(.VSS(VSS),.VDD(VDD),.Y(g23269),.A(I30260));
  NOT NOT1_8517(.VSS(VSS),.VDD(VDD),.Y(I30263),.A(g22768));
  NOT NOT1_8518(.VSS(VSS),.VDD(VDD),.Y(g23270),.A(I30263));
  NOT NOT1_8519(.VSS(VSS),.VDD(VDD),.Y(I30266),.A(g22744));
  NOT NOT1_8520(.VSS(VSS),.VDD(VDD),.Y(g23271),.A(I30266));
  NOT NOT1_8521(.VSS(VSS),.VDD(VDD),.Y(I30269),.A(g22769));
  NOT NOT1_8522(.VSS(VSS),.VDD(VDD),.Y(g23272),.A(I30269));
  NOT NOT1_8523(.VSS(VSS),.VDD(VDD),.Y(I30272),.A(g22797));
  NOT NOT1_8524(.VSS(VSS),.VDD(VDD),.Y(g23273),.A(I30272));
  NOT NOT1_8525(.VSS(VSS),.VDD(VDD),.Y(I30275),.A(g22156));
  NOT NOT1_8526(.VSS(VSS),.VDD(VDD),.Y(g23274),.A(I30275));
  NOT NOT1_8527(.VSS(VSS),.VDD(VDD),.Y(I30278),.A(g22691));
  NOT NOT1_8528(.VSS(VSS),.VDD(VDD),.Y(g23275),.A(I30278));
  NOT NOT1_8529(.VSS(VSS),.VDD(VDD),.Y(I30281),.A(g22635));
  NOT NOT1_8530(.VSS(VSS),.VDD(VDD),.Y(g23276),.A(I30281));
  NOT NOT1_8531(.VSS(VSS),.VDD(VDD),.Y(I30284),.A(g22662));
  NOT NOT1_8532(.VSS(VSS),.VDD(VDD),.Y(g23277),.A(I30284));
  NOT NOT1_8533(.VSS(VSS),.VDD(VDD),.Y(I30287),.A(g22692));
  NOT NOT1_8534(.VSS(VSS),.VDD(VDD),.Y(g23278),.A(I30287));
  NOT NOT1_8535(.VSS(VSS),.VDD(VDD),.Y(I30290),.A(g22663));
  NOT NOT1_8536(.VSS(VSS),.VDD(VDD),.Y(g23279),.A(I30290));
  NOT NOT1_8537(.VSS(VSS),.VDD(VDD),.Y(I30293),.A(g22693));
  NOT NOT1_8538(.VSS(VSS),.VDD(VDD),.Y(g23280),.A(I30293));
  NOT NOT1_8539(.VSS(VSS),.VDD(VDD),.Y(I30296),.A(g22723));
  NOT NOT1_8540(.VSS(VSS),.VDD(VDD),.Y(g23281),.A(I30296));
  NOT NOT1_8541(.VSS(VSS),.VDD(VDD),.Y(I30299),.A(g22694));
  NOT NOT1_8542(.VSS(VSS),.VDD(VDD),.Y(g23282),.A(I30299));
  NOT NOT1_8543(.VSS(VSS),.VDD(VDD),.Y(I30302),.A(g22724));
  NOT NOT1_8544(.VSS(VSS),.VDD(VDD),.Y(g23283),.A(I30302));
  NOT NOT1_8545(.VSS(VSS),.VDD(VDD),.Y(I30305),.A(g22746));
  NOT NOT1_8546(.VSS(VSS),.VDD(VDD),.Y(g23284),.A(I30305));
  NOT NOT1_8547(.VSS(VSS),.VDD(VDD),.Y(I30308),.A(g22725));
  NOT NOT1_8548(.VSS(VSS),.VDD(VDD),.Y(g23285),.A(I30308));
  NOT NOT1_8549(.VSS(VSS),.VDD(VDD),.Y(I30311),.A(g22747));
  NOT NOT1_8550(.VSS(VSS),.VDD(VDD),.Y(g23286),.A(I30311));
  NOT NOT1_8551(.VSS(VSS),.VDD(VDD),.Y(I30314),.A(g22772));
  NOT NOT1_8552(.VSS(VSS),.VDD(VDD),.Y(g23287),.A(I30314));
  NOT NOT1_8553(.VSS(VSS),.VDD(VDD),.Y(I30317),.A(g22748));
  NOT NOT1_8554(.VSS(VSS),.VDD(VDD),.Y(g23288),.A(I30317));
  NOT NOT1_8555(.VSS(VSS),.VDD(VDD),.Y(I30320),.A(g22773));
  NOT NOT1_8556(.VSS(VSS),.VDD(VDD),.Y(g23289),.A(I30320));
  NOT NOT1_8557(.VSS(VSS),.VDD(VDD),.Y(I30323),.A(g22799));
  NOT NOT1_8558(.VSS(VSS),.VDD(VDD),.Y(g23290),.A(I30323));
  NOT NOT1_8559(.VSS(VSS),.VDD(VDD),.Y(I30326),.A(g22774));
  NOT NOT1_8560(.VSS(VSS),.VDD(VDD),.Y(g23291),.A(I30326));
  NOT NOT1_8561(.VSS(VSS),.VDD(VDD),.Y(I30329),.A(g22800));
  NOT NOT1_8562(.VSS(VSS),.VDD(VDD),.Y(g23292),.A(I30329));
  NOT NOT1_8563(.VSS(VSS),.VDD(VDD),.Y(I30332),.A(g22836));
  NOT NOT1_8564(.VSS(VSS),.VDD(VDD),.Y(g23293),.A(I30332));
  NOT NOT1_8565(.VSS(VSS),.VDD(VDD),.Y(I30335),.A(g22801));
  NOT NOT1_8566(.VSS(VSS),.VDD(VDD),.Y(g23294),.A(I30335));
  NOT NOT1_8567(.VSS(VSS),.VDD(VDD),.Y(I30338),.A(g22837));
  NOT NOT1_8568(.VSS(VSS),.VDD(VDD),.Y(g23295),.A(I30338));
  NOT NOT1_8569(.VSS(VSS),.VDD(VDD),.Y(I30341),.A(g22871));
  NOT NOT1_8570(.VSS(VSS),.VDD(VDD),.Y(g23296),.A(I30341));
  NOT NOT1_8571(.VSS(VSS),.VDD(VDD),.Y(I30344),.A(g22838));
  NOT NOT1_8572(.VSS(VSS),.VDD(VDD),.Y(g23297),.A(I30344));
  NOT NOT1_8573(.VSS(VSS),.VDD(VDD),.Y(I30347),.A(g22872));
  NOT NOT1_8574(.VSS(VSS),.VDD(VDD),.Y(g23298),.A(I30347));
  NOT NOT1_8575(.VSS(VSS),.VDD(VDD),.Y(I30350),.A(g22901));
  NOT NOT1_8576(.VSS(VSS),.VDD(VDD),.Y(g23299),.A(I30350));
  NOT NOT1_8577(.VSS(VSS),.VDD(VDD),.Y(I30353),.A(g22873));
  NOT NOT1_8578(.VSS(VSS),.VDD(VDD),.Y(g23300),.A(I30353));
  NOT NOT1_8579(.VSS(VSS),.VDD(VDD),.Y(I30356),.A(g22902));
  NOT NOT1_8580(.VSS(VSS),.VDD(VDD),.Y(g23301),.A(I30356));
  NOT NOT1_8581(.VSS(VSS),.VDD(VDD),.Y(I30359),.A(g22934));
  NOT NOT1_8582(.VSS(VSS),.VDD(VDD),.Y(g23302),.A(I30359));
  NOT NOT1_8583(.VSS(VSS),.VDD(VDD),.Y(I30362),.A(g22636));
  NOT NOT1_8584(.VSS(VSS),.VDD(VDD),.Y(g23303),.A(I30362));
  NOT NOT1_8585(.VSS(VSS),.VDD(VDD),.Y(I30365),.A(g22664));
  NOT NOT1_8586(.VSS(VSS),.VDD(VDD),.Y(g23304),.A(I30365));
  NOT NOT1_8587(.VSS(VSS),.VDD(VDD),.Y(I30368),.A(g22695));
  NOT NOT1_8588(.VSS(VSS),.VDD(VDD),.Y(g23305),.A(I30368));
  NOT NOT1_8589(.VSS(VSS),.VDD(VDD),.Y(I30371),.A(g22749));
  NOT NOT1_8590(.VSS(VSS),.VDD(VDD),.Y(g23306),.A(I30371));
  NOT NOT1_8591(.VSS(VSS),.VDD(VDD),.Y(I30374),.A(g22775));
  NOT NOT1_8592(.VSS(VSS),.VDD(VDD),.Y(g23307),.A(I30374));
  NOT NOT1_8593(.VSS(VSS),.VDD(VDD),.Y(I30377),.A(g22802));
  NOT NOT1_8594(.VSS(VSS),.VDD(VDD),.Y(g23308),.A(I30377));
  NOT NOT1_8595(.VSS(VSS),.VDD(VDD),.Y(I30380),.A(g22776));
  NOT NOT1_8596(.VSS(VSS),.VDD(VDD),.Y(g23309),.A(I30380));
  NOT NOT1_8597(.VSS(VSS),.VDD(VDD),.Y(I30383),.A(g22803));
  NOT NOT1_8598(.VSS(VSS),.VDD(VDD),.Y(g23310),.A(I30383));
  NOT NOT1_8599(.VSS(VSS),.VDD(VDD),.Y(I30386),.A(g22839));
  NOT NOT1_8600(.VSS(VSS),.VDD(VDD),.Y(g23311),.A(I30386));
  NOT NOT1_8601(.VSS(VSS),.VDD(VDD),.Y(I30389),.A(g22225));
  NOT NOT1_8602(.VSS(VSS),.VDD(VDD),.Y(g23312),.A(I30389));
  NOT NOT1_8603(.VSS(VSS),.VDD(VDD),.Y(I30392),.A(g22226));
  NOT NOT1_8604(.VSS(VSS),.VDD(VDD),.Y(g23313),.A(I30392));
  NOT NOT1_8605(.VSS(VSS),.VDD(VDD),.Y(I30395),.A(g22253));
  NOT NOT1_8606(.VSS(VSS),.VDD(VDD),.Y(g23314),.A(I30395));
  NOT NOT1_8607(.VSS(VSS),.VDD(VDD),.Y(I30398),.A(g22840));
  NOT NOT1_8608(.VSS(VSS),.VDD(VDD),.Y(g23315),.A(I30398));
  NOT NOT1_8609(.VSS(VSS),.VDD(VDD),.Y(I30401),.A(g22444));
  NOT NOT1_8610(.VSS(VSS),.VDD(VDD),.Y(g23316),.A(I30401));
  NOT NOT1_8611(.VSS(VSS),.VDD(VDD),.Y(I30404),.A(g22948));
  NOT NOT1_8612(.VSS(VSS),.VDD(VDD),.Y(g23317),.A(I30404));
  NOT NOT1_8613(.VSS(VSS),.VDD(VDD),.Y(I30407),.A(g22970));
  NOT NOT1_8614(.VSS(VSS),.VDD(VDD),.Y(g23318),.A(I30407));
  NOT NOT1_8615(.VSS(VSS),.VDD(VDD),.Y(g23403),.A(g23052));
  NOT NOT1_8616(.VSS(VSS),.VDD(VDD),.Y(g23410),.A(g23071));
  NOT NOT1_8617(.VSS(VSS),.VDD(VDD),.Y(g23415),.A(g23084));
  NOT NOT1_8618(.VSS(VSS),.VDD(VDD),.Y(g23420),.A(g23089));
  NOT NOT1_8619(.VSS(VSS),.VDD(VDD),.Y(g23424),.A(g23100));
  NOT NOT1_8620(.VSS(VSS),.VDD(VDD),.Y(g23429),.A(g23107));
  NOT NOT1_8621(.VSS(VSS),.VDD(VDD),.Y(g23435),.A(g23120));
  NOT NOT1_8622(.VSS(VSS),.VDD(VDD),.Y(I30467),.A(g23000));
  NOT NOT1_8623(.VSS(VSS),.VDD(VDD),.Y(g23438),.A(I30467));
  NOT NOT1_8624(.VSS(VSS),.VDD(VDD),.Y(I30470),.A(g23117));
  NOT NOT1_8625(.VSS(VSS),.VDD(VDD),.Y(g23439),.A(I30470));
  NOT NOT1_8626(.VSS(VSS),.VDD(VDD),.Y(g23441),.A(g23129));
  NOT NOT1_8627(.VSS(VSS),.VDD(VDD),.Y(g23444),.A(g22945));
  NOT NOT1_8628(.VSS(VSS),.VDD(VDD),.Y(I30476),.A(g22876));
  NOT NOT1_8629(.VSS(VSS),.VDD(VDD),.Y(g23448),.A(I30476));
  NOT NOT1_8630(.VSS(VSS),.VDD(VDD),.Y(I30480),.A(g23014));
  NOT NOT1_8631(.VSS(VSS),.VDD(VDD),.Y(g23452),.A(I30480));
  NOT NOT1_8632(.VSS(VSS),.VDD(VDD),.Y(I30483),.A(g23126));
  NOT NOT1_8633(.VSS(VSS),.VDD(VDD),.Y(g23453),.A(I30483));
  NOT NOT1_8634(.VSS(VSS),.VDD(VDD),.Y(I30486),.A(g23022));
  NOT NOT1_8635(.VSS(VSS),.VDD(VDD),.Y(g23454),.A(I30486));
  NOT NOT1_8636(.VSS(VSS),.VDD(VDD),.Y(I30489),.A(g22911));
  NOT NOT1_8637(.VSS(VSS),.VDD(VDD),.Y(g23455),.A(I30489));
  NOT NOT1_8638(.VSS(VSS),.VDD(VDD),.Y(I30493),.A(g23030));
  NOT NOT1_8639(.VSS(VSS),.VDD(VDD),.Y(g23459),.A(I30493));
  NOT NOT1_8640(.VSS(VSS),.VDD(VDD),.Y(I30496),.A(g23137));
  NOT NOT1_8641(.VSS(VSS),.VDD(VDD),.Y(g23460),.A(I30496));
  NOT NOT1_8642(.VSS(VSS),.VDD(VDD),.Y(I30501),.A(g23039));
  NOT NOT1_8643(.VSS(VSS),.VDD(VDD),.Y(g23463),.A(I30501));
  NOT NOT1_8644(.VSS(VSS),.VDD(VDD),.Y(I30504),.A(g22936));
  NOT NOT1_8645(.VSS(VSS),.VDD(VDD),.Y(g23464),.A(I30504));
  NOT NOT1_8646(.VSS(VSS),.VDD(VDD),.Y(I30508),.A(g23047));
  NOT NOT1_8647(.VSS(VSS),.VDD(VDD),.Y(g23468),.A(I30508));
  NOT NOT1_8648(.VSS(VSS),.VDD(VDD),.Y(I30511),.A(g21970));
  NOT NOT1_8649(.VSS(VSS),.VDD(VDD),.Y(g23469),.A(I30511));
  NOT NOT1_8650(.VSS(VSS),.VDD(VDD),.Y(g23470),.A(g22188));
  NOT NOT1_8651(.VSS(VSS),.VDD(VDD),.Y(I30516),.A(g23058));
  NOT NOT1_8652(.VSS(VSS),.VDD(VDD),.Y(g23472),.A(I30516));
  NOT NOT1_8653(.VSS(VSS),.VDD(VDD),.Y(I30519),.A(g22942));
  NOT NOT1_8654(.VSS(VSS),.VDD(VDD),.Y(g23473),.A(I30519));
  NOT NOT1_8655(.VSS(VSS),.VDD(VDD),.Y(I30525),.A(g23067));
  NOT NOT1_8656(.VSS(VSS),.VDD(VDD),.Y(g23481),.A(I30525));
  NOT NOT1_8657(.VSS(VSS),.VDD(VDD),.Y(g23482),.A(g22197));
  NOT NOT1_8658(.VSS(VSS),.VDD(VDD),.Y(I30531),.A(g23076));
  NOT NOT1_8659(.VSS(VSS),.VDD(VDD),.Y(g23485),.A(I30531));
  NOT NOT1_8660(.VSS(VSS),.VDD(VDD),.Y(I30536),.A(g23081));
  NOT NOT1_8661(.VSS(VSS),.VDD(VDD),.Y(g23492),.A(I30536));
  NOT NOT1_8662(.VSS(VSS),.VDD(VDD),.Y(g23493),.A(g22203));
  NOT NOT1_8663(.VSS(VSS),.VDD(VDD),.Y(I30544),.A(g23092));
  NOT NOT1_8664(.VSS(VSS),.VDD(VDD),.Y(g23500),.A(I30544));
  NOT NOT1_8665(.VSS(VSS),.VDD(VDD),.Y(I30547),.A(g23093));
  NOT NOT1_8666(.VSS(VSS),.VDD(VDD),.Y(g23501),.A(I30547));
  NOT NOT1_8667(.VSS(VSS),.VDD(VDD),.Y(I30552),.A(g23097));
  NOT NOT1_8668(.VSS(VSS),.VDD(VDD),.Y(g23508),.A(I30552));
  NOT NOT1_8669(.VSS(VSS),.VDD(VDD),.Y(g23509),.A(g22209));
  NOT NOT1_8670(.VSS(VSS),.VDD(VDD),.Y(I30560),.A(g23110));
  NOT NOT1_8671(.VSS(VSS),.VDD(VDD),.Y(g23516),.A(I30560));
  NOT NOT1_8672(.VSS(VSS),.VDD(VDD),.Y(I30563),.A(g23111));
  NOT NOT1_8673(.VSS(VSS),.VDD(VDD),.Y(g23517),.A(I30563));
  NOT NOT1_8674(.VSS(VSS),.VDD(VDD),.Y(I30568),.A(g23114));
  NOT NOT1_8675(.VSS(VSS),.VDD(VDD),.Y(g23524),.A(I30568));
  NOT NOT1_8676(.VSS(VSS),.VDD(VDD),.Y(I30575),.A(g23123));
  NOT NOT1_8677(.VSS(VSS),.VDD(VDD),.Y(g23531),.A(I30575));
  NOT NOT1_8678(.VSS(VSS),.VDD(VDD),.Y(I30578),.A(g23124));
  NOT NOT1_8679(.VSS(VSS),.VDD(VDD),.Y(g23532),.A(I30578));
  NOT NOT1_8680(.VSS(VSS),.VDD(VDD),.Y(I30586),.A(g23132));
  NOT NOT1_8681(.VSS(VSS),.VDD(VDD),.Y(g23542),.A(I30586));
  NOT NOT1_8682(.VSS(VSS),.VDD(VDD),.Y(I30589),.A(g23133));
  NOT NOT1_8683(.VSS(VSS),.VDD(VDD),.Y(g23543),.A(I30589));
  NOT NOT1_8684(.VSS(VSS),.VDD(VDD),.Y(I30594),.A(g22025));
  NOT NOT1_8685(.VSS(VSS),.VDD(VDD),.Y(g23546),.A(I30594));
  NOT NOT1_8686(.VSS(VSS),.VDD(VDD),.Y(I30598),.A(g22027));
  NOT NOT1_8687(.VSS(VSS),.VDD(VDD),.Y(g23548),.A(I30598));
  NOT NOT1_8688(.VSS(VSS),.VDD(VDD),.Y(I30601),.A(g22028));
  NOT NOT1_8689(.VSS(VSS),.VDD(VDD),.Y(g23549),.A(I30601));
  NOT NOT1_8690(.VSS(VSS),.VDD(VDD),.Y(I30607),.A(g22029));
  NOT NOT1_8691(.VSS(VSS),.VDD(VDD),.Y(g23553),.A(I30607));
  NOT NOT1_8692(.VSS(VSS),.VDD(VDD),.Y(I30611),.A(g22030));
  NOT NOT1_8693(.VSS(VSS),.VDD(VDD),.Y(g23555),.A(I30611));
  NOT NOT1_8694(.VSS(VSS),.VDD(VDD),.Y(I30614),.A(g22031));
  NOT NOT1_8695(.VSS(VSS),.VDD(VDD),.Y(g23556),.A(I30614));
  NOT NOT1_8696(.VSS(VSS),.VDD(VDD),.Y(I30617),.A(g22032));
  NOT NOT1_8697(.VSS(VSS),.VDD(VDD),.Y(g23557),.A(I30617));
  NOT NOT1_8698(.VSS(VSS),.VDD(VDD),.Y(I30623),.A(g22033));
  NOT NOT1_8699(.VSS(VSS),.VDD(VDD),.Y(g23561),.A(I30623));
  NOT NOT1_8700(.VSS(VSS),.VDD(VDD),.Y(I30626),.A(g22034));
  NOT NOT1_8701(.VSS(VSS),.VDD(VDD),.Y(g23562),.A(I30626));
  NOT NOT1_8702(.VSS(VSS),.VDD(VDD),.Y(I30632),.A(g22035));
  NOT NOT1_8703(.VSS(VSS),.VDD(VDD),.Y(g23566),.A(I30632));
  NOT NOT1_8704(.VSS(VSS),.VDD(VDD),.Y(I30636),.A(g22037));
  NOT NOT1_8705(.VSS(VSS),.VDD(VDD),.Y(g23568),.A(I30636));
  NOT NOT1_8706(.VSS(VSS),.VDD(VDD),.Y(I30639),.A(g22038));
  NOT NOT1_8707(.VSS(VSS),.VDD(VDD),.Y(g23569),.A(I30639));
  NOT NOT1_8708(.VSS(VSS),.VDD(VDD),.Y(I30642),.A(g22039));
  NOT NOT1_8709(.VSS(VSS),.VDD(VDD),.Y(g23570),.A(I30642));
  NOT NOT1_8710(.VSS(VSS),.VDD(VDD),.Y(I30648),.A(g22040));
  NOT NOT1_8711(.VSS(VSS),.VDD(VDD),.Y(g23574),.A(I30648));
  NOT NOT1_8712(.VSS(VSS),.VDD(VDD),.Y(I30651),.A(g22041));
  NOT NOT1_8713(.VSS(VSS),.VDD(VDD),.Y(g23575),.A(I30651));
  NOT NOT1_8714(.VSS(VSS),.VDD(VDD),.Y(I30654),.A(g22042));
  NOT NOT1_8715(.VSS(VSS),.VDD(VDD),.Y(g23576),.A(I30654));
  NOT NOT1_8716(.VSS(VSS),.VDD(VDD),.Y(I30660),.A(g22043));
  NOT NOT1_8717(.VSS(VSS),.VDD(VDD),.Y(g23580),.A(I30660));
  NOT NOT1_8718(.VSS(VSS),.VDD(VDD),.Y(I30663),.A(g22044));
  NOT NOT1_8719(.VSS(VSS),.VDD(VDD),.Y(g23581),.A(I30663));
  NOT NOT1_8720(.VSS(VSS),.VDD(VDD),.Y(I30669),.A(g22045));
  NOT NOT1_8721(.VSS(VSS),.VDD(VDD),.Y(g23585),.A(I30669));
  NOT NOT1_8722(.VSS(VSS),.VDD(VDD),.Y(I30673),.A(g22047));
  NOT NOT1_8723(.VSS(VSS),.VDD(VDD),.Y(g23587),.A(I30673));
  NOT NOT1_8724(.VSS(VSS),.VDD(VDD),.Y(I30676),.A(g22048));
  NOT NOT1_8725(.VSS(VSS),.VDD(VDD),.Y(g23588),.A(I30676));
  NOT NOT1_8726(.VSS(VSS),.VDD(VDD),.Y(I30679),.A(g22049));
  NOT NOT1_8727(.VSS(VSS),.VDD(VDD),.Y(g23589),.A(I30679));
  NOT NOT1_8728(.VSS(VSS),.VDD(VDD),.Y(I30686),.A(g23136));
  NOT NOT1_8729(.VSS(VSS),.VDD(VDD),.Y(g23594),.A(I30686));
  NOT NOT1_8730(.VSS(VSS),.VDD(VDD),.Y(I30689),.A(g22054));
  NOT NOT1_8731(.VSS(VSS),.VDD(VDD),.Y(g23595),.A(I30689));
  NOT NOT1_8732(.VSS(VSS),.VDD(VDD),.Y(I30692),.A(g22055));
  NOT NOT1_8733(.VSS(VSS),.VDD(VDD),.Y(g23596),.A(I30692));
  NOT NOT1_8734(.VSS(VSS),.VDD(VDD),.Y(I30695),.A(g22056));
  NOT NOT1_8735(.VSS(VSS),.VDD(VDD),.Y(g23597),.A(I30695));
  NOT NOT1_8736(.VSS(VSS),.VDD(VDD),.Y(I30701),.A(g22057));
  NOT NOT1_8737(.VSS(VSS),.VDD(VDD),.Y(g23601),.A(I30701));
  NOT NOT1_8738(.VSS(VSS),.VDD(VDD),.Y(I30704),.A(g22058));
  NOT NOT1_8739(.VSS(VSS),.VDD(VDD),.Y(g23602),.A(I30704));
  NOT NOT1_8740(.VSS(VSS),.VDD(VDD),.Y(I30707),.A(g22059));
  NOT NOT1_8741(.VSS(VSS),.VDD(VDD),.Y(g23603),.A(I30707));
  NOT NOT1_8742(.VSS(VSS),.VDD(VDD),.Y(I30713),.A(g22060));
  NOT NOT1_8743(.VSS(VSS),.VDD(VDD),.Y(g23607),.A(I30713));
  NOT NOT1_8744(.VSS(VSS),.VDD(VDD),.Y(I30716),.A(g22061));
  NOT NOT1_8745(.VSS(VSS),.VDD(VDD),.Y(g23608),.A(I30716));
  NOT NOT1_8746(.VSS(VSS),.VDD(VDD),.Y(I30722),.A(g22063));
  NOT NOT1_8747(.VSS(VSS),.VDD(VDD),.Y(g23612),.A(I30722));
  NOT NOT1_8748(.VSS(VSS),.VDD(VDD),.Y(I30725),.A(g22064));
  NOT NOT1_8749(.VSS(VSS),.VDD(VDD),.Y(g23613),.A(I30725));
  NOT NOT1_8750(.VSS(VSS),.VDD(VDD),.Y(I30728),.A(g22065));
  NOT NOT1_8751(.VSS(VSS),.VDD(VDD),.Y(g23614),.A(I30728));
  NOT NOT1_8752(.VSS(VSS),.VDD(VDD),.Y(I30735),.A(g22066));
  NOT NOT1_8753(.VSS(VSS),.VDD(VDD),.Y(g23619),.A(I30735));
  NOT NOT1_8754(.VSS(VSS),.VDD(VDD),.Y(I30738),.A(g22067));
  NOT NOT1_8755(.VSS(VSS),.VDD(VDD),.Y(g23620),.A(I30738));
  NOT NOT1_8756(.VSS(VSS),.VDD(VDD),.Y(I30741),.A(g22068));
  NOT NOT1_8757(.VSS(VSS),.VDD(VDD),.Y(g23621),.A(I30741));
  NOT NOT1_8758(.VSS(VSS),.VDD(VDD),.Y(I30748),.A(g21969));
  NOT NOT1_8759(.VSS(VSS),.VDD(VDD),.Y(g23626),.A(I30748));
  NOT NOT1_8760(.VSS(VSS),.VDD(VDD),.Y(I30751),.A(g22073));
  NOT NOT1_8761(.VSS(VSS),.VDD(VDD),.Y(g23627),.A(I30751));
  NOT NOT1_8762(.VSS(VSS),.VDD(VDD),.Y(I30754),.A(g22074));
  NOT NOT1_8763(.VSS(VSS),.VDD(VDD),.Y(g23628),.A(I30754));
  NOT NOT1_8764(.VSS(VSS),.VDD(VDD),.Y(I30757),.A(g22075));
  NOT NOT1_8765(.VSS(VSS),.VDD(VDD),.Y(g23629),.A(I30757));
  NOT NOT1_8766(.VSS(VSS),.VDD(VDD),.Y(I30763),.A(g22076));
  NOT NOT1_8767(.VSS(VSS),.VDD(VDD),.Y(g23633),.A(I30763));
  NOT NOT1_8768(.VSS(VSS),.VDD(VDD),.Y(I30766),.A(g22077));
  NOT NOT1_8769(.VSS(VSS),.VDD(VDD),.Y(g23634),.A(I30766));
  NOT NOT1_8770(.VSS(VSS),.VDD(VDD),.Y(I30769),.A(g22078));
  NOT NOT1_8771(.VSS(VSS),.VDD(VDD),.Y(g23635),.A(I30769));
  NOT NOT1_8772(.VSS(VSS),.VDD(VDD),.Y(I30776),.A(g22079));
  NOT NOT1_8773(.VSS(VSS),.VDD(VDD),.Y(g23640),.A(I30776));
  NOT NOT1_8774(.VSS(VSS),.VDD(VDD),.Y(I30779),.A(g22080));
  NOT NOT1_8775(.VSS(VSS),.VDD(VDD),.Y(g23641),.A(I30779));
  NOT NOT1_8776(.VSS(VSS),.VDD(VDD),.Y(I30782),.A(g22081));
  NOT NOT1_8777(.VSS(VSS),.VDD(VDD),.Y(g23642),.A(I30782));
  NOT NOT1_8778(.VSS(VSS),.VDD(VDD),.Y(I30786),.A(g22454));
  NOT NOT1_8779(.VSS(VSS),.VDD(VDD),.Y(g23644),.A(I30786));
  NOT NOT1_8780(.VSS(VSS),.VDD(VDD),.Y(I30797),.A(g22087));
  NOT NOT1_8781(.VSS(VSS),.VDD(VDD),.Y(g23661),.A(I30797));
  NOT NOT1_8782(.VSS(VSS),.VDD(VDD),.Y(I30800),.A(g22088));
  NOT NOT1_8783(.VSS(VSS),.VDD(VDD),.Y(g23662),.A(I30800));
  NOT NOT1_8784(.VSS(VSS),.VDD(VDD),.Y(I30803),.A(g22089));
  NOT NOT1_8785(.VSS(VSS),.VDD(VDD),.Y(g23663),.A(I30803));
  NOT NOT1_8786(.VSS(VSS),.VDD(VDD),.Y(I30810),.A(g22090));
  NOT NOT1_8787(.VSS(VSS),.VDD(VDD),.Y(g23668),.A(I30810));
  NOT NOT1_8788(.VSS(VSS),.VDD(VDD),.Y(I30813),.A(g22091));
  NOT NOT1_8789(.VSS(VSS),.VDD(VDD),.Y(g23669),.A(I30813));
  NOT NOT1_8790(.VSS(VSS),.VDD(VDD),.Y(I30816),.A(g22092));
  NOT NOT1_8791(.VSS(VSS),.VDD(VDD),.Y(g23670),.A(I30816));
  NOT NOT1_8792(.VSS(VSS),.VDD(VDD),.Y(I30823),.A(g21972));
  NOT NOT1_8793(.VSS(VSS),.VDD(VDD),.Y(g23675),.A(I30823));
  NOT NOT1_8794(.VSS(VSS),.VDD(VDD),.Y(I30826),.A(g22097));
  NOT NOT1_8795(.VSS(VSS),.VDD(VDD),.Y(g23676),.A(I30826));
  NOT NOT1_8796(.VSS(VSS),.VDD(VDD),.Y(I30829),.A(g22098));
  NOT NOT1_8797(.VSS(VSS),.VDD(VDD),.Y(g23677),.A(I30829));
  NOT NOT1_8798(.VSS(VSS),.VDD(VDD),.Y(I30832),.A(g22099));
  NOT NOT1_8799(.VSS(VSS),.VDD(VDD),.Y(g23678),.A(I30832));
  NOT NOT1_8800(.VSS(VSS),.VDD(VDD),.Y(I30838),.A(g22100));
  NOT NOT1_8801(.VSS(VSS),.VDD(VDD),.Y(g23682),.A(I30838));
  NOT NOT1_8802(.VSS(VSS),.VDD(VDD),.Y(I30841),.A(g22101));
  NOT NOT1_8803(.VSS(VSS),.VDD(VDD),.Y(g23683),.A(I30841));
  NOT NOT1_8804(.VSS(VSS),.VDD(VDD),.Y(I30844),.A(g22102));
  NOT NOT1_8805(.VSS(VSS),.VDD(VDD),.Y(g23684),.A(I30844));
  NOT NOT1_8806(.VSS(VSS),.VDD(VDD),.Y(I30847),.A(g22103));
  NOT NOT1_8807(.VSS(VSS),.VDD(VDD),.Y(g23685),.A(I30847));
  NOT NOT1_8808(.VSS(VSS),.VDD(VDD),.Y(I30854),.A(g22104));
  NOT NOT1_8809(.VSS(VSS),.VDD(VDD),.Y(g23690),.A(I30854));
  NOT NOT1_8810(.VSS(VSS),.VDD(VDD),.Y(I30857),.A(g22105));
  NOT NOT1_8811(.VSS(VSS),.VDD(VDD),.Y(g23691),.A(I30857));
  NOT NOT1_8812(.VSS(VSS),.VDD(VDD),.Y(I30860),.A(g22106));
  NOT NOT1_8813(.VSS(VSS),.VDD(VDD),.Y(g23692),.A(I30860));
  NOT NOT1_8814(.VSS(VSS),.VDD(VDD),.Y(I30864),.A(g22493));
  NOT NOT1_8815(.VSS(VSS),.VDD(VDD),.Y(g23694),.A(I30864));
  NOT NOT1_8816(.VSS(VSS),.VDD(VDD),.Y(I30875),.A(g22112));
  NOT NOT1_8817(.VSS(VSS),.VDD(VDD),.Y(g23711),.A(I30875));
  NOT NOT1_8818(.VSS(VSS),.VDD(VDD),.Y(I30878),.A(g22113));
  NOT NOT1_8819(.VSS(VSS),.VDD(VDD),.Y(g23712),.A(I30878));
  NOT NOT1_8820(.VSS(VSS),.VDD(VDD),.Y(I30881),.A(g22114));
  NOT NOT1_8821(.VSS(VSS),.VDD(VDD),.Y(g23713),.A(I30881));
  NOT NOT1_8822(.VSS(VSS),.VDD(VDD),.Y(I30888),.A(g22115));
  NOT NOT1_8823(.VSS(VSS),.VDD(VDD),.Y(g23718),.A(I30888));
  NOT NOT1_8824(.VSS(VSS),.VDD(VDD),.Y(I30891),.A(g22116));
  NOT NOT1_8825(.VSS(VSS),.VDD(VDD),.Y(g23719),.A(I30891));
  NOT NOT1_8826(.VSS(VSS),.VDD(VDD),.Y(I30894),.A(g22117));
  NOT NOT1_8827(.VSS(VSS),.VDD(VDD),.Y(g23720),.A(I30894));
  NOT NOT1_8828(.VSS(VSS),.VDD(VDD),.Y(I30901),.A(g21974));
  NOT NOT1_8829(.VSS(VSS),.VDD(VDD),.Y(g23725),.A(I30901));
  NOT NOT1_8830(.VSS(VSS),.VDD(VDD),.Y(I30905),.A(g22122));
  NOT NOT1_8831(.VSS(VSS),.VDD(VDD),.Y(g23727),.A(I30905));
  NOT NOT1_8832(.VSS(VSS),.VDD(VDD),.Y(I30908),.A(g22123));
  NOT NOT1_8833(.VSS(VSS),.VDD(VDD),.Y(g23728),.A(I30908));
  NOT NOT1_8834(.VSS(VSS),.VDD(VDD),.Y(I30911),.A(g22124));
  NOT NOT1_8835(.VSS(VSS),.VDD(VDD),.Y(g23729),.A(I30911));
  NOT NOT1_8836(.VSS(VSS),.VDD(VDD),.Y(I30914),.A(g22125));
  NOT NOT1_8837(.VSS(VSS),.VDD(VDD),.Y(g23730),.A(I30914));
  NOT NOT1_8838(.VSS(VSS),.VDD(VDD),.Y(I30917),.A(g22806));
  NOT NOT1_8839(.VSS(VSS),.VDD(VDD),.Y(g23731),.A(I30917));
  NOT NOT1_8840(.VSS(VSS),.VDD(VDD),.Y(I30922),.A(g22126));
  NOT NOT1_8841(.VSS(VSS),.VDD(VDD),.Y(g23736),.A(I30922));
  NOT NOT1_8842(.VSS(VSS),.VDD(VDD),.Y(I30925),.A(g22127));
  NOT NOT1_8843(.VSS(VSS),.VDD(VDD),.Y(g23737),.A(I30925));
  NOT NOT1_8844(.VSS(VSS),.VDD(VDD),.Y(I30928),.A(g22128));
  NOT NOT1_8845(.VSS(VSS),.VDD(VDD),.Y(g23738),.A(I30928));
  NOT NOT1_8846(.VSS(VSS),.VDD(VDD),.Y(I30931),.A(g22129));
  NOT NOT1_8847(.VSS(VSS),.VDD(VDD),.Y(g23739),.A(I30931));
  NOT NOT1_8848(.VSS(VSS),.VDD(VDD),.Y(I30938),.A(g22130));
  NOT NOT1_8849(.VSS(VSS),.VDD(VDD),.Y(g23744),.A(I30938));
  NOT NOT1_8850(.VSS(VSS),.VDD(VDD),.Y(I30941),.A(g22131));
  NOT NOT1_8851(.VSS(VSS),.VDD(VDD),.Y(g23745),.A(I30941));
  NOT NOT1_8852(.VSS(VSS),.VDD(VDD),.Y(I30944),.A(g22132));
  NOT NOT1_8853(.VSS(VSS),.VDD(VDD),.Y(g23746),.A(I30944));
  NOT NOT1_8854(.VSS(VSS),.VDD(VDD),.Y(I30948),.A(g22536));
  NOT NOT1_8855(.VSS(VSS),.VDD(VDD),.Y(g23748),.A(I30948));
  NOT NOT1_8856(.VSS(VSS),.VDD(VDD),.Y(I30959),.A(g22138));
  NOT NOT1_8857(.VSS(VSS),.VDD(VDD),.Y(g23765),.A(I30959));
  NOT NOT1_8858(.VSS(VSS),.VDD(VDD),.Y(I30962),.A(g22139));
  NOT NOT1_8859(.VSS(VSS),.VDD(VDD),.Y(g23766),.A(I30962));
  NOT NOT1_8860(.VSS(VSS),.VDD(VDD),.Y(I30965),.A(g22140));
  NOT NOT1_8861(.VSS(VSS),.VDD(VDD),.Y(g23767),.A(I30965));
  NOT NOT1_8862(.VSS(VSS),.VDD(VDD),.Y(I30973),.A(g22141));
  NOT NOT1_8863(.VSS(VSS),.VDD(VDD),.Y(g23773),.A(I30973));
  NOT NOT1_8864(.VSS(VSS),.VDD(VDD),.Y(I30976),.A(g22142));
  NOT NOT1_8865(.VSS(VSS),.VDD(VDD),.Y(g23774),.A(I30976));
  NOT NOT1_8866(.VSS(VSS),.VDD(VDD),.Y(I30979),.A(g22143));
  NOT NOT1_8867(.VSS(VSS),.VDD(VDD),.Y(g23775),.A(I30979));
  NOT NOT1_8868(.VSS(VSS),.VDD(VDD),.Y(I30985),.A(g22992));
  NOT NOT1_8869(.VSS(VSS),.VDD(VDD),.Y(g23779),.A(I30985));
  NOT NOT1_8870(.VSS(VSS),.VDD(VDD),.Y(I30988),.A(g22145));
  NOT NOT1_8871(.VSS(VSS),.VDD(VDD),.Y(g23782),.A(I30988));
  NOT NOT1_8872(.VSS(VSS),.VDD(VDD),.Y(I30991),.A(g22146));
  NOT NOT1_8873(.VSS(VSS),.VDD(VDD),.Y(g23783),.A(I30991));
  NOT NOT1_8874(.VSS(VSS),.VDD(VDD),.Y(I30994),.A(g22147));
  NOT NOT1_8875(.VSS(VSS),.VDD(VDD),.Y(g23784),.A(I30994));
  NOT NOT1_8876(.VSS(VSS),.VDD(VDD),.Y(I30997),.A(g22148));
  NOT NOT1_8877(.VSS(VSS),.VDD(VDD),.Y(g23785),.A(I30997));
  NOT NOT1_8878(.VSS(VSS),.VDD(VDD),.Y(I31000),.A(g22847));
  NOT NOT1_8879(.VSS(VSS),.VDD(VDD),.Y(g23786),.A(I31000));
  NOT NOT1_8880(.VSS(VSS),.VDD(VDD),.Y(I31005),.A(g22149));
  NOT NOT1_8881(.VSS(VSS),.VDD(VDD),.Y(g23791),.A(I31005));
  NOT NOT1_8882(.VSS(VSS),.VDD(VDD),.Y(I31008),.A(g22150));
  NOT NOT1_8883(.VSS(VSS),.VDD(VDD),.Y(g23792),.A(I31008));
  NOT NOT1_8884(.VSS(VSS),.VDD(VDD),.Y(I31011),.A(g22151));
  NOT NOT1_8885(.VSS(VSS),.VDD(VDD),.Y(g23793),.A(I31011));
  NOT NOT1_8886(.VSS(VSS),.VDD(VDD),.Y(I31014),.A(g22152));
  NOT NOT1_8887(.VSS(VSS),.VDD(VDD),.Y(g23794),.A(I31014));
  NOT NOT1_8888(.VSS(VSS),.VDD(VDD),.Y(I31021),.A(g22153));
  NOT NOT1_8889(.VSS(VSS),.VDD(VDD),.Y(g23799),.A(I31021));
  NOT NOT1_8890(.VSS(VSS),.VDD(VDD),.Y(I31024),.A(g22154));
  NOT NOT1_8891(.VSS(VSS),.VDD(VDD),.Y(g23800),.A(I31024));
  NOT NOT1_8892(.VSS(VSS),.VDD(VDD),.Y(I31027),.A(g22155));
  NOT NOT1_8893(.VSS(VSS),.VDD(VDD),.Y(g23801),.A(I31027));
  NOT NOT1_8894(.VSS(VSS),.VDD(VDD),.Y(I31031),.A(g22576));
  NOT NOT1_8895(.VSS(VSS),.VDD(VDD),.Y(g23803),.A(I31031));
  NOT NOT1_8896(.VSS(VSS),.VDD(VDD),.Y(I31043),.A(g22161));
  NOT NOT1_8897(.VSS(VSS),.VDD(VDD),.Y(g23821),.A(I31043));
  NOT NOT1_8898(.VSS(VSS),.VDD(VDD),.Y(I31050),.A(g22162));
  NOT NOT1_8899(.VSS(VSS),.VDD(VDD),.Y(g23826),.A(I31050));
  NOT NOT1_8900(.VSS(VSS),.VDD(VDD),.Y(I31053),.A(g22163));
  NOT NOT1_8901(.VSS(VSS),.VDD(VDD),.Y(g23827),.A(I31053));
  NOT NOT1_8902(.VSS(VSS),.VDD(VDD),.Y(I31056),.A(g22164));
  NOT NOT1_8903(.VSS(VSS),.VDD(VDD),.Y(g23828),.A(I31056));
  NOT NOT1_8904(.VSS(VSS),.VDD(VDD),.Y(I31062),.A(g23003));
  NOT NOT1_8905(.VSS(VSS),.VDD(VDD),.Y(g23832),.A(I31062));
  NOT NOT1_8906(.VSS(VSS),.VDD(VDD),.Y(I31065),.A(g22166));
  NOT NOT1_8907(.VSS(VSS),.VDD(VDD),.Y(g23835),.A(I31065));
  NOT NOT1_8908(.VSS(VSS),.VDD(VDD),.Y(I31068),.A(g22167));
  NOT NOT1_8909(.VSS(VSS),.VDD(VDD),.Y(g23836),.A(I31068));
  NOT NOT1_8910(.VSS(VSS),.VDD(VDD),.Y(I31071),.A(g22168));
  NOT NOT1_8911(.VSS(VSS),.VDD(VDD),.Y(g23837),.A(I31071));
  NOT NOT1_8912(.VSS(VSS),.VDD(VDD),.Y(I31074),.A(g22169));
  NOT NOT1_8913(.VSS(VSS),.VDD(VDD),.Y(g23838),.A(I31074));
  NOT NOT1_8914(.VSS(VSS),.VDD(VDD),.Y(I31077),.A(g22882));
  NOT NOT1_8915(.VSS(VSS),.VDD(VDD),.Y(g23839),.A(I31077));
  NOT NOT1_8916(.VSS(VSS),.VDD(VDD),.Y(I31082),.A(g22170));
  NOT NOT1_8917(.VSS(VSS),.VDD(VDD),.Y(g23844),.A(I31082));
  NOT NOT1_8918(.VSS(VSS),.VDD(VDD),.Y(I31085),.A(g22171));
  NOT NOT1_8919(.VSS(VSS),.VDD(VDD),.Y(g23845),.A(I31085));
  NOT NOT1_8920(.VSS(VSS),.VDD(VDD),.Y(I31088),.A(g22172));
  NOT NOT1_8921(.VSS(VSS),.VDD(VDD),.Y(g23846),.A(I31088));
  NOT NOT1_8922(.VSS(VSS),.VDD(VDD),.Y(I31091),.A(g22173));
  NOT NOT1_8923(.VSS(VSS),.VDD(VDD),.Y(g23847),.A(I31091));
  NOT NOT1_8924(.VSS(VSS),.VDD(VDD),.Y(g23853),.A(g22300));
  NOT NOT1_8925(.VSS(VSS),.VDD(VDD),.Y(I31102),.A(g22177));
  NOT NOT1_8926(.VSS(VSS),.VDD(VDD),.Y(g23856),.A(I31102));
  NOT NOT1_8927(.VSS(VSS),.VDD(VDD),.Y(I31109),.A(g22178));
  NOT NOT1_8928(.VSS(VSS),.VDD(VDD),.Y(g23861),.A(I31109));
  NOT NOT1_8929(.VSS(VSS),.VDD(VDD),.Y(I31112),.A(g22179));
  NOT NOT1_8930(.VSS(VSS),.VDD(VDD),.Y(g23862),.A(I31112));
  NOT NOT1_8931(.VSS(VSS),.VDD(VDD),.Y(I31115),.A(g22180));
  NOT NOT1_8932(.VSS(VSS),.VDD(VDD),.Y(g23863),.A(I31115));
  NOT NOT1_8933(.VSS(VSS),.VDD(VDD),.Y(I31121),.A(g23017));
  NOT NOT1_8934(.VSS(VSS),.VDD(VDD),.Y(g23867),.A(I31121));
  NOT NOT1_8935(.VSS(VSS),.VDD(VDD),.Y(I31124),.A(g22182));
  NOT NOT1_8936(.VSS(VSS),.VDD(VDD),.Y(g23870),.A(I31124));
  NOT NOT1_8937(.VSS(VSS),.VDD(VDD),.Y(I31127),.A(g22183));
  NOT NOT1_8938(.VSS(VSS),.VDD(VDD),.Y(g23871),.A(I31127));
  NOT NOT1_8939(.VSS(VSS),.VDD(VDD),.Y(I31130),.A(g22184));
  NOT NOT1_8940(.VSS(VSS),.VDD(VDD),.Y(g23872),.A(I31130));
  NOT NOT1_8941(.VSS(VSS),.VDD(VDD),.Y(I31133),.A(g22185));
  NOT NOT1_8942(.VSS(VSS),.VDD(VDD),.Y(g23873),.A(I31133));
  NOT NOT1_8943(.VSS(VSS),.VDD(VDD),.Y(I31136),.A(g22917));
  NOT NOT1_8944(.VSS(VSS),.VDD(VDD),.Y(g23874),.A(I31136));
  NOT NOT1_8945(.VSS(VSS),.VDD(VDD),.Y(I31141),.A(g22777));
  NOT NOT1_8946(.VSS(VSS),.VDD(VDD),.Y(g23879),.A(I31141));
  NOT NOT1_8947(.VSS(VSS),.VDD(VDD),.Y(I31144),.A(g22935));
  NOT NOT1_8948(.VSS(VSS),.VDD(VDD),.Y(g23882),.A(I31144));
  NOT NOT1_8949(.VSS(VSS),.VDD(VDD),.Y(g23885),.A(g22062));
  NOT NOT1_8950(.VSS(VSS),.VDD(VDD),.Y(g23887),.A(g22328));
  NOT NOT1_8951(.VSS(VSS),.VDD(VDD),.Y(I31152),.A(g22191));
  NOT NOT1_8952(.VSS(VSS),.VDD(VDD),.Y(g23890),.A(I31152));
  NOT NOT1_8953(.VSS(VSS),.VDD(VDD),.Y(I31159),.A(g22192));
  NOT NOT1_8954(.VSS(VSS),.VDD(VDD),.Y(g23895),.A(I31159));
  NOT NOT1_8955(.VSS(VSS),.VDD(VDD),.Y(I31162),.A(g22193));
  NOT NOT1_8956(.VSS(VSS),.VDD(VDD),.Y(g23896),.A(I31162));
  NOT NOT1_8957(.VSS(VSS),.VDD(VDD),.Y(I31165),.A(g22194));
  NOT NOT1_8958(.VSS(VSS),.VDD(VDD),.Y(g23897),.A(I31165));
  NOT NOT1_8959(.VSS(VSS),.VDD(VDD),.Y(I31171),.A(g23033));
  NOT NOT1_8960(.VSS(VSS),.VDD(VDD),.Y(g23901),.A(I31171));
  NOT NOT1_8961(.VSS(VSS),.VDD(VDD),.Y(g23905),.A(g22046));
  NOT NOT1_8962(.VSS(VSS),.VDD(VDD),.Y(g23908),.A(g22353));
  NOT NOT1_8963(.VSS(VSS),.VDD(VDD),.Y(I31181),.A(g22200));
  NOT NOT1_8964(.VSS(VSS),.VDD(VDD),.Y(g23911),.A(I31181));
  NOT NOT1_8965(.VSS(VSS),.VDD(VDD),.Y(I31188),.A(g21989));
  NOT NOT1_8966(.VSS(VSS),.VDD(VDD),.Y(g23916),.A(I31188));
  NOT NOT1_8967(.VSS(VSS),.VDD(VDD),.Y(g23918),.A(g22036));
  NOT NOT1_8968(.VSS(VSS),.VDD(VDD),.Y(I31195),.A(g22578));
  NOT NOT1_8969(.VSS(VSS),.VDD(VDD),.Y(g23923),.A(I31195));
  NOT NOT1_8970(.VSS(VSS),.VDD(VDD),.Y(g23940),.A(g22376));
  NOT NOT1_8971(.VSS(VSS),.VDD(VDD),.Y(I31205),.A(g22002));
  NOT NOT1_8972(.VSS(VSS),.VDD(VDD),.Y(g23943),.A(I31205));
  NOT NOT1_8973(.VSS(VSS),.VDD(VDD),.Y(I31213),.A(g22615));
  NOT NOT1_8974(.VSS(VSS),.VDD(VDD),.Y(g23955),.A(I31213));
  NOT NOT1_8975(.VSS(VSS),.VDD(VDD),.Y(I31226),.A(g22651));
  NOT NOT1_8976(.VSS(VSS),.VDD(VDD),.Y(g23984),.A(I31226));
  NOT NOT1_8977(.VSS(VSS),.VDD(VDD),.Y(I31232),.A(g22026));
  NOT NOT1_8978(.VSS(VSS),.VDD(VDD),.Y(g24000),.A(I31232));
  NOT NOT1_8979(.VSS(VSS),.VDD(VDD),.Y(I31235),.A(g22218));
  NOT NOT1_8980(.VSS(VSS),.VDD(VDD),.Y(g24001),.A(I31235));
  NOT NOT1_8981(.VSS(VSS),.VDD(VDD),.Y(I31244),.A(g22687));
  NOT NOT1_8982(.VSS(VSS),.VDD(VDD),.Y(g24014),.A(I31244));
  NOT NOT1_8983(.VSS(VSS),.VDD(VDD),.Y(I31250),.A(g22953));
  NOT NOT1_8984(.VSS(VSS),.VDD(VDD),.Y(g24030),.A(I31250));
  NOT NOT1_8985(.VSS(VSS),.VDD(VDD),.Y(I31253),.A(g22231));
  NOT NOT1_8986(.VSS(VSS),.VDD(VDD),.Y(g24033),.A(I31253));
  NOT NOT1_8987(.VSS(VSS),.VDD(VDD),.Y(I31257),.A(g22234));
  NOT NOT1_8988(.VSS(VSS),.VDD(VDD),.Y(g24035),.A(I31257));
  NOT NOT1_8989(.VSS(VSS),.VDD(VDD),.Y(g24047),.A(g23023));
  NOT NOT1_8990(.VSS(VSS),.VDD(VDD),.Y(I31266),.A(g22242));
  NOT NOT1_8991(.VSS(VSS),.VDD(VDD),.Y(g24051),.A(I31266));
  NOT NOT1_8992(.VSS(VSS),.VDD(VDD),.Y(I31270),.A(g22247));
  NOT NOT1_8993(.VSS(VSS),.VDD(VDD),.Y(g24053),.A(I31270));
  NOT NOT1_8994(.VSS(VSS),.VDD(VDD),.Y(I31274),.A(g22249));
  NOT NOT1_8995(.VSS(VSS),.VDD(VDD),.Y(g24055),.A(I31274));
  NOT NOT1_8996(.VSS(VSS),.VDD(VDD),.Y(g24060),.A(g23040));
  NOT NOT1_8997(.VSS(VSS),.VDD(VDD),.Y(I31282),.A(g22263));
  NOT NOT1_8998(.VSS(VSS),.VDD(VDD),.Y(g24064),.A(I31282));
  NOT NOT1_8999(.VSS(VSS),.VDD(VDD),.Y(I31286),.A(g22267));
  NOT NOT1_9000(.VSS(VSS),.VDD(VDD),.Y(g24066),.A(I31286));
  NOT NOT1_9001(.VSS(VSS),.VDD(VDD),.Y(I31290),.A(g22269));
  NOT NOT1_9002(.VSS(VSS),.VDD(VDD),.Y(g24068),.A(I31290));
  NOT NOT1_9003(.VSS(VSS),.VDD(VDD),.Y(g24073),.A(g23059));
  NOT NOT1_9004(.VSS(VSS),.VDD(VDD),.Y(I31298),.A(g22280));
  NOT NOT1_9005(.VSS(VSS),.VDD(VDD),.Y(g24077),.A(I31298));
  NOT NOT1_9006(.VSS(VSS),.VDD(VDD),.Y(I31302),.A(g22284));
  NOT NOT1_9007(.VSS(VSS),.VDD(VDD),.Y(g24079),.A(I31302));
  NOT NOT1_9008(.VSS(VSS),.VDD(VDD),.Y(g24084),.A(g23077));
  NOT NOT1_9009(.VSS(VSS),.VDD(VDD),.Y(I31310),.A(g22299));
  NOT NOT1_9010(.VSS(VSS),.VDD(VDD),.Y(g24088),.A(I31310));
  NOT NOT1_9011(.VSS(VSS),.VDD(VDD),.Y(g24094),.A(g22339));
  NOT NOT1_9012(.VSS(VSS),.VDD(VDD),.Y(g24095),.A(g22362));
  NOT NOT1_9013(.VSS(VSS),.VDD(VDD),.Y(g24096),.A(g22405));
  NOT NOT1_9014(.VSS(VSS),.VDD(VDD),.Y(g24097),.A(g22382));
  NOT NOT1_9015(.VSS(VSS),.VDD(VDD),.Y(g24098),.A(g22409));
  NOT NOT1_9016(.VSS(VSS),.VDD(VDD),.Y(g24099),.A(g22412));
  NOT NOT1_9017(.VSS(VSS),.VDD(VDD),.Y(g24101),.A(g22415));
  NOT NOT1_9018(.VSS(VSS),.VDD(VDD),.Y(g24102),.A(g22418));
  NOT NOT1_9019(.VSS(VSS),.VDD(VDD),.Y(g24103),.A(g22397));
  NOT NOT1_9020(.VSS(VSS),.VDD(VDD),.Y(g24104),.A(g22422));
  NOT NOT1_9021(.VSS(VSS),.VDD(VDD),.Y(g24105),.A(g22425));
  NOT NOT1_9022(.VSS(VSS),.VDD(VDD),.Y(g24106),.A(g22428));
  NOT NOT1_9023(.VSS(VSS),.VDD(VDD),.Y(g24107),.A(g22431));
  NOT NOT1_9024(.VSS(VSS),.VDD(VDD),.Y(g24108),.A(g22434));
  NOT NOT1_9025(.VSS(VSS),.VDD(VDD),.Y(g24110),.A(g22437));
  NOT NOT1_9026(.VSS(VSS),.VDD(VDD),.Y(g24111),.A(g22440));
  NOT NOT1_9027(.VSS(VSS),.VDD(VDD),.Y(g24112),.A(g22445));
  NOT NOT1_9028(.VSS(VSS),.VDD(VDD),.Y(g24113),.A(g22448));
  NOT NOT1_9029(.VSS(VSS),.VDD(VDD),.Y(g24114),.A(g22451));
  NOT NOT1_9030(.VSS(VSS),.VDD(VDD),.Y(g24115),.A(g22381));
  NOT NOT1_9031(.VSS(VSS),.VDD(VDD),.Y(g24121),.A(g22455));
  NOT NOT1_9032(.VSS(VSS),.VDD(VDD),.Y(g24122),.A(g22458));
  NOT NOT1_9033(.VSS(VSS),.VDD(VDD),.Y(g24123),.A(g22461));
  NOT NOT1_9034(.VSS(VSS),.VDD(VDD),.Y(g24124),.A(g22464));
  NOT NOT1_9035(.VSS(VSS),.VDD(VDD),.Y(g24125),.A(g22467));
  NOT NOT1_9036(.VSS(VSS),.VDD(VDD),.Y(g24127),.A(g22470));
  NOT NOT1_9037(.VSS(VSS),.VDD(VDD),.Y(g24128),.A(g22473));
  NOT NOT1_9038(.VSS(VSS),.VDD(VDD),.Y(g24129),.A(g22477));
  NOT NOT1_9039(.VSS(VSS),.VDD(VDD),.Y(g24130),.A(g22480));
  NOT NOT1_9040(.VSS(VSS),.VDD(VDD),.Y(g24131),.A(g22484));
  NOT NOT1_9041(.VSS(VSS),.VDD(VDD),.Y(g24132),.A(g22487));
  NOT NOT1_9042(.VSS(VSS),.VDD(VDD),.Y(g24133),.A(g22490));
  NOT NOT1_9043(.VSS(VSS),.VDD(VDD),.Y(g24134),.A(g22396));
  NOT NOT1_9044(.VSS(VSS),.VDD(VDD),.Y(g24140),.A(g22494));
  NOT NOT1_9045(.VSS(VSS),.VDD(VDD),.Y(g24141),.A(g22497));
  NOT NOT1_9046(.VSS(VSS),.VDD(VDD),.Y(g24142),.A(g22500));
  NOT NOT1_9047(.VSS(VSS),.VDD(VDD),.Y(g24143),.A(g22503));
  NOT NOT1_9048(.VSS(VSS),.VDD(VDD),.Y(g24144),.A(g22506));
  NOT NOT1_9049(.VSS(VSS),.VDD(VDD),.Y(g24146),.A(g22509));
  NOT NOT1_9050(.VSS(VSS),.VDD(VDD),.Y(g24147),.A(g22512));
  NOT NOT1_9051(.VSS(VSS),.VDD(VDD),.Y(g24148),.A(g22520));
  NOT NOT1_9052(.VSS(VSS),.VDD(VDD),.Y(g24149),.A(g22523));
  NOT NOT1_9053(.VSS(VSS),.VDD(VDD),.Y(g24150),.A(g22527));
  NOT NOT1_9054(.VSS(VSS),.VDD(VDD),.Y(g24151),.A(g22530));
  NOT NOT1_9055(.VSS(VSS),.VDD(VDD),.Y(g24152),.A(g22533));
  NOT NOT1_9056(.VSS(VSS),.VDD(VDD),.Y(g24153),.A(g22399));
  NOT NOT1_9057(.VSS(VSS),.VDD(VDD),.Y(g24159),.A(g22537));
  NOT NOT1_9058(.VSS(VSS),.VDD(VDD),.Y(g24160),.A(g22540));
  NOT NOT1_9059(.VSS(VSS),.VDD(VDD),.Y(g24161),.A(g22543));
  NOT NOT1_9060(.VSS(VSS),.VDD(VDD),.Y(g24162),.A(g22552));
  NOT NOT1_9061(.VSS(VSS),.VDD(VDD),.Y(g24163),.A(g22560));
  NOT NOT1_9062(.VSS(VSS),.VDD(VDD),.Y(g24164),.A(g22563));
  NOT NOT1_9063(.VSS(VSS),.VDD(VDD),.Y(g24165),.A(g22567));
  NOT NOT1_9064(.VSS(VSS),.VDD(VDD),.Y(g24166),.A(g22570));
  NOT NOT1_9065(.VSS(VSS),.VDD(VDD),.Y(g24167),.A(g22573));
  NOT NOT1_9066(.VSS(VSS),.VDD(VDD),.Y(g24168),.A(g22400));
  NOT NOT1_9067(.VSS(VSS),.VDD(VDD),.Y(g24175),.A(g22592));
  NOT NOT1_9068(.VSS(VSS),.VDD(VDD),.Y(g24176),.A(g22600));
  NOT NOT1_9069(.VSS(VSS),.VDD(VDD),.Y(g24177),.A(g22603));
  NOT NOT1_9070(.VSS(VSS),.VDD(VDD),.Y(g24180),.A(g22629));
  NOT NOT1_9071(.VSS(VSS),.VDD(VDD),.Y(I31387),.A(g22811));
  NOT NOT1_9072(.VSS(VSS),.VDD(VDD),.Y(g24183),.A(I31387));
  NOT NOT1_9073(.VSS(VSS),.VDD(VDD),.Y(g24210),.A(g22696));
  NOT NOT1_9074(.VSS(VSS),.VDD(VDD),.Y(g24220),.A(g22750));
  NOT NOT1_9075(.VSS(VSS),.VDD(VDD),.Y(I31417),.A(g22578));
  NOT NOT1_9076(.VSS(VSS),.VDD(VDD),.Y(g24233),.A(I31417));
  NOT NOT1_9077(.VSS(VSS),.VDD(VDD),.Y(I31426),.A(g22615));
  NOT NOT1_9078(.VSS(VSS),.VDD(VDD),.Y(g24240),.A(I31426));
  NOT NOT1_9079(.VSS(VSS),.VDD(VDD),.Y(I31436),.A(g22651));
  NOT NOT1_9080(.VSS(VSS),.VDD(VDD),.Y(g24248),.A(I31436));
  NOT NOT1_9081(.VSS(VSS),.VDD(VDD),.Y(g24251),.A(g22903));
  NOT NOT1_9082(.VSS(VSS),.VDD(VDD),.Y(I31445),.A(g22687));
  NOT NOT1_9083(.VSS(VSS),.VDD(VDD),.Y(g24255),.A(I31445));
  NOT NOT1_9084(.VSS(VSS),.VDD(VDD),.Y(I31451),.A(g23682));
  NOT NOT1_9085(.VSS(VSS),.VDD(VDD),.Y(g24259),.A(I31451));
  NOT NOT1_9086(.VSS(VSS),.VDD(VDD),.Y(I31454),.A(g23727));
  NOT NOT1_9087(.VSS(VSS),.VDD(VDD),.Y(g24260),.A(I31454));
  NOT NOT1_9088(.VSS(VSS),.VDD(VDD),.Y(I31457),.A(g23773));
  NOT NOT1_9089(.VSS(VSS),.VDD(VDD),.Y(g24261),.A(I31457));
  NOT NOT1_9090(.VSS(VSS),.VDD(VDD),.Y(I31460),.A(g23728));
  NOT NOT1_9091(.VSS(VSS),.VDD(VDD),.Y(g24262),.A(I31460));
  NOT NOT1_9092(.VSS(VSS),.VDD(VDD),.Y(I31463),.A(g23774));
  NOT NOT1_9093(.VSS(VSS),.VDD(VDD),.Y(g24263),.A(I31463));
  NOT NOT1_9094(.VSS(VSS),.VDD(VDD),.Y(I31466),.A(g23821));
  NOT NOT1_9095(.VSS(VSS),.VDD(VDD),.Y(g24264),.A(I31466));
  NOT NOT1_9096(.VSS(VSS),.VDD(VDD),.Y(I31469),.A(g23546));
  NOT NOT1_9097(.VSS(VSS),.VDD(VDD),.Y(g24265),.A(I31469));
  NOT NOT1_9098(.VSS(VSS),.VDD(VDD),.Y(I31472),.A(g23548));
  NOT NOT1_9099(.VSS(VSS),.VDD(VDD),.Y(g24266),.A(I31472));
  NOT NOT1_9100(.VSS(VSS),.VDD(VDD),.Y(I31475),.A(g23555));
  NOT NOT1_9101(.VSS(VSS),.VDD(VDD),.Y(g24267),.A(I31475));
  NOT NOT1_9102(.VSS(VSS),.VDD(VDD),.Y(I31478),.A(g23549));
  NOT NOT1_9103(.VSS(VSS),.VDD(VDD),.Y(g24268),.A(I31478));
  NOT NOT1_9104(.VSS(VSS),.VDD(VDD),.Y(I31481),.A(g23556));
  NOT NOT1_9105(.VSS(VSS),.VDD(VDD),.Y(g24269),.A(I31481));
  NOT NOT1_9106(.VSS(VSS),.VDD(VDD),.Y(I31484),.A(g23568));
  NOT NOT1_9107(.VSS(VSS),.VDD(VDD),.Y(g24270),.A(I31484));
  NOT NOT1_9108(.VSS(VSS),.VDD(VDD),.Y(I31487),.A(g23557));
  NOT NOT1_9109(.VSS(VSS),.VDD(VDD),.Y(g24271),.A(I31487));
  NOT NOT1_9110(.VSS(VSS),.VDD(VDD),.Y(I31490),.A(g23569));
  NOT NOT1_9111(.VSS(VSS),.VDD(VDD),.Y(g24272),.A(I31490));
  NOT NOT1_9112(.VSS(VSS),.VDD(VDD),.Y(I31493),.A(g23587));
  NOT NOT1_9113(.VSS(VSS),.VDD(VDD),.Y(g24273),.A(I31493));
  NOT NOT1_9114(.VSS(VSS),.VDD(VDD),.Y(I31496),.A(g23570));
  NOT NOT1_9115(.VSS(VSS),.VDD(VDD),.Y(g24274),.A(I31496));
  NOT NOT1_9116(.VSS(VSS),.VDD(VDD),.Y(I31499),.A(g23588));
  NOT NOT1_9117(.VSS(VSS),.VDD(VDD),.Y(g24275),.A(I31499));
  NOT NOT1_9118(.VSS(VSS),.VDD(VDD),.Y(I31502),.A(g23612));
  NOT NOT1_9119(.VSS(VSS),.VDD(VDD),.Y(g24276),.A(I31502));
  NOT NOT1_9120(.VSS(VSS),.VDD(VDD),.Y(I31505),.A(g23589));
  NOT NOT1_9121(.VSS(VSS),.VDD(VDD),.Y(g24277),.A(I31505));
  NOT NOT1_9122(.VSS(VSS),.VDD(VDD),.Y(I31508),.A(g23613));
  NOT NOT1_9123(.VSS(VSS),.VDD(VDD),.Y(g24278),.A(I31508));
  NOT NOT1_9124(.VSS(VSS),.VDD(VDD),.Y(I31511),.A(g23640));
  NOT NOT1_9125(.VSS(VSS),.VDD(VDD),.Y(g24279),.A(I31511));
  NOT NOT1_9126(.VSS(VSS),.VDD(VDD),.Y(I31514),.A(g23614));
  NOT NOT1_9127(.VSS(VSS),.VDD(VDD),.Y(g24280),.A(I31514));
  NOT NOT1_9128(.VSS(VSS),.VDD(VDD),.Y(I31517),.A(g23641));
  NOT NOT1_9129(.VSS(VSS),.VDD(VDD),.Y(g24281),.A(I31517));
  NOT NOT1_9130(.VSS(VSS),.VDD(VDD),.Y(I31520),.A(g23683));
  NOT NOT1_9131(.VSS(VSS),.VDD(VDD),.Y(g24282),.A(I31520));
  NOT NOT1_9132(.VSS(VSS),.VDD(VDD),.Y(I31523),.A(g23642));
  NOT NOT1_9133(.VSS(VSS),.VDD(VDD),.Y(g24283),.A(I31523));
  NOT NOT1_9134(.VSS(VSS),.VDD(VDD),.Y(I31526),.A(g23684));
  NOT NOT1_9135(.VSS(VSS),.VDD(VDD),.Y(g24284),.A(I31526));
  NOT NOT1_9136(.VSS(VSS),.VDD(VDD),.Y(I31529),.A(g23729));
  NOT NOT1_9137(.VSS(VSS),.VDD(VDD),.Y(g24285),.A(I31529));
  NOT NOT1_9138(.VSS(VSS),.VDD(VDD),.Y(I31532),.A(g23685));
  NOT NOT1_9139(.VSS(VSS),.VDD(VDD),.Y(g24286),.A(I31532));
  NOT NOT1_9140(.VSS(VSS),.VDD(VDD),.Y(I31535),.A(g23730));
  NOT NOT1_9141(.VSS(VSS),.VDD(VDD),.Y(g24287),.A(I31535));
  NOT NOT1_9142(.VSS(VSS),.VDD(VDD),.Y(I31538),.A(g23775));
  NOT NOT1_9143(.VSS(VSS),.VDD(VDD),.Y(g24288),.A(I31538));
  NOT NOT1_9144(.VSS(VSS),.VDD(VDD),.Y(I31541),.A(g23500));
  NOT NOT1_9145(.VSS(VSS),.VDD(VDD),.Y(g24289),.A(I31541));
  NOT NOT1_9146(.VSS(VSS),.VDD(VDD),.Y(I31544),.A(g23438));
  NOT NOT1_9147(.VSS(VSS),.VDD(VDD),.Y(g24290),.A(I31544));
  NOT NOT1_9148(.VSS(VSS),.VDD(VDD),.Y(I31547),.A(g23454));
  NOT NOT1_9149(.VSS(VSS),.VDD(VDD),.Y(g24291),.A(I31547));
  NOT NOT1_9150(.VSS(VSS),.VDD(VDD),.Y(I31550),.A(g23481));
  NOT NOT1_9151(.VSS(VSS),.VDD(VDD),.Y(g24292),.A(I31550));
  NOT NOT1_9152(.VSS(VSS),.VDD(VDD),.Y(I31553),.A(g23501));
  NOT NOT1_9153(.VSS(VSS),.VDD(VDD),.Y(g24293),.A(I31553));
  NOT NOT1_9154(.VSS(VSS),.VDD(VDD),.Y(I31556),.A(g23439));
  NOT NOT1_9155(.VSS(VSS),.VDD(VDD),.Y(g24294),.A(I31556));
  NOT NOT1_9156(.VSS(VSS),.VDD(VDD),.Y(I31559),.A(g24233));
  NOT NOT1_9157(.VSS(VSS),.VDD(VDD),.Y(g24295),.A(I31559));
  NOT NOT1_9158(.VSS(VSS),.VDD(VDD),.Y(I31562),.A(g23594));
  NOT NOT1_9159(.VSS(VSS),.VDD(VDD),.Y(g24296),.A(I31562));
  NOT NOT1_9160(.VSS(VSS),.VDD(VDD),.Y(I31565),.A(g24001));
  NOT NOT1_9161(.VSS(VSS),.VDD(VDD),.Y(g24297),.A(I31565));
  NOT NOT1_9162(.VSS(VSS),.VDD(VDD),.Y(I31568),.A(g24033));
  NOT NOT1_9163(.VSS(VSS),.VDD(VDD),.Y(g24298),.A(I31568));
  NOT NOT1_9164(.VSS(VSS),.VDD(VDD),.Y(I31571),.A(g24051));
  NOT NOT1_9165(.VSS(VSS),.VDD(VDD),.Y(g24299),.A(I31571));
  NOT NOT1_9166(.VSS(VSS),.VDD(VDD),.Y(I31574),.A(g23736));
  NOT NOT1_9167(.VSS(VSS),.VDD(VDD),.Y(g24300),.A(I31574));
  NOT NOT1_9168(.VSS(VSS),.VDD(VDD),.Y(I31577),.A(g23782));
  NOT NOT1_9169(.VSS(VSS),.VDD(VDD),.Y(g24301),.A(I31577));
  NOT NOT1_9170(.VSS(VSS),.VDD(VDD),.Y(I31580),.A(g23826));
  NOT NOT1_9171(.VSS(VSS),.VDD(VDD),.Y(g24302),.A(I31580));
  NOT NOT1_9172(.VSS(VSS),.VDD(VDD),.Y(I31583),.A(g23783));
  NOT NOT1_9173(.VSS(VSS),.VDD(VDD),.Y(g24303),.A(I31583));
  NOT NOT1_9174(.VSS(VSS),.VDD(VDD),.Y(I31586),.A(g23827));
  NOT NOT1_9175(.VSS(VSS),.VDD(VDD),.Y(g24304),.A(I31586));
  NOT NOT1_9176(.VSS(VSS),.VDD(VDD),.Y(I31589),.A(g23856));
  NOT NOT1_9177(.VSS(VSS),.VDD(VDD),.Y(g24305),.A(I31589));
  NOT NOT1_9178(.VSS(VSS),.VDD(VDD),.Y(I31592),.A(g23553));
  NOT NOT1_9179(.VSS(VSS),.VDD(VDD),.Y(g24306),.A(I31592));
  NOT NOT1_9180(.VSS(VSS),.VDD(VDD),.Y(I31595),.A(g23561));
  NOT NOT1_9181(.VSS(VSS),.VDD(VDD),.Y(g24307),.A(I31595));
  NOT NOT1_9182(.VSS(VSS),.VDD(VDD),.Y(I31598),.A(g23574));
  NOT NOT1_9183(.VSS(VSS),.VDD(VDD),.Y(g24308),.A(I31598));
  NOT NOT1_9184(.VSS(VSS),.VDD(VDD),.Y(I31601),.A(g23562));
  NOT NOT1_9185(.VSS(VSS),.VDD(VDD),.Y(g24309),.A(I31601));
  NOT NOT1_9186(.VSS(VSS),.VDD(VDD),.Y(I31604),.A(g23575));
  NOT NOT1_9187(.VSS(VSS),.VDD(VDD),.Y(g24310),.A(I31604));
  NOT NOT1_9188(.VSS(VSS),.VDD(VDD),.Y(I31607),.A(g23595));
  NOT NOT1_9189(.VSS(VSS),.VDD(VDD),.Y(g24311),.A(I31607));
  NOT NOT1_9190(.VSS(VSS),.VDD(VDD),.Y(I31610),.A(g23576));
  NOT NOT1_9191(.VSS(VSS),.VDD(VDD),.Y(g24312),.A(I31610));
  NOT NOT1_9192(.VSS(VSS),.VDD(VDD),.Y(I31613),.A(g23596));
  NOT NOT1_9193(.VSS(VSS),.VDD(VDD),.Y(g24313),.A(I31613));
  NOT NOT1_9194(.VSS(VSS),.VDD(VDD),.Y(I31616),.A(g23619));
  NOT NOT1_9195(.VSS(VSS),.VDD(VDD),.Y(g24314),.A(I31616));
  NOT NOT1_9196(.VSS(VSS),.VDD(VDD),.Y(I31619),.A(g23597));
  NOT NOT1_9197(.VSS(VSS),.VDD(VDD),.Y(g24315),.A(I31619));
  NOT NOT1_9198(.VSS(VSS),.VDD(VDD),.Y(I31622),.A(g23620));
  NOT NOT1_9199(.VSS(VSS),.VDD(VDD),.Y(g24316),.A(I31622));
  NOT NOT1_9200(.VSS(VSS),.VDD(VDD),.Y(I31625),.A(g23661));
  NOT NOT1_9201(.VSS(VSS),.VDD(VDD),.Y(g24317),.A(I31625));
  NOT NOT1_9202(.VSS(VSS),.VDD(VDD),.Y(I31628),.A(g23621));
  NOT NOT1_9203(.VSS(VSS),.VDD(VDD),.Y(g24318),.A(I31628));
  NOT NOT1_9204(.VSS(VSS),.VDD(VDD),.Y(I31631),.A(g23662));
  NOT NOT1_9205(.VSS(VSS),.VDD(VDD),.Y(g24319),.A(I31631));
  NOT NOT1_9206(.VSS(VSS),.VDD(VDD),.Y(I31634),.A(g23690));
  NOT NOT1_9207(.VSS(VSS),.VDD(VDD),.Y(g24320),.A(I31634));
  NOT NOT1_9208(.VSS(VSS),.VDD(VDD),.Y(I31637),.A(g23663));
  NOT NOT1_9209(.VSS(VSS),.VDD(VDD),.Y(g24321),.A(I31637));
  NOT NOT1_9210(.VSS(VSS),.VDD(VDD),.Y(I31640),.A(g23691));
  NOT NOT1_9211(.VSS(VSS),.VDD(VDD),.Y(g24322),.A(I31640));
  NOT NOT1_9212(.VSS(VSS),.VDD(VDD),.Y(I31643),.A(g23737));
  NOT NOT1_9213(.VSS(VSS),.VDD(VDD),.Y(g24323),.A(I31643));
  NOT NOT1_9214(.VSS(VSS),.VDD(VDD),.Y(I31646),.A(g23692));
  NOT NOT1_9215(.VSS(VSS),.VDD(VDD),.Y(g24324),.A(I31646));
  NOT NOT1_9216(.VSS(VSS),.VDD(VDD),.Y(I31649),.A(g23738));
  NOT NOT1_9217(.VSS(VSS),.VDD(VDD),.Y(g24325),.A(I31649));
  NOT NOT1_9218(.VSS(VSS),.VDD(VDD),.Y(I31652),.A(g23784));
  NOT NOT1_9219(.VSS(VSS),.VDD(VDD),.Y(g24326),.A(I31652));
  NOT NOT1_9220(.VSS(VSS),.VDD(VDD),.Y(I31655),.A(g23739));
  NOT NOT1_9221(.VSS(VSS),.VDD(VDD),.Y(g24327),.A(I31655));
  NOT NOT1_9222(.VSS(VSS),.VDD(VDD),.Y(I31658),.A(g23785));
  NOT NOT1_9223(.VSS(VSS),.VDD(VDD),.Y(g24328),.A(I31658));
  NOT NOT1_9224(.VSS(VSS),.VDD(VDD),.Y(I31661),.A(g23828));
  NOT NOT1_9225(.VSS(VSS),.VDD(VDD),.Y(g24329),.A(I31661));
  NOT NOT1_9226(.VSS(VSS),.VDD(VDD),.Y(I31664),.A(g23516));
  NOT NOT1_9227(.VSS(VSS),.VDD(VDD),.Y(g24330),.A(I31664));
  NOT NOT1_9228(.VSS(VSS),.VDD(VDD),.Y(I31667),.A(g23452));
  NOT NOT1_9229(.VSS(VSS),.VDD(VDD),.Y(g24331),.A(I31667));
  NOT NOT1_9230(.VSS(VSS),.VDD(VDD),.Y(I31670),.A(g23463));
  NOT NOT1_9231(.VSS(VSS),.VDD(VDD),.Y(g24332),.A(I31670));
  NOT NOT1_9232(.VSS(VSS),.VDD(VDD),.Y(I31673),.A(g23492));
  NOT NOT1_9233(.VSS(VSS),.VDD(VDD),.Y(g24333),.A(I31673));
  NOT NOT1_9234(.VSS(VSS),.VDD(VDD),.Y(I31676),.A(g23517));
  NOT NOT1_9235(.VSS(VSS),.VDD(VDD),.Y(g24334),.A(I31676));
  NOT NOT1_9236(.VSS(VSS),.VDD(VDD),.Y(I31679),.A(g23453));
  NOT NOT1_9237(.VSS(VSS),.VDD(VDD),.Y(g24335),.A(I31679));
  NOT NOT1_9238(.VSS(VSS),.VDD(VDD),.Y(I31682),.A(g24240));
  NOT NOT1_9239(.VSS(VSS),.VDD(VDD),.Y(g24336),.A(I31682));
  NOT NOT1_9240(.VSS(VSS),.VDD(VDD),.Y(I31685),.A(g23626));
  NOT NOT1_9241(.VSS(VSS),.VDD(VDD),.Y(g24337),.A(I31685));
  NOT NOT1_9242(.VSS(VSS),.VDD(VDD),.Y(I31688),.A(g24035));
  NOT NOT1_9243(.VSS(VSS),.VDD(VDD),.Y(g24338),.A(I31688));
  NOT NOT1_9244(.VSS(VSS),.VDD(VDD),.Y(I31691),.A(g24053));
  NOT NOT1_9245(.VSS(VSS),.VDD(VDD),.Y(g24339),.A(I31691));
  NOT NOT1_9246(.VSS(VSS),.VDD(VDD),.Y(I31694),.A(g24064));
  NOT NOT1_9247(.VSS(VSS),.VDD(VDD),.Y(g24340),.A(I31694));
  NOT NOT1_9248(.VSS(VSS),.VDD(VDD),.Y(I31697),.A(g23791));
  NOT NOT1_9249(.VSS(VSS),.VDD(VDD),.Y(g24341),.A(I31697));
  NOT NOT1_9250(.VSS(VSS),.VDD(VDD),.Y(I31700),.A(g23835));
  NOT NOT1_9251(.VSS(VSS),.VDD(VDD),.Y(g24342),.A(I31700));
  NOT NOT1_9252(.VSS(VSS),.VDD(VDD),.Y(I31703),.A(g23861));
  NOT NOT1_9253(.VSS(VSS),.VDD(VDD),.Y(g24343),.A(I31703));
  NOT NOT1_9254(.VSS(VSS),.VDD(VDD),.Y(I31706),.A(g23836));
  NOT NOT1_9255(.VSS(VSS),.VDD(VDD),.Y(g24344),.A(I31706));
  NOT NOT1_9256(.VSS(VSS),.VDD(VDD),.Y(I31709),.A(g23862));
  NOT NOT1_9257(.VSS(VSS),.VDD(VDD),.Y(g24345),.A(I31709));
  NOT NOT1_9258(.VSS(VSS),.VDD(VDD),.Y(I31712),.A(g23890));
  NOT NOT1_9259(.VSS(VSS),.VDD(VDD),.Y(g24346),.A(I31712));
  NOT NOT1_9260(.VSS(VSS),.VDD(VDD),.Y(I31715),.A(g23566));
  NOT NOT1_9261(.VSS(VSS),.VDD(VDD),.Y(g24347),.A(I31715));
  NOT NOT1_9262(.VSS(VSS),.VDD(VDD),.Y(I31718),.A(g23580));
  NOT NOT1_9263(.VSS(VSS),.VDD(VDD),.Y(g24348),.A(I31718));
  NOT NOT1_9264(.VSS(VSS),.VDD(VDD),.Y(I31721),.A(g23601));
  NOT NOT1_9265(.VSS(VSS),.VDD(VDD),.Y(g24349),.A(I31721));
  NOT NOT1_9266(.VSS(VSS),.VDD(VDD),.Y(I31724),.A(g23581));
  NOT NOT1_9267(.VSS(VSS),.VDD(VDD),.Y(g24350),.A(I31724));
  NOT NOT1_9268(.VSS(VSS),.VDD(VDD),.Y(I31727),.A(g23602));
  NOT NOT1_9269(.VSS(VSS),.VDD(VDD),.Y(g24351),.A(I31727));
  NOT NOT1_9270(.VSS(VSS),.VDD(VDD),.Y(I31730),.A(g23627));
  NOT NOT1_9271(.VSS(VSS),.VDD(VDD),.Y(g24352),.A(I31730));
  NOT NOT1_9272(.VSS(VSS),.VDD(VDD),.Y(I31733),.A(g23603));
  NOT NOT1_9273(.VSS(VSS),.VDD(VDD),.Y(g24353),.A(I31733));
  NOT NOT1_9274(.VSS(VSS),.VDD(VDD),.Y(I31736),.A(g23628));
  NOT NOT1_9275(.VSS(VSS),.VDD(VDD),.Y(g24354),.A(I31736));
  NOT NOT1_9276(.VSS(VSS),.VDD(VDD),.Y(I31739),.A(g23668));
  NOT NOT1_9277(.VSS(VSS),.VDD(VDD),.Y(g24355),.A(I31739));
  NOT NOT1_9278(.VSS(VSS),.VDD(VDD),.Y(I31742),.A(g23629));
  NOT NOT1_9279(.VSS(VSS),.VDD(VDD),.Y(g24356),.A(I31742));
  NOT NOT1_9280(.VSS(VSS),.VDD(VDD),.Y(I31745),.A(g23669));
  NOT NOT1_9281(.VSS(VSS),.VDD(VDD),.Y(g24357),.A(I31745));
  NOT NOT1_9282(.VSS(VSS),.VDD(VDD),.Y(I31748),.A(g23711));
  NOT NOT1_9283(.VSS(VSS),.VDD(VDD),.Y(g24358),.A(I31748));
  NOT NOT1_9284(.VSS(VSS),.VDD(VDD),.Y(I31751),.A(g23670));
  NOT NOT1_9285(.VSS(VSS),.VDD(VDD),.Y(g24359),.A(I31751));
  NOT NOT1_9286(.VSS(VSS),.VDD(VDD),.Y(I31754),.A(g23712));
  NOT NOT1_9287(.VSS(VSS),.VDD(VDD),.Y(g24360),.A(I31754));
  NOT NOT1_9288(.VSS(VSS),.VDD(VDD),.Y(I31757),.A(g23744));
  NOT NOT1_9289(.VSS(VSS),.VDD(VDD),.Y(g24361),.A(I31757));
  NOT NOT1_9290(.VSS(VSS),.VDD(VDD),.Y(I31760),.A(g23713));
  NOT NOT1_9291(.VSS(VSS),.VDD(VDD),.Y(g24362),.A(I31760));
  NOT NOT1_9292(.VSS(VSS),.VDD(VDD),.Y(I31763),.A(g23745));
  NOT NOT1_9293(.VSS(VSS),.VDD(VDD),.Y(g24363),.A(I31763));
  NOT NOT1_9294(.VSS(VSS),.VDD(VDD),.Y(I31766),.A(g23792));
  NOT NOT1_9295(.VSS(VSS),.VDD(VDD),.Y(g24364),.A(I31766));
  NOT NOT1_9296(.VSS(VSS),.VDD(VDD),.Y(I31769),.A(g23746));
  NOT NOT1_9297(.VSS(VSS),.VDD(VDD),.Y(g24365),.A(I31769));
  NOT NOT1_9298(.VSS(VSS),.VDD(VDD),.Y(I31772),.A(g23793));
  NOT NOT1_9299(.VSS(VSS),.VDD(VDD),.Y(g24366),.A(I31772));
  NOT NOT1_9300(.VSS(VSS),.VDD(VDD),.Y(I31775),.A(g23837));
  NOT NOT1_9301(.VSS(VSS),.VDD(VDD),.Y(g24367),.A(I31775));
  NOT NOT1_9302(.VSS(VSS),.VDD(VDD),.Y(I31778),.A(g23794));
  NOT NOT1_9303(.VSS(VSS),.VDD(VDD),.Y(g24368),.A(I31778));
  NOT NOT1_9304(.VSS(VSS),.VDD(VDD),.Y(I31781),.A(g23838));
  NOT NOT1_9305(.VSS(VSS),.VDD(VDD),.Y(g24369),.A(I31781));
  NOT NOT1_9306(.VSS(VSS),.VDD(VDD),.Y(I31784),.A(g23863));
  NOT NOT1_9307(.VSS(VSS),.VDD(VDD),.Y(g24370),.A(I31784));
  NOT NOT1_9308(.VSS(VSS),.VDD(VDD),.Y(I31787),.A(g23531));
  NOT NOT1_9309(.VSS(VSS),.VDD(VDD),.Y(g24371),.A(I31787));
  NOT NOT1_9310(.VSS(VSS),.VDD(VDD),.Y(I31790),.A(g23459));
  NOT NOT1_9311(.VSS(VSS),.VDD(VDD),.Y(g24372),.A(I31790));
  NOT NOT1_9312(.VSS(VSS),.VDD(VDD),.Y(I31793),.A(g23472));
  NOT NOT1_9313(.VSS(VSS),.VDD(VDD),.Y(g24373),.A(I31793));
  NOT NOT1_9314(.VSS(VSS),.VDD(VDD),.Y(I31796),.A(g23508));
  NOT NOT1_9315(.VSS(VSS),.VDD(VDD),.Y(g24374),.A(I31796));
  NOT NOT1_9316(.VSS(VSS),.VDD(VDD),.Y(I31799),.A(g23532));
  NOT NOT1_9317(.VSS(VSS),.VDD(VDD),.Y(g24375),.A(I31799));
  NOT NOT1_9318(.VSS(VSS),.VDD(VDD),.Y(I31802),.A(g23460));
  NOT NOT1_9319(.VSS(VSS),.VDD(VDD),.Y(g24376),.A(I31802));
  NOT NOT1_9320(.VSS(VSS),.VDD(VDD),.Y(I31805),.A(g24248));
  NOT NOT1_9321(.VSS(VSS),.VDD(VDD),.Y(g24377),.A(I31805));
  NOT NOT1_9322(.VSS(VSS),.VDD(VDD),.Y(I31808),.A(g23675));
  NOT NOT1_9323(.VSS(VSS),.VDD(VDD),.Y(g24378),.A(I31808));
  NOT NOT1_9324(.VSS(VSS),.VDD(VDD),.Y(I31811),.A(g24055));
  NOT NOT1_9325(.VSS(VSS),.VDD(VDD),.Y(g24379),.A(I31811));
  NOT NOT1_9326(.VSS(VSS),.VDD(VDD),.Y(I31814),.A(g24066));
  NOT NOT1_9327(.VSS(VSS),.VDD(VDD),.Y(g24380),.A(I31814));
  NOT NOT1_9328(.VSS(VSS),.VDD(VDD),.Y(I31817),.A(g24077));
  NOT NOT1_9329(.VSS(VSS),.VDD(VDD),.Y(g24381),.A(I31817));
  NOT NOT1_9330(.VSS(VSS),.VDD(VDD),.Y(I31820),.A(g23844));
  NOT NOT1_9331(.VSS(VSS),.VDD(VDD),.Y(g24382),.A(I31820));
  NOT NOT1_9332(.VSS(VSS),.VDD(VDD),.Y(I31823),.A(g23870));
  NOT NOT1_9333(.VSS(VSS),.VDD(VDD),.Y(g24383),.A(I31823));
  NOT NOT1_9334(.VSS(VSS),.VDD(VDD),.Y(I31826),.A(g23895));
  NOT NOT1_9335(.VSS(VSS),.VDD(VDD),.Y(g24384),.A(I31826));
  NOT NOT1_9336(.VSS(VSS),.VDD(VDD),.Y(I31829),.A(g23871));
  NOT NOT1_9337(.VSS(VSS),.VDD(VDD),.Y(g24385),.A(I31829));
  NOT NOT1_9338(.VSS(VSS),.VDD(VDD),.Y(I31832),.A(g23896));
  NOT NOT1_9339(.VSS(VSS),.VDD(VDD),.Y(g24386),.A(I31832));
  NOT NOT1_9340(.VSS(VSS),.VDD(VDD),.Y(I31835),.A(g23911));
  NOT NOT1_9341(.VSS(VSS),.VDD(VDD),.Y(g24387),.A(I31835));
  NOT NOT1_9342(.VSS(VSS),.VDD(VDD),.Y(I31838),.A(g23585));
  NOT NOT1_9343(.VSS(VSS),.VDD(VDD),.Y(g24388),.A(I31838));
  NOT NOT1_9344(.VSS(VSS),.VDD(VDD),.Y(I31841),.A(g23607));
  NOT NOT1_9345(.VSS(VSS),.VDD(VDD),.Y(g24389),.A(I31841));
  NOT NOT1_9346(.VSS(VSS),.VDD(VDD),.Y(I31844),.A(g23633));
  NOT NOT1_9347(.VSS(VSS),.VDD(VDD),.Y(g24390),.A(I31844));
  NOT NOT1_9348(.VSS(VSS),.VDD(VDD),.Y(I31847),.A(g23608));
  NOT NOT1_9349(.VSS(VSS),.VDD(VDD),.Y(g24391),.A(I31847));
  NOT NOT1_9350(.VSS(VSS),.VDD(VDD),.Y(I31850),.A(g23634));
  NOT NOT1_9351(.VSS(VSS),.VDD(VDD),.Y(g24392),.A(I31850));
  NOT NOT1_9352(.VSS(VSS),.VDD(VDD),.Y(I31853),.A(g23676));
  NOT NOT1_9353(.VSS(VSS),.VDD(VDD),.Y(g24393),.A(I31853));
  NOT NOT1_9354(.VSS(VSS),.VDD(VDD),.Y(I31856),.A(g23635));
  NOT NOT1_9355(.VSS(VSS),.VDD(VDD),.Y(g24394),.A(I31856));
  NOT NOT1_9356(.VSS(VSS),.VDD(VDD),.Y(I31859),.A(g23677));
  NOT NOT1_9357(.VSS(VSS),.VDD(VDD),.Y(g24395),.A(I31859));
  NOT NOT1_9358(.VSS(VSS),.VDD(VDD),.Y(I31862),.A(g23718));
  NOT NOT1_9359(.VSS(VSS),.VDD(VDD),.Y(g24396),.A(I31862));
  NOT NOT1_9360(.VSS(VSS),.VDD(VDD),.Y(I31865),.A(g23678));
  NOT NOT1_9361(.VSS(VSS),.VDD(VDD),.Y(g24397),.A(I31865));
  NOT NOT1_9362(.VSS(VSS),.VDD(VDD),.Y(I31868),.A(g23719));
  NOT NOT1_9363(.VSS(VSS),.VDD(VDD),.Y(g24398),.A(I31868));
  NOT NOT1_9364(.VSS(VSS),.VDD(VDD),.Y(I31871),.A(g23765));
  NOT NOT1_9365(.VSS(VSS),.VDD(VDD),.Y(g24399),.A(I31871));
  NOT NOT1_9366(.VSS(VSS),.VDD(VDD),.Y(I31874),.A(g23720));
  NOT NOT1_9367(.VSS(VSS),.VDD(VDD),.Y(g24400),.A(I31874));
  NOT NOT1_9368(.VSS(VSS),.VDD(VDD),.Y(I31877),.A(g23766));
  NOT NOT1_9369(.VSS(VSS),.VDD(VDD),.Y(g24401),.A(I31877));
  NOT NOT1_9370(.VSS(VSS),.VDD(VDD),.Y(I31880),.A(g23799));
  NOT NOT1_9371(.VSS(VSS),.VDD(VDD),.Y(g24402),.A(I31880));
  NOT NOT1_9372(.VSS(VSS),.VDD(VDD),.Y(I31883),.A(g23767));
  NOT NOT1_9373(.VSS(VSS),.VDD(VDD),.Y(g24403),.A(I31883));
  NOT NOT1_9374(.VSS(VSS),.VDD(VDD),.Y(I31886),.A(g23800));
  NOT NOT1_9375(.VSS(VSS),.VDD(VDD),.Y(g24404),.A(I31886));
  NOT NOT1_9376(.VSS(VSS),.VDD(VDD),.Y(I31889),.A(g23845));
  NOT NOT1_9377(.VSS(VSS),.VDD(VDD),.Y(g24405),.A(I31889));
  NOT NOT1_9378(.VSS(VSS),.VDD(VDD),.Y(I31892),.A(g23801));
  NOT NOT1_9379(.VSS(VSS),.VDD(VDD),.Y(g24406),.A(I31892));
  NOT NOT1_9380(.VSS(VSS),.VDD(VDD),.Y(I31895),.A(g23846));
  NOT NOT1_9381(.VSS(VSS),.VDD(VDD),.Y(g24407),.A(I31895));
  NOT NOT1_9382(.VSS(VSS),.VDD(VDD),.Y(I31898),.A(g23872));
  NOT NOT1_9383(.VSS(VSS),.VDD(VDD),.Y(g24408),.A(I31898));
  NOT NOT1_9384(.VSS(VSS),.VDD(VDD),.Y(I31901),.A(g23847));
  NOT NOT1_9385(.VSS(VSS),.VDD(VDD),.Y(g24409),.A(I31901));
  NOT NOT1_9386(.VSS(VSS),.VDD(VDD),.Y(I31904),.A(g23873));
  NOT NOT1_9387(.VSS(VSS),.VDD(VDD),.Y(g24410),.A(I31904));
  NOT NOT1_9388(.VSS(VSS),.VDD(VDD),.Y(I31907),.A(g23897));
  NOT NOT1_9389(.VSS(VSS),.VDD(VDD),.Y(g24411),.A(I31907));
  NOT NOT1_9390(.VSS(VSS),.VDD(VDD),.Y(I31910),.A(g23542));
  NOT NOT1_9391(.VSS(VSS),.VDD(VDD),.Y(g24412),.A(I31910));
  NOT NOT1_9392(.VSS(VSS),.VDD(VDD),.Y(I31913),.A(g23468));
  NOT NOT1_9393(.VSS(VSS),.VDD(VDD),.Y(g24413),.A(I31913));
  NOT NOT1_9394(.VSS(VSS),.VDD(VDD),.Y(I31916),.A(g23485));
  NOT NOT1_9395(.VSS(VSS),.VDD(VDD),.Y(g24414),.A(I31916));
  NOT NOT1_9396(.VSS(VSS),.VDD(VDD),.Y(I31919),.A(g23524));
  NOT NOT1_9397(.VSS(VSS),.VDD(VDD),.Y(g24415),.A(I31919));
  NOT NOT1_9398(.VSS(VSS),.VDD(VDD),.Y(I31922),.A(g23543));
  NOT NOT1_9399(.VSS(VSS),.VDD(VDD),.Y(g24416),.A(I31922));
  NOT NOT1_9400(.VSS(VSS),.VDD(VDD),.Y(I31925),.A(g23469));
  NOT NOT1_9401(.VSS(VSS),.VDD(VDD),.Y(g24417),.A(I31925));
  NOT NOT1_9402(.VSS(VSS),.VDD(VDD),.Y(I31928),.A(g24255));
  NOT NOT1_9403(.VSS(VSS),.VDD(VDD),.Y(g24418),.A(I31928));
  NOT NOT1_9404(.VSS(VSS),.VDD(VDD),.Y(I31931),.A(g23725));
  NOT NOT1_9405(.VSS(VSS),.VDD(VDD),.Y(g24419),.A(I31931));
  NOT NOT1_9406(.VSS(VSS),.VDD(VDD),.Y(I31934),.A(g24068));
  NOT NOT1_9407(.VSS(VSS),.VDD(VDD),.Y(g24420),.A(I31934));
  NOT NOT1_9408(.VSS(VSS),.VDD(VDD),.Y(I31937),.A(g24079));
  NOT NOT1_9409(.VSS(VSS),.VDD(VDD),.Y(g24421),.A(I31937));
  NOT NOT1_9410(.VSS(VSS),.VDD(VDD),.Y(I31940),.A(g24088));
  NOT NOT1_9411(.VSS(VSS),.VDD(VDD),.Y(g24422),.A(I31940));
  NOT NOT1_9412(.VSS(VSS),.VDD(VDD),.Y(I31943),.A(g24000));
  NOT NOT1_9413(.VSS(VSS),.VDD(VDD),.Y(g24423),.A(I31943));
  NOT NOT1_9414(.VSS(VSS),.VDD(VDD),.Y(I31946),.A(g23916));
  NOT NOT1_9415(.VSS(VSS),.VDD(VDD),.Y(g24424),.A(I31946));
  NOT NOT1_9416(.VSS(VSS),.VDD(VDD),.Y(I31949),.A(g23943));
  NOT NOT1_9417(.VSS(VSS),.VDD(VDD),.Y(g24425),.A(I31949));
  NOT NOT1_9418(.VSS(VSS),.VDD(VDD),.Y(g24482),.A(g24183));
  NOT NOT1_9419(.VSS(VSS),.VDD(VDD),.Y(I32042),.A(g23399));
  NOT NOT1_9420(.VSS(VSS),.VDD(VDD),.Y(g24518),.A(I32042));
  NOT NOT1_9421(.VSS(VSS),.VDD(VDD),.Y(I32057),.A(g23406));
  NOT NOT1_9422(.VSS(VSS),.VDD(VDD),.Y(g24531),.A(I32057));
  NOT NOT1_9423(.VSS(VSS),.VDD(VDD),.Y(I32067),.A(g24174));
  NOT NOT1_9424(.VSS(VSS),.VDD(VDD),.Y(g24539),.A(I32067));
  NOT NOT1_9425(.VSS(VSS),.VDD(VDD),.Y(I32074),.A(g23413));
  NOT NOT1_9426(.VSS(VSS),.VDD(VDD),.Y(g24544),.A(I32074));
  NOT NOT1_9427(.VSS(VSS),.VDD(VDD),.Y(I32081),.A(g24178));
  NOT NOT1_9428(.VSS(VSS),.VDD(VDD),.Y(g24549),.A(I32081));
  NOT NOT1_9429(.VSS(VSS),.VDD(VDD),.Y(I32085),.A(g24179));
  NOT NOT1_9430(.VSS(VSS),.VDD(VDD),.Y(g24551),.A(I32085));
  NOT NOT1_9431(.VSS(VSS),.VDD(VDD),.Y(I32092),.A(g23418));
  NOT NOT1_9432(.VSS(VSS),.VDD(VDD),.Y(g24556),.A(I32092));
  NOT NOT1_9433(.VSS(VSS),.VDD(VDD),.Y(I32098),.A(g24181));
  NOT NOT1_9434(.VSS(VSS),.VDD(VDD),.Y(g24560),.A(I32098));
  NOT NOT1_9435(.VSS(VSS),.VDD(VDD),.Y(I32102),.A(g24182));
  NOT NOT1_9436(.VSS(VSS),.VDD(VDD),.Y(g24562),.A(I32102));
  NOT NOT1_9437(.VSS(VSS),.VDD(VDD),.Y(I32109),.A(g24206));
  NOT NOT1_9438(.VSS(VSS),.VDD(VDD),.Y(g24567),.A(I32109));
  NOT NOT1_9439(.VSS(VSS),.VDD(VDD),.Y(I32112),.A(g24207));
  NOT NOT1_9440(.VSS(VSS),.VDD(VDD),.Y(g24568),.A(I32112));
  NOT NOT1_9441(.VSS(VSS),.VDD(VDD),.Y(I32116),.A(g24208));
  NOT NOT1_9442(.VSS(VSS),.VDD(VDD),.Y(g24570),.A(I32116));
  NOT NOT1_9443(.VSS(VSS),.VDD(VDD),.Y(I32120),.A(g24209));
  NOT NOT1_9444(.VSS(VSS),.VDD(VDD),.Y(g24572),.A(I32120));
  NOT NOT1_9445(.VSS(VSS),.VDD(VDD),.Y(I32126),.A(g24212));
  NOT NOT1_9446(.VSS(VSS),.VDD(VDD),.Y(g24576),.A(I32126));
  NOT NOT1_9447(.VSS(VSS),.VDD(VDD),.Y(I32129),.A(g24213));
  NOT NOT1_9448(.VSS(VSS),.VDD(VDD),.Y(g24577),.A(I32129));
  NOT NOT1_9449(.VSS(VSS),.VDD(VDD),.Y(I32133),.A(g24214));
  NOT NOT1_9450(.VSS(VSS),.VDD(VDD),.Y(g24579),.A(I32133));
  NOT NOT1_9451(.VSS(VSS),.VDD(VDD),.Y(I32137),.A(g24215));
  NOT NOT1_9452(.VSS(VSS),.VDD(VDD),.Y(g24581),.A(I32137));
  NOT NOT1_9453(.VSS(VSS),.VDD(VDD),.Y(I32140),.A(g24216));
  NOT NOT1_9454(.VSS(VSS),.VDD(VDD),.Y(g24582),.A(I32140));
  NOT NOT1_9455(.VSS(VSS),.VDD(VDD),.Y(I32143),.A(g24218));
  NOT NOT1_9456(.VSS(VSS),.VDD(VDD),.Y(g24583),.A(I32143));
  NOT NOT1_9457(.VSS(VSS),.VDD(VDD),.Y(I32146),.A(g24219));
  NOT NOT1_9458(.VSS(VSS),.VDD(VDD),.Y(g24584),.A(I32146));
  NOT NOT1_9459(.VSS(VSS),.VDD(VDD),.Y(I32150),.A(g24222));
  NOT NOT1_9460(.VSS(VSS),.VDD(VDD),.Y(g24586),.A(I32150));
  NOT NOT1_9461(.VSS(VSS),.VDD(VDD),.Y(I32153),.A(g24223));
  NOT NOT1_9462(.VSS(VSS),.VDD(VDD),.Y(g24587),.A(I32153));
  NOT NOT1_9463(.VSS(VSS),.VDD(VDD),.Y(I32156),.A(g24225));
  NOT NOT1_9464(.VSS(VSS),.VDD(VDD),.Y(g24588),.A(I32156));
  NOT NOT1_9465(.VSS(VSS),.VDD(VDD),.Y(I32159),.A(g24226));
  NOT NOT1_9466(.VSS(VSS),.VDD(VDD),.Y(g24589),.A(I32159));
  NOT NOT1_9467(.VSS(VSS),.VDD(VDD),.Y(I32164),.A(g24228));
  NOT NOT1_9468(.VSS(VSS),.VDD(VDD),.Y(g24592),.A(I32164));
  NOT NOT1_9469(.VSS(VSS),.VDD(VDD),.Y(I32167),.A(g24230));
  NOT NOT1_9470(.VSS(VSS),.VDD(VDD),.Y(g24593),.A(I32167));
  NOT NOT1_9471(.VSS(VSS),.VDD(VDD),.Y(I32170),.A(g24231));
  NOT NOT1_9472(.VSS(VSS),.VDD(VDD),.Y(g24594),.A(I32170));
  NOT NOT1_9473(.VSS(VSS),.VDD(VDD),.Y(I32175),.A(g24235));
  NOT NOT1_9474(.VSS(VSS),.VDD(VDD),.Y(g24597),.A(I32175));
  NOT NOT1_9475(.VSS(VSS),.VDD(VDD),.Y(I32178),.A(g24237));
  NOT NOT1_9476(.VSS(VSS),.VDD(VDD),.Y(g24598),.A(I32178));
  NOT NOT1_9477(.VSS(VSS),.VDD(VDD),.Y(I32181),.A(g24238));
  NOT NOT1_9478(.VSS(VSS),.VDD(VDD),.Y(g24599),.A(I32181));
  NOT NOT1_9479(.VSS(VSS),.VDD(VDD),.Y(I32184),.A(g23497));
  NOT NOT1_9480(.VSS(VSS),.VDD(VDD),.Y(g24600),.A(I32184));
  NOT NOT1_9481(.VSS(VSS),.VDD(VDD),.Y(I32189),.A(g24243));
  NOT NOT1_9482(.VSS(VSS),.VDD(VDD),.Y(g24605),.A(I32189));
  NOT NOT1_9483(.VSS(VSS),.VDD(VDD),.Y(I32193),.A(g23513));
  NOT NOT1_9484(.VSS(VSS),.VDD(VDD),.Y(g24607),.A(I32193));
  NOT NOT1_9485(.VSS(VSS),.VDD(VDD),.Y(I32198),.A(g24250));
  NOT NOT1_9486(.VSS(VSS),.VDD(VDD),.Y(g24612),.A(I32198));
  NOT NOT1_9487(.VSS(VSS),.VDD(VDD),.Y(I32203),.A(g23528));
  NOT NOT1_9488(.VSS(VSS),.VDD(VDD),.Y(g24619),.A(I32203));
  NOT NOT1_9489(.VSS(VSS),.VDD(VDD),.Y(I32210),.A(g23539));
  NOT NOT1_9490(.VSS(VSS),.VDD(VDD),.Y(g24630),.A(I32210));
  NOT NOT1_9491(.VSS(VSS),.VDD(VDD),.Y(g24648),.A(g23470));
  NOT NOT1_9492(.VSS(VSS),.VDD(VDD),.Y(g24668),.A(g23482));
  NOT NOT1_9493(.VSS(VSS),.VDD(VDD),.Y(g24687),.A(g23493));
  NOT NOT1_9494(.VSS(VSS),.VDD(VDD),.Y(g24704),.A(g23509));
  NOT NOT1_9495(.VSS(VSS),.VDD(VDD),.Y(I32248),.A(g23919));
  NOT NOT1_9496(.VSS(VSS),.VDD(VDD),.Y(g24734),.A(I32248));
  NOT NOT1_9497(.VSS(VSS),.VDD(VDD),.Y(I32251),.A(g23919));
  NOT NOT1_9498(.VSS(VSS),.VDD(VDD),.Y(g24735),.A(I32251));
  NOT NOT1_9499(.VSS(VSS),.VDD(VDD),.Y(I32281),.A(g23950));
  NOT NOT1_9500(.VSS(VSS),.VDD(VDD),.Y(g24763),.A(I32281));
  NOT NOT1_9501(.VSS(VSS),.VDD(VDD),.Y(I32320),.A(g23979));
  NOT NOT1_9502(.VSS(VSS),.VDD(VDD),.Y(g24784),.A(I32320));
  NOT NOT1_9503(.VSS(VSS),.VDD(VDD),.Y(I32365),.A(g24009));
  NOT NOT1_9504(.VSS(VSS),.VDD(VDD),.Y(g24805),.A(I32365));
  NOT NOT1_9505(.VSS(VSS),.VDD(VDD),.Y(g24815),.A(g23448));
  NOT NOT1_9506(.VSS(VSS),.VDD(VDD),.Y(I32388),.A(g23385));
  NOT NOT1_9507(.VSS(VSS),.VDD(VDD),.Y(g24816),.A(I32388));
  NOT NOT1_9508(.VSS(VSS),.VDD(VDD),.Y(I32419),.A(g24043));
  NOT NOT1_9509(.VSS(VSS),.VDD(VDD),.Y(g24827),.A(I32419));
  NOT NOT1_9510(.VSS(VSS),.VDD(VDD),.Y(g24834),.A(g23455));
  NOT NOT1_9511(.VSS(VSS),.VDD(VDD),.Y(I32439),.A(g23392));
  NOT NOT1_9512(.VSS(VSS),.VDD(VDD),.Y(g24835),.A(I32439));
  NOT NOT1_9513(.VSS(VSS),.VDD(VDD),.Y(g24850),.A(g23464));
  NOT NOT1_9514(.VSS(VSS),.VDD(VDD),.Y(I32487),.A(g23400));
  NOT NOT1_9515(.VSS(VSS),.VDD(VDD),.Y(g24851),.A(I32487));
  NOT NOT1_9516(.VSS(VSS),.VDD(VDD),.Y(I32506),.A(g23324));
  NOT NOT1_9517(.VSS(VSS),.VDD(VDD),.Y(g24856),.A(I32506));
  NOT NOT1_9518(.VSS(VSS),.VDD(VDD),.Y(g24864),.A(g23473));
  NOT NOT1_9519(.VSS(VSS),.VDD(VDD),.Y(I32535),.A(g23407));
  NOT NOT1_9520(.VSS(VSS),.VDD(VDD),.Y(g24865),.A(I32535));
  NOT NOT1_9521(.VSS(VSS),.VDD(VDD),.Y(I32556),.A(g23329));
  NOT NOT1_9522(.VSS(VSS),.VDD(VDD),.Y(g24872),.A(I32556));
  NOT NOT1_9523(.VSS(VSS),.VDD(VDD),.Y(I32583),.A(g23330));
  NOT NOT1_9524(.VSS(VSS),.VDD(VDD),.Y(g24879),.A(I32583));
  NOT NOT1_9525(.VSS(VSS),.VDD(VDD),.Y(I32604),.A(g23339));
  NOT NOT1_9526(.VSS(VSS),.VDD(VDD),.Y(g24886),.A(I32604));
  NOT NOT1_9527(.VSS(VSS),.VDD(VDD),.Y(g24893),.A(g23486));
  NOT NOT1_9528(.VSS(VSS),.VDD(VDD),.Y(I32642),.A(g23348));
  NOT NOT1_9529(.VSS(VSS),.VDD(VDD),.Y(g24903),.A(I32642));
  NOT NOT1_9530(.VSS(VSS),.VDD(VDD),.Y(g24912),.A(g23495));
  NOT NOT1_9531(.VSS(VSS),.VDD(VDD),.Y(g24916),.A(g23502));
  NOT NOT1_9532(.VSS(VSS),.VDD(VDD),.Y(g24929),.A(g23511));
  NOT NOT1_9533(.VSS(VSS),.VDD(VDD),.Y(g24933),.A(g23518));
  NOT NOT1_9534(.VSS(VSS),.VDD(VDD),.Y(g24939),.A(g23660));
  NOT NOT1_9535(.VSS(VSS),.VDD(VDD),.Y(g24941),.A(g23526));
  NOT NOT1_9536(.VSS(VSS),.VDD(VDD),.Y(g24945),.A(g23533));
  NOT NOT1_9537(.VSS(VSS),.VDD(VDD),.Y(I32704),.A(g23357));
  NOT NOT1_9538(.VSS(VSS),.VDD(VDD),.Y(g24949),.A(I32704));
  NOT NOT1_9539(.VSS(VSS),.VDD(VDD),.Y(g24950),.A(g23710));
  NOT NOT1_9540(.VSS(VSS),.VDD(VDD),.Y(g24952),.A(g23537));
  NOT NOT1_9541(.VSS(VSS),.VDD(VDD),.Y(I32716),.A(g23358));
  NOT NOT1_9542(.VSS(VSS),.VDD(VDD),.Y(g24956),.A(I32716));
  NOT NOT1_9543(.VSS(VSS),.VDD(VDD),.Y(I32719),.A(g23359));
  NOT NOT1_9544(.VSS(VSS),.VDD(VDD),.Y(g24957),.A(I32719));
  NOT NOT1_9545(.VSS(VSS),.VDD(VDD),.Y(g24958),.A(g23478));
  NOT NOT1_9546(.VSS(VSS),.VDD(VDD),.Y(g24962),.A(g23764));
  NOT NOT1_9547(.VSS(VSS),.VDD(VDD),.Y(g24969),.A(g23489));
  NOT NOT1_9548(.VSS(VSS),.VDD(VDD),.Y(g24973),.A(g23819));
  NOT NOT1_9549(.VSS(VSS),.VDD(VDD),.Y(g24982),.A(g23505));
  NOT NOT1_9550(.VSS(VSS),.VDD(VDD),.Y(g24993),.A(g23521));
  NOT NOT1_9551(.VSS(VSS),.VDD(VDD),.Y(g25087),.A(g23731));
  NOT NOT1_9552(.VSS(VSS),.VDD(VDD),.Y(g25094),.A(g23779));
  NOT NOT1_9553(.VSS(VSS),.VDD(VDD),.Y(g25095),.A(g23786));
  NOT NOT1_9554(.VSS(VSS),.VDD(VDD),.Y(I32829),.A(g24059));
  NOT NOT1_9555(.VSS(VSS),.VDD(VDD),.Y(g25103),.A(I32829));
  NOT NOT1_9556(.VSS(VSS),.VDD(VDD),.Y(g25104),.A(g23832));
  NOT NOT1_9557(.VSS(VSS),.VDD(VDD),.Y(g25105),.A(g23839));
  NOT NOT1_9558(.VSS(VSS),.VDD(VDD),.Y(I32835),.A(g24072));
  NOT NOT1_9559(.VSS(VSS),.VDD(VDD),.Y(g25109),.A(I32835));
  NOT NOT1_9560(.VSS(VSS),.VDD(VDD),.Y(g25110),.A(g23867));
  NOT NOT1_9561(.VSS(VSS),.VDD(VDD),.Y(g25111),.A(g23874));
  NOT NOT1_9562(.VSS(VSS),.VDD(VDD),.Y(g25115),.A(g23879));
  NOT NOT1_9563(.VSS(VSS),.VDD(VDD),.Y(g25116),.A(g23882));
  NOT NOT1_9564(.VSS(VSS),.VDD(VDD),.Y(I32844),.A(g23644));
  NOT NOT1_9565(.VSS(VSS),.VDD(VDD),.Y(g25118),.A(I32844));
  NOT NOT1_9566(.VSS(VSS),.VDD(VDD),.Y(I32847),.A(g24083));
  NOT NOT1_9567(.VSS(VSS),.VDD(VDD),.Y(g25119),.A(I32847));
  NOT NOT1_9568(.VSS(VSS),.VDD(VDD),.Y(g25120),.A(g23901));
  NOT NOT1_9569(.VSS(VSS),.VDD(VDD),.Y(I32851),.A(g23694));
  NOT NOT1_9570(.VSS(VSS),.VDD(VDD),.Y(g25121),.A(I32851));
  NOT NOT1_9571(.VSS(VSS),.VDD(VDD),.Y(I32854),.A(g24092));
  NOT NOT1_9572(.VSS(VSS),.VDD(VDD),.Y(g25122),.A(I32854));
  NOT NOT1_9573(.VSS(VSS),.VDD(VDD),.Y(I32857),.A(g23748));
  NOT NOT1_9574(.VSS(VSS),.VDD(VDD),.Y(g25123),.A(I32857));
  NOT NOT1_9575(.VSS(VSS),.VDD(VDD),.Y(I32860),.A(g23803));
  NOT NOT1_9576(.VSS(VSS),.VDD(VDD),.Y(g25124),.A(I32860));
  NOT NOT1_9577(.VSS(VSS),.VDD(VDD),.Y(g25126),.A(g24030));
  NOT NOT1_9578(.VSS(VSS),.VDD(VDD),.Y(I32868),.A(g25118));
  NOT NOT1_9579(.VSS(VSS),.VDD(VDD),.Y(g25130),.A(I32868));
  NOT NOT1_9580(.VSS(VSS),.VDD(VDD),.Y(I32871),.A(g24518));
  NOT NOT1_9581(.VSS(VSS),.VDD(VDD),.Y(g25131),.A(I32871));
  NOT NOT1_9582(.VSS(VSS),.VDD(VDD),.Y(I32874),.A(g24539));
  NOT NOT1_9583(.VSS(VSS),.VDD(VDD),.Y(g25132),.A(I32874));
  NOT NOT1_9584(.VSS(VSS),.VDD(VDD),.Y(I32877),.A(g24567));
  NOT NOT1_9585(.VSS(VSS),.VDD(VDD),.Y(g25133),.A(I32877));
  NOT NOT1_9586(.VSS(VSS),.VDD(VDD),.Y(I32880),.A(g24581));
  NOT NOT1_9587(.VSS(VSS),.VDD(VDD),.Y(g25134),.A(I32880));
  NOT NOT1_9588(.VSS(VSS),.VDD(VDD),.Y(I32883),.A(g24592));
  NOT NOT1_9589(.VSS(VSS),.VDD(VDD),.Y(g25135),.A(I32883));
  NOT NOT1_9590(.VSS(VSS),.VDD(VDD),.Y(I32886),.A(g24549));
  NOT NOT1_9591(.VSS(VSS),.VDD(VDD),.Y(g25136),.A(I32886));
  NOT NOT1_9592(.VSS(VSS),.VDD(VDD),.Y(I32889),.A(g24568));
  NOT NOT1_9593(.VSS(VSS),.VDD(VDD),.Y(g25137),.A(I32889));
  NOT NOT1_9594(.VSS(VSS),.VDD(VDD),.Y(I32892),.A(g24582));
  NOT NOT1_9595(.VSS(VSS),.VDD(VDD),.Y(g25138),.A(I32892));
  NOT NOT1_9596(.VSS(VSS),.VDD(VDD),.Y(I32895),.A(g24816));
  NOT NOT1_9597(.VSS(VSS),.VDD(VDD),.Y(g25139),.A(I32895));
  NOT NOT1_9598(.VSS(VSS),.VDD(VDD),.Y(I32898),.A(g24856));
  NOT NOT1_9599(.VSS(VSS),.VDD(VDD),.Y(g25140),.A(I32898));
  NOT NOT1_9600(.VSS(VSS),.VDD(VDD),.Y(I32901),.A(g25121));
  NOT NOT1_9601(.VSS(VSS),.VDD(VDD),.Y(g25141),.A(I32901));
  NOT NOT1_9602(.VSS(VSS),.VDD(VDD),.Y(I32904),.A(g24531));
  NOT NOT1_9603(.VSS(VSS),.VDD(VDD),.Y(g25142),.A(I32904));
  NOT NOT1_9604(.VSS(VSS),.VDD(VDD),.Y(I32907),.A(g24551));
  NOT NOT1_9605(.VSS(VSS),.VDD(VDD),.Y(g25143),.A(I32907));
  NOT NOT1_9606(.VSS(VSS),.VDD(VDD),.Y(I32910),.A(g24576));
  NOT NOT1_9607(.VSS(VSS),.VDD(VDD),.Y(g25144),.A(I32910));
  NOT NOT1_9608(.VSS(VSS),.VDD(VDD),.Y(I32913),.A(g24586));
  NOT NOT1_9609(.VSS(VSS),.VDD(VDD),.Y(g25145),.A(I32913));
  NOT NOT1_9610(.VSS(VSS),.VDD(VDD),.Y(I32916),.A(g24597));
  NOT NOT1_9611(.VSS(VSS),.VDD(VDD),.Y(g25146),.A(I32916));
  NOT NOT1_9612(.VSS(VSS),.VDD(VDD),.Y(I32919),.A(g24560));
  NOT NOT1_9613(.VSS(VSS),.VDD(VDD),.Y(g25147),.A(I32919));
  NOT NOT1_9614(.VSS(VSS),.VDD(VDD),.Y(I32922),.A(g24577));
  NOT NOT1_9615(.VSS(VSS),.VDD(VDD),.Y(g25148),.A(I32922));
  NOT NOT1_9616(.VSS(VSS),.VDD(VDD),.Y(I32925),.A(g24587));
  NOT NOT1_9617(.VSS(VSS),.VDD(VDD),.Y(g25149),.A(I32925));
  NOT NOT1_9618(.VSS(VSS),.VDD(VDD),.Y(I32928),.A(g24835));
  NOT NOT1_9619(.VSS(VSS),.VDD(VDD),.Y(g25150),.A(I32928));
  NOT NOT1_9620(.VSS(VSS),.VDD(VDD),.Y(I32931),.A(g24872));
  NOT NOT1_9621(.VSS(VSS),.VDD(VDD),.Y(g25151),.A(I32931));
  NOT NOT1_9622(.VSS(VSS),.VDD(VDD),.Y(I32934),.A(g25123));
  NOT NOT1_9623(.VSS(VSS),.VDD(VDD),.Y(g25152),.A(I32934));
  NOT NOT1_9624(.VSS(VSS),.VDD(VDD),.Y(I32937),.A(g24544));
  NOT NOT1_9625(.VSS(VSS),.VDD(VDD),.Y(g25153),.A(I32937));
  NOT NOT1_9626(.VSS(VSS),.VDD(VDD),.Y(I32940),.A(g24562));
  NOT NOT1_9627(.VSS(VSS),.VDD(VDD),.Y(g25154),.A(I32940));
  NOT NOT1_9628(.VSS(VSS),.VDD(VDD),.Y(I32943),.A(g24583));
  NOT NOT1_9629(.VSS(VSS),.VDD(VDD),.Y(g25155),.A(I32943));
  NOT NOT1_9630(.VSS(VSS),.VDD(VDD),.Y(I32946),.A(g24593));
  NOT NOT1_9631(.VSS(VSS),.VDD(VDD),.Y(g25156),.A(I32946));
  NOT NOT1_9632(.VSS(VSS),.VDD(VDD),.Y(I32949),.A(g24605));
  NOT NOT1_9633(.VSS(VSS),.VDD(VDD),.Y(g25157),.A(I32949));
  NOT NOT1_9634(.VSS(VSS),.VDD(VDD),.Y(I32952),.A(g24570));
  NOT NOT1_9635(.VSS(VSS),.VDD(VDD),.Y(g25158),.A(I32952));
  NOT NOT1_9636(.VSS(VSS),.VDD(VDD),.Y(I32955),.A(g24584));
  NOT NOT1_9637(.VSS(VSS),.VDD(VDD),.Y(g25159),.A(I32955));
  NOT NOT1_9638(.VSS(VSS),.VDD(VDD),.Y(I32958),.A(g24594));
  NOT NOT1_9639(.VSS(VSS),.VDD(VDD),.Y(g25160),.A(I32958));
  NOT NOT1_9640(.VSS(VSS),.VDD(VDD),.Y(I32961),.A(g24851));
  NOT NOT1_9641(.VSS(VSS),.VDD(VDD),.Y(g25161),.A(I32961));
  NOT NOT1_9642(.VSS(VSS),.VDD(VDD),.Y(I32964),.A(g24886));
  NOT NOT1_9643(.VSS(VSS),.VDD(VDD),.Y(g25162),.A(I32964));
  NOT NOT1_9644(.VSS(VSS),.VDD(VDD),.Y(I32967),.A(g25124));
  NOT NOT1_9645(.VSS(VSS),.VDD(VDD),.Y(g25163),.A(I32967));
  NOT NOT1_9646(.VSS(VSS),.VDD(VDD),.Y(I32970),.A(g24556));
  NOT NOT1_9647(.VSS(VSS),.VDD(VDD),.Y(g25164),.A(I32970));
  NOT NOT1_9648(.VSS(VSS),.VDD(VDD),.Y(I32973),.A(g24572));
  NOT NOT1_9649(.VSS(VSS),.VDD(VDD),.Y(g25165),.A(I32973));
  NOT NOT1_9650(.VSS(VSS),.VDD(VDD),.Y(I32976),.A(g24588));
  NOT NOT1_9651(.VSS(VSS),.VDD(VDD),.Y(g25166),.A(I32976));
  NOT NOT1_9652(.VSS(VSS),.VDD(VDD),.Y(I32979),.A(g24598));
  NOT NOT1_9653(.VSS(VSS),.VDD(VDD),.Y(g25167),.A(I32979));
  NOT NOT1_9654(.VSS(VSS),.VDD(VDD),.Y(I32982),.A(g24612));
  NOT NOT1_9655(.VSS(VSS),.VDD(VDD),.Y(g25168),.A(I32982));
  NOT NOT1_9656(.VSS(VSS),.VDD(VDD),.Y(I32985),.A(g24579));
  NOT NOT1_9657(.VSS(VSS),.VDD(VDD),.Y(g25169),.A(I32985));
  NOT NOT1_9658(.VSS(VSS),.VDD(VDD),.Y(I32988),.A(g24589));
  NOT NOT1_9659(.VSS(VSS),.VDD(VDD),.Y(g25170),.A(I32988));
  NOT NOT1_9660(.VSS(VSS),.VDD(VDD),.Y(I32991),.A(g24599));
  NOT NOT1_9661(.VSS(VSS),.VDD(VDD),.Y(g25171),.A(I32991));
  NOT NOT1_9662(.VSS(VSS),.VDD(VDD),.Y(I32994),.A(g24865));
  NOT NOT1_9663(.VSS(VSS),.VDD(VDD),.Y(g25172),.A(I32994));
  NOT NOT1_9664(.VSS(VSS),.VDD(VDD),.Y(I32997),.A(g24903));
  NOT NOT1_9665(.VSS(VSS),.VDD(VDD),.Y(g25173),.A(I32997));
  NOT NOT1_9666(.VSS(VSS),.VDD(VDD),.Y(I33000),.A(g24949));
  NOT NOT1_9667(.VSS(VSS),.VDD(VDD),.Y(g25174),.A(I33000));
  NOT NOT1_9668(.VSS(VSS),.VDD(VDD),.Y(I33003),.A(g24956));
  NOT NOT1_9669(.VSS(VSS),.VDD(VDD),.Y(g25175),.A(I33003));
  NOT NOT1_9670(.VSS(VSS),.VDD(VDD),.Y(I33006),.A(g24957));
  NOT NOT1_9671(.VSS(VSS),.VDD(VDD),.Y(g25176),.A(I33006));
  NOT NOT1_9672(.VSS(VSS),.VDD(VDD),.Y(I33009),.A(g24879));
  NOT NOT1_9673(.VSS(VSS),.VDD(VDD),.Y(g25177),.A(I33009));
  NOT NOT1_9674(.VSS(VSS),.VDD(VDD),.Y(I33013),.A(g25119));
  NOT NOT1_9675(.VSS(VSS),.VDD(VDD),.Y(g25179),.A(I33013));
  NOT NOT1_9676(.VSS(VSS),.VDD(VDD),.Y(I33016),.A(g25122));
  NOT NOT1_9677(.VSS(VSS),.VDD(VDD),.Y(g25180),.A(I33016));
  NOT NOT1_9678(.VSS(VSS),.VDD(VDD),.Y(g25274),.A(g24912));
  NOT NOT1_9679(.VSS(VSS),.VDD(VDD),.Y(g25283),.A(g24929));
  NOT NOT1_9680(.VSS(VSS),.VDD(VDD),.Y(g25291),.A(g24941));
  NOT NOT1_9681(.VSS(VSS),.VDD(VDD),.Y(I33128),.A(g24975));
  NOT NOT1_9682(.VSS(VSS),.VDD(VDD),.Y(g25296),.A(I33128));
  NOT NOT1_9683(.VSS(VSS),.VDD(VDD),.Y(g25301),.A(g24952));
  NOT NOT1_9684(.VSS(VSS),.VDD(VDD),.Y(g25305),.A(g24880));
  NOT NOT1_9685(.VSS(VSS),.VDD(VDD),.Y(I33136),.A(g24986));
  NOT NOT1_9686(.VSS(VSS),.VDD(VDD),.Y(g25306),.A(I33136));
  NOT NOT1_9687(.VSS(VSS),.VDD(VDD),.Y(g25313),.A(g24868));
  NOT NOT1_9688(.VSS(VSS),.VDD(VDD),.Y(g25314),.A(g24897));
  NOT NOT1_9689(.VSS(VSS),.VDD(VDD),.Y(I33145),.A(g24997));
  NOT NOT1_9690(.VSS(VSS),.VDD(VDD),.Y(g25315),.A(I33145));
  NOT NOT1_9691(.VSS(VSS),.VDD(VDD),.Y(g25319),.A(g24857));
  NOT NOT1_9692(.VSS(VSS),.VDD(VDD),.Y(g25322),.A(g24883));
  NOT NOT1_9693(.VSS(VSS),.VDD(VDD),.Y(g25323),.A(g24920));
  NOT NOT1_9694(.VSS(VSS),.VDD(VDD),.Y(I33154),.A(g25005));
  NOT NOT1_9695(.VSS(VSS),.VDD(VDD),.Y(g25324),.A(I33154));
  NOT NOT1_9696(.VSS(VSS),.VDD(VDD),.Y(I33157),.A(g25027));
  NOT NOT1_9697(.VSS(VSS),.VDD(VDD),.Y(g25327),.A(I33157));
  NOT NOT1_9698(.VSS(VSS),.VDD(VDD),.Y(g25329),.A(g24844));
  NOT NOT1_9699(.VSS(VSS),.VDD(VDD),.Y(g25330),.A(g24873));
  NOT NOT1_9700(.VSS(VSS),.VDD(VDD),.Y(g25332),.A(g24900));
  NOT NOT1_9701(.VSS(VSS),.VDD(VDD),.Y(g25333),.A(g24937));
  NOT NOT1_9702(.VSS(VSS),.VDD(VDD),.Y(g25335),.A(g24832));
  NOT NOT1_9703(.VSS(VSS),.VDD(VDD),.Y(I33168),.A(g25042));
  NOT NOT1_9704(.VSS(VSS),.VDD(VDD),.Y(g25336),.A(I33168));
  NOT NOT1_9705(.VSS(VSS),.VDD(VDD),.Y(g25338),.A(g24860));
  NOT NOT1_9706(.VSS(VSS),.VDD(VDD),.Y(g25339),.A(g24887));
  NOT NOT1_9707(.VSS(VSS),.VDD(VDD),.Y(g25341),.A(g24923));
  NOT NOT1_9708(.VSS(VSS),.VDD(VDD),.Y(g25347),.A(g24817));
  NOT NOT1_9709(.VSS(VSS),.VDD(VDD),.Y(g25349),.A(g24848));
  NOT NOT1_9710(.VSS(VSS),.VDD(VDD),.Y(I33182),.A(g25056));
  NOT NOT1_9711(.VSS(VSS),.VDD(VDD),.Y(g25350),.A(I33182));
  NOT NOT1_9712(.VSS(VSS),.VDD(VDD),.Y(g25352),.A(g24875));
  NOT NOT1_9713(.VSS(VSS),.VDD(VDD),.Y(g25353),.A(g24904));
  NOT NOT1_9714(.VSS(VSS),.VDD(VDD),.Y(I33188),.A(g24814));
  NOT NOT1_9715(.VSS(VSS),.VDD(VDD),.Y(g25354),.A(I33188));
  NOT NOT1_9716(.VSS(VSS),.VDD(VDD),.Y(g25355),.A(g24797));
  NOT NOT1_9717(.VSS(VSS),.VDD(VDD),.Y(g25361),.A(g24837));
  NOT NOT1_9718(.VSS(VSS),.VDD(VDD),.Y(g25363),.A(g24862));
  NOT NOT1_9719(.VSS(VSS),.VDD(VDD),.Y(I33198),.A(g25067));
  NOT NOT1_9720(.VSS(VSS),.VDD(VDD),.Y(g25364),.A(I33198));
  NOT NOT1_9721(.VSS(VSS),.VDD(VDD),.Y(g25366),.A(g24889));
  NOT NOT1_9722(.VSS(VSS),.VDD(VDD),.Y(g25367),.A(g24676));
  NOT NOT1_9723(.VSS(VSS),.VDD(VDD),.Y(g25368),.A(g24778));
  NOT NOT1_9724(.VSS(VSS),.VDD(VDD),.Y(I33205),.A(g24833));
  NOT NOT1_9725(.VSS(VSS),.VDD(VDD),.Y(g25369),.A(I33205));
  NOT NOT1_9726(.VSS(VSS),.VDD(VDD),.Y(g25370),.A(g24820));
  NOT NOT1_9727(.VSS(VSS),.VDD(VDD),.Y(g25376),.A(g24852));
  NOT NOT1_9728(.VSS(VSS),.VDD(VDD),.Y(g25378),.A(g24877));
  NOT NOT1_9729(.VSS(VSS),.VDD(VDD),.Y(g25379),.A(g24893));
  NOT NOT1_9730(.VSS(VSS),.VDD(VDD),.Y(g25383),.A(g24766));
  NOT NOT1_9731(.VSS(VSS),.VDD(VDD),.Y(g25384),.A(g24695));
  NOT NOT1_9732(.VSS(VSS),.VDD(VDD),.Y(g25385),.A(g24801));
  NOT NOT1_9733(.VSS(VSS),.VDD(VDD),.Y(I33219),.A(g24849));
  NOT NOT1_9734(.VSS(VSS),.VDD(VDD),.Y(g25386),.A(I33219));
  NOT NOT1_9735(.VSS(VSS),.VDD(VDD),.Y(g25387),.A(g24839));
  NOT NOT1_9736(.VSS(VSS),.VDD(VDD),.Y(g25393),.A(g24866));
  NOT NOT1_9737(.VSS(VSS),.VDD(VDD),.Y(g25394),.A(g24753));
  NOT NOT1_9738(.VSS(VSS),.VDD(VDD),.Y(g25395),.A(g24916));
  NOT NOT1_9739(.VSS(VSS),.VDD(VDD),.Y(g25399),.A(g24787));
  NOT NOT1_9740(.VSS(VSS),.VDD(VDD),.Y(g25400),.A(g24712));
  NOT NOT1_9741(.VSS(VSS),.VDD(VDD),.Y(g25401),.A(g24823));
  NOT NOT1_9742(.VSS(VSS),.VDD(VDD),.Y(I33232),.A(g24863));
  NOT NOT1_9743(.VSS(VSS),.VDD(VDD),.Y(g25402),.A(I33232));
  NOT NOT1_9744(.VSS(VSS),.VDD(VDD),.Y(g25403),.A(g24854));
  NOT NOT1_9745(.VSS(VSS),.VDD(VDD),.Y(g25404),.A(g24771));
  NOT NOT1_9746(.VSS(VSS),.VDD(VDD),.Y(g25405),.A(g24933));
  NOT NOT1_9747(.VSS(VSS),.VDD(VDD),.Y(g25409),.A(g24808));
  NOT NOT1_9748(.VSS(VSS),.VDD(VDD),.Y(g25410),.A(g24723));
  NOT NOT1_9749(.VSS(VSS),.VDD(VDD),.Y(g25411),.A(g24842));
  NOT NOT1_9750(.VSS(VSS),.VDD(VDD),.Y(g25412),.A(g24791));
  NOT NOT1_9751(.VSS(VSS),.VDD(VDD),.Y(g25413),.A(g24945));
  NOT NOT1_9752(.VSS(VSS),.VDD(VDD),.Y(g25417),.A(g24830));
  NOT NOT1_9753(.VSS(VSS),.VDD(VDD),.Y(g25419),.A(g24812));
  NOT NOT1_9754(.VSS(VSS),.VDD(VDD),.Y(I33246),.A(g24890));
  NOT NOT1_9755(.VSS(VSS),.VDD(VDD),.Y(g25420),.A(I33246));
  NOT NOT1_9756(.VSS(VSS),.VDD(VDD),.Y(I33249),.A(g24890));
  NOT NOT1_9757(.VSS(VSS),.VDD(VDD),.Y(g25421),.A(I33249));
  NOT NOT1_9758(.VSS(VSS),.VDD(VDD),.Y(g25422),.A(g24958));
  NOT NOT1_9759(.VSS(VSS),.VDD(VDD),.Y(g25430),.A(g24616));
  NOT NOT1_9760(.VSS(VSS),.VDD(VDD),.Y(g25431),.A(g24969));
  NOT NOT1_9761(.VSS(VSS),.VDD(VDD),.Y(I33257),.A(g24909));
  NOT NOT1_9762(.VSS(VSS),.VDD(VDD),.Y(g25435),.A(I33257));
  NOT NOT1_9763(.VSS(VSS),.VDD(VDD),.Y(I33260),.A(g24909));
  NOT NOT1_9764(.VSS(VSS),.VDD(VDD),.Y(g25436),.A(I33260));
  NOT NOT1_9765(.VSS(VSS),.VDD(VDD),.Y(g25437),.A(g24627));
  NOT NOT1_9766(.VSS(VSS),.VDD(VDD),.Y(g25438),.A(g24982));
  NOT NOT1_9767(.VSS(VSS),.VDD(VDD),.Y(I33265),.A(g24925));
  NOT NOT1_9768(.VSS(VSS),.VDD(VDD),.Y(g25442),.A(I33265));
  NOT NOT1_9769(.VSS(VSS),.VDD(VDD),.Y(I33268),.A(g24925));
  NOT NOT1_9770(.VSS(VSS),.VDD(VDD),.Y(g25443),.A(I33268));
  NOT NOT1_9771(.VSS(VSS),.VDD(VDD),.Y(g25444),.A(g24641));
  NOT NOT1_9772(.VSS(VSS),.VDD(VDD),.Y(g25445),.A(g24993));
  NOT NOT1_9773(.VSS(VSS),.VDD(VDD),.Y(g25449),.A(g24660));
  NOT NOT1_9774(.VSS(VSS),.VDD(VDD),.Y(I33278),.A(g25088));
  NOT NOT1_9775(.VSS(VSS),.VDD(VDD),.Y(g25454),.A(I33278));
  NOT NOT1_9776(.VSS(VSS),.VDD(VDD),.Y(I33282),.A(g25096));
  NOT NOT1_9777(.VSS(VSS),.VDD(VDD),.Y(g25458),.A(I33282));
  NOT NOT1_9778(.VSS(VSS),.VDD(VDD),.Y(I33286),.A(g24426));
  NOT NOT1_9779(.VSS(VSS),.VDD(VDD),.Y(g25462),.A(I33286));
  NOT NOT1_9780(.VSS(VSS),.VDD(VDD),.Y(I33289),.A(g25106));
  NOT NOT1_9781(.VSS(VSS),.VDD(VDD),.Y(g25463),.A(I33289));
  NOT NOT1_9782(.VSS(VSS),.VDD(VDD),.Y(I33293),.A(g25008));
  NOT NOT1_9783(.VSS(VSS),.VDD(VDD),.Y(g25467),.A(I33293));
  NOT NOT1_9784(.VSS(VSS),.VDD(VDD),.Y(I33297),.A(g24430));
  NOT NOT1_9785(.VSS(VSS),.VDD(VDD),.Y(g25471),.A(I33297));
  NOT NOT1_9786(.VSS(VSS),.VDD(VDD),.Y(I33300),.A(g25112));
  NOT NOT1_9787(.VSS(VSS),.VDD(VDD),.Y(g25472),.A(I33300));
  NOT NOT1_9788(.VSS(VSS),.VDD(VDD),.Y(I33304),.A(g25004));
  NOT NOT1_9789(.VSS(VSS),.VDD(VDD),.Y(g25476),.A(I33304));
  NOT NOT1_9790(.VSS(VSS),.VDD(VDD),.Y(I33307),.A(g25011));
  NOT NOT1_9791(.VSS(VSS),.VDD(VDD),.Y(g25479),.A(I33307));
  NOT NOT1_9792(.VSS(VSS),.VDD(VDD),.Y(I33312),.A(g25014));
  NOT NOT1_9793(.VSS(VSS),.VDD(VDD),.Y(g25484),.A(I33312));
  NOT NOT1_9794(.VSS(VSS),.VDD(VDD),.Y(I33316),.A(g24434));
  NOT NOT1_9795(.VSS(VSS),.VDD(VDD),.Y(g25488),.A(I33316));
  NOT NOT1_9796(.VSS(VSS),.VDD(VDD),.Y(I33321),.A(g24442));
  NOT NOT1_9797(.VSS(VSS),.VDD(VDD),.Y(g25493),.A(I33321));
  NOT NOT1_9798(.VSS(VSS),.VDD(VDD),.Y(I33324),.A(g25009));
  NOT NOT1_9799(.VSS(VSS),.VDD(VDD),.Y(g25496),.A(I33324));
  NOT NOT1_9800(.VSS(VSS),.VDD(VDD),.Y(I33327),.A(g25017));
  NOT NOT1_9801(.VSS(VSS),.VDD(VDD),.Y(g25499),.A(I33327));
  NOT NOT1_9802(.VSS(VSS),.VDD(VDD),.Y(I33330),.A(g25019));
  NOT NOT1_9803(.VSS(VSS),.VDD(VDD),.Y(g25502),.A(I33330));
  NOT NOT1_9804(.VSS(VSS),.VDD(VDD),.Y(I33335),.A(g25010));
  NOT NOT1_9805(.VSS(VSS),.VDD(VDD),.Y(g25507),.A(I33335));
  NOT NOT1_9806(.VSS(VSS),.VDD(VDD),.Y(I33338),.A(g25021));
  NOT NOT1_9807(.VSS(VSS),.VDD(VDD),.Y(g25510),.A(I33338));
  NOT NOT1_9808(.VSS(VSS),.VDD(VDD),.Y(I33343),.A(g25024));
  NOT NOT1_9809(.VSS(VSS),.VDD(VDD),.Y(g25515),.A(I33343));
  NOT NOT1_9810(.VSS(VSS),.VDD(VDD),.Y(I33347),.A(g24438));
  NOT NOT1_9811(.VSS(VSS),.VDD(VDD),.Y(g25519),.A(I33347));
  NOT NOT1_9812(.VSS(VSS),.VDD(VDD),.Y(I33352),.A(g24443));
  NOT NOT1_9813(.VSS(VSS),.VDD(VDD),.Y(g25524),.A(I33352));
  NOT NOT1_9814(.VSS(VSS),.VDD(VDD),.Y(I33355),.A(g25012));
  NOT NOT1_9815(.VSS(VSS),.VDD(VDD),.Y(g25527),.A(I33355));
  NOT NOT1_9816(.VSS(VSS),.VDD(VDD),.Y(I33358),.A(g25028));
  NOT NOT1_9817(.VSS(VSS),.VDD(VDD),.Y(g25530),.A(I33358));
  NOT NOT1_9818(.VSS(VSS),.VDD(VDD),.Y(I33361),.A(g25013));
  NOT NOT1_9819(.VSS(VSS),.VDD(VDD),.Y(g25533),.A(I33361));
  NOT NOT1_9820(.VSS(VSS),.VDD(VDD),.Y(I33364),.A(g25029));
  NOT NOT1_9821(.VSS(VSS),.VDD(VDD),.Y(g25536),.A(I33364));
  NOT NOT1_9822(.VSS(VSS),.VDD(VDD),.Y(I33368),.A(g24444));
  NOT NOT1_9823(.VSS(VSS),.VDD(VDD),.Y(g25540),.A(I33368));
  NOT NOT1_9824(.VSS(VSS),.VDD(VDD),.Y(I33371),.A(g25015));
  NOT NOT1_9825(.VSS(VSS),.VDD(VDD),.Y(g25543),.A(I33371));
  NOT NOT1_9826(.VSS(VSS),.VDD(VDD),.Y(I33374),.A(g25031));
  NOT NOT1_9827(.VSS(VSS),.VDD(VDD),.Y(g25546),.A(I33374));
  NOT NOT1_9828(.VSS(VSS),.VDD(VDD),.Y(I33377),.A(g25033));
  NOT NOT1_9829(.VSS(VSS),.VDD(VDD),.Y(g25549),.A(I33377));
  NOT NOT1_9830(.VSS(VSS),.VDD(VDD),.Y(I33382),.A(g25016));
  NOT NOT1_9831(.VSS(VSS),.VDD(VDD),.Y(g25554),.A(I33382));
  NOT NOT1_9832(.VSS(VSS),.VDD(VDD),.Y(I33385),.A(g25035));
  NOT NOT1_9833(.VSS(VSS),.VDD(VDD),.Y(g25557),.A(I33385));
  NOT NOT1_9834(.VSS(VSS),.VDD(VDD),.Y(I33390),.A(g25038));
  NOT NOT1_9835(.VSS(VSS),.VDD(VDD),.Y(g25562),.A(I33390));
  NOT NOT1_9836(.VSS(VSS),.VDD(VDD),.Y(I33396),.A(g24447));
  NOT NOT1_9837(.VSS(VSS),.VDD(VDD),.Y(g25573),.A(I33396));
  NOT NOT1_9838(.VSS(VSS),.VDD(VDD),.Y(I33399),.A(g25018));
  NOT NOT1_9839(.VSS(VSS),.VDD(VDD),.Y(g25576),.A(I33399));
  NOT NOT1_9840(.VSS(VSS),.VDD(VDD),.Y(I33402),.A(g24448));
  NOT NOT1_9841(.VSS(VSS),.VDD(VDD),.Y(g25579),.A(I33402));
  NOT NOT1_9842(.VSS(VSS),.VDD(VDD),.Y(I33405),.A(g25020));
  NOT NOT1_9843(.VSS(VSS),.VDD(VDD),.Y(g25582),.A(I33405));
  NOT NOT1_9844(.VSS(VSS),.VDD(VDD),.Y(I33408),.A(g25040));
  NOT NOT1_9845(.VSS(VSS),.VDD(VDD),.Y(g25585),.A(I33408));
  NOT NOT1_9846(.VSS(VSS),.VDD(VDD),.Y(I33411),.A(g24491));
  NOT NOT1_9847(.VSS(VSS),.VDD(VDD),.Y(g25588),.A(I33411));
  NOT NOT1_9848(.VSS(VSS),.VDD(VDD),.Y(I33415),.A(g24449));
  NOT NOT1_9849(.VSS(VSS),.VDD(VDD),.Y(g25590),.A(I33415));
  NOT NOT1_9850(.VSS(VSS),.VDD(VDD),.Y(I33418),.A(g25022));
  NOT NOT1_9851(.VSS(VSS),.VDD(VDD),.Y(g25593),.A(I33418));
  NOT NOT1_9852(.VSS(VSS),.VDD(VDD),.Y(I33421),.A(g25043));
  NOT NOT1_9853(.VSS(VSS),.VDD(VDD),.Y(g25596),.A(I33421));
  NOT NOT1_9854(.VSS(VSS),.VDD(VDD),.Y(I33424),.A(g25023));
  NOT NOT1_9855(.VSS(VSS),.VDD(VDD),.Y(g25599),.A(I33424));
  NOT NOT1_9856(.VSS(VSS),.VDD(VDD),.Y(I33427),.A(g25044));
  NOT NOT1_9857(.VSS(VSS),.VDD(VDD),.Y(g25602),.A(I33427));
  NOT NOT1_9858(.VSS(VSS),.VDD(VDD),.Y(I33431),.A(g24450));
  NOT NOT1_9859(.VSS(VSS),.VDD(VDD),.Y(g25606),.A(I33431));
  NOT NOT1_9860(.VSS(VSS),.VDD(VDD),.Y(I33434),.A(g25025));
  NOT NOT1_9861(.VSS(VSS),.VDD(VDD),.Y(g25609),.A(I33434));
  NOT NOT1_9862(.VSS(VSS),.VDD(VDD),.Y(I33437),.A(g25046));
  NOT NOT1_9863(.VSS(VSS),.VDD(VDD),.Y(g25612),.A(I33437));
  NOT NOT1_9864(.VSS(VSS),.VDD(VDD),.Y(I33440),.A(g25048));
  NOT NOT1_9865(.VSS(VSS),.VDD(VDD),.Y(g25615),.A(I33440));
  NOT NOT1_9866(.VSS(VSS),.VDD(VDD),.Y(I33445),.A(g25026));
  NOT NOT1_9867(.VSS(VSS),.VDD(VDD),.Y(g25620),.A(I33445));
  NOT NOT1_9868(.VSS(VSS),.VDD(VDD),.Y(I33448),.A(g25050));
  NOT NOT1_9869(.VSS(VSS),.VDD(VDD),.Y(g25623),.A(I33448));
  NOT NOT1_9870(.VSS(VSS),.VDD(VDD),.Y(g25630),.A(g24478));
  NOT NOT1_9871(.VSS(VSS),.VDD(VDD),.Y(I33457),.A(g24451));
  NOT NOT1_9872(.VSS(VSS),.VDD(VDD),.Y(g25634),.A(I33457));
  NOT NOT1_9873(.VSS(VSS),.VDD(VDD),.Y(I33460),.A(g24452));
  NOT NOT1_9874(.VSS(VSS),.VDD(VDD),.Y(g25637),.A(I33460));
  NOT NOT1_9875(.VSS(VSS),.VDD(VDD),.Y(I33463),.A(g25030));
  NOT NOT1_9876(.VSS(VSS),.VDD(VDD),.Y(g25640),.A(I33463));
  NOT NOT1_9877(.VSS(VSS),.VDD(VDD),.Y(I33466),.A(g25053));
  NOT NOT1_9878(.VSS(VSS),.VDD(VDD),.Y(g25643),.A(I33466));
  NOT NOT1_9879(.VSS(VSS),.VDD(VDD),.Y(I33469),.A(g24498));
  NOT NOT1_9880(.VSS(VSS),.VDD(VDD),.Y(g25646),.A(I33469));
  NOT NOT1_9881(.VSS(VSS),.VDD(VDD),.Y(I33472),.A(g24499));
  NOT NOT1_9882(.VSS(VSS),.VDD(VDD),.Y(g25647),.A(I33472));
  NOT NOT1_9883(.VSS(VSS),.VDD(VDD),.Y(I33476),.A(g24453));
  NOT NOT1_9884(.VSS(VSS),.VDD(VDD),.Y(g25652),.A(I33476));
  NOT NOT1_9885(.VSS(VSS),.VDD(VDD),.Y(I33479),.A(g25032));
  NOT NOT1_9886(.VSS(VSS),.VDD(VDD),.Y(g25655),.A(I33479));
  NOT NOT1_9887(.VSS(VSS),.VDD(VDD),.Y(I33482),.A(g24454));
  NOT NOT1_9888(.VSS(VSS),.VDD(VDD),.Y(g25658),.A(I33482));
  NOT NOT1_9889(.VSS(VSS),.VDD(VDD),.Y(I33485),.A(g25034));
  NOT NOT1_9890(.VSS(VSS),.VDD(VDD),.Y(g25661),.A(I33485));
  NOT NOT1_9891(.VSS(VSS),.VDD(VDD),.Y(I33488),.A(g25054));
  NOT NOT1_9892(.VSS(VSS),.VDD(VDD),.Y(g25664),.A(I33488));
  NOT NOT1_9893(.VSS(VSS),.VDD(VDD),.Y(I33491),.A(g24501));
  NOT NOT1_9894(.VSS(VSS),.VDD(VDD),.Y(g25667),.A(I33491));
  NOT NOT1_9895(.VSS(VSS),.VDD(VDD),.Y(I33495),.A(g24455));
  NOT NOT1_9896(.VSS(VSS),.VDD(VDD),.Y(g25669),.A(I33495));
  NOT NOT1_9897(.VSS(VSS),.VDD(VDD),.Y(I33498),.A(g25036));
  NOT NOT1_9898(.VSS(VSS),.VDD(VDD),.Y(g25672),.A(I33498));
  NOT NOT1_9899(.VSS(VSS),.VDD(VDD),.Y(I33501),.A(g25057));
  NOT NOT1_9900(.VSS(VSS),.VDD(VDD),.Y(g25675),.A(I33501));
  NOT NOT1_9901(.VSS(VSS),.VDD(VDD),.Y(I33504),.A(g25037));
  NOT NOT1_9902(.VSS(VSS),.VDD(VDD),.Y(g25678),.A(I33504));
  NOT NOT1_9903(.VSS(VSS),.VDD(VDD),.Y(I33507),.A(g25058));
  NOT NOT1_9904(.VSS(VSS),.VDD(VDD),.Y(g25681),.A(I33507));
  NOT NOT1_9905(.VSS(VSS),.VDD(VDD),.Y(I33511),.A(g24456));
  NOT NOT1_9906(.VSS(VSS),.VDD(VDD),.Y(g25685),.A(I33511));
  NOT NOT1_9907(.VSS(VSS),.VDD(VDD),.Y(I33514),.A(g25039));
  NOT NOT1_9908(.VSS(VSS),.VDD(VDD),.Y(g25688),.A(I33514));
  NOT NOT1_9909(.VSS(VSS),.VDD(VDD),.Y(I33517),.A(g25060));
  NOT NOT1_9910(.VSS(VSS),.VDD(VDD),.Y(g25691),.A(I33517));
  NOT NOT1_9911(.VSS(VSS),.VDD(VDD),.Y(I33520),.A(g25062));
  NOT NOT1_9912(.VSS(VSS),.VDD(VDD),.Y(g25694),.A(I33520));
  NOT NOT1_9913(.VSS(VSS),.VDD(VDD),.Y(g25698),.A(g24600));
  NOT NOT1_9914(.VSS(VSS),.VDD(VDD),.Y(I33526),.A(g24457));
  NOT NOT1_9915(.VSS(VSS),.VDD(VDD),.Y(g25700),.A(I33526));
  NOT NOT1_9916(.VSS(VSS),.VDD(VDD),.Y(I33529),.A(g25041));
  NOT NOT1_9917(.VSS(VSS),.VDD(VDD),.Y(g25703),.A(I33529));
  NOT NOT1_9918(.VSS(VSS),.VDD(VDD),.Y(I33532),.A(g24507));
  NOT NOT1_9919(.VSS(VSS),.VDD(VDD),.Y(g25706),.A(I33532));
  NOT NOT1_9920(.VSS(VSS),.VDD(VDD),.Y(I33535),.A(g24508));
  NOT NOT1_9921(.VSS(VSS),.VDD(VDD),.Y(g25707),.A(I33535));
  NOT NOT1_9922(.VSS(VSS),.VDD(VDD),.Y(I33539),.A(g24458));
  NOT NOT1_9923(.VSS(VSS),.VDD(VDD),.Y(g25711),.A(I33539));
  NOT NOT1_9924(.VSS(VSS),.VDD(VDD),.Y(I33542),.A(g24459));
  NOT NOT1_9925(.VSS(VSS),.VDD(VDD),.Y(g25714),.A(I33542));
  NOT NOT1_9926(.VSS(VSS),.VDD(VDD),.Y(I33545),.A(g25045));
  NOT NOT1_9927(.VSS(VSS),.VDD(VDD),.Y(g25717),.A(I33545));
  NOT NOT1_9928(.VSS(VSS),.VDD(VDD),.Y(I33548),.A(g25064));
  NOT NOT1_9929(.VSS(VSS),.VDD(VDD),.Y(g25720),.A(I33548));
  NOT NOT1_9930(.VSS(VSS),.VDD(VDD),.Y(I33551),.A(g24510));
  NOT NOT1_9931(.VSS(VSS),.VDD(VDD),.Y(g25723),.A(I33551));
  NOT NOT1_9932(.VSS(VSS),.VDD(VDD),.Y(I33554),.A(g24511));
  NOT NOT1_9933(.VSS(VSS),.VDD(VDD),.Y(g25724),.A(I33554));
  NOT NOT1_9934(.VSS(VSS),.VDD(VDD),.Y(I33558),.A(g24460));
  NOT NOT1_9935(.VSS(VSS),.VDD(VDD),.Y(g25729),.A(I33558));
  NOT NOT1_9936(.VSS(VSS),.VDD(VDD),.Y(I33561),.A(g25047));
  NOT NOT1_9937(.VSS(VSS),.VDD(VDD),.Y(g25732),.A(I33561));
  NOT NOT1_9938(.VSS(VSS),.VDD(VDD),.Y(I33564),.A(g24461));
  NOT NOT1_9939(.VSS(VSS),.VDD(VDD),.Y(g25735),.A(I33564));
  NOT NOT1_9940(.VSS(VSS),.VDD(VDD),.Y(I33567),.A(g25049));
  NOT NOT1_9941(.VSS(VSS),.VDD(VDD),.Y(g25738),.A(I33567));
  NOT NOT1_9942(.VSS(VSS),.VDD(VDD),.Y(I33570),.A(g25065));
  NOT NOT1_9943(.VSS(VSS),.VDD(VDD),.Y(g25741),.A(I33570));
  NOT NOT1_9944(.VSS(VSS),.VDD(VDD),.Y(I33573),.A(g24513));
  NOT NOT1_9945(.VSS(VSS),.VDD(VDD),.Y(g25744),.A(I33573));
  NOT NOT1_9946(.VSS(VSS),.VDD(VDD),.Y(I33577),.A(g24462));
  NOT NOT1_9947(.VSS(VSS),.VDD(VDD),.Y(g25746),.A(I33577));
  NOT NOT1_9948(.VSS(VSS),.VDD(VDD),.Y(I33580),.A(g25051));
  NOT NOT1_9949(.VSS(VSS),.VDD(VDD),.Y(g25749),.A(I33580));
  NOT NOT1_9950(.VSS(VSS),.VDD(VDD),.Y(I33583),.A(g25068));
  NOT NOT1_9951(.VSS(VSS),.VDD(VDD),.Y(g25752),.A(I33583));
  NOT NOT1_9952(.VSS(VSS),.VDD(VDD),.Y(I33586),.A(g25052));
  NOT NOT1_9953(.VSS(VSS),.VDD(VDD),.Y(g25755),.A(I33586));
  NOT NOT1_9954(.VSS(VSS),.VDD(VDD),.Y(I33589),.A(g25069));
  NOT NOT1_9955(.VSS(VSS),.VDD(VDD),.Y(g25758),.A(I33589));
  NOT NOT1_9956(.VSS(VSS),.VDD(VDD),.Y(I33593),.A(g24445));
  NOT NOT1_9957(.VSS(VSS),.VDD(VDD),.Y(g25762),.A(I33593));
  NOT NOT1_9958(.VSS(VSS),.VDD(VDD),.Y(I33596),.A(g24446));
  NOT NOT1_9959(.VSS(VSS),.VDD(VDD),.Y(g25763),.A(I33596));
  NOT NOT1_9960(.VSS(VSS),.VDD(VDD),.Y(I33600),.A(g24463));
  NOT NOT1_9961(.VSS(VSS),.VDD(VDD),.Y(g25767),.A(I33600));
  NOT NOT1_9962(.VSS(VSS),.VDD(VDD),.Y(I33603),.A(g24519));
  NOT NOT1_9963(.VSS(VSS),.VDD(VDD),.Y(g25770),.A(I33603));
  NOT NOT1_9964(.VSS(VSS),.VDD(VDD),.Y(g25771),.A(g24607));
  NOT NOT1_9965(.VSS(VSS),.VDD(VDD),.Y(I33608),.A(g24464));
  NOT NOT1_9966(.VSS(VSS),.VDD(VDD),.Y(g25773),.A(I33608));
  NOT NOT1_9967(.VSS(VSS),.VDD(VDD),.Y(I33611),.A(g25055));
  NOT NOT1_9968(.VSS(VSS),.VDD(VDD),.Y(g25776),.A(I33611));
  NOT NOT1_9969(.VSS(VSS),.VDD(VDD),.Y(I33614),.A(g24521));
  NOT NOT1_9970(.VSS(VSS),.VDD(VDD),.Y(g25779),.A(I33614));
  NOT NOT1_9971(.VSS(VSS),.VDD(VDD),.Y(I33617),.A(g24522));
  NOT NOT1_9972(.VSS(VSS),.VDD(VDD),.Y(g25780),.A(I33617));
  NOT NOT1_9973(.VSS(VSS),.VDD(VDD),.Y(I33621),.A(g24465));
  NOT NOT1_9974(.VSS(VSS),.VDD(VDD),.Y(g25784),.A(I33621));
  NOT NOT1_9975(.VSS(VSS),.VDD(VDD),.Y(I33624),.A(g24466));
  NOT NOT1_9976(.VSS(VSS),.VDD(VDD),.Y(g25787),.A(I33624));
  NOT NOT1_9977(.VSS(VSS),.VDD(VDD),.Y(I33627),.A(g25059));
  NOT NOT1_9978(.VSS(VSS),.VDD(VDD),.Y(g25790),.A(I33627));
  NOT NOT1_9979(.VSS(VSS),.VDD(VDD),.Y(I33630),.A(g25071));
  NOT NOT1_9980(.VSS(VSS),.VDD(VDD),.Y(g25793),.A(I33630));
  NOT NOT1_9981(.VSS(VSS),.VDD(VDD),.Y(I33633),.A(g24524));
  NOT NOT1_9982(.VSS(VSS),.VDD(VDD),.Y(g25796),.A(I33633));
  NOT NOT1_9983(.VSS(VSS),.VDD(VDD),.Y(I33636),.A(g24525));
  NOT NOT1_9984(.VSS(VSS),.VDD(VDD),.Y(g25797),.A(I33636));
  NOT NOT1_9985(.VSS(VSS),.VDD(VDD),.Y(I33640),.A(g24467));
  NOT NOT1_9986(.VSS(VSS),.VDD(VDD),.Y(g25802),.A(I33640));
  NOT NOT1_9987(.VSS(VSS),.VDD(VDD),.Y(I33643),.A(g25061));
  NOT NOT1_9988(.VSS(VSS),.VDD(VDD),.Y(g25805),.A(I33643));
  NOT NOT1_9989(.VSS(VSS),.VDD(VDD),.Y(I33646),.A(g24468));
  NOT NOT1_9990(.VSS(VSS),.VDD(VDD),.Y(g25808),.A(I33646));
  NOT NOT1_9991(.VSS(VSS),.VDD(VDD),.Y(I33649),.A(g25063));
  NOT NOT1_9992(.VSS(VSS),.VDD(VDD),.Y(g25811),.A(I33649));
  NOT NOT1_9993(.VSS(VSS),.VDD(VDD),.Y(I33652),.A(g25072));
  NOT NOT1_9994(.VSS(VSS),.VDD(VDD),.Y(g25814),.A(I33652));
  NOT NOT1_9995(.VSS(VSS),.VDD(VDD),.Y(I33655),.A(g24527));
  NOT NOT1_9996(.VSS(VSS),.VDD(VDD),.Y(g25817),.A(I33655));
  NOT NOT1_9997(.VSS(VSS),.VDD(VDD),.Y(I33659),.A(g24469));
  NOT NOT1_9998(.VSS(VSS),.VDD(VDD),.Y(g25821),.A(I33659));
  NOT NOT1_9999(.VSS(VSS),.VDD(VDD),.Y(I33662),.A(g24532));
  NOT NOT1_10000(.VSS(VSS),.VDD(VDD),.Y(g25824),.A(I33662));
  NOT NOT1_10001(.VSS(VSS),.VDD(VDD),.Y(g25825),.A(g24619));
  NOT NOT1_10002(.VSS(VSS),.VDD(VDD),.Y(I33667),.A(g24470));
  NOT NOT1_10003(.VSS(VSS),.VDD(VDD),.Y(g25827),.A(I33667));
  NOT NOT1_10004(.VSS(VSS),.VDD(VDD),.Y(I33670),.A(g25066));
  NOT NOT1_10005(.VSS(VSS),.VDD(VDD),.Y(g25830),.A(I33670));
  NOT NOT1_10006(.VSS(VSS),.VDD(VDD),.Y(I33673),.A(g24534));
  NOT NOT1_10007(.VSS(VSS),.VDD(VDD),.Y(g25833),.A(I33673));
  NOT NOT1_10008(.VSS(VSS),.VDD(VDD),.Y(I33676),.A(g24535));
  NOT NOT1_10009(.VSS(VSS),.VDD(VDD),.Y(g25834),.A(I33676));
  NOT NOT1_10010(.VSS(VSS),.VDD(VDD),.Y(I33680),.A(g24471));
  NOT NOT1_10011(.VSS(VSS),.VDD(VDD),.Y(g25838),.A(I33680));
  NOT NOT1_10012(.VSS(VSS),.VDD(VDD),.Y(I33683),.A(g24472));
  NOT NOT1_10013(.VSS(VSS),.VDD(VDD),.Y(g25841),.A(I33683));
  NOT NOT1_10014(.VSS(VSS),.VDD(VDD),.Y(I33686),.A(g25070));
  NOT NOT1_10015(.VSS(VSS),.VDD(VDD),.Y(g25844),.A(I33686));
  NOT NOT1_10016(.VSS(VSS),.VDD(VDD),.Y(I33689),.A(g25074));
  NOT NOT1_10017(.VSS(VSS),.VDD(VDD),.Y(g25847),.A(I33689));
  NOT NOT1_10018(.VSS(VSS),.VDD(VDD),.Y(I33692),.A(g24537));
  NOT NOT1_10019(.VSS(VSS),.VDD(VDD),.Y(g25850),.A(I33692));
  NOT NOT1_10020(.VSS(VSS),.VDD(VDD),.Y(I33695),.A(g24538));
  NOT NOT1_10021(.VSS(VSS),.VDD(VDD),.Y(g25851),.A(I33695));
  NOT NOT1_10022(.VSS(VSS),.VDD(VDD),.Y(I33700),.A(g24474));
  NOT NOT1_10023(.VSS(VSS),.VDD(VDD),.Y(g25856),.A(I33700));
  NOT NOT1_10024(.VSS(VSS),.VDD(VDD),.Y(I33703),.A(g24545));
  NOT NOT1_10025(.VSS(VSS),.VDD(VDD),.Y(g25859),.A(I33703));
  NOT NOT1_10026(.VSS(VSS),.VDD(VDD),.Y(g25860),.A(g24630));
  NOT NOT1_10027(.VSS(VSS),.VDD(VDD),.Y(I33708),.A(g24475));
  NOT NOT1_10028(.VSS(VSS),.VDD(VDD),.Y(g25862),.A(I33708));
  NOT NOT1_10029(.VSS(VSS),.VDD(VDD),.Y(I33711),.A(g25073));
  NOT NOT1_10030(.VSS(VSS),.VDD(VDD),.Y(g25865),.A(I33711));
  NOT NOT1_10031(.VSS(VSS),.VDD(VDD),.Y(I33714),.A(g24547));
  NOT NOT1_10032(.VSS(VSS),.VDD(VDD),.Y(g25868),.A(I33714));
  NOT NOT1_10033(.VSS(VSS),.VDD(VDD),.Y(I33717),.A(g24548));
  NOT NOT1_10034(.VSS(VSS),.VDD(VDD),.Y(g25869),.A(I33717));
  NOT NOT1_10035(.VSS(VSS),.VDD(VDD),.Y(I33723),.A(g24477));
  NOT NOT1_10036(.VSS(VSS),.VDD(VDD),.Y(g25877),.A(I33723));
  NOT NOT1_10037(.VSS(VSS),.VDD(VDD),.Y(I33726),.A(g24557));
  NOT NOT1_10038(.VSS(VSS),.VDD(VDD),.Y(g25880),.A(I33726));
  NOT NOT1_10039(.VSS(VSS),.VDD(VDD),.Y(I33732),.A(g24473));
  NOT NOT1_10040(.VSS(VSS),.VDD(VDD),.Y(g25886),.A(I33732));
  NOT NOT1_10041(.VSS(VSS),.VDD(VDD),.Y(I33737),.A(g24476));
  NOT NOT1_10042(.VSS(VSS),.VDD(VDD),.Y(g25891),.A(I33737));
  NOT NOT1_10043(.VSS(VSS),.VDD(VDD),.Y(g25895),.A(g24939));
  NOT NOT1_10044(.VSS(VSS),.VDD(VDD),.Y(g25899),.A(g24928));
  NOT NOT1_10045(.VSS(VSS),.VDD(VDD),.Y(g25903),.A(g24950));
  NOT NOT1_10046(.VSS(VSS),.VDD(VDD),.Y(g25907),.A(g24940));
  NOT NOT1_10047(.VSS(VSS),.VDD(VDD),.Y(g25911),.A(g24962));
  NOT NOT1_10048(.VSS(VSS),.VDD(VDD),.Y(g25915),.A(g24951));
  NOT NOT1_10049(.VSS(VSS),.VDD(VDD),.Y(g25919),.A(g24973));
  NOT NOT1_10050(.VSS(VSS),.VDD(VDD),.Y(g25923),.A(g24963));
  NOT NOT1_10051(.VSS(VSS),.VDD(VDD),.Y(g25937),.A(g24763));
  NOT NOT1_10052(.VSS(VSS),.VDD(VDD),.Y(g25939),.A(g24784));
  NOT NOT1_10053(.VSS(VSS),.VDD(VDD),.Y(g25942),.A(g24805));
  NOT NOT1_10054(.VSS(VSS),.VDD(VDD),.Y(g25945),.A(g24827));
  NOT NOT1_10055(.VSS(VSS),.VDD(VDD),.Y(g25952),.A(g24735));
  NOT NOT1_10056(.VSS(VSS),.VDD(VDD),.Y(I33790),.A(g25103));
  NOT NOT1_10057(.VSS(VSS),.VDD(VDD),.Y(g25976),.A(I33790));
  NOT NOT1_10058(.VSS(VSS),.VDD(VDD),.Y(I33798),.A(g25109));
  NOT NOT1_10059(.VSS(VSS),.VDD(VDD),.Y(g25982),.A(I33798));
  NOT NOT1_10060(.VSS(VSS),.VDD(VDD),.Y(I33801),.A(g25327));
  NOT NOT1_10061(.VSS(VSS),.VDD(VDD),.Y(g25983),.A(I33801));
  NOT NOT1_10062(.VSS(VSS),.VDD(VDD),.Y(I33804),.A(g25976));
  NOT NOT1_10063(.VSS(VSS),.VDD(VDD),.Y(g25984),.A(I33804));
  NOT NOT1_10064(.VSS(VSS),.VDD(VDD),.Y(I33807),.A(g25588));
  NOT NOT1_10065(.VSS(VSS),.VDD(VDD),.Y(g25985),.A(I33807));
  NOT NOT1_10066(.VSS(VSS),.VDD(VDD),.Y(I33810),.A(g25646));
  NOT NOT1_10067(.VSS(VSS),.VDD(VDD),.Y(g25986),.A(I33810));
  NOT NOT1_10068(.VSS(VSS),.VDD(VDD),.Y(I33813),.A(g25706));
  NOT NOT1_10069(.VSS(VSS),.VDD(VDD),.Y(g25987),.A(I33813));
  NOT NOT1_10070(.VSS(VSS),.VDD(VDD),.Y(I33816),.A(g25647));
  NOT NOT1_10071(.VSS(VSS),.VDD(VDD),.Y(g25988),.A(I33816));
  NOT NOT1_10072(.VSS(VSS),.VDD(VDD),.Y(I33819),.A(g25707));
  NOT NOT1_10073(.VSS(VSS),.VDD(VDD),.Y(g25989),.A(I33819));
  NOT NOT1_10074(.VSS(VSS),.VDD(VDD),.Y(I33822),.A(g25770));
  NOT NOT1_10075(.VSS(VSS),.VDD(VDD),.Y(g25990),.A(I33822));
  NOT NOT1_10076(.VSS(VSS),.VDD(VDD),.Y(I33825),.A(g25462));
  NOT NOT1_10077(.VSS(VSS),.VDD(VDD),.Y(g25991),.A(I33825));
  NOT NOT1_10078(.VSS(VSS),.VDD(VDD),.Y(I33828),.A(g25336));
  NOT NOT1_10079(.VSS(VSS),.VDD(VDD),.Y(g25992),.A(I33828));
  NOT NOT1_10080(.VSS(VSS),.VDD(VDD),.Y(I33831),.A(g25982));
  NOT NOT1_10081(.VSS(VSS),.VDD(VDD),.Y(g25993),.A(I33831));
  NOT NOT1_10082(.VSS(VSS),.VDD(VDD),.Y(I33834),.A(g25667));
  NOT NOT1_10083(.VSS(VSS),.VDD(VDD),.Y(g25994),.A(I33834));
  NOT NOT1_10084(.VSS(VSS),.VDD(VDD),.Y(I33837),.A(g25723));
  NOT NOT1_10085(.VSS(VSS),.VDD(VDD),.Y(g25995),.A(I33837));
  NOT NOT1_10086(.VSS(VSS),.VDD(VDD),.Y(I33840),.A(g25779));
  NOT NOT1_10087(.VSS(VSS),.VDD(VDD),.Y(g25996),.A(I33840));
  NOT NOT1_10088(.VSS(VSS),.VDD(VDD),.Y(I33843),.A(g25724));
  NOT NOT1_10089(.VSS(VSS),.VDD(VDD),.Y(g25997),.A(I33843));
  NOT NOT1_10090(.VSS(VSS),.VDD(VDD),.Y(I33846),.A(g25780));
  NOT NOT1_10091(.VSS(VSS),.VDD(VDD),.Y(g25998),.A(I33846));
  NOT NOT1_10092(.VSS(VSS),.VDD(VDD),.Y(I33849),.A(g25824));
  NOT NOT1_10093(.VSS(VSS),.VDD(VDD),.Y(g25999),.A(I33849));
  NOT NOT1_10094(.VSS(VSS),.VDD(VDD),.Y(I33852),.A(g25471));
  NOT NOT1_10095(.VSS(VSS),.VDD(VDD),.Y(g26000),.A(I33852));
  NOT NOT1_10096(.VSS(VSS),.VDD(VDD),.Y(I33855),.A(g25350));
  NOT NOT1_10097(.VSS(VSS),.VDD(VDD),.Y(g26001),.A(I33855));
  NOT NOT1_10098(.VSS(VSS),.VDD(VDD),.Y(I33858),.A(g25179));
  NOT NOT1_10099(.VSS(VSS),.VDD(VDD),.Y(g26002),.A(I33858));
  NOT NOT1_10100(.VSS(VSS),.VDD(VDD),.Y(I33861),.A(g25744));
  NOT NOT1_10101(.VSS(VSS),.VDD(VDD),.Y(g26003),.A(I33861));
  NOT NOT1_10102(.VSS(VSS),.VDD(VDD),.Y(I33864),.A(g25796));
  NOT NOT1_10103(.VSS(VSS),.VDD(VDD),.Y(g26004),.A(I33864));
  NOT NOT1_10104(.VSS(VSS),.VDD(VDD),.Y(I33867),.A(g25833));
  NOT NOT1_10105(.VSS(VSS),.VDD(VDD),.Y(g26005),.A(I33867));
  NOT NOT1_10106(.VSS(VSS),.VDD(VDD),.Y(I33870),.A(g25797));
  NOT NOT1_10107(.VSS(VSS),.VDD(VDD),.Y(g26006),.A(I33870));
  NOT NOT1_10108(.VSS(VSS),.VDD(VDD),.Y(I33873),.A(g25834));
  NOT NOT1_10109(.VSS(VSS),.VDD(VDD),.Y(g26007),.A(I33873));
  NOT NOT1_10110(.VSS(VSS),.VDD(VDD),.Y(I33876),.A(g25859));
  NOT NOT1_10111(.VSS(VSS),.VDD(VDD),.Y(g26008),.A(I33876));
  NOT NOT1_10112(.VSS(VSS),.VDD(VDD),.Y(I33879),.A(g25488));
  NOT NOT1_10113(.VSS(VSS),.VDD(VDD),.Y(g26009),.A(I33879));
  NOT NOT1_10114(.VSS(VSS),.VDD(VDD),.Y(I33882),.A(g25364));
  NOT NOT1_10115(.VSS(VSS),.VDD(VDD),.Y(g26010),.A(I33882));
  NOT NOT1_10116(.VSS(VSS),.VDD(VDD),.Y(I33885),.A(g25180));
  NOT NOT1_10117(.VSS(VSS),.VDD(VDD),.Y(g26011),.A(I33885));
  NOT NOT1_10118(.VSS(VSS),.VDD(VDD),.Y(I33888),.A(g25817));
  NOT NOT1_10119(.VSS(VSS),.VDD(VDD),.Y(g26012),.A(I33888));
  NOT NOT1_10120(.VSS(VSS),.VDD(VDD),.Y(I33891),.A(g25850));
  NOT NOT1_10121(.VSS(VSS),.VDD(VDD),.Y(g26013),.A(I33891));
  NOT NOT1_10122(.VSS(VSS),.VDD(VDD),.Y(I33894),.A(g25868));
  NOT NOT1_10123(.VSS(VSS),.VDD(VDD),.Y(g26014),.A(I33894));
  NOT NOT1_10124(.VSS(VSS),.VDD(VDD),.Y(I33897),.A(g25851));
  NOT NOT1_10125(.VSS(VSS),.VDD(VDD),.Y(g26015),.A(I33897));
  NOT NOT1_10126(.VSS(VSS),.VDD(VDD),.Y(I33900),.A(g25869));
  NOT NOT1_10127(.VSS(VSS),.VDD(VDD),.Y(g26016),.A(I33900));
  NOT NOT1_10128(.VSS(VSS),.VDD(VDD),.Y(I33903),.A(g25880));
  NOT NOT1_10129(.VSS(VSS),.VDD(VDD),.Y(g26017),.A(I33903));
  NOT NOT1_10130(.VSS(VSS),.VDD(VDD),.Y(I33906),.A(g25519));
  NOT NOT1_10131(.VSS(VSS),.VDD(VDD),.Y(g26018),.A(I33906));
  NOT NOT1_10132(.VSS(VSS),.VDD(VDD),.Y(I33909),.A(g25886));
  NOT NOT1_10133(.VSS(VSS),.VDD(VDD),.Y(g26019),.A(I33909));
  NOT NOT1_10134(.VSS(VSS),.VDD(VDD),.Y(I33912),.A(g25891));
  NOT NOT1_10135(.VSS(VSS),.VDD(VDD),.Y(g26020),.A(I33912));
  NOT NOT1_10136(.VSS(VSS),.VDD(VDD),.Y(I33915),.A(g25762));
  NOT NOT1_10137(.VSS(VSS),.VDD(VDD),.Y(g26021),.A(I33915));
  NOT NOT1_10138(.VSS(VSS),.VDD(VDD),.Y(I33918),.A(g25763));
  NOT NOT1_10139(.VSS(VSS),.VDD(VDD),.Y(g26022),.A(I33918));
  NOT NOT1_10140(.VSS(VSS),.VDD(VDD),.Y(I33954),.A(g25343));
  NOT NOT1_10141(.VSS(VSS),.VDD(VDD),.Y(g26056),.A(I33954));
  NOT NOT1_10142(.VSS(VSS),.VDD(VDD),.Y(I33961),.A(g25357));
  NOT NOT1_10143(.VSS(VSS),.VDD(VDD),.Y(g26063),.A(I33961));
  NOT NOT1_10144(.VSS(VSS),.VDD(VDD),.Y(I33968),.A(g25372));
  NOT NOT1_10145(.VSS(VSS),.VDD(VDD),.Y(g26070),.A(I33968));
  NOT NOT1_10146(.VSS(VSS),.VDD(VDD),.Y(I33974),.A(g25389));
  NOT NOT1_10147(.VSS(VSS),.VDD(VDD),.Y(g26076),.A(I33974));
  NOT NOT1_10148(.VSS(VSS),.VDD(VDD),.Y(I33984),.A(g25932));
  NOT NOT1_10149(.VSS(VSS),.VDD(VDD),.Y(g26086),.A(I33984));
  NOT NOT1_10150(.VSS(VSS),.VDD(VDD),.Y(I33990),.A(g25870));
  NOT NOT1_10151(.VSS(VSS),.VDD(VDD),.Y(g26092),.A(I33990));
  NOT NOT1_10152(.VSS(VSS),.VDD(VDD),.Y(I33995),.A(g25935));
  NOT NOT1_10153(.VSS(VSS),.VDD(VDD),.Y(g26102),.A(I33995));
  NOT NOT1_10154(.VSS(VSS),.VDD(VDD),.Y(I33999),.A(g25490));
  NOT NOT1_10155(.VSS(VSS),.VDD(VDD),.Y(g26104),.A(I33999));
  NOT NOT1_10156(.VSS(VSS),.VDD(VDD),.Y(I34002),.A(g25490));
  NOT NOT1_10157(.VSS(VSS),.VDD(VDD),.Y(g26105),.A(I34002));
  NOT NOT1_10158(.VSS(VSS),.VDD(VDD),.Y(I34009),.A(g25882));
  NOT NOT1_10159(.VSS(VSS),.VDD(VDD),.Y(g26114),.A(I34009));
  NOT NOT1_10160(.VSS(VSS),.VDD(VDD),.Y(I34012),.A(g25938));
  NOT NOT1_10161(.VSS(VSS),.VDD(VDD),.Y(g26118),.A(I34012));
  NOT NOT1_10162(.VSS(VSS),.VDD(VDD),.Y(I34017),.A(g25887));
  NOT NOT1_10163(.VSS(VSS),.VDD(VDD),.Y(g26121),.A(I34017));
  NOT NOT1_10164(.VSS(VSS),.VDD(VDD),.Y(I34020),.A(g25940));
  NOT NOT1_10165(.VSS(VSS),.VDD(VDD),.Y(g26125),.A(I34020));
  NOT NOT1_10166(.VSS(VSS),.VDD(VDD),.Y(I34026),.A(g25892));
  NOT NOT1_10167(.VSS(VSS),.VDD(VDD),.Y(g26131),.A(I34026));
  NOT NOT1_10168(.VSS(VSS),.VDD(VDD),.Y(I34029),.A(g25520));
  NOT NOT1_10169(.VSS(VSS),.VDD(VDD),.Y(g26135),.A(I34029));
  NOT NOT1_10170(.VSS(VSS),.VDD(VDD),.Y(I34032),.A(g25520));
  NOT NOT1_10171(.VSS(VSS),.VDD(VDD),.Y(g26136),.A(I34032));
  NOT NOT1_10172(.VSS(VSS),.VDD(VDD),.Y(I34041),.A(g25566));
  NOT NOT1_10173(.VSS(VSS),.VDD(VDD),.Y(g26149),.A(I34041));
  NOT NOT1_10174(.VSS(VSS),.VDD(VDD),.Y(I34044),.A(g25566));
  NOT NOT1_10175(.VSS(VSS),.VDD(VDD),.Y(g26150),.A(I34044));
  NOT NOT1_10176(.VSS(VSS),.VDD(VDD),.Y(I34051),.A(g25204));
  NOT NOT1_10177(.VSS(VSS),.VDD(VDD),.Y(g26159),.A(I34051));
  NOT NOT1_10178(.VSS(VSS),.VDD(VDD),.Y(I34056),.A(g25206));
  NOT NOT1_10179(.VSS(VSS),.VDD(VDD),.Y(g26164),.A(I34056));
  NOT NOT1_10180(.VSS(VSS),.VDD(VDD),.Y(I34059),.A(g25207));
  NOT NOT1_10181(.VSS(VSS),.VDD(VDD),.Y(g26165),.A(I34059));
  NOT NOT1_10182(.VSS(VSS),.VDD(VDD),.Y(I34063),.A(g25209));
  NOT NOT1_10183(.VSS(VSS),.VDD(VDD),.Y(g26167),.A(I34063));
  NOT NOT1_10184(.VSS(VSS),.VDD(VDD),.Y(I34068),.A(g25211));
  NOT NOT1_10185(.VSS(VSS),.VDD(VDD),.Y(g26172),.A(I34068));
  NOT NOT1_10186(.VSS(VSS),.VDD(VDD),.Y(I34071),.A(g25212));
  NOT NOT1_10187(.VSS(VSS),.VDD(VDD),.Y(g26173),.A(I34071));
  NOT NOT1_10188(.VSS(VSS),.VDD(VDD),.Y(I34074),.A(g25213));
  NOT NOT1_10189(.VSS(VSS),.VDD(VDD),.Y(g26174),.A(I34074));
  NOT NOT1_10190(.VSS(VSS),.VDD(VDD),.Y(I34077),.A(g25954));
  NOT NOT1_10191(.VSS(VSS),.VDD(VDD),.Y(g26175),.A(I34077));
  NOT NOT1_10192(.VSS(VSS),.VDD(VDD),.Y(I34080),.A(g25539));
  NOT NOT1_10193(.VSS(VSS),.VDD(VDD),.Y(g26178),.A(I34080));
  NOT NOT1_10194(.VSS(VSS),.VDD(VDD),.Y(I34083),.A(g25214));
  NOT NOT1_10195(.VSS(VSS),.VDD(VDD),.Y(g26181),.A(I34083));
  NOT NOT1_10196(.VSS(VSS),.VDD(VDD),.Y(I34086),.A(g25215));
  NOT NOT1_10197(.VSS(VSS),.VDD(VDD),.Y(g26182),.A(I34086));
  NOT NOT1_10198(.VSS(VSS),.VDD(VDD),.Y(I34091),.A(g25217));
  NOT NOT1_10199(.VSS(VSS),.VDD(VDD),.Y(g26187),.A(I34091));
  NOT NOT1_10200(.VSS(VSS),.VDD(VDD),.Y(g26189),.A(g25952));
  NOT NOT1_10201(.VSS(VSS),.VDD(VDD),.Y(I34096),.A(g25218));
  NOT NOT1_10202(.VSS(VSS),.VDD(VDD),.Y(g26190),.A(I34096));
  NOT NOT1_10203(.VSS(VSS),.VDD(VDD),.Y(I34099),.A(g25219));
  NOT NOT1_10204(.VSS(VSS),.VDD(VDD),.Y(g26191),.A(I34099));
  NOT NOT1_10205(.VSS(VSS),.VDD(VDD),.Y(I34102),.A(g25220));
  NOT NOT1_10206(.VSS(VSS),.VDD(VDD),.Y(g26192),.A(I34102));
  NOT NOT1_10207(.VSS(VSS),.VDD(VDD),.Y(I34105),.A(g25221));
  NOT NOT1_10208(.VSS(VSS),.VDD(VDD),.Y(g26193),.A(I34105));
  NOT NOT1_10209(.VSS(VSS),.VDD(VDD),.Y(I34108),.A(g25222));
  NOT NOT1_10210(.VSS(VSS),.VDD(VDD),.Y(g26194),.A(I34108));
  NOT NOT1_10211(.VSS(VSS),.VDD(VDD),.Y(I34111),.A(g25223));
  NOT NOT1_10212(.VSS(VSS),.VDD(VDD),.Y(g26195),.A(I34111));
  NOT NOT1_10213(.VSS(VSS),.VDD(VDD),.Y(I34114),.A(g25958));
  NOT NOT1_10214(.VSS(VSS),.VDD(VDD),.Y(g26196),.A(I34114));
  NOT NOT1_10215(.VSS(VSS),.VDD(VDD),.Y(I34118),.A(g25605));
  NOT NOT1_10216(.VSS(VSS),.VDD(VDD),.Y(g26202),.A(I34118));
  NOT NOT1_10217(.VSS(VSS),.VDD(VDD),.Y(I34121),.A(g25224));
  NOT NOT1_10218(.VSS(VSS),.VDD(VDD),.Y(g26205),.A(I34121));
  NOT NOT1_10219(.VSS(VSS),.VDD(VDD),.Y(I34124),.A(g25225));
  NOT NOT1_10220(.VSS(VSS),.VDD(VDD),.Y(g26206),.A(I34124));
  NOT NOT1_10221(.VSS(VSS),.VDD(VDD),.Y(I34128),.A(g25227));
  NOT NOT1_10222(.VSS(VSS),.VDD(VDD),.Y(g26208),.A(I34128));
  NOT NOT1_10223(.VSS(VSS),.VDD(VDD),.Y(g26209),.A(g25296));
  NOT NOT1_10224(.VSS(VSS),.VDD(VDD),.Y(I34132),.A(g25228));
  NOT NOT1_10225(.VSS(VSS),.VDD(VDD),.Y(g26210),.A(I34132));
  NOT NOT1_10226(.VSS(VSS),.VDD(VDD),.Y(I34135),.A(g25229));
  NOT NOT1_10227(.VSS(VSS),.VDD(VDD),.Y(g26211),.A(I34135));
  NOT NOT1_10228(.VSS(VSS),.VDD(VDD),.Y(I34140),.A(g25230));
  NOT NOT1_10229(.VSS(VSS),.VDD(VDD),.Y(g26214),.A(I34140));
  NOT NOT1_10230(.VSS(VSS),.VDD(VDD),.Y(I34143),.A(g25231));
  NOT NOT1_10231(.VSS(VSS),.VDD(VDD),.Y(g26215),.A(I34143));
  NOT NOT1_10232(.VSS(VSS),.VDD(VDD),.Y(I34146),.A(g25232));
  NOT NOT1_10233(.VSS(VSS),.VDD(VDD),.Y(g26216),.A(I34146));
  NOT NOT1_10234(.VSS(VSS),.VDD(VDD),.Y(I34150),.A(g25233));
  NOT NOT1_10235(.VSS(VSS),.VDD(VDD),.Y(g26220),.A(I34150));
  NOT NOT1_10236(.VSS(VSS),.VDD(VDD),.Y(I34153),.A(g25234));
  NOT NOT1_10237(.VSS(VSS),.VDD(VDD),.Y(g26221),.A(I34153));
  NOT NOT1_10238(.VSS(VSS),.VDD(VDD),.Y(I34156),.A(g25235));
  NOT NOT1_10239(.VSS(VSS),.VDD(VDD),.Y(g26222),.A(I34156));
  NOT NOT1_10240(.VSS(VSS),.VDD(VDD),.Y(I34159),.A(g25964));
  NOT NOT1_10241(.VSS(VSS),.VDD(VDD),.Y(g26223),.A(I34159));
  NOT NOT1_10242(.VSS(VSS),.VDD(VDD),.Y(I34162),.A(g25684));
  NOT NOT1_10243(.VSS(VSS),.VDD(VDD),.Y(g26226),.A(I34162));
  NOT NOT1_10244(.VSS(VSS),.VDD(VDD),.Y(I34165),.A(g25236));
  NOT NOT1_10245(.VSS(VSS),.VDD(VDD),.Y(g26229),.A(I34165));
  NOT NOT1_10246(.VSS(VSS),.VDD(VDD),.Y(I34168),.A(g25237));
  NOT NOT1_10247(.VSS(VSS),.VDD(VDD),.Y(g26230),.A(I34168));
  NOT NOT1_10248(.VSS(VSS),.VDD(VDD),.Y(I34172),.A(g25239));
  NOT NOT1_10249(.VSS(VSS),.VDD(VDD),.Y(g26232),.A(I34172));
  NOT NOT1_10250(.VSS(VSS),.VDD(VDD),.Y(g26237),.A(g25306));
  NOT NOT1_10251(.VSS(VSS),.VDD(VDD),.Y(I34180),.A(g25240));
  NOT NOT1_10252(.VSS(VSS),.VDD(VDD),.Y(g26238),.A(I34180));
  NOT NOT1_10253(.VSS(VSS),.VDD(VDD),.Y(I34183),.A(g25241));
  NOT NOT1_10254(.VSS(VSS),.VDD(VDD),.Y(g26239),.A(I34183));
  NOT NOT1_10255(.VSS(VSS),.VDD(VDD),.Y(I34189),.A(g25242));
  NOT NOT1_10256(.VSS(VSS),.VDD(VDD),.Y(g26245),.A(I34189));
  NOT NOT1_10257(.VSS(VSS),.VDD(VDD),.Y(I34192),.A(g25243));
  NOT NOT1_10258(.VSS(VSS),.VDD(VDD),.Y(g26246),.A(I34192));
  NOT NOT1_10259(.VSS(VSS),.VDD(VDD),.Y(I34195),.A(g25244));
  NOT NOT1_10260(.VSS(VSS),.VDD(VDD),.Y(g26247),.A(I34195));
  NOT NOT1_10261(.VSS(VSS),.VDD(VDD),.Y(I34198),.A(g25245));
  NOT NOT1_10262(.VSS(VSS),.VDD(VDD),.Y(g26248),.A(I34198));
  NOT NOT1_10263(.VSS(VSS),.VDD(VDD),.Y(I34201),.A(g25246));
  NOT NOT1_10264(.VSS(VSS),.VDD(VDD),.Y(g26249),.A(I34201));
  NOT NOT1_10265(.VSS(VSS),.VDD(VDD),.Y(I34204),.A(g25247));
  NOT NOT1_10266(.VSS(VSS),.VDD(VDD),.Y(g26250),.A(I34204));
  NOT NOT1_10267(.VSS(VSS),.VDD(VDD),.Y(I34207),.A(g25969));
  NOT NOT1_10268(.VSS(VSS),.VDD(VDD),.Y(g26251),.A(I34207));
  NOT NOT1_10269(.VSS(VSS),.VDD(VDD),.Y(I34210),.A(g25761));
  NOT NOT1_10270(.VSS(VSS),.VDD(VDD),.Y(g26254),.A(I34210));
  NOT NOT1_10271(.VSS(VSS),.VDD(VDD),.Y(I34220),.A(g25248));
  NOT NOT1_10272(.VSS(VSS),.VDD(VDD),.Y(g26264),.A(I34220));
  NOT NOT1_10273(.VSS(VSS),.VDD(VDD),.Y(g26275),.A(g25315));
  NOT NOT1_10274(.VSS(VSS),.VDD(VDD),.Y(I34230),.A(g25249));
  NOT NOT1_10275(.VSS(VSS),.VDD(VDD),.Y(g26276),.A(I34230));
  NOT NOT1_10276(.VSS(VSS),.VDD(VDD),.Y(I34233),.A(g25250));
  NOT NOT1_10277(.VSS(VSS),.VDD(VDD),.Y(g26277),.A(I34233));
  NOT NOT1_10278(.VSS(VSS),.VDD(VDD),.Y(I34238),.A(g25251));
  NOT NOT1_10279(.VSS(VSS),.VDD(VDD),.Y(g26280),.A(I34238));
  NOT NOT1_10280(.VSS(VSS),.VDD(VDD),.Y(I34241),.A(g25252));
  NOT NOT1_10281(.VSS(VSS),.VDD(VDD),.Y(g26281),.A(I34241));
  NOT NOT1_10282(.VSS(VSS),.VDD(VDD),.Y(I34244),.A(g25253));
  NOT NOT1_10283(.VSS(VSS),.VDD(VDD),.Y(g26282),.A(I34244));
  NOT NOT1_10284(.VSS(VSS),.VDD(VDD),.Y(I34254),.A(g25185));
  NOT NOT1_10285(.VSS(VSS),.VDD(VDD),.Y(g26294),.A(I34254));
  NOT NOT1_10286(.VSS(VSS),.VDD(VDD),.Y(I34266),.A(g25255));
  NOT NOT1_10287(.VSS(VSS),.VDD(VDD),.Y(g26308),.A(I34266));
  NOT NOT1_10288(.VSS(VSS),.VDD(VDD),.Y(g26313),.A(g25324));
  NOT NOT1_10289(.VSS(VSS),.VDD(VDD),.Y(I34274),.A(g25256));
  NOT NOT1_10290(.VSS(VSS),.VDD(VDD),.Y(g26314),.A(I34274));
  NOT NOT1_10291(.VSS(VSS),.VDD(VDD),.Y(I34277),.A(g25257));
  NOT NOT1_10292(.VSS(VSS),.VDD(VDD),.Y(g26315),.A(I34277));
  NOT NOT1_10293(.VSS(VSS),.VDD(VDD),.Y(I34296),.A(g25189));
  NOT NOT1_10294(.VSS(VSS),.VDD(VDD),.Y(g26341),.A(I34296));
  NOT NOT1_10295(.VSS(VSS),.VDD(VDD),.Y(I34306),.A(g25259));
  NOT NOT1_10296(.VSS(VSS),.VDD(VDD),.Y(g26349),.A(I34306));
  NOT NOT1_10297(.VSS(VSS),.VDD(VDD),.Y(I34313),.A(g25265));
  NOT NOT1_10298(.VSS(VSS),.VDD(VDD),.Y(g26354),.A(I34313));
  NOT NOT1_10299(.VSS(VSS),.VDD(VDD),.Y(I34316),.A(g25191));
  NOT NOT1_10300(.VSS(VSS),.VDD(VDD),.Y(g26355),.A(I34316));
  NOT NOT1_10301(.VSS(VSS),.VDD(VDD),.Y(I34321),.A(g25928));
  NOT NOT1_10302(.VSS(VSS),.VDD(VDD),.Y(g26358),.A(I34321));
  NOT NOT1_10303(.VSS(VSS),.VDD(VDD),.Y(I34327),.A(g25260));
  NOT NOT1_10304(.VSS(VSS),.VDD(VDD),.Y(g26364),.A(I34327));
  NOT NOT1_10305(.VSS(VSS),.VDD(VDD),.Y(I34343),.A(g25194));
  NOT NOT1_10306(.VSS(VSS),.VDD(VDD),.Y(g26385),.A(I34343));
  NOT NOT1_10307(.VSS(VSS),.VDD(VDD),.Y(I34353),.A(g25927));
  NOT NOT1_10308(.VSS(VSS),.VDD(VDD),.Y(g26393),.A(I34353));
  NOT NOT1_10309(.VSS(VSS),.VDD(VDD),.Y(I34358),.A(g25262));
  NOT NOT1_10310(.VSS(VSS),.VDD(VDD),.Y(g26398),.A(I34358));
  NOT NOT1_10311(.VSS(VSS),.VDD(VDD),.Y(I34363),.A(g25930));
  NOT NOT1_10312(.VSS(VSS),.VDD(VDD),.Y(g26401),.A(I34363));
  NOT NOT1_10313(.VSS(VSS),.VDD(VDD),.Y(I34369),.A(g25263));
  NOT NOT1_10314(.VSS(VSS),.VDD(VDD),.Y(g26407),.A(I34369));
  NOT NOT1_10315(.VSS(VSS),.VDD(VDD),.Y(I34385),.A(g25197));
  NOT NOT1_10316(.VSS(VSS),.VDD(VDD),.Y(g26428),.A(I34385));
  NOT NOT1_10317(.VSS(VSS),.VDD(VDD),.Y(I34388),.A(g25200));
  NOT NOT1_10318(.VSS(VSS),.VDD(VDD),.Y(g26429),.A(I34388));
  NOT NOT1_10319(.VSS(VSS),.VDD(VDD),.Y(I34392),.A(g25266));
  NOT NOT1_10320(.VSS(VSS),.VDD(VDD),.Y(g26433),.A(I34392));
  NOT NOT1_10321(.VSS(VSS),.VDD(VDD),.Y(I34395),.A(g25929));
  NOT NOT1_10322(.VSS(VSS),.VDD(VDD),.Y(g26434),.A(I34395));
  NOT NOT1_10323(.VSS(VSS),.VDD(VDD),.Y(I34400),.A(g25267));
  NOT NOT1_10324(.VSS(VSS),.VDD(VDD),.Y(g26439),.A(I34400));
  NOT NOT1_10325(.VSS(VSS),.VDD(VDD),.Y(I34405),.A(g25933));
  NOT NOT1_10326(.VSS(VSS),.VDD(VDD),.Y(g26442),.A(I34405));
  NOT NOT1_10327(.VSS(VSS),.VDD(VDD),.Y(I34411),.A(g25268));
  NOT NOT1_10328(.VSS(VSS),.VDD(VDD),.Y(g26448),.A(I34411));
  NOT NOT1_10329(.VSS(VSS),.VDD(VDD),.Y(I34421),.A(g25203));
  NOT NOT1_10330(.VSS(VSS),.VDD(VDD),.Y(g26461),.A(I34421));
  NOT NOT1_10331(.VSS(VSS),.VDD(VDD),.Y(I34425),.A(g25270));
  NOT NOT1_10332(.VSS(VSS),.VDD(VDD),.Y(g26465),.A(I34425));
  NOT NOT1_10333(.VSS(VSS),.VDD(VDD),.Y(I34428),.A(g25931));
  NOT NOT1_10334(.VSS(VSS),.VDD(VDD),.Y(g26466),.A(I34428));
  NOT NOT1_10335(.VSS(VSS),.VDD(VDD),.Y(I34433),.A(g25271));
  NOT NOT1_10336(.VSS(VSS),.VDD(VDD),.Y(g26471),.A(I34433));
  NOT NOT1_10337(.VSS(VSS),.VDD(VDD),.Y(I34438),.A(g25936));
  NOT NOT1_10338(.VSS(VSS),.VDD(VDD),.Y(g26474),.A(I34438));
  NOT NOT1_10339(.VSS(VSS),.VDD(VDD),.Y(I34444),.A(g25272));
  NOT NOT1_10340(.VSS(VSS),.VDD(VDD),.Y(g26480),.A(I34444));
  NOT NOT1_10341(.VSS(VSS),.VDD(VDD),.Y(g26481),.A(g25764));
  NOT NOT1_10342(.VSS(VSS),.VDD(VDD),.Y(I34449),.A(g25205));
  NOT NOT1_10343(.VSS(VSS),.VDD(VDD),.Y(g26485),.A(I34449));
  NOT NOT1_10344(.VSS(VSS),.VDD(VDD),.Y(I34453),.A(g25279));
  NOT NOT1_10345(.VSS(VSS),.VDD(VDD),.Y(g26489),.A(I34453));
  NOT NOT1_10346(.VSS(VSS),.VDD(VDD),.Y(I34456),.A(g25934));
  NOT NOT1_10347(.VSS(VSS),.VDD(VDD),.Y(g26490),.A(I34456));
  NOT NOT1_10348(.VSS(VSS),.VDD(VDD),.Y(I34461),.A(g25280));
  NOT NOT1_10349(.VSS(VSS),.VDD(VDD),.Y(g26495),.A(I34461));
  NOT NOT1_10350(.VSS(VSS),.VDD(VDD),.Y(I34464),.A(g25199));
  NOT NOT1_10351(.VSS(VSS),.VDD(VDD),.Y(g26496),.A(I34464));
  NOT NOT1_10352(.VSS(VSS),.VDD(VDD),.Y(g26497),.A(g25818));
  NOT NOT1_10353(.VSS(VSS),.VDD(VDD),.Y(I34469),.A(g25210));
  NOT NOT1_10354(.VSS(VSS),.VDD(VDD),.Y(g26501),.A(I34469));
  NOT NOT1_10355(.VSS(VSS),.VDD(VDD),.Y(I34473),.A(g25288));
  NOT NOT1_10356(.VSS(VSS),.VDD(VDD),.Y(g26505),.A(I34473));
  NOT NOT1_10357(.VSS(VSS),.VDD(VDD),.Y(I34476),.A(g25201));
  NOT NOT1_10358(.VSS(VSS),.VDD(VDD),.Y(g26506),.A(I34476));
  NOT NOT1_10359(.VSS(VSS),.VDD(VDD),.Y(I34479),.A(g25202));
  NOT NOT1_10360(.VSS(VSS),.VDD(VDD),.Y(g26507),.A(I34479));
  NOT NOT1_10361(.VSS(VSS),.VDD(VDD),.Y(g26508),.A(g25312));
  NOT NOT1_10362(.VSS(VSS),.VDD(VDD),.Y(g26512),.A(g25853));
  NOT NOT1_10363(.VSS(VSS),.VDD(VDD),.Y(g26516),.A(g25320));
  NOT NOT1_10364(.VSS(VSS),.VDD(VDD),.Y(g26520),.A(g25874));
  NOT NOT1_10365(.VSS(VSS),.VDD(VDD),.Y(g26521),.A(g25331));
  NOT NOT1_10366(.VSS(VSS),.VDD(VDD),.Y(g26525),.A(g25340));
  NOT NOT1_10367(.VSS(VSS),.VDD(VDD),.Y(g26533),.A(g25454));
  NOT NOT1_10368(.VSS(VSS),.VDD(VDD),.Y(g26538),.A(g25458));
  NOT NOT1_10369(.VSS(VSS),.VDD(VDD),.Y(g26539),.A(g25463));
  NOT NOT1_10370(.VSS(VSS),.VDD(VDD),.Y(g26540),.A(g25467));
  NOT NOT1_10371(.VSS(VSS),.VDD(VDD),.Y(g26542),.A(g25472));
  NOT NOT1_10372(.VSS(VSS),.VDD(VDD),.Y(g26543),.A(g25476));
  NOT NOT1_10373(.VSS(VSS),.VDD(VDD),.Y(g26544),.A(g25479));
  NOT NOT1_10374(.VSS(VSS),.VDD(VDD),.Y(g26546),.A(g25484));
  NOT NOT1_10375(.VSS(VSS),.VDD(VDD),.Y(I34505),.A(g25450));
  NOT NOT1_10376(.VSS(VSS),.VDD(VDD),.Y(g26548),.A(I34505));
  NOT NOT1_10377(.VSS(VSS),.VDD(VDD),.Y(g26549),.A(g25421));
  NOT NOT1_10378(.VSS(VSS),.VDD(VDD),.Y(g26550),.A(g25493));
  NOT NOT1_10379(.VSS(VSS),.VDD(VDD),.Y(g26551),.A(g25496));
  NOT NOT1_10380(.VSS(VSS),.VDD(VDD),.Y(g26552),.A(g25499));
  NOT NOT1_10381(.VSS(VSS),.VDD(VDD),.Y(g26554),.A(g25502));
  NOT NOT1_10382(.VSS(VSS),.VDD(VDD),.Y(g26555),.A(g25507));
  NOT NOT1_10383(.VSS(VSS),.VDD(VDD),.Y(g26556),.A(g25510));
  NOT NOT1_10384(.VSS(VSS),.VDD(VDD),.Y(g26558),.A(g25515));
  NOT NOT1_10385(.VSS(VSS),.VDD(VDD),.Y(g26561),.A(g25524));
  NOT NOT1_10386(.VSS(VSS),.VDD(VDD),.Y(g26562),.A(g25527));
  NOT NOT1_10387(.VSS(VSS),.VDD(VDD),.Y(g26563),.A(g25530));
  NOT NOT1_10388(.VSS(VSS),.VDD(VDD),.Y(g26564),.A(g25533));
  NOT NOT1_10389(.VSS(VSS),.VDD(VDD),.Y(g26565),.A(g25536));
  NOT NOT1_10390(.VSS(VSS),.VDD(VDD),.Y(g26566),.A(g25540));
  NOT NOT1_10391(.VSS(VSS),.VDD(VDD),.Y(g26567),.A(g25543));
  NOT NOT1_10392(.VSS(VSS),.VDD(VDD),.Y(g26568),.A(g25546));
  NOT NOT1_10393(.VSS(VSS),.VDD(VDD),.Y(g26570),.A(g25549));
  NOT NOT1_10394(.VSS(VSS),.VDD(VDD),.Y(g26571),.A(g25554));
  NOT NOT1_10395(.VSS(VSS),.VDD(VDD),.Y(g26572),.A(g25557));
  NOT NOT1_10396(.VSS(VSS),.VDD(VDD),.Y(g26574),.A(g25562));
  NOT NOT1_10397(.VSS(VSS),.VDD(VDD),.Y(I34535),.A(g25451));
  NOT NOT1_10398(.VSS(VSS),.VDD(VDD),.Y(g26576),.A(I34535));
  NOT NOT1_10399(.VSS(VSS),.VDD(VDD),.Y(g26577),.A(g25436));
  NOT NOT1_10400(.VSS(VSS),.VDD(VDD),.Y(g26578),.A(g25573));
  NOT NOT1_10401(.VSS(VSS),.VDD(VDD),.Y(g26579),.A(g25576));
  NOT NOT1_10402(.VSS(VSS),.VDD(VDD),.Y(g26580),.A(g25579));
  NOT NOT1_10403(.VSS(VSS),.VDD(VDD),.Y(g26581),.A(g25582));
  NOT NOT1_10404(.VSS(VSS),.VDD(VDD),.Y(g26582),.A(g25585));
  NOT NOT1_10405(.VSS(VSS),.VDD(VDD),.Y(g26584),.A(g25590));
  NOT NOT1_10406(.VSS(VSS),.VDD(VDD),.Y(g26585),.A(g25593));
  NOT NOT1_10407(.VSS(VSS),.VDD(VDD),.Y(g26586),.A(g25596));
  NOT NOT1_10408(.VSS(VSS),.VDD(VDD),.Y(g26587),.A(g25599));
  NOT NOT1_10409(.VSS(VSS),.VDD(VDD),.Y(g26588),.A(g25602));
  NOT NOT1_10410(.VSS(VSS),.VDD(VDD),.Y(g26589),.A(g25606));
  NOT NOT1_10411(.VSS(VSS),.VDD(VDD),.Y(g26590),.A(g25609));
  NOT NOT1_10412(.VSS(VSS),.VDD(VDD),.Y(g26591),.A(g25612));
  NOT NOT1_10413(.VSS(VSS),.VDD(VDD),.Y(g26593),.A(g25615));
  NOT NOT1_10414(.VSS(VSS),.VDD(VDD),.Y(g26594),.A(g25620));
  NOT NOT1_10415(.VSS(VSS),.VDD(VDD),.Y(g26595),.A(g25623));
  NOT NOT1_10416(.VSS(VSS),.VDD(VDD),.Y(g26597),.A(g25443));
  NOT NOT1_10417(.VSS(VSS),.VDD(VDD),.Y(g26598),.A(g25634));
  NOT NOT1_10418(.VSS(VSS),.VDD(VDD),.Y(g26599),.A(g25637));
  NOT NOT1_10419(.VSS(VSS),.VDD(VDD),.Y(g26600),.A(g25640));
  NOT NOT1_10420(.VSS(VSS),.VDD(VDD),.Y(g26601),.A(g25643));
  NOT NOT1_10421(.VSS(VSS),.VDD(VDD),.Y(g26602),.A(g25652));
  NOT NOT1_10422(.VSS(VSS),.VDD(VDD),.Y(g26603),.A(g25655));
  NOT NOT1_10423(.VSS(VSS),.VDD(VDD),.Y(g26604),.A(g25658));
  NOT NOT1_10424(.VSS(VSS),.VDD(VDD),.Y(g26605),.A(g25661));
  NOT NOT1_10425(.VSS(VSS),.VDD(VDD),.Y(g26606),.A(g25664));
  NOT NOT1_10426(.VSS(VSS),.VDD(VDD),.Y(g26608),.A(g25669));
  NOT NOT1_10427(.VSS(VSS),.VDD(VDD),.Y(g26609),.A(g25672));
  NOT NOT1_10428(.VSS(VSS),.VDD(VDD),.Y(g26610),.A(g25675));
  NOT NOT1_10429(.VSS(VSS),.VDD(VDD),.Y(g26611),.A(g25678));
  NOT NOT1_10430(.VSS(VSS),.VDD(VDD),.Y(g26612),.A(g25681));
  NOT NOT1_10431(.VSS(VSS),.VDD(VDD),.Y(g26613),.A(g25685));
  NOT NOT1_10432(.VSS(VSS),.VDD(VDD),.Y(g26614),.A(g25688));
  NOT NOT1_10433(.VSS(VSS),.VDD(VDD),.Y(g26615),.A(g25691));
  NOT NOT1_10434(.VSS(VSS),.VDD(VDD),.Y(g26617),.A(g25694));
  NOT NOT1_10435(.VSS(VSS),.VDD(VDD),.Y(I34579),.A(g25452));
  NOT NOT1_10436(.VSS(VSS),.VDD(VDD),.Y(g26618),.A(I34579));
  NOT NOT1_10437(.VSS(VSS),.VDD(VDD),.Y(g26619),.A(g25700));
  NOT NOT1_10438(.VSS(VSS),.VDD(VDD),.Y(g26620),.A(g25703));
  NOT NOT1_10439(.VSS(VSS),.VDD(VDD),.Y(g26621),.A(g25711));
  NOT NOT1_10440(.VSS(VSS),.VDD(VDD),.Y(g26622),.A(g25714));
  NOT NOT1_10441(.VSS(VSS),.VDD(VDD),.Y(g26623),.A(g25717));
  NOT NOT1_10442(.VSS(VSS),.VDD(VDD),.Y(g26624),.A(g25720));
  NOT NOT1_10443(.VSS(VSS),.VDD(VDD),.Y(g26625),.A(g25729));
  NOT NOT1_10444(.VSS(VSS),.VDD(VDD),.Y(g26626),.A(g25732));
  NOT NOT1_10445(.VSS(VSS),.VDD(VDD),.Y(g26627),.A(g25735));
  NOT NOT1_10446(.VSS(VSS),.VDD(VDD),.Y(g26628),.A(g25738));
  NOT NOT1_10447(.VSS(VSS),.VDD(VDD),.Y(g26629),.A(g25741));
  NOT NOT1_10448(.VSS(VSS),.VDD(VDD),.Y(g26631),.A(g25746));
  NOT NOT1_10449(.VSS(VSS),.VDD(VDD),.Y(g26632),.A(g25749));
  NOT NOT1_10450(.VSS(VSS),.VDD(VDD),.Y(g26633),.A(g25752));
  NOT NOT1_10451(.VSS(VSS),.VDD(VDD),.Y(g26634),.A(g25755));
  NOT NOT1_10452(.VSS(VSS),.VDD(VDD),.Y(g26635),.A(g25758));
  NOT NOT1_10453(.VSS(VSS),.VDD(VDD),.Y(g26636),.A(g25767));
  NOT NOT1_10454(.VSS(VSS),.VDD(VDD),.Y(g26637),.A(g25773));
  NOT NOT1_10455(.VSS(VSS),.VDD(VDD),.Y(g26638),.A(g25776));
  NOT NOT1_10456(.VSS(VSS),.VDD(VDD),.Y(g26639),.A(g25784));
  NOT NOT1_10457(.VSS(VSS),.VDD(VDD),.Y(g26640),.A(g25787));
  NOT NOT1_10458(.VSS(VSS),.VDD(VDD),.Y(g26641),.A(g25790));
  NOT NOT1_10459(.VSS(VSS),.VDD(VDD),.Y(g26642),.A(g25793));
  NOT NOT1_10460(.VSS(VSS),.VDD(VDD),.Y(g26643),.A(g25802));
  NOT NOT1_10461(.VSS(VSS),.VDD(VDD),.Y(g26644),.A(g25805));
  NOT NOT1_10462(.VSS(VSS),.VDD(VDD),.Y(g26645),.A(g25808));
  NOT NOT1_10463(.VSS(VSS),.VDD(VDD),.Y(g26646),.A(g25811));
  NOT NOT1_10464(.VSS(VSS),.VDD(VDD),.Y(g26647),.A(g25814));
  NOT NOT1_10465(.VSS(VSS),.VDD(VDD),.Y(g26648),.A(g25821));
  NOT NOT1_10466(.VSS(VSS),.VDD(VDD),.Y(g26649),.A(g25827));
  NOT NOT1_10467(.VSS(VSS),.VDD(VDD),.Y(g26650),.A(g25830));
  NOT NOT1_10468(.VSS(VSS),.VDD(VDD),.Y(g26651),.A(g25838));
  NOT NOT1_10469(.VSS(VSS),.VDD(VDD),.Y(g26652),.A(g25841));
  NOT NOT1_10470(.VSS(VSS),.VDD(VDD),.Y(g26653),.A(g25844));
  NOT NOT1_10471(.VSS(VSS),.VDD(VDD),.Y(g26654),.A(g25847));
  NOT NOT1_10472(.VSS(VSS),.VDD(VDD),.Y(g26656),.A(g25856));
  NOT NOT1_10473(.VSS(VSS),.VDD(VDD),.Y(g26657),.A(g25862));
  NOT NOT1_10474(.VSS(VSS),.VDD(VDD),.Y(g26658),.A(g25865));
  NOT NOT1_10475(.VSS(VSS),.VDD(VDD),.Y(g26662),.A(g25877));
  NOT NOT1_10476(.VSS(VSS),.VDD(VDD),.Y(I34641),.A(g26086));
  NOT NOT1_10477(.VSS(VSS),.VDD(VDD),.Y(g26678),.A(I34641));
  NOT NOT1_10478(.VSS(VSS),.VDD(VDD),.Y(I34644),.A(g26159));
  NOT NOT1_10479(.VSS(VSS),.VDD(VDD),.Y(g26679),.A(I34644));
  NOT NOT1_10480(.VSS(VSS),.VDD(VDD),.Y(I34647),.A(g26164));
  NOT NOT1_10481(.VSS(VSS),.VDD(VDD),.Y(g26680),.A(I34647));
  NOT NOT1_10482(.VSS(VSS),.VDD(VDD),.Y(I34650),.A(g26172));
  NOT NOT1_10483(.VSS(VSS),.VDD(VDD),.Y(g26681),.A(I34650));
  NOT NOT1_10484(.VSS(VSS),.VDD(VDD),.Y(I34653),.A(g26165));
  NOT NOT1_10485(.VSS(VSS),.VDD(VDD),.Y(g26682),.A(I34653));
  NOT NOT1_10486(.VSS(VSS),.VDD(VDD),.Y(I34656),.A(g26173));
  NOT NOT1_10487(.VSS(VSS),.VDD(VDD),.Y(g26683),.A(I34656));
  NOT NOT1_10488(.VSS(VSS),.VDD(VDD),.Y(I34659),.A(g26190));
  NOT NOT1_10489(.VSS(VSS),.VDD(VDD),.Y(g26684),.A(I34659));
  NOT NOT1_10490(.VSS(VSS),.VDD(VDD),.Y(I34662),.A(g26174));
  NOT NOT1_10491(.VSS(VSS),.VDD(VDD),.Y(g26685),.A(I34662));
  NOT NOT1_10492(.VSS(VSS),.VDD(VDD),.Y(I34665),.A(g26191));
  NOT NOT1_10493(.VSS(VSS),.VDD(VDD),.Y(g26686),.A(I34665));
  NOT NOT1_10494(.VSS(VSS),.VDD(VDD),.Y(I34668),.A(g26210));
  NOT NOT1_10495(.VSS(VSS),.VDD(VDD),.Y(g26687),.A(I34668));
  NOT NOT1_10496(.VSS(VSS),.VDD(VDD),.Y(I34671),.A(g26192));
  NOT NOT1_10497(.VSS(VSS),.VDD(VDD),.Y(g26688),.A(I34671));
  NOT NOT1_10498(.VSS(VSS),.VDD(VDD),.Y(I34674),.A(g26211));
  NOT NOT1_10499(.VSS(VSS),.VDD(VDD),.Y(g26689),.A(I34674));
  NOT NOT1_10500(.VSS(VSS),.VDD(VDD),.Y(I34677),.A(g26232));
  NOT NOT1_10501(.VSS(VSS),.VDD(VDD),.Y(g26690),.A(I34677));
  NOT NOT1_10502(.VSS(VSS),.VDD(VDD),.Y(I34680),.A(g26294));
  NOT NOT1_10503(.VSS(VSS),.VDD(VDD),.Y(g26691),.A(I34680));
  NOT NOT1_10504(.VSS(VSS),.VDD(VDD),.Y(I34683),.A(g26364));
  NOT NOT1_10505(.VSS(VSS),.VDD(VDD),.Y(g26692),.A(I34683));
  NOT NOT1_10506(.VSS(VSS),.VDD(VDD),.Y(I34686),.A(g26398));
  NOT NOT1_10507(.VSS(VSS),.VDD(VDD),.Y(g26693),.A(I34686));
  NOT NOT1_10508(.VSS(VSS),.VDD(VDD),.Y(I34689),.A(g26433));
  NOT NOT1_10509(.VSS(VSS),.VDD(VDD),.Y(g26694),.A(I34689));
  NOT NOT1_10510(.VSS(VSS),.VDD(VDD),.Y(I34692),.A(g26102));
  NOT NOT1_10511(.VSS(VSS),.VDD(VDD),.Y(g26695),.A(I34692));
  NOT NOT1_10512(.VSS(VSS),.VDD(VDD),.Y(I34695),.A(g26167));
  NOT NOT1_10513(.VSS(VSS),.VDD(VDD),.Y(g26696),.A(I34695));
  NOT NOT1_10514(.VSS(VSS),.VDD(VDD),.Y(I34698),.A(g26181));
  NOT NOT1_10515(.VSS(VSS),.VDD(VDD),.Y(g26697),.A(I34698));
  NOT NOT1_10516(.VSS(VSS),.VDD(VDD),.Y(I34701),.A(g26193));
  NOT NOT1_10517(.VSS(VSS),.VDD(VDD),.Y(g26698),.A(I34701));
  NOT NOT1_10518(.VSS(VSS),.VDD(VDD),.Y(I34704),.A(g26182));
  NOT NOT1_10519(.VSS(VSS),.VDD(VDD),.Y(g26699),.A(I34704));
  NOT NOT1_10520(.VSS(VSS),.VDD(VDD),.Y(I34707),.A(g26194));
  NOT NOT1_10521(.VSS(VSS),.VDD(VDD),.Y(g26700),.A(I34707));
  NOT NOT1_10522(.VSS(VSS),.VDD(VDD),.Y(I34710),.A(g26214));
  NOT NOT1_10523(.VSS(VSS),.VDD(VDD),.Y(g26701),.A(I34710));
  NOT NOT1_10524(.VSS(VSS),.VDD(VDD),.Y(I34713),.A(g26195));
  NOT NOT1_10525(.VSS(VSS),.VDD(VDD),.Y(g26702),.A(I34713));
  NOT NOT1_10526(.VSS(VSS),.VDD(VDD),.Y(I34716),.A(g26215));
  NOT NOT1_10527(.VSS(VSS),.VDD(VDD),.Y(g26703),.A(I34716));
  NOT NOT1_10528(.VSS(VSS),.VDD(VDD),.Y(I34719),.A(g26238));
  NOT NOT1_10529(.VSS(VSS),.VDD(VDD),.Y(g26704),.A(I34719));
  NOT NOT1_10530(.VSS(VSS),.VDD(VDD),.Y(I34722),.A(g26216));
  NOT NOT1_10531(.VSS(VSS),.VDD(VDD),.Y(g26705),.A(I34722));
  NOT NOT1_10532(.VSS(VSS),.VDD(VDD),.Y(I34725),.A(g26239));
  NOT NOT1_10533(.VSS(VSS),.VDD(VDD),.Y(g26706),.A(I34725));
  NOT NOT1_10534(.VSS(VSS),.VDD(VDD),.Y(I34728),.A(g26264));
  NOT NOT1_10535(.VSS(VSS),.VDD(VDD),.Y(g26707),.A(I34728));
  NOT NOT1_10536(.VSS(VSS),.VDD(VDD),.Y(I34731),.A(g26341));
  NOT NOT1_10537(.VSS(VSS),.VDD(VDD),.Y(g26708),.A(I34731));
  NOT NOT1_10538(.VSS(VSS),.VDD(VDD),.Y(I34734),.A(g26407));
  NOT NOT1_10539(.VSS(VSS),.VDD(VDD),.Y(g26709),.A(I34734));
  NOT NOT1_10540(.VSS(VSS),.VDD(VDD),.Y(I34737),.A(g26439));
  NOT NOT1_10541(.VSS(VSS),.VDD(VDD),.Y(g26710),.A(I34737));
  NOT NOT1_10542(.VSS(VSS),.VDD(VDD),.Y(I34740),.A(g26465));
  NOT NOT1_10543(.VSS(VSS),.VDD(VDD),.Y(g26711),.A(I34740));
  NOT NOT1_10544(.VSS(VSS),.VDD(VDD),.Y(I34743),.A(g26118));
  NOT NOT1_10545(.VSS(VSS),.VDD(VDD),.Y(g26712),.A(I34743));
  NOT NOT1_10546(.VSS(VSS),.VDD(VDD),.Y(I34746),.A(g26187));
  NOT NOT1_10547(.VSS(VSS),.VDD(VDD),.Y(g26713),.A(I34746));
  NOT NOT1_10548(.VSS(VSS),.VDD(VDD),.Y(I34749),.A(g26205));
  NOT NOT1_10549(.VSS(VSS),.VDD(VDD),.Y(g26714),.A(I34749));
  NOT NOT1_10550(.VSS(VSS),.VDD(VDD),.Y(I34752),.A(g26220));
  NOT NOT1_10551(.VSS(VSS),.VDD(VDD),.Y(g26715),.A(I34752));
  NOT NOT1_10552(.VSS(VSS),.VDD(VDD),.Y(I34755),.A(g26206));
  NOT NOT1_10553(.VSS(VSS),.VDD(VDD),.Y(g26716),.A(I34755));
  NOT NOT1_10554(.VSS(VSS),.VDD(VDD),.Y(I34758),.A(g26221));
  NOT NOT1_10555(.VSS(VSS),.VDD(VDD),.Y(g26717),.A(I34758));
  NOT NOT1_10556(.VSS(VSS),.VDD(VDD),.Y(I34761),.A(g26245));
  NOT NOT1_10557(.VSS(VSS),.VDD(VDD),.Y(g26718),.A(I34761));
  NOT NOT1_10558(.VSS(VSS),.VDD(VDD),.Y(I34764),.A(g26222));
  NOT NOT1_10559(.VSS(VSS),.VDD(VDD),.Y(g26719),.A(I34764));
  NOT NOT1_10560(.VSS(VSS),.VDD(VDD),.Y(I34767),.A(g26246));
  NOT NOT1_10561(.VSS(VSS),.VDD(VDD),.Y(g26720),.A(I34767));
  NOT NOT1_10562(.VSS(VSS),.VDD(VDD),.Y(I34770),.A(g26276));
  NOT NOT1_10563(.VSS(VSS),.VDD(VDD),.Y(g26721),.A(I34770));
  NOT NOT1_10564(.VSS(VSS),.VDD(VDD),.Y(I34773),.A(g26247));
  NOT NOT1_10565(.VSS(VSS),.VDD(VDD),.Y(g26722),.A(I34773));
  NOT NOT1_10566(.VSS(VSS),.VDD(VDD),.Y(I34776),.A(g26277));
  NOT NOT1_10567(.VSS(VSS),.VDD(VDD),.Y(g26723),.A(I34776));
  NOT NOT1_10568(.VSS(VSS),.VDD(VDD),.Y(I34779),.A(g26308));
  NOT NOT1_10569(.VSS(VSS),.VDD(VDD),.Y(g26724),.A(I34779));
  NOT NOT1_10570(.VSS(VSS),.VDD(VDD),.Y(I34782),.A(g26385));
  NOT NOT1_10571(.VSS(VSS),.VDD(VDD),.Y(g26725),.A(I34782));
  NOT NOT1_10572(.VSS(VSS),.VDD(VDD),.Y(I34785),.A(g26448));
  NOT NOT1_10573(.VSS(VSS),.VDD(VDD),.Y(g26726),.A(I34785));
  NOT NOT1_10574(.VSS(VSS),.VDD(VDD),.Y(I34788),.A(g26471));
  NOT NOT1_10575(.VSS(VSS),.VDD(VDD),.Y(g26727),.A(I34788));
  NOT NOT1_10576(.VSS(VSS),.VDD(VDD),.Y(I34791),.A(g26489));
  NOT NOT1_10577(.VSS(VSS),.VDD(VDD),.Y(g26728),.A(I34791));
  NOT NOT1_10578(.VSS(VSS),.VDD(VDD),.Y(I34794),.A(g26125));
  NOT NOT1_10579(.VSS(VSS),.VDD(VDD),.Y(g26729),.A(I34794));
  NOT NOT1_10580(.VSS(VSS),.VDD(VDD),.Y(I34797),.A(g26208));
  NOT NOT1_10581(.VSS(VSS),.VDD(VDD),.Y(g26730),.A(I34797));
  NOT NOT1_10582(.VSS(VSS),.VDD(VDD),.Y(I34800),.A(g26229));
  NOT NOT1_10583(.VSS(VSS),.VDD(VDD),.Y(g26731),.A(I34800));
  NOT NOT1_10584(.VSS(VSS),.VDD(VDD),.Y(I34803),.A(g26248));
  NOT NOT1_10585(.VSS(VSS),.VDD(VDD),.Y(g26732),.A(I34803));
  NOT NOT1_10586(.VSS(VSS),.VDD(VDD),.Y(I34806),.A(g26230));
  NOT NOT1_10587(.VSS(VSS),.VDD(VDD),.Y(g26733),.A(I34806));
  NOT NOT1_10588(.VSS(VSS),.VDD(VDD),.Y(I34809),.A(g26249));
  NOT NOT1_10589(.VSS(VSS),.VDD(VDD),.Y(g26734),.A(I34809));
  NOT NOT1_10590(.VSS(VSS),.VDD(VDD),.Y(I34812),.A(g26280));
  NOT NOT1_10591(.VSS(VSS),.VDD(VDD),.Y(g26735),.A(I34812));
  NOT NOT1_10592(.VSS(VSS),.VDD(VDD),.Y(I34815),.A(g26250));
  NOT NOT1_10593(.VSS(VSS),.VDD(VDD),.Y(g26736),.A(I34815));
  NOT NOT1_10594(.VSS(VSS),.VDD(VDD),.Y(I34818),.A(g26281));
  NOT NOT1_10595(.VSS(VSS),.VDD(VDD),.Y(g26737),.A(I34818));
  NOT NOT1_10596(.VSS(VSS),.VDD(VDD),.Y(I34821),.A(g26314));
  NOT NOT1_10597(.VSS(VSS),.VDD(VDD),.Y(g26738),.A(I34821));
  NOT NOT1_10598(.VSS(VSS),.VDD(VDD),.Y(I34824),.A(g26282));
  NOT NOT1_10599(.VSS(VSS),.VDD(VDD),.Y(g26739),.A(I34824));
  NOT NOT1_10600(.VSS(VSS),.VDD(VDD),.Y(I34827),.A(g26315));
  NOT NOT1_10601(.VSS(VSS),.VDD(VDD),.Y(g26740),.A(I34827));
  NOT NOT1_10602(.VSS(VSS),.VDD(VDD),.Y(I34830),.A(g26349));
  NOT NOT1_10603(.VSS(VSS),.VDD(VDD),.Y(g26741),.A(I34830));
  NOT NOT1_10604(.VSS(VSS),.VDD(VDD),.Y(I34833),.A(g26428));
  NOT NOT1_10605(.VSS(VSS),.VDD(VDD),.Y(g26742),.A(I34833));
  NOT NOT1_10606(.VSS(VSS),.VDD(VDD),.Y(I34836),.A(g26480));
  NOT NOT1_10607(.VSS(VSS),.VDD(VDD),.Y(g26743),.A(I34836));
  NOT NOT1_10608(.VSS(VSS),.VDD(VDD),.Y(I34839),.A(g26495));
  NOT NOT1_10609(.VSS(VSS),.VDD(VDD),.Y(g26744),.A(I34839));
  NOT NOT1_10610(.VSS(VSS),.VDD(VDD),.Y(I34842),.A(g26505));
  NOT NOT1_10611(.VSS(VSS),.VDD(VDD),.Y(g26745),.A(I34842));
  NOT NOT1_10612(.VSS(VSS),.VDD(VDD),.Y(I34845),.A(g26496));
  NOT NOT1_10613(.VSS(VSS),.VDD(VDD),.Y(g26746),.A(I34845));
  NOT NOT1_10614(.VSS(VSS),.VDD(VDD),.Y(I34848),.A(g26506));
  NOT NOT1_10615(.VSS(VSS),.VDD(VDD),.Y(g26747),.A(I34848));
  NOT NOT1_10616(.VSS(VSS),.VDD(VDD),.Y(I34851),.A(g26354));
  NOT NOT1_10617(.VSS(VSS),.VDD(VDD),.Y(g26748),.A(I34851));
  NOT NOT1_10618(.VSS(VSS),.VDD(VDD),.Y(I34854),.A(g26507));
  NOT NOT1_10619(.VSS(VSS),.VDD(VDD),.Y(g26749),.A(I34854));
  NOT NOT1_10620(.VSS(VSS),.VDD(VDD),.Y(I34857),.A(g26355));
  NOT NOT1_10621(.VSS(VSS),.VDD(VDD),.Y(g26750),.A(I34857));
  NOT NOT1_10622(.VSS(VSS),.VDD(VDD),.Y(I34860),.A(g26548));
  NOT NOT1_10623(.VSS(VSS),.VDD(VDD),.Y(g26751),.A(I34860));
  NOT NOT1_10624(.VSS(VSS),.VDD(VDD),.Y(I34863),.A(g26576));
  NOT NOT1_10625(.VSS(VSS),.VDD(VDD),.Y(g26752),.A(I34863));
  NOT NOT1_10626(.VSS(VSS),.VDD(VDD),.Y(I34866),.A(g26618));
  NOT NOT1_10627(.VSS(VSS),.VDD(VDD),.Y(g26753),.A(I34866));
  NOT NOT1_10628(.VSS(VSS),.VDD(VDD),.Y(I34872),.A(g26217));
  NOT NOT1_10629(.VSS(VSS),.VDD(VDD),.Y(g26757),.A(I34872));
  NOT NOT1_10630(.VSS(VSS),.VDD(VDD),.Y(I34879),.A(g26240));
  NOT NOT1_10631(.VSS(VSS),.VDD(VDD),.Y(g26762),.A(I34879));
  NOT NOT1_10632(.VSS(VSS),.VDD(VDD),.Y(I34901),.A(g26295));
  NOT NOT1_10633(.VSS(VSS),.VDD(VDD),.Y(g26782),.A(I34901));
  NOT NOT1_10634(.VSS(VSS),.VDD(VDD),.Y(I34909),.A(g26265));
  NOT NOT1_10635(.VSS(VSS),.VDD(VDD),.Y(g26788),.A(I34909));
  NOT NOT1_10636(.VSS(VSS),.VDD(VDD),.Y(I34916),.A(g26240));
  NOT NOT1_10637(.VSS(VSS),.VDD(VDD),.Y(g26793),.A(I34916));
  NOT NOT1_10638(.VSS(VSS),.VDD(VDD),.Y(I34921),.A(g26217));
  NOT NOT1_10639(.VSS(VSS),.VDD(VDD),.Y(g26796),.A(I34921));
  NOT NOT1_10640(.VSS(VSS),.VDD(VDD),.Y(I34946),.A(g26534));
  NOT NOT1_10641(.VSS(VSS),.VDD(VDD),.Y(g26819),.A(I34946));
  NOT NOT1_10642(.VSS(VSS),.VDD(VDD),.Y(I34957),.A(g26541));
  NOT NOT1_10643(.VSS(VSS),.VDD(VDD),.Y(g26828),.A(I34957));
  NOT NOT1_10644(.VSS(VSS),.VDD(VDD),.Y(I34961),.A(g26545));
  NOT NOT1_10645(.VSS(VSS),.VDD(VDD),.Y(g26830),.A(I34961));
  NOT NOT1_10646(.VSS(VSS),.VDD(VDD),.Y(I34964),.A(g26547));
  NOT NOT1_10647(.VSS(VSS),.VDD(VDD),.Y(g26831),.A(I34964));
  NOT NOT1_10648(.VSS(VSS),.VDD(VDD),.Y(I34967),.A(g26553));
  NOT NOT1_10649(.VSS(VSS),.VDD(VDD),.Y(g26832),.A(I34967));
  NOT NOT1_10650(.VSS(VSS),.VDD(VDD),.Y(I34971),.A(g26557));
  NOT NOT1_10651(.VSS(VSS),.VDD(VDD),.Y(g26834),.A(I34971));
  NOT NOT1_10652(.VSS(VSS),.VDD(VDD),.Y(I34974),.A(g26168));
  NOT NOT1_10653(.VSS(VSS),.VDD(VDD),.Y(g26835),.A(I34974));
  NOT NOT1_10654(.VSS(VSS),.VDD(VDD),.Y(I34977),.A(g26559));
  NOT NOT1_10655(.VSS(VSS),.VDD(VDD),.Y(g26836),.A(I34977));
  NOT NOT1_10656(.VSS(VSS),.VDD(VDD),.Y(I34980),.A(g26458));
  NOT NOT1_10657(.VSS(VSS),.VDD(VDD),.Y(g26837),.A(I34980));
  NOT NOT1_10658(.VSS(VSS),.VDD(VDD),.Y(I34983),.A(g26569));
  NOT NOT1_10659(.VSS(VSS),.VDD(VDD),.Y(g26840),.A(I34983));
  NOT NOT1_10660(.VSS(VSS),.VDD(VDD),.Y(I34986),.A(g26160));
  NOT NOT1_10661(.VSS(VSS),.VDD(VDD),.Y(g26841),.A(I34986));
  NOT NOT1_10662(.VSS(VSS),.VDD(VDD),.Y(I34990),.A(g26573));
  NOT NOT1_10663(.VSS(VSS),.VDD(VDD),.Y(g26843),.A(I34990));
  NOT NOT1_10664(.VSS(VSS),.VDD(VDD),.Y(I34993),.A(g26575));
  NOT NOT1_10665(.VSS(VSS),.VDD(VDD),.Y(g26844),.A(I34993));
  NOT NOT1_10666(.VSS(VSS),.VDD(VDD),.Y(I34997),.A(g26482));
  NOT NOT1_10667(.VSS(VSS),.VDD(VDD),.Y(g26846),.A(I34997));
  NOT NOT1_10668(.VSS(VSS),.VDD(VDD),.Y(I35000),.A(g26336));
  NOT NOT1_10669(.VSS(VSS),.VDD(VDD),.Y(g26849),.A(I35000));
  NOT NOT1_10670(.VSS(VSS),.VDD(VDD),.Y(I35003),.A(g26592));
  NOT NOT1_10671(.VSS(VSS),.VDD(VDD),.Y(g26850),.A(I35003));
  NOT NOT1_10672(.VSS(VSS),.VDD(VDD),.Y(I35007),.A(g26596));
  NOT NOT1_10673(.VSS(VSS),.VDD(VDD),.Y(g26852),.A(I35007));
  NOT NOT1_10674(.VSS(VSS),.VDD(VDD),.Y(I35011),.A(g26304));
  NOT NOT1_10675(.VSS(VSS),.VDD(VDD),.Y(g26854),.A(I35011));
  NOT NOT1_10676(.VSS(VSS),.VDD(VDD),.Y(I35014),.A(g26498));
  NOT NOT1_10677(.VSS(VSS),.VDD(VDD),.Y(g26855),.A(I35014));
  NOT NOT1_10678(.VSS(VSS),.VDD(VDD),.Y(I35017),.A(g26616));
  NOT NOT1_10679(.VSS(VSS),.VDD(VDD),.Y(g26858),.A(I35017));
  NOT NOT1_10680(.VSS(VSS),.VDD(VDD),.Y(I35028),.A(g26513));
  NOT NOT1_10681(.VSS(VSS),.VDD(VDD),.Y(g26861),.A(I35028));
  NOT NOT1_10682(.VSS(VSS),.VDD(VDD),.Y(I35031),.A(g26529));
  NOT NOT1_10683(.VSS(VSS),.VDD(VDD),.Y(g26864),.A(I35031));
  NOT NOT1_10684(.VSS(VSS),.VDD(VDD),.Y(I35049),.A(g26530));
  NOT NOT1_10685(.VSS(VSS),.VDD(VDD),.Y(g26868),.A(I35049));
  NOT NOT1_10686(.VSS(VSS),.VDD(VDD),.Y(I35053),.A(g26655));
  NOT NOT1_10687(.VSS(VSS),.VDD(VDD),.Y(g26872),.A(I35053));
  NOT NOT1_10688(.VSS(VSS),.VDD(VDD),.Y(I35064),.A(g26531));
  NOT NOT1_10689(.VSS(VSS),.VDD(VDD),.Y(g26875),.A(I35064));
  NOT NOT1_10690(.VSS(VSS),.VDD(VDD),.Y(I35067),.A(g26659));
  NOT NOT1_10691(.VSS(VSS),.VDD(VDD),.Y(g26876),.A(I35067));
  NOT NOT1_10692(.VSS(VSS),.VDD(VDD),.Y(I35072),.A(g26661));
  NOT NOT1_10693(.VSS(VSS),.VDD(VDD),.Y(g26881),.A(I35072));
  NOT NOT1_10694(.VSS(VSS),.VDD(VDD),.Y(I35076),.A(g26532));
  NOT NOT1_10695(.VSS(VSS),.VDD(VDD),.Y(g26883),.A(I35076));
  NOT NOT1_10696(.VSS(VSS),.VDD(VDD),.Y(I35079),.A(g26664));
  NOT NOT1_10697(.VSS(VSS),.VDD(VDD),.Y(g26884),.A(I35079));
  NOT NOT1_10698(.VSS(VSS),.VDD(VDD),.Y(I35083),.A(g26665));
  NOT NOT1_10699(.VSS(VSS),.VDD(VDD),.Y(g26886),.A(I35083));
  NOT NOT1_10700(.VSS(VSS),.VDD(VDD),.Y(I35087),.A(g26667));
  NOT NOT1_10701(.VSS(VSS),.VDD(VDD),.Y(g26890),.A(I35087));
  NOT NOT1_10702(.VSS(VSS),.VDD(VDD),.Y(I35092),.A(g26669));
  NOT NOT1_10703(.VSS(VSS),.VDD(VDD),.Y(g26895),.A(I35092));
  NOT NOT1_10704(.VSS(VSS),.VDD(VDD),.Y(I35095),.A(g26670));
  NOT NOT1_10705(.VSS(VSS),.VDD(VDD),.Y(g26896),.A(I35095));
  NOT NOT1_10706(.VSS(VSS),.VDD(VDD),.Y(I35099),.A(g26672));
  NOT NOT1_10707(.VSS(VSS),.VDD(VDD),.Y(g26900),.A(I35099));
  NOT NOT1_10708(.VSS(VSS),.VDD(VDD),.Y(I35106),.A(g26675));
  NOT NOT1_10709(.VSS(VSS),.VDD(VDD),.Y(g26909),.A(I35106));
  NOT NOT1_10710(.VSS(VSS),.VDD(VDD),.Y(I35109),.A(g26676));
  NOT NOT1_10711(.VSS(VSS),.VDD(VDD),.Y(g26910),.A(I35109));
  NOT NOT1_10712(.VSS(VSS),.VDD(VDD),.Y(I35116),.A(g26025));
  NOT NOT1_10713(.VSS(VSS),.VDD(VDD),.Y(g26921),.A(I35116));
  NOT NOT1_10714(.VSS(VSS),.VDD(VDD),.Y(g26922),.A(g26283));
  NOT NOT1_10715(.VSS(VSS),.VDD(VDD),.Y(g26935),.A(g26327));
  NOT NOT1_10716(.VSS(VSS),.VDD(VDD),.Y(g26944),.A(g26374));
  NOT NOT1_10717(.VSS(VSS),.VDD(VDD),.Y(g26950),.A(g26417));
  NOT NOT1_10718(.VSS(VSS),.VDD(VDD),.Y(I35136),.A(g26660));
  NOT NOT1_10719(.VSS(VSS),.VDD(VDD),.Y(g26953),.A(I35136));
  NOT NOT1_10720(.VSS(VSS),.VDD(VDD),.Y(g26954),.A(g26549));
  NOT NOT1_10721(.VSS(VSS),.VDD(VDD),.Y(I35141),.A(g26666));
  NOT NOT1_10722(.VSS(VSS),.VDD(VDD),.Y(g26956),.A(I35141));
  NOT NOT1_10723(.VSS(VSS),.VDD(VDD),.Y(g26957),.A(g26577));
  NOT NOT1_10724(.VSS(VSS),.VDD(VDD),.Y(I35146),.A(g26671));
  NOT NOT1_10725(.VSS(VSS),.VDD(VDD),.Y(g26959),.A(I35146));
  NOT NOT1_10726(.VSS(VSS),.VDD(VDD),.Y(g26960),.A(g26597));
  NOT NOT1_10727(.VSS(VSS),.VDD(VDD),.Y(I35153),.A(g26677));
  NOT NOT1_10728(.VSS(VSS),.VDD(VDD),.Y(g26964),.A(I35153));
  NOT NOT1_10729(.VSS(VSS),.VDD(VDD),.Y(I35172),.A(g26272));
  NOT NOT1_10730(.VSS(VSS),.VDD(VDD),.Y(g26983),.A(I35172));
  NOT NOT1_10731(.VSS(VSS),.VDD(VDD),.Y(g26987),.A(g26056));
  NOT NOT1_10732(.VSS(VSS),.VDD(VDD),.Y(g27010),.A(g26063));
  NOT NOT1_10733(.VSS(VSS),.VDD(VDD),.Y(g27036),.A(g26070));
  NOT NOT1_10734(.VSS(VSS),.VDD(VDD),.Y(g27064),.A(g26076));
  NOT NOT1_10735(.VSS(VSS),.VDD(VDD),.Y(I35254),.A(g26048));
  NOT NOT1_10736(.VSS(VSS),.VDD(VDD),.Y(g27075),.A(I35254));
  NOT NOT1_10737(.VSS(VSS),.VDD(VDD),.Y(I35283),.A(g26031));
  NOT NOT1_10738(.VSS(VSS),.VDD(VDD),.Y(g27102),.A(I35283));
  NOT NOT1_10739(.VSS(VSS),.VDD(VDD),.Y(I35297),.A(g26199));
  NOT NOT1_10740(.VSS(VSS),.VDD(VDD),.Y(g27114),.A(I35297));
  NOT NOT1_10741(.VSS(VSS),.VDD(VDD),.Y(I35301),.A(g26037));
  NOT NOT1_10742(.VSS(VSS),.VDD(VDD),.Y(g27116),.A(I35301));
  NOT NOT1_10743(.VSS(VSS),.VDD(VDD),.Y(I35313),.A(g26534));
  NOT NOT1_10744(.VSS(VSS),.VDD(VDD),.Y(g27126),.A(I35313));
  NOT NOT1_10745(.VSS(VSS),.VDD(VDD),.Y(I35319),.A(g26183));
  NOT NOT1_10746(.VSS(VSS),.VDD(VDD),.Y(g27132),.A(I35319));
  NOT NOT1_10747(.VSS(VSS),.VDD(VDD),.Y(g27133),.A(g26105));
  NOT NOT1_10748(.VSS(VSS),.VDD(VDD),.Y(g27134),.A(g26175));
  NOT NOT1_10749(.VSS(VSS),.VDD(VDD),.Y(g27135),.A(g26178));
  NOT NOT1_10750(.VSS(VSS),.VDD(VDD),.Y(g27136),.A(g26196));
  NOT NOT1_10751(.VSS(VSS),.VDD(VDD),.Y(g27137),.A(g26202));
  NOT NOT1_10752(.VSS(VSS),.VDD(VDD),.Y(g27138),.A(g26223));
  NOT NOT1_10753(.VSS(VSS),.VDD(VDD),.Y(g27139),.A(g26226));
  NOT NOT1_10754(.VSS(VSS),.VDD(VDD),.Y(g27140),.A(g26136));
  NOT NOT1_10755(.VSS(VSS),.VDD(VDD),.Y(g27141),.A(g26251));
  NOT NOT1_10756(.VSS(VSS),.VDD(VDD),.Y(g27142),.A(g26254));
  NOT NOT1_10757(.VSS(VSS),.VDD(VDD),.Y(g27143),.A(g26150));
  NOT NOT1_10758(.VSS(VSS),.VDD(VDD),.Y(I35334),.A(g26106));
  NOT NOT1_10759(.VSS(VSS),.VDD(VDD),.Y(g27145),.A(I35334));
  NOT NOT1_10760(.VSS(VSS),.VDD(VDD),.Y(g27146),.A(g26358));
  NOT NOT1_10761(.VSS(VSS),.VDD(VDD),.Y(g27148),.A(g26393));
  NOT NOT1_10762(.VSS(VSS),.VDD(VDD),.Y(I35341),.A(g26120));
  NOT NOT1_10763(.VSS(VSS),.VDD(VDD),.Y(g27150),.A(I35341));
  NOT NOT1_10764(.VSS(VSS),.VDD(VDD),.Y(g27151),.A(g26401));
  NOT NOT1_10765(.VSS(VSS),.VDD(VDD),.Y(g27153),.A(g26429));
  NOT NOT1_10766(.VSS(VSS),.VDD(VDD),.Y(I35347),.A(g26265));
  NOT NOT1_10767(.VSS(VSS),.VDD(VDD),.Y(g27154),.A(I35347));
  NOT NOT1_10768(.VSS(VSS),.VDD(VDD),.Y(g27155),.A(g26434));
  NOT NOT1_10769(.VSS(VSS),.VDD(VDD),.Y(I35351),.A(g26272));
  NOT NOT1_10770(.VSS(VSS),.VDD(VDD),.Y(g27156),.A(I35351));
  NOT NOT1_10771(.VSS(VSS),.VDD(VDD),.Y(I35355),.A(g26130));
  NOT NOT1_10772(.VSS(VSS),.VDD(VDD),.Y(g27158),.A(I35355));
  NOT NOT1_10773(.VSS(VSS),.VDD(VDD),.Y(g27159),.A(g26442));
  NOT NOT1_10774(.VSS(VSS),.VDD(VDD),.Y(I35360),.A(g26295));
  NOT NOT1_10775(.VSS(VSS),.VDD(VDD),.Y(g27161),.A(I35360));
  NOT NOT1_10776(.VSS(VSS),.VDD(VDD),.Y(g27162),.A(g26461));
  NOT NOT1_10777(.VSS(VSS),.VDD(VDD),.Y(I35364),.A(g26304));
  NOT NOT1_10778(.VSS(VSS),.VDD(VDD),.Y(g27163),.A(I35364));
  NOT NOT1_10779(.VSS(VSS),.VDD(VDD),.Y(g27164),.A(g26466));
  NOT NOT1_10780(.VSS(VSS),.VDD(VDD),.Y(I35369),.A(g26144));
  NOT NOT1_10781(.VSS(VSS),.VDD(VDD),.Y(g27166),.A(I35369));
  NOT NOT1_10782(.VSS(VSS),.VDD(VDD),.Y(g27167),.A(g26474));
  NOT NOT1_10783(.VSS(VSS),.VDD(VDD),.Y(I35373),.A(g26189));
  NOT NOT1_10784(.VSS(VSS),.VDD(VDD),.Y(g27168),.A(I35373));
  NOT NOT1_10785(.VSS(VSS),.VDD(VDD),.Y(I35376),.A(g26336));
  NOT NOT1_10786(.VSS(VSS),.VDD(VDD),.Y(g27171),.A(I35376));
  NOT NOT1_10787(.VSS(VSS),.VDD(VDD),.Y(g27172),.A(g26485));
  NOT NOT1_10788(.VSS(VSS),.VDD(VDD),.Y(g27173),.A(g26490));
  NOT NOT1_10789(.VSS(VSS),.VDD(VDD),.Y(I35383),.A(g26160));
  NOT NOT1_10790(.VSS(VSS),.VDD(VDD),.Y(g27176),.A(I35383));
  NOT NOT1_10791(.VSS(VSS),.VDD(VDD),.Y(g27177),.A(g26501));
  NOT NOT1_10792(.VSS(VSS),.VDD(VDD),.Y(I35389),.A(g26168));
  NOT NOT1_10793(.VSS(VSS),.VDD(VDD),.Y(g27180),.A(I35389));
  NOT NOT1_10794(.VSS(VSS),.VDD(VDD),.Y(I35394),.A(g26183));
  NOT NOT1_10795(.VSS(VSS),.VDD(VDD),.Y(g27183),.A(I35394));
  NOT NOT1_10796(.VSS(VSS),.VDD(VDD),.Y(I35399),.A(g26199));
  NOT NOT1_10797(.VSS(VSS),.VDD(VDD),.Y(g27186),.A(I35399));
  NOT NOT1_10798(.VSS(VSS),.VDD(VDD),.Y(I35404),.A(g26864));
  NOT NOT1_10799(.VSS(VSS),.VDD(VDD),.Y(g27189),.A(I35404));
  NOT NOT1_10800(.VSS(VSS),.VDD(VDD),.Y(I35407),.A(g27145));
  NOT NOT1_10801(.VSS(VSS),.VDD(VDD),.Y(g27190),.A(I35407));
  NOT NOT1_10802(.VSS(VSS),.VDD(VDD),.Y(I35410),.A(g26872));
  NOT NOT1_10803(.VSS(VSS),.VDD(VDD),.Y(g27191),.A(I35410));
  NOT NOT1_10804(.VSS(VSS),.VDD(VDD),.Y(I35413),.A(g26876));
  NOT NOT1_10805(.VSS(VSS),.VDD(VDD),.Y(g27192),.A(I35413));
  NOT NOT1_10806(.VSS(VSS),.VDD(VDD),.Y(I35416),.A(g26884));
  NOT NOT1_10807(.VSS(VSS),.VDD(VDD),.Y(g27193),.A(I35416));
  NOT NOT1_10808(.VSS(VSS),.VDD(VDD),.Y(I35419),.A(g26828));
  NOT NOT1_10809(.VSS(VSS),.VDD(VDD),.Y(g27194),.A(I35419));
  NOT NOT1_10810(.VSS(VSS),.VDD(VDD),.Y(I35422),.A(g26830));
  NOT NOT1_10811(.VSS(VSS),.VDD(VDD),.Y(g27195),.A(I35422));
  NOT NOT1_10812(.VSS(VSS),.VDD(VDD),.Y(I35425),.A(g26832));
  NOT NOT1_10813(.VSS(VSS),.VDD(VDD),.Y(g27196),.A(I35425));
  NOT NOT1_10814(.VSS(VSS),.VDD(VDD),.Y(I35428),.A(g26953));
  NOT NOT1_10815(.VSS(VSS),.VDD(VDD),.Y(g27197),.A(I35428));
  NOT NOT1_10816(.VSS(VSS),.VDD(VDD),.Y(I35431),.A(g26868));
  NOT NOT1_10817(.VSS(VSS),.VDD(VDD),.Y(g27198),.A(I35431));
  NOT NOT1_10818(.VSS(VSS),.VDD(VDD),.Y(I35434),.A(g27150));
  NOT NOT1_10819(.VSS(VSS),.VDD(VDD),.Y(g27199),.A(I35434));
  NOT NOT1_10820(.VSS(VSS),.VDD(VDD),.Y(I35437),.A(g27183));
  NOT NOT1_10821(.VSS(VSS),.VDD(VDD),.Y(g27200),.A(I35437));
  NOT NOT1_10822(.VSS(VSS),.VDD(VDD),.Y(I35440),.A(g27186));
  NOT NOT1_10823(.VSS(VSS),.VDD(VDD),.Y(g27201),.A(I35440));
  NOT NOT1_10824(.VSS(VSS),.VDD(VDD),.Y(I35443),.A(g26757));
  NOT NOT1_10825(.VSS(VSS),.VDD(VDD),.Y(g27202),.A(I35443));
  NOT NOT1_10826(.VSS(VSS),.VDD(VDD),.Y(I35446),.A(g26762));
  NOT NOT1_10827(.VSS(VSS),.VDD(VDD),.Y(g27203),.A(I35446));
  NOT NOT1_10828(.VSS(VSS),.VDD(VDD),.Y(I35449),.A(g27154));
  NOT NOT1_10829(.VSS(VSS),.VDD(VDD),.Y(g27204),.A(I35449));
  NOT NOT1_10830(.VSS(VSS),.VDD(VDD),.Y(I35452),.A(g27161));
  NOT NOT1_10831(.VSS(VSS),.VDD(VDD),.Y(g27205),.A(I35452));
  NOT NOT1_10832(.VSS(VSS),.VDD(VDD),.Y(I35455),.A(g26881));
  NOT NOT1_10833(.VSS(VSS),.VDD(VDD),.Y(g27206),.A(I35455));
  NOT NOT1_10834(.VSS(VSS),.VDD(VDD),.Y(I35458),.A(g26886));
  NOT NOT1_10835(.VSS(VSS),.VDD(VDD),.Y(g27207),.A(I35458));
  NOT NOT1_10836(.VSS(VSS),.VDD(VDD),.Y(I35461),.A(g26895));
  NOT NOT1_10837(.VSS(VSS),.VDD(VDD),.Y(g27208),.A(I35461));
  NOT NOT1_10838(.VSS(VSS),.VDD(VDD),.Y(I35464),.A(g26831));
  NOT NOT1_10839(.VSS(VSS),.VDD(VDD),.Y(g27209),.A(I35464));
  NOT NOT1_10840(.VSS(VSS),.VDD(VDD),.Y(I35467),.A(g26834));
  NOT NOT1_10841(.VSS(VSS),.VDD(VDD),.Y(g27210),.A(I35467));
  NOT NOT1_10842(.VSS(VSS),.VDD(VDD),.Y(I35470),.A(g26840));
  NOT NOT1_10843(.VSS(VSS),.VDD(VDD),.Y(g27211),.A(I35470));
  NOT NOT1_10844(.VSS(VSS),.VDD(VDD),.Y(I35473),.A(g27156));
  NOT NOT1_10845(.VSS(VSS),.VDD(VDD),.Y(g27212),.A(I35473));
  NOT NOT1_10846(.VSS(VSS),.VDD(VDD),.Y(I35476),.A(g27163));
  NOT NOT1_10847(.VSS(VSS),.VDD(VDD),.Y(g27213),.A(I35476));
  NOT NOT1_10848(.VSS(VSS),.VDD(VDD),.Y(I35479),.A(g27171));
  NOT NOT1_10849(.VSS(VSS),.VDD(VDD),.Y(g27214),.A(I35479));
  NOT NOT1_10850(.VSS(VSS),.VDD(VDD),.Y(I35482),.A(g27176));
  NOT NOT1_10851(.VSS(VSS),.VDD(VDD),.Y(g27215),.A(I35482));
  NOT NOT1_10852(.VSS(VSS),.VDD(VDD),.Y(I35485),.A(g27180));
  NOT NOT1_10853(.VSS(VSS),.VDD(VDD),.Y(g27216),.A(I35485));
  NOT NOT1_10854(.VSS(VSS),.VDD(VDD),.Y(I35488),.A(g26819));
  NOT NOT1_10855(.VSS(VSS),.VDD(VDD),.Y(g27217),.A(I35488));
  NOT NOT1_10856(.VSS(VSS),.VDD(VDD),.Y(I35491),.A(g26956));
  NOT NOT1_10857(.VSS(VSS),.VDD(VDD),.Y(g27218),.A(I35491));
  NOT NOT1_10858(.VSS(VSS),.VDD(VDD),.Y(I35494),.A(g26875));
  NOT NOT1_10859(.VSS(VSS),.VDD(VDD),.Y(g27219),.A(I35494));
  NOT NOT1_10860(.VSS(VSS),.VDD(VDD),.Y(I35497),.A(g27158));
  NOT NOT1_10861(.VSS(VSS),.VDD(VDD),.Y(g27220),.A(I35497));
  NOT NOT1_10862(.VSS(VSS),.VDD(VDD),.Y(I35500),.A(g26890));
  NOT NOT1_10863(.VSS(VSS),.VDD(VDD),.Y(g27221),.A(I35500));
  NOT NOT1_10864(.VSS(VSS),.VDD(VDD),.Y(I35503),.A(g26896));
  NOT NOT1_10865(.VSS(VSS),.VDD(VDD),.Y(g27222),.A(I35503));
  NOT NOT1_10866(.VSS(VSS),.VDD(VDD),.Y(I35506),.A(g26909));
  NOT NOT1_10867(.VSS(VSS),.VDD(VDD),.Y(g27223),.A(I35506));
  NOT NOT1_10868(.VSS(VSS),.VDD(VDD),.Y(I35509),.A(g26836));
  NOT NOT1_10869(.VSS(VSS),.VDD(VDD),.Y(g27224),.A(I35509));
  NOT NOT1_10870(.VSS(VSS),.VDD(VDD),.Y(I35512),.A(g26843));
  NOT NOT1_10871(.VSS(VSS),.VDD(VDD),.Y(g27225),.A(I35512));
  NOT NOT1_10872(.VSS(VSS),.VDD(VDD),.Y(I35515),.A(g26850));
  NOT NOT1_10873(.VSS(VSS),.VDD(VDD),.Y(g27226),.A(I35515));
  NOT NOT1_10874(.VSS(VSS),.VDD(VDD),.Y(I35518),.A(g26959));
  NOT NOT1_10875(.VSS(VSS),.VDD(VDD),.Y(g27227),.A(I35518));
  NOT NOT1_10876(.VSS(VSS),.VDD(VDD),.Y(I35521),.A(g26883));
  NOT NOT1_10877(.VSS(VSS),.VDD(VDD),.Y(g27228),.A(I35521));
  NOT NOT1_10878(.VSS(VSS),.VDD(VDD),.Y(I35524),.A(g27166));
  NOT NOT1_10879(.VSS(VSS),.VDD(VDD),.Y(g27229),.A(I35524));
  NOT NOT1_10880(.VSS(VSS),.VDD(VDD),.Y(I35527),.A(g26900));
  NOT NOT1_10881(.VSS(VSS),.VDD(VDD),.Y(g27230),.A(I35527));
  NOT NOT1_10882(.VSS(VSS),.VDD(VDD),.Y(I35530),.A(g26910));
  NOT NOT1_10883(.VSS(VSS),.VDD(VDD),.Y(g27231),.A(I35530));
  NOT NOT1_10884(.VSS(VSS),.VDD(VDD),.Y(I35533),.A(g26921));
  NOT NOT1_10885(.VSS(VSS),.VDD(VDD),.Y(g27232),.A(I35533));
  NOT NOT1_10886(.VSS(VSS),.VDD(VDD),.Y(I35536),.A(g26844));
  NOT NOT1_10887(.VSS(VSS),.VDD(VDD),.Y(g27233),.A(I35536));
  NOT NOT1_10888(.VSS(VSS),.VDD(VDD),.Y(I35539),.A(g26852));
  NOT NOT1_10889(.VSS(VSS),.VDD(VDD),.Y(g27234),.A(I35539));
  NOT NOT1_10890(.VSS(VSS),.VDD(VDD),.Y(I35542),.A(g26858));
  NOT NOT1_10891(.VSS(VSS),.VDD(VDD),.Y(g27235),.A(I35542));
  NOT NOT1_10892(.VSS(VSS),.VDD(VDD),.Y(I35545),.A(g26964));
  NOT NOT1_10893(.VSS(VSS),.VDD(VDD),.Y(g27236),.A(I35545));
  NOT NOT1_10894(.VSS(VSS),.VDD(VDD),.Y(I35548),.A(g27116));
  NOT NOT1_10895(.VSS(VSS),.VDD(VDD),.Y(g27237),.A(I35548));
  NOT NOT1_10896(.VSS(VSS),.VDD(VDD),.Y(I35551),.A(g27075));
  NOT NOT1_10897(.VSS(VSS),.VDD(VDD),.Y(g27238),.A(I35551));
  NOT NOT1_10898(.VSS(VSS),.VDD(VDD),.Y(I35554),.A(g27102));
  NOT NOT1_10899(.VSS(VSS),.VDD(VDD),.Y(g27239),.A(I35554));
  NOT NOT1_10900(.VSS(VSS),.VDD(VDD),.Y(g27349),.A(g27126));
  NOT NOT1_10901(.VSS(VSS),.VDD(VDD),.Y(I35667),.A(g27120));
  NOT NOT1_10902(.VSS(VSS),.VDD(VDD),.Y(g27353),.A(I35667));
  NOT NOT1_10903(.VSS(VSS),.VDD(VDD),.Y(I35673),.A(g27123));
  NOT NOT1_10904(.VSS(VSS),.VDD(VDD),.Y(g27357),.A(I35673));
  NOT NOT1_10905(.VSS(VSS),.VDD(VDD),.Y(I35678),.A(g27129));
  NOT NOT1_10906(.VSS(VSS),.VDD(VDD),.Y(g27360),.A(I35678));
  NOT NOT1_10907(.VSS(VSS),.VDD(VDD),.Y(I35681),.A(g26869));
  NOT NOT1_10908(.VSS(VSS),.VDD(VDD),.Y(g27361),.A(I35681));
  NOT NOT1_10909(.VSS(VSS),.VDD(VDD),.Y(I35686),.A(g27131));
  NOT NOT1_10910(.VSS(VSS),.VDD(VDD),.Y(g27366),.A(I35686));
  NOT NOT1_10911(.VSS(VSS),.VDD(VDD),.Y(I35689),.A(g26878));
  NOT NOT1_10912(.VSS(VSS),.VDD(VDD),.Y(g27367),.A(I35689));
  NOT NOT1_10913(.VSS(VSS),.VDD(VDD),.Y(I35695),.A(g26887));
  NOT NOT1_10914(.VSS(VSS),.VDD(VDD),.Y(g27373),.A(I35695));
  NOT NOT1_10915(.VSS(VSS),.VDD(VDD),.Y(I35698),.A(g26897));
  NOT NOT1_10916(.VSS(VSS),.VDD(VDD),.Y(g27376),.A(I35698));
  NOT NOT1_10917(.VSS(VSS),.VDD(VDD),.Y(I35708),.A(g26974));
  NOT NOT1_10918(.VSS(VSS),.VDD(VDD),.Y(g27380),.A(I35708));
  NOT NOT1_10919(.VSS(VSS),.VDD(VDD),.Y(I35711),.A(g26974));
  NOT NOT1_10920(.VSS(VSS),.VDD(VDD),.Y(g27381),.A(I35711));
  NOT NOT1_10921(.VSS(VSS),.VDD(VDD),.Y(g27383),.A(g27133));
  NOT NOT1_10922(.VSS(VSS),.VDD(VDD),.Y(g27384),.A(g27140));
  NOT NOT1_10923(.VSS(VSS),.VDD(VDD),.Y(I35723),.A(g27168));
  NOT NOT1_10924(.VSS(VSS),.VDD(VDD),.Y(g27385),.A(I35723));
  NOT NOT1_10925(.VSS(VSS),.VDD(VDD),.Y(g27386),.A(g27143));
  NOT NOT1_10926(.VSS(VSS),.VDD(VDD),.Y(I35727),.A(g26902));
  NOT NOT1_10927(.VSS(VSS),.VDD(VDD),.Y(g27387),.A(I35727));
  NOT NOT1_10928(.VSS(VSS),.VDD(VDD),.Y(I35731),.A(g26892));
  NOT NOT1_10929(.VSS(VSS),.VDD(VDD),.Y(g27391),.A(I35731));
  NOT NOT1_10930(.VSS(VSS),.VDD(VDD),.Y(I35737),.A(g26915));
  NOT NOT1_10931(.VSS(VSS),.VDD(VDD),.Y(g27397),.A(I35737));
  NOT NOT1_10932(.VSS(VSS),.VDD(VDD),.Y(I35741),.A(g27118));
  NOT NOT1_10933(.VSS(VSS),.VDD(VDD),.Y(g27401),.A(I35741));
  NOT NOT1_10934(.VSS(VSS),.VDD(VDD),.Y(I35744),.A(g26906));
  NOT NOT1_10935(.VSS(VSS),.VDD(VDD),.Y(g27404),.A(I35744));
  NOT NOT1_10936(.VSS(VSS),.VDD(VDD),.Y(I35750),.A(g26928));
  NOT NOT1_10937(.VSS(VSS),.VDD(VDD),.Y(g27410),.A(I35750));
  NOT NOT1_10938(.VSS(VSS),.VDD(VDD),.Y(I35756),.A(g27117));
  NOT NOT1_10939(.VSS(VSS),.VDD(VDD),.Y(g27416),.A(I35756));
  NOT NOT1_10940(.VSS(VSS),.VDD(VDD),.Y(I35759),.A(g27121));
  NOT NOT1_10941(.VSS(VSS),.VDD(VDD),.Y(g27419),.A(I35759));
  NOT NOT1_10942(.VSS(VSS),.VDD(VDD),.Y(I35762),.A(g26918));
  NOT NOT1_10943(.VSS(VSS),.VDD(VDD),.Y(g27422),.A(I35762));
  NOT NOT1_10944(.VSS(VSS),.VDD(VDD),.Y(I35768),.A(g26941));
  NOT NOT1_10945(.VSS(VSS),.VDD(VDD),.Y(g27428),.A(I35768));
  NOT NOT1_10946(.VSS(VSS),.VDD(VDD),.Y(I35772),.A(g26772));
  NOT NOT1_10947(.VSS(VSS),.VDD(VDD),.Y(g27432),.A(I35772));
  NOT NOT1_10948(.VSS(VSS),.VDD(VDD),.Y(I35777),.A(g27119));
  NOT NOT1_10949(.VSS(VSS),.VDD(VDD),.Y(g27437),.A(I35777));
  NOT NOT1_10950(.VSS(VSS),.VDD(VDD),.Y(I35780),.A(g27124));
  NOT NOT1_10951(.VSS(VSS),.VDD(VDD),.Y(g27440),.A(I35780));
  NOT NOT1_10952(.VSS(VSS),.VDD(VDD),.Y(I35783),.A(g26931));
  NOT NOT1_10953(.VSS(VSS),.VDD(VDD),.Y(g27443),.A(I35783));
  NOT NOT1_10954(.VSS(VSS),.VDD(VDD),.Y(g27449),.A(g26837));
  NOT NOT1_10955(.VSS(VSS),.VDD(VDD),.Y(I35791),.A(g26779));
  NOT NOT1_10956(.VSS(VSS),.VDD(VDD),.Y(g27451),.A(I35791));
  NOT NOT1_10957(.VSS(VSS),.VDD(VDD),.Y(I35796),.A(g27122));
  NOT NOT1_10958(.VSS(VSS),.VDD(VDD),.Y(g27456),.A(I35796));
  NOT NOT1_10959(.VSS(VSS),.VDD(VDD),.Y(I35799),.A(g27130));
  NOT NOT1_10960(.VSS(VSS),.VDD(VDD),.Y(g27459),.A(I35799));
  NOT NOT1_10961(.VSS(VSS),.VDD(VDD),.Y(I35803),.A(g26803));
  NOT NOT1_10962(.VSS(VSS),.VDD(VDD),.Y(g27463),.A(I35803));
  NOT NOT1_10963(.VSS(VSS),.VDD(VDD),.Y(g27465),.A(g26846));
  NOT NOT1_10964(.VSS(VSS),.VDD(VDD),.Y(I35809),.A(g26785));
  NOT NOT1_10965(.VSS(VSS),.VDD(VDD),.Y(g27467),.A(I35809));
  NOT NOT1_10966(.VSS(VSS),.VDD(VDD),.Y(I35814),.A(g27125));
  NOT NOT1_10967(.VSS(VSS),.VDD(VDD),.Y(g27472),.A(I35814));
  NOT NOT1_10968(.VSS(VSS),.VDD(VDD),.Y(I35817),.A(g26922));
  NOT NOT1_10969(.VSS(VSS),.VDD(VDD),.Y(g27475),.A(I35817));
  NOT NOT1_10970(.VSS(VSS),.VDD(VDD),.Y(I35821),.A(g26804));
  NOT NOT1_10971(.VSS(VSS),.VDD(VDD),.Y(g27479),.A(I35821));
  NOT NOT1_10972(.VSS(VSS),.VDD(VDD),.Y(I35824),.A(g26805));
  NOT NOT1_10973(.VSS(VSS),.VDD(VDD),.Y(g27480),.A(I35824));
  NOT NOT1_10974(.VSS(VSS),.VDD(VDD),.Y(I35829),.A(g26806));
  NOT NOT1_10975(.VSS(VSS),.VDD(VDD),.Y(g27483),.A(I35829));
  NOT NOT1_10976(.VSS(VSS),.VDD(VDD),.Y(g27484),.A(g26855));
  NOT NOT1_10977(.VSS(VSS),.VDD(VDD),.Y(I35834),.A(g26792));
  NOT NOT1_10978(.VSS(VSS),.VDD(VDD),.Y(g27486),.A(I35834));
  NOT NOT1_10979(.VSS(VSS),.VDD(VDD),.Y(I35837),.A(g26911));
  NOT NOT1_10980(.VSS(VSS),.VDD(VDD),.Y(g27489),.A(I35837));
  NOT NOT1_10981(.VSS(VSS),.VDD(VDD),.Y(I35841),.A(g26807));
  NOT NOT1_10982(.VSS(VSS),.VDD(VDD),.Y(g27493),.A(I35841));
  NOT NOT1_10983(.VSS(VSS),.VDD(VDD),.Y(I35844),.A(g26808));
  NOT NOT1_10984(.VSS(VSS),.VDD(VDD),.Y(g27494),.A(I35844));
  NOT NOT1_10985(.VSS(VSS),.VDD(VDD),.Y(I35849),.A(g26776));
  NOT NOT1_10986(.VSS(VSS),.VDD(VDD),.Y(g27497),.A(I35849));
  NOT NOT1_10987(.VSS(VSS),.VDD(VDD),.Y(I35852),.A(g26935));
  NOT NOT1_10988(.VSS(VSS),.VDD(VDD),.Y(g27498),.A(I35852));
  NOT NOT1_10989(.VSS(VSS),.VDD(VDD),.Y(I35856),.A(g26809));
  NOT NOT1_10990(.VSS(VSS),.VDD(VDD),.Y(g27502),.A(I35856));
  NOT NOT1_10991(.VSS(VSS),.VDD(VDD),.Y(I35859),.A(g26810));
  NOT NOT1_10992(.VSS(VSS),.VDD(VDD),.Y(g27503),.A(I35859));
  NOT NOT1_10993(.VSS(VSS),.VDD(VDD),.Y(I35863),.A(g26811));
  NOT NOT1_10994(.VSS(VSS),.VDD(VDD),.Y(g27505),.A(I35863));
  NOT NOT1_10995(.VSS(VSS),.VDD(VDD),.Y(g27506),.A(g26861));
  NOT NOT1_10996(.VSS(VSS),.VDD(VDD),.Y(I35868),.A(g26812));
  NOT NOT1_10997(.VSS(VSS),.VDD(VDD),.Y(g27508),.A(I35868));
  NOT NOT1_10998(.VSS(VSS),.VDD(VDD),.Y(I35872),.A(g26925));
  NOT NOT1_10999(.VSS(VSS),.VDD(VDD),.Y(g27510),.A(I35872));
  NOT NOT1_11000(.VSS(VSS),.VDD(VDD),.Y(I35876),.A(g26813));
  NOT NOT1_11001(.VSS(VSS),.VDD(VDD),.Y(g27514),.A(I35876));
  NOT NOT1_11002(.VSS(VSS),.VDD(VDD),.Y(I35879),.A(g26814));
  NOT NOT1_11003(.VSS(VSS),.VDD(VDD),.Y(g27515),.A(I35879));
  NOT NOT1_11004(.VSS(VSS),.VDD(VDD),.Y(I35883),.A(g26781));
  NOT NOT1_11005(.VSS(VSS),.VDD(VDD),.Y(g27517),.A(I35883));
  NOT NOT1_11006(.VSS(VSS),.VDD(VDD),.Y(I35886),.A(g26944));
  NOT NOT1_11007(.VSS(VSS),.VDD(VDD),.Y(g27518),.A(I35886));
  NOT NOT1_11008(.VSS(VSS),.VDD(VDD),.Y(I35890),.A(g26815));
  NOT NOT1_11009(.VSS(VSS),.VDD(VDD),.Y(g27522),.A(I35890));
  NOT NOT1_11010(.VSS(VSS),.VDD(VDD),.Y(I35893),.A(g26816));
  NOT NOT1_11011(.VSS(VSS),.VDD(VDD),.Y(g27523),.A(I35893));
  NOT NOT1_11012(.VSS(VSS),.VDD(VDD),.Y(I35897),.A(g26817));
  NOT NOT1_11013(.VSS(VSS),.VDD(VDD),.Y(g27525),.A(I35897));
  NOT NOT1_11014(.VSS(VSS),.VDD(VDD),.Y(I35900),.A(g26786));
  NOT NOT1_11015(.VSS(VSS),.VDD(VDD),.Y(g27526),.A(I35900));
  NOT NOT1_11016(.VSS(VSS),.VDD(VDD),.Y(I35915),.A(g26818));
  NOT NOT1_11017(.VSS(VSS),.VDD(VDD),.Y(g27533),.A(I35915));
  NOT NOT1_11018(.VSS(VSS),.VDD(VDD),.Y(I35919),.A(g26938));
  NOT NOT1_11019(.VSS(VSS),.VDD(VDD),.Y(g27535),.A(I35919));
  NOT NOT1_11020(.VSS(VSS),.VDD(VDD),.Y(I35923),.A(g26820));
  NOT NOT1_11021(.VSS(VSS),.VDD(VDD),.Y(g27539),.A(I35923));
  NOT NOT1_11022(.VSS(VSS),.VDD(VDD),.Y(I35926),.A(g26821));
  NOT NOT1_11023(.VSS(VSS),.VDD(VDD),.Y(g27540),.A(I35926));
  NOT NOT1_11024(.VSS(VSS),.VDD(VDD),.Y(I35930),.A(g26789));
  NOT NOT1_11025(.VSS(VSS),.VDD(VDD),.Y(g27542),.A(I35930));
  NOT NOT1_11026(.VSS(VSS),.VDD(VDD),.Y(I35933),.A(g26950));
  NOT NOT1_11027(.VSS(VSS),.VDD(VDD),.Y(g27543),.A(I35933));
  NOT NOT1_11028(.VSS(VSS),.VDD(VDD),.Y(I35937),.A(g26822));
  NOT NOT1_11029(.VSS(VSS),.VDD(VDD),.Y(g27547),.A(I35937));
  NOT NOT1_11030(.VSS(VSS),.VDD(VDD),.Y(I35940),.A(g26823));
  NOT NOT1_11031(.VSS(VSS),.VDD(VDD),.Y(g27548),.A(I35940));
  NOT NOT1_11032(.VSS(VSS),.VDD(VDD),.Y(I35953),.A(g26824));
  NOT NOT1_11033(.VSS(VSS),.VDD(VDD),.Y(g27553),.A(I35953));
  NOT NOT1_11034(.VSS(VSS),.VDD(VDD),.Y(I35957),.A(g26947));
  NOT NOT1_11035(.VSS(VSS),.VDD(VDD),.Y(g27555),.A(I35957));
  NOT NOT1_11036(.VSS(VSS),.VDD(VDD),.Y(I35961),.A(g26825));
  NOT NOT1_11037(.VSS(VSS),.VDD(VDD),.Y(g27559),.A(I35961));
  NOT NOT1_11038(.VSS(VSS),.VDD(VDD),.Y(I35964),.A(g26826));
  NOT NOT1_11039(.VSS(VSS),.VDD(VDD),.Y(g27560),.A(I35964));
  NOT NOT1_11040(.VSS(VSS),.VDD(VDD),.Y(I35968),.A(g26795));
  NOT NOT1_11041(.VSS(VSS),.VDD(VDD),.Y(g27562),.A(I35968));
  NOT NOT1_11042(.VSS(VSS),.VDD(VDD),.Y(I35983),.A(g26827));
  NOT NOT1_11043(.VSS(VSS),.VDD(VDD),.Y(g27569),.A(I35983));
  NOT NOT1_11044(.VSS(VSS),.VDD(VDD),.Y(I36008),.A(g26798));
  NOT NOT1_11045(.VSS(VSS),.VDD(VDD),.Y(g27586),.A(I36008));
  NOT NOT1_11046(.VSS(VSS),.VDD(VDD),.Y(g27589),.A(g27168));
  NOT NOT1_11047(.VSS(VSS),.VDD(VDD),.Y(g27590),.A(g27144));
  NOT NOT1_11048(.VSS(VSS),.VDD(VDD),.Y(g27595),.A(g27149));
  NOT NOT1_11049(.VSS(VSS),.VDD(VDD),.Y(g27599),.A(g27147));
  NOT NOT1_11050(.VSS(VSS),.VDD(VDD),.Y(g27604),.A(g27157));
  NOT NOT1_11051(.VSS(VSS),.VDD(VDD),.Y(g27608),.A(g27152));
  NOT NOT1_11052(.VSS(VSS),.VDD(VDD),.Y(g27613),.A(g27165));
  NOT NOT1_11053(.VSS(VSS),.VDD(VDD),.Y(g27617),.A(g27160));
  NOT NOT1_11054(.VSS(VSS),.VDD(VDD),.Y(g27622),.A(g27174));
  NOT NOT1_11055(.VSS(VSS),.VDD(VDD),.Y(I36032),.A(g27113));
  NOT NOT1_11056(.VSS(VSS),.VDD(VDD),.Y(g27632),.A(I36032));
  NOT NOT1_11057(.VSS(VSS),.VDD(VDD),.Y(I36042),.A(g26960));
  NOT NOT1_11058(.VSS(VSS),.VDD(VDD),.Y(g27662),.A(I36042));
  NOT NOT1_11059(.VSS(VSS),.VDD(VDD),.Y(I36046),.A(g26957));
  NOT NOT1_11060(.VSS(VSS),.VDD(VDD),.Y(g27667),.A(I36046));
  NOT NOT1_11061(.VSS(VSS),.VDD(VDD),.Y(I36052),.A(g26954));
  NOT NOT1_11062(.VSS(VSS),.VDD(VDD),.Y(g27674),.A(I36052));
  NOT NOT1_11063(.VSS(VSS),.VDD(VDD),.Y(I36060),.A(g27353));
  NOT NOT1_11064(.VSS(VSS),.VDD(VDD),.Y(g27683),.A(I36060));
  NOT NOT1_11065(.VSS(VSS),.VDD(VDD),.Y(I36063),.A(g27463));
  NOT NOT1_11066(.VSS(VSS),.VDD(VDD),.Y(g27684),.A(I36063));
  NOT NOT1_11067(.VSS(VSS),.VDD(VDD),.Y(I36066),.A(g27479));
  NOT NOT1_11068(.VSS(VSS),.VDD(VDD),.Y(g27685),.A(I36066));
  NOT NOT1_11069(.VSS(VSS),.VDD(VDD),.Y(I36069),.A(g27493));
  NOT NOT1_11070(.VSS(VSS),.VDD(VDD),.Y(g27686),.A(I36069));
  NOT NOT1_11071(.VSS(VSS),.VDD(VDD),.Y(I36072),.A(g27480));
  NOT NOT1_11072(.VSS(VSS),.VDD(VDD),.Y(g27687),.A(I36072));
  NOT NOT1_11073(.VSS(VSS),.VDD(VDD),.Y(I36075),.A(g27494));
  NOT NOT1_11074(.VSS(VSS),.VDD(VDD),.Y(g27688),.A(I36075));
  NOT NOT1_11075(.VSS(VSS),.VDD(VDD),.Y(I36078),.A(g27508));
  NOT NOT1_11076(.VSS(VSS),.VDD(VDD),.Y(g27689),.A(I36078));
  NOT NOT1_11077(.VSS(VSS),.VDD(VDD),.Y(I36081),.A(g27497));
  NOT NOT1_11078(.VSS(VSS),.VDD(VDD),.Y(g27690),.A(I36081));
  NOT NOT1_11079(.VSS(VSS),.VDD(VDD),.Y(I36084),.A(g27357));
  NOT NOT1_11080(.VSS(VSS),.VDD(VDD),.Y(g27691),.A(I36084));
  NOT NOT1_11081(.VSS(VSS),.VDD(VDD),.Y(I36087),.A(g27483));
  NOT NOT1_11082(.VSS(VSS),.VDD(VDD),.Y(g27692),.A(I36087));
  NOT NOT1_11083(.VSS(VSS),.VDD(VDD),.Y(I36090),.A(g27502));
  NOT NOT1_11084(.VSS(VSS),.VDD(VDD),.Y(g27693),.A(I36090));
  NOT NOT1_11085(.VSS(VSS),.VDD(VDD),.Y(I36093),.A(g27514));
  NOT NOT1_11086(.VSS(VSS),.VDD(VDD),.Y(g27694),.A(I36093));
  NOT NOT1_11087(.VSS(VSS),.VDD(VDD),.Y(I36096),.A(g27503));
  NOT NOT1_11088(.VSS(VSS),.VDD(VDD),.Y(g27695),.A(I36096));
  NOT NOT1_11089(.VSS(VSS),.VDD(VDD),.Y(I36099),.A(g27515));
  NOT NOT1_11090(.VSS(VSS),.VDD(VDD),.Y(g27696),.A(I36099));
  NOT NOT1_11091(.VSS(VSS),.VDD(VDD),.Y(I36102),.A(g27533));
  NOT NOT1_11092(.VSS(VSS),.VDD(VDD),.Y(g27697),.A(I36102));
  NOT NOT1_11093(.VSS(VSS),.VDD(VDD),.Y(I36105),.A(g27517));
  NOT NOT1_11094(.VSS(VSS),.VDD(VDD),.Y(g27698),.A(I36105));
  NOT NOT1_11095(.VSS(VSS),.VDD(VDD),.Y(I36108),.A(g27360));
  NOT NOT1_11096(.VSS(VSS),.VDD(VDD),.Y(g27699),.A(I36108));
  NOT NOT1_11097(.VSS(VSS),.VDD(VDD),.Y(I36111),.A(g27505));
  NOT NOT1_11098(.VSS(VSS),.VDD(VDD),.Y(g27700),.A(I36111));
  NOT NOT1_11099(.VSS(VSS),.VDD(VDD),.Y(I36114),.A(g27522));
  NOT NOT1_11100(.VSS(VSS),.VDD(VDD),.Y(g27701),.A(I36114));
  NOT NOT1_11101(.VSS(VSS),.VDD(VDD),.Y(I36117),.A(g27539));
  NOT NOT1_11102(.VSS(VSS),.VDD(VDD),.Y(g27702),.A(I36117));
  NOT NOT1_11103(.VSS(VSS),.VDD(VDD),.Y(I36120),.A(g27523));
  NOT NOT1_11104(.VSS(VSS),.VDD(VDD),.Y(g27703),.A(I36120));
  NOT NOT1_11105(.VSS(VSS),.VDD(VDD),.Y(I36123),.A(g27540));
  NOT NOT1_11106(.VSS(VSS),.VDD(VDD),.Y(g27704),.A(I36123));
  NOT NOT1_11107(.VSS(VSS),.VDD(VDD),.Y(I36126),.A(g27553));
  NOT NOT1_11108(.VSS(VSS),.VDD(VDD),.Y(g27705),.A(I36126));
  NOT NOT1_11109(.VSS(VSS),.VDD(VDD),.Y(I36129),.A(g27542));
  NOT NOT1_11110(.VSS(VSS),.VDD(VDD),.Y(g27706),.A(I36129));
  NOT NOT1_11111(.VSS(VSS),.VDD(VDD),.Y(I36132),.A(g27366));
  NOT NOT1_11112(.VSS(VSS),.VDD(VDD),.Y(g27707),.A(I36132));
  NOT NOT1_11113(.VSS(VSS),.VDD(VDD),.Y(I36135),.A(g27525));
  NOT NOT1_11114(.VSS(VSS),.VDD(VDD),.Y(g27708),.A(I36135));
  NOT NOT1_11115(.VSS(VSS),.VDD(VDD),.Y(I36138),.A(g27547));
  NOT NOT1_11116(.VSS(VSS),.VDD(VDD),.Y(g27709),.A(I36138));
  NOT NOT1_11117(.VSS(VSS),.VDD(VDD),.Y(I36141),.A(g27559));
  NOT NOT1_11118(.VSS(VSS),.VDD(VDD),.Y(g27710),.A(I36141));
  NOT NOT1_11119(.VSS(VSS),.VDD(VDD),.Y(I36144),.A(g27548));
  NOT NOT1_11120(.VSS(VSS),.VDD(VDD),.Y(g27711),.A(I36144));
  NOT NOT1_11121(.VSS(VSS),.VDD(VDD),.Y(I36147),.A(g27560));
  NOT NOT1_11122(.VSS(VSS),.VDD(VDD),.Y(g27712),.A(I36147));
  NOT NOT1_11123(.VSS(VSS),.VDD(VDD),.Y(I36150),.A(g27569));
  NOT NOT1_11124(.VSS(VSS),.VDD(VDD),.Y(g27713),.A(I36150));
  NOT NOT1_11125(.VSS(VSS),.VDD(VDD),.Y(I36153),.A(g27562));
  NOT NOT1_11126(.VSS(VSS),.VDD(VDD),.Y(g27714),.A(I36153));
  NOT NOT1_11127(.VSS(VSS),.VDD(VDD),.Y(I36156),.A(g27586));
  NOT NOT1_11128(.VSS(VSS),.VDD(VDD),.Y(g27715),.A(I36156));
  NOT NOT1_11129(.VSS(VSS),.VDD(VDD),.Y(I36159),.A(g27526));
  NOT NOT1_11130(.VSS(VSS),.VDD(VDD),.Y(g27716),.A(I36159));
  NOT NOT1_11131(.VSS(VSS),.VDD(VDD),.Y(I36162),.A(g27385));
  NOT NOT1_11132(.VSS(VSS),.VDD(VDD),.Y(g27717),.A(I36162));
  NOT NOT1_11133(.VSS(VSS),.VDD(VDD),.Y(g27748),.A(g27632));
  NOT NOT1_11134(.VSS(VSS),.VDD(VDD),.Y(I36213),.A(g27571));
  NOT NOT1_11135(.VSS(VSS),.VDD(VDD),.Y(g27776),.A(I36213));
  NOT NOT1_11136(.VSS(VSS),.VDD(VDD),.Y(I36217),.A(g27580));
  NOT NOT1_11137(.VSS(VSS),.VDD(VDD),.Y(g27780),.A(I36217));
  NOT NOT1_11138(.VSS(VSS),.VDD(VDD),.Y(I36221),.A(g27662));
  NOT NOT1_11139(.VSS(VSS),.VDD(VDD),.Y(g27784),.A(I36221));
  NOT NOT1_11140(.VSS(VSS),.VDD(VDD),.Y(I36224),.A(g27589));
  NOT NOT1_11141(.VSS(VSS),.VDD(VDD),.Y(g27785),.A(I36224));
  NOT NOT1_11142(.VSS(VSS),.VDD(VDD),.Y(I36227),.A(g27594));
  NOT NOT1_11143(.VSS(VSS),.VDD(VDD),.Y(g27786),.A(I36227));
  NOT NOT1_11144(.VSS(VSS),.VDD(VDD),.Y(I36230),.A(g27583));
  NOT NOT1_11145(.VSS(VSS),.VDD(VDD),.Y(g27787),.A(I36230));
  NOT NOT1_11146(.VSS(VSS),.VDD(VDD),.Y(I36234),.A(g27667));
  NOT NOT1_11147(.VSS(VSS),.VDD(VDD),.Y(g27791),.A(I36234));
  NOT NOT1_11148(.VSS(VSS),.VDD(VDD),.Y(I36237),.A(g27662));
  NOT NOT1_11149(.VSS(VSS),.VDD(VDD),.Y(g27792),.A(I36237));
  NOT NOT1_11150(.VSS(VSS),.VDD(VDD),.Y(I36240),.A(g27603));
  NOT NOT1_11151(.VSS(VSS),.VDD(VDD),.Y(g27793),.A(I36240));
  NOT NOT1_11152(.VSS(VSS),.VDD(VDD),.Y(I36243),.A(g27587));
  NOT NOT1_11153(.VSS(VSS),.VDD(VDD),.Y(g27794),.A(I36243));
  NOT NOT1_11154(.VSS(VSS),.VDD(VDD),.Y(I36246),.A(g27674));
  NOT NOT1_11155(.VSS(VSS),.VDD(VDD),.Y(g27797),.A(I36246));
  NOT NOT1_11156(.VSS(VSS),.VDD(VDD),.Y(I36250),.A(g27612));
  NOT NOT1_11157(.VSS(VSS),.VDD(VDD),.Y(g27799),.A(I36250));
  NOT NOT1_11158(.VSS(VSS),.VDD(VDD),.Y(I36253),.A(g27674));
  NOT NOT1_11159(.VSS(VSS),.VDD(VDD),.Y(g27800),.A(I36253));
  NOT NOT1_11160(.VSS(VSS),.VDD(VDD),.Y(I36264),.A(g27621));
  NOT NOT1_11161(.VSS(VSS),.VDD(VDD),.Y(g27805),.A(I36264));
  NOT NOT1_11162(.VSS(VSS),.VDD(VDD),.Y(I36267),.A(g27395));
  NOT NOT1_11163(.VSS(VSS),.VDD(VDD),.Y(g27806),.A(I36267));
  NOT NOT1_11164(.VSS(VSS),.VDD(VDD),.Y(I36280),.A(g27390));
  NOT NOT1_11165(.VSS(VSS),.VDD(VDD),.Y(g27817),.A(I36280));
  NOT NOT1_11166(.VSS(VSS),.VDD(VDD),.Y(I36283),.A(g27408));
  NOT NOT1_11167(.VSS(VSS),.VDD(VDD),.Y(g27820),.A(I36283));
  NOT NOT1_11168(.VSS(VSS),.VDD(VDD),.Y(I36296),.A(g27626));
  NOT NOT1_11169(.VSS(VSS),.VDD(VDD),.Y(g27831),.A(I36296));
  NOT NOT1_11170(.VSS(VSS),.VDD(VDD),.Y(I36307),.A(g27400));
  NOT NOT1_11171(.VSS(VSS),.VDD(VDD),.Y(g27839),.A(I36307));
  NOT NOT1_11172(.VSS(VSS),.VDD(VDD),.Y(I36311),.A(g27426));
  NOT NOT1_11173(.VSS(VSS),.VDD(VDD),.Y(g27843),.A(I36311));
  NOT NOT1_11174(.VSS(VSS),.VDD(VDD),.Y(I36321),.A(g27627));
  NOT NOT1_11175(.VSS(VSS),.VDD(VDD),.Y(g27847),.A(I36321));
  NOT NOT1_11176(.VSS(VSS),.VDD(VDD),.Y(I36327),.A(g27413));
  NOT NOT1_11177(.VSS(VSS),.VDD(VDD),.Y(g27858),.A(I36327));
  NOT NOT1_11178(.VSS(VSS),.VDD(VDD),.Y(I36330),.A(g27447));
  NOT NOT1_11179(.VSS(VSS),.VDD(VDD),.Y(g27861),.A(I36330));
  NOT NOT1_11180(.VSS(VSS),.VDD(VDD),.Y(I36337),.A(g27628));
  NOT NOT1_11181(.VSS(VSS),.VDD(VDD),.Y(g27872),.A(I36337));
  NOT NOT1_11182(.VSS(VSS),.VDD(VDD),.Y(I36341),.A(g27431));
  NOT NOT1_11183(.VSS(VSS),.VDD(VDD),.Y(g27879),.A(I36341));
  NOT NOT1_11184(.VSS(VSS),.VDD(VDD),.Y(I36347),.A(g27630));
  NOT NOT1_11185(.VSS(VSS),.VDD(VDD),.Y(g27889),.A(I36347));
  NOT NOT1_11186(.VSS(VSS),.VDD(VDD),.Y(I36354),.A(g27662));
  NOT NOT1_11187(.VSS(VSS),.VDD(VDD),.Y(g27903),.A(I36354));
  NOT NOT1_11188(.VSS(VSS),.VDD(VDD),.Y(I36358),.A(g27672));
  NOT NOT1_11189(.VSS(VSS),.VDD(VDD),.Y(g27905),.A(I36358));
  NOT NOT1_11190(.VSS(VSS),.VDD(VDD),.Y(I36362),.A(g27667));
  NOT NOT1_11191(.VSS(VSS),.VDD(VDD),.Y(g27907),.A(I36362));
  NOT NOT1_11192(.VSS(VSS),.VDD(VDD),.Y(I36367),.A(g27678));
  NOT NOT1_11193(.VSS(VSS),.VDD(VDD),.Y(g27910),.A(I36367));
  NOT NOT1_11194(.VSS(VSS),.VDD(VDD),.Y(I36371),.A(g27674));
  NOT NOT1_11195(.VSS(VSS),.VDD(VDD),.Y(g27912),.A(I36371));
  NOT NOT1_11196(.VSS(VSS),.VDD(VDD),.Y(I36379),.A(g27682));
  NOT NOT1_11197(.VSS(VSS),.VDD(VDD),.Y(g27918),.A(I36379));
  NOT NOT1_11198(.VSS(VSS),.VDD(VDD),.Y(I36382),.A(g27563));
  NOT NOT1_11199(.VSS(VSS),.VDD(VDD),.Y(g27919),.A(I36382));
  NOT NOT1_11200(.VSS(VSS),.VDD(VDD),.Y(I36390),.A(g27243));
  NOT NOT1_11201(.VSS(VSS),.VDD(VDD),.Y(g27927),.A(I36390));
  NOT NOT1_11202(.VSS(VSS),.VDD(VDD),.Y(I36393),.A(g27572));
  NOT NOT1_11203(.VSS(VSS),.VDD(VDD),.Y(g27928),.A(I36393));
  NOT NOT1_11204(.VSS(VSS),.VDD(VDD),.Y(I36397),.A(g27574));
  NOT NOT1_11205(.VSS(VSS),.VDD(VDD),.Y(g27932),.A(I36397));
  NOT NOT1_11206(.VSS(VSS),.VDD(VDD),.Y(I36404),.A(g27450));
  NOT NOT1_11207(.VSS(VSS),.VDD(VDD),.Y(g27939),.A(I36404));
  NOT NOT1_11208(.VSS(VSS),.VDD(VDD),.Y(I36407),.A(g27581));
  NOT NOT1_11209(.VSS(VSS),.VDD(VDD),.Y(g27942),.A(I36407));
  NOT NOT1_11210(.VSS(VSS),.VDD(VDD),.Y(I36411),.A(g27582));
  NOT NOT1_11211(.VSS(VSS),.VDD(VDD),.Y(g27946),.A(I36411));
  NOT NOT1_11212(.VSS(VSS),.VDD(VDD),.Y(I36417),.A(g27462));
  NOT NOT1_11213(.VSS(VSS),.VDD(VDD),.Y(g27952),.A(I36417));
  NOT NOT1_11214(.VSS(VSS),.VDD(VDD),.Y(I36420),.A(g27253));
  NOT NOT1_11215(.VSS(VSS),.VDD(VDD),.Y(g27955),.A(I36420));
  NOT NOT1_11216(.VSS(VSS),.VDD(VDD),.Y(I36423),.A(g27466));
  NOT NOT1_11217(.VSS(VSS),.VDD(VDD),.Y(g27956),.A(I36423));
  NOT NOT1_11218(.VSS(VSS),.VDD(VDD),.Y(I36426),.A(g27584));
  NOT NOT1_11219(.VSS(VSS),.VDD(VDD),.Y(g27959),.A(I36426));
  NOT NOT1_11220(.VSS(VSS),.VDD(VDD),.Y(I36432),.A(g27585));
  NOT NOT1_11221(.VSS(VSS),.VDD(VDD),.Y(g27965),.A(I36432));
  NOT NOT1_11222(.VSS(VSS),.VDD(VDD),.Y(g27969),.A(g27361));
  NOT NOT1_11223(.VSS(VSS),.VDD(VDD),.Y(I36438),.A(g27255));
  NOT NOT1_11224(.VSS(VSS),.VDD(VDD),.Y(g27971),.A(I36438));
  NOT NOT1_11225(.VSS(VSS),.VDD(VDD),.Y(I36441),.A(g27256));
  NOT NOT1_11226(.VSS(VSS),.VDD(VDD),.Y(g27972),.A(I36441));
  NOT NOT1_11227(.VSS(VSS),.VDD(VDD),.Y(I36444),.A(g27482));
  NOT NOT1_11228(.VSS(VSS),.VDD(VDD),.Y(g27973),.A(I36444));
  NOT NOT1_11229(.VSS(VSS),.VDD(VDD),.Y(I36447),.A(g27257));
  NOT NOT1_11230(.VSS(VSS),.VDD(VDD),.Y(g27976),.A(I36447));
  NOT NOT1_11231(.VSS(VSS),.VDD(VDD),.Y(I36450),.A(g27485));
  NOT NOT1_11232(.VSS(VSS),.VDD(VDD),.Y(g27977),.A(I36450));
  NOT NOT1_11233(.VSS(VSS),.VDD(VDD),.Y(I36454),.A(g27588));
  NOT NOT1_11234(.VSS(VSS),.VDD(VDD),.Y(g27981),.A(I36454));
  NOT NOT1_11235(.VSS(VSS),.VDD(VDD),.Y(I36459),.A(g27258));
  NOT NOT1_11236(.VSS(VSS),.VDD(VDD),.Y(g27986),.A(I36459));
  NOT NOT1_11237(.VSS(VSS),.VDD(VDD),.Y(I36462),.A(g27259));
  NOT NOT1_11238(.VSS(VSS),.VDD(VDD),.Y(g27987),.A(I36462));
  NOT NOT1_11239(.VSS(VSS),.VDD(VDD),.Y(I36465),.A(g27260));
  NOT NOT1_11240(.VSS(VSS),.VDD(VDD),.Y(g27988),.A(I36465));
  NOT NOT1_11241(.VSS(VSS),.VDD(VDD),.Y(I36468),.A(g27261));
  NOT NOT1_11242(.VSS(VSS),.VDD(VDD),.Y(g27989),.A(I36468));
  NOT NOT1_11243(.VSS(VSS),.VDD(VDD),.Y(g27990),.A(g27367));
  NOT NOT1_11244(.VSS(VSS),.VDD(VDD),.Y(I36473),.A(g27262));
  NOT NOT1_11245(.VSS(VSS),.VDD(VDD),.Y(g27992),.A(I36473));
  NOT NOT1_11246(.VSS(VSS),.VDD(VDD),.Y(I36476),.A(g27263));
  NOT NOT1_11247(.VSS(VSS),.VDD(VDD),.Y(g27993),.A(I36476));
  NOT NOT1_11248(.VSS(VSS),.VDD(VDD),.Y(I36479),.A(g27504));
  NOT NOT1_11249(.VSS(VSS),.VDD(VDD),.Y(g27994),.A(I36479));
  NOT NOT1_11250(.VSS(VSS),.VDD(VDD),.Y(I36483),.A(g27264));
  NOT NOT1_11251(.VSS(VSS),.VDD(VDD),.Y(g27998),.A(I36483));
  NOT NOT1_11252(.VSS(VSS),.VDD(VDD),.Y(I36486),.A(g27507));
  NOT NOT1_11253(.VSS(VSS),.VDD(VDD),.Y(g27999),.A(I36486));
  NOT NOT1_11254(.VSS(VSS),.VDD(VDD),.Y(I36490),.A(g27265));
  NOT NOT1_11255(.VSS(VSS),.VDD(VDD),.Y(g28003),.A(I36490));
  NOT NOT1_11256(.VSS(VSS),.VDD(VDD),.Y(I36493),.A(g27266));
  NOT NOT1_11257(.VSS(VSS),.VDD(VDD),.Y(g28004),.A(I36493));
  NOT NOT1_11258(.VSS(VSS),.VDD(VDD),.Y(I36496),.A(g27267));
  NOT NOT1_11259(.VSS(VSS),.VDD(VDD),.Y(g28005),.A(I36496));
  NOT NOT1_11260(.VSS(VSS),.VDD(VDD),.Y(I36499),.A(g27268));
  NOT NOT1_11261(.VSS(VSS),.VDD(VDD),.Y(g28006),.A(I36499));
  NOT NOT1_11262(.VSS(VSS),.VDD(VDD),.Y(I36502),.A(g27269));
  NOT NOT1_11263(.VSS(VSS),.VDD(VDD),.Y(g28007),.A(I36502));
  NOT NOT1_11264(.VSS(VSS),.VDD(VDD),.Y(I36507),.A(g27270));
  NOT NOT1_11265(.VSS(VSS),.VDD(VDD),.Y(g28010),.A(I36507));
  NOT NOT1_11266(.VSS(VSS),.VDD(VDD),.Y(I36510),.A(g27271));
  NOT NOT1_11267(.VSS(VSS),.VDD(VDD),.Y(g28011),.A(I36510));
  NOT NOT1_11268(.VSS(VSS),.VDD(VDD),.Y(I36513),.A(g27272));
  NOT NOT1_11269(.VSS(VSS),.VDD(VDD),.Y(g28012),.A(I36513));
  NOT NOT1_11270(.VSS(VSS),.VDD(VDD),.Y(I36516),.A(g27273));
  NOT NOT1_11271(.VSS(VSS),.VDD(VDD),.Y(g28013),.A(I36516));
  NOT NOT1_11272(.VSS(VSS),.VDD(VDD),.Y(g28014),.A(g27373));
  NOT NOT1_11273(.VSS(VSS),.VDD(VDD),.Y(I36521),.A(g27274));
  NOT NOT1_11274(.VSS(VSS),.VDD(VDD),.Y(g28016),.A(I36521));
  NOT NOT1_11275(.VSS(VSS),.VDD(VDD),.Y(I36524),.A(g27275));
  NOT NOT1_11276(.VSS(VSS),.VDD(VDD),.Y(g28017),.A(I36524));
  NOT NOT1_11277(.VSS(VSS),.VDD(VDD),.Y(I36527),.A(g27524));
  NOT NOT1_11278(.VSS(VSS),.VDD(VDD),.Y(g28018),.A(I36527));
  NOT NOT1_11279(.VSS(VSS),.VDD(VDD),.Y(I36530),.A(g27276));
  NOT NOT1_11280(.VSS(VSS),.VDD(VDD),.Y(g28021),.A(I36530));
  NOT NOT1_11281(.VSS(VSS),.VDD(VDD),.Y(I36533),.A(g27277));
  NOT NOT1_11282(.VSS(VSS),.VDD(VDD),.Y(g28022),.A(I36533));
  NOT NOT1_11283(.VSS(VSS),.VDD(VDD),.Y(I36536),.A(g27278));
  NOT NOT1_11284(.VSS(VSS),.VDD(VDD),.Y(g28023),.A(I36536));
  NOT NOT1_11285(.VSS(VSS),.VDD(VDD),.Y(I36539),.A(g27279));
  NOT NOT1_11286(.VSS(VSS),.VDD(VDD),.Y(g28024),.A(I36539));
  NOT NOT1_11287(.VSS(VSS),.VDD(VDD),.Y(I36542),.A(g27280));
  NOT NOT1_11288(.VSS(VSS),.VDD(VDD),.Y(g28025),.A(I36542));
  NOT NOT1_11289(.VSS(VSS),.VDD(VDD),.Y(I36545),.A(g27281));
  NOT NOT1_11290(.VSS(VSS),.VDD(VDD),.Y(g28026),.A(I36545));
  NOT NOT1_11291(.VSS(VSS),.VDD(VDD),.Y(I36551),.A(g27282));
  NOT NOT1_11292(.VSS(VSS),.VDD(VDD),.Y(g28030),.A(I36551));
  NOT NOT1_11293(.VSS(VSS),.VDD(VDD),.Y(I36554),.A(g27283));
  NOT NOT1_11294(.VSS(VSS),.VDD(VDD),.Y(g28031),.A(I36554));
  NOT NOT1_11295(.VSS(VSS),.VDD(VDD),.Y(I36557),.A(g27284));
  NOT NOT1_11296(.VSS(VSS),.VDD(VDD),.Y(g28032),.A(I36557));
  NOT NOT1_11297(.VSS(VSS),.VDD(VDD),.Y(I36560),.A(g27285));
  NOT NOT1_11298(.VSS(VSS),.VDD(VDD),.Y(g28033),.A(I36560));
  NOT NOT1_11299(.VSS(VSS),.VDD(VDD),.Y(I36563),.A(g27286));
  NOT NOT1_11300(.VSS(VSS),.VDD(VDD),.Y(g28034),.A(I36563));
  NOT NOT1_11301(.VSS(VSS),.VDD(VDD),.Y(I36568),.A(g27287));
  NOT NOT1_11302(.VSS(VSS),.VDD(VDD),.Y(g28037),.A(I36568));
  NOT NOT1_11303(.VSS(VSS),.VDD(VDD),.Y(I36571),.A(g27288));
  NOT NOT1_11304(.VSS(VSS),.VDD(VDD),.Y(g28038),.A(I36571));
  NOT NOT1_11305(.VSS(VSS),.VDD(VDD),.Y(I36574),.A(g27289));
  NOT NOT1_11306(.VSS(VSS),.VDD(VDD),.Y(g28039),.A(I36574));
  NOT NOT1_11307(.VSS(VSS),.VDD(VDD),.Y(I36577),.A(g27290));
  NOT NOT1_11308(.VSS(VSS),.VDD(VDD),.Y(g28040),.A(I36577));
  NOT NOT1_11309(.VSS(VSS),.VDD(VDD),.Y(g28041),.A(g27376));
  NOT NOT1_11310(.VSS(VSS),.VDD(VDD),.Y(I36582),.A(g27291));
  NOT NOT1_11311(.VSS(VSS),.VDD(VDD),.Y(g28043),.A(I36582));
  NOT NOT1_11312(.VSS(VSS),.VDD(VDD),.Y(I36585),.A(g27292));
  NOT NOT1_11313(.VSS(VSS),.VDD(VDD),.Y(g28044),.A(I36585));
  NOT NOT1_11314(.VSS(VSS),.VDD(VDD),.Y(I36588),.A(g27293));
  NOT NOT1_11315(.VSS(VSS),.VDD(VDD),.Y(g28045),.A(I36588));
  NOT NOT1_11316(.VSS(VSS),.VDD(VDD),.Y(I36598),.A(g27294));
  NOT NOT1_11317(.VSS(VSS),.VDD(VDD),.Y(g28047),.A(I36598));
  NOT NOT1_11318(.VSS(VSS),.VDD(VDD),.Y(I36601),.A(g27295));
  NOT NOT1_11319(.VSS(VSS),.VDD(VDD),.Y(g28048),.A(I36601));
  NOT NOT1_11320(.VSS(VSS),.VDD(VDD),.Y(I36604),.A(g27296));
  NOT NOT1_11321(.VSS(VSS),.VDD(VDD),.Y(g28049),.A(I36604));
  NOT NOT1_11322(.VSS(VSS),.VDD(VDD),.Y(I36609),.A(g27297));
  NOT NOT1_11323(.VSS(VSS),.VDD(VDD),.Y(g28052),.A(I36609));
  NOT NOT1_11324(.VSS(VSS),.VDD(VDD),.Y(I36612),.A(g27298));
  NOT NOT1_11325(.VSS(VSS),.VDD(VDD),.Y(g28053),.A(I36612));
  NOT NOT1_11326(.VSS(VSS),.VDD(VDD),.Y(I36615),.A(g27299));
  NOT NOT1_11327(.VSS(VSS),.VDD(VDD),.Y(g28054),.A(I36615));
  NOT NOT1_11328(.VSS(VSS),.VDD(VDD),.Y(I36618),.A(g27300));
  NOT NOT1_11329(.VSS(VSS),.VDD(VDD),.Y(g28055),.A(I36618));
  NOT NOT1_11330(.VSS(VSS),.VDD(VDD),.Y(I36621),.A(g27301));
  NOT NOT1_11331(.VSS(VSS),.VDD(VDD),.Y(g28056),.A(I36621));
  NOT NOT1_11332(.VSS(VSS),.VDD(VDD),.Y(I36627),.A(g27302));
  NOT NOT1_11333(.VSS(VSS),.VDD(VDD),.Y(g28060),.A(I36627));
  NOT NOT1_11334(.VSS(VSS),.VDD(VDD),.Y(I36630),.A(g27303));
  NOT NOT1_11335(.VSS(VSS),.VDD(VDD),.Y(g28061),.A(I36630));
  NOT NOT1_11336(.VSS(VSS),.VDD(VDD),.Y(I36633),.A(g27304));
  NOT NOT1_11337(.VSS(VSS),.VDD(VDD),.Y(g28062),.A(I36633));
  NOT NOT1_11338(.VSS(VSS),.VDD(VDD),.Y(I36636),.A(g27305));
  NOT NOT1_11339(.VSS(VSS),.VDD(VDD),.Y(g28063),.A(I36636));
  NOT NOT1_11340(.VSS(VSS),.VDD(VDD),.Y(I36639),.A(g27306));
  NOT NOT1_11341(.VSS(VSS),.VDD(VDD),.Y(g28064),.A(I36639));
  NOT NOT1_11342(.VSS(VSS),.VDD(VDD),.Y(I36644),.A(g27307));
  NOT NOT1_11343(.VSS(VSS),.VDD(VDD),.Y(g28067),.A(I36644));
  NOT NOT1_11344(.VSS(VSS),.VDD(VDD),.Y(I36647),.A(g27308));
  NOT NOT1_11345(.VSS(VSS),.VDD(VDD),.Y(g28068),.A(I36647));
  NOT NOT1_11346(.VSS(VSS),.VDD(VDD),.Y(I36650),.A(g27309));
  NOT NOT1_11347(.VSS(VSS),.VDD(VDD),.Y(g28069),.A(I36650));
  NOT NOT1_11348(.VSS(VSS),.VDD(VDD),.Y(I36653),.A(g27310));
  NOT NOT1_11349(.VSS(VSS),.VDD(VDD),.Y(g28070),.A(I36653));
  NOT NOT1_11350(.VSS(VSS),.VDD(VDD),.Y(I36656),.A(g27311));
  NOT NOT1_11351(.VSS(VSS),.VDD(VDD),.Y(g28071),.A(I36656));
  NOT NOT1_11352(.VSS(VSS),.VDD(VDD),.Y(I36659),.A(g27312));
  NOT NOT1_11353(.VSS(VSS),.VDD(VDD),.Y(g28072),.A(I36659));
  NOT NOT1_11354(.VSS(VSS),.VDD(VDD),.Y(I36663),.A(g27313));
  NOT NOT1_11355(.VSS(VSS),.VDD(VDD),.Y(g28074),.A(I36663));
  NOT NOT1_11356(.VSS(VSS),.VDD(VDD),.Y(I36673),.A(g27314));
  NOT NOT1_11357(.VSS(VSS),.VDD(VDD),.Y(g28076),.A(I36673));
  NOT NOT1_11358(.VSS(VSS),.VDD(VDD),.Y(I36676),.A(g27315));
  NOT NOT1_11359(.VSS(VSS),.VDD(VDD),.Y(g28077),.A(I36676));
  NOT NOT1_11360(.VSS(VSS),.VDD(VDD),.Y(I36679),.A(g27316));
  NOT NOT1_11361(.VSS(VSS),.VDD(VDD),.Y(g28078),.A(I36679));
  NOT NOT1_11362(.VSS(VSS),.VDD(VDD),.Y(I36684),.A(g27317));
  NOT NOT1_11363(.VSS(VSS),.VDD(VDD),.Y(g28081),.A(I36684));
  NOT NOT1_11364(.VSS(VSS),.VDD(VDD),.Y(I36687),.A(g27318));
  NOT NOT1_11365(.VSS(VSS),.VDD(VDD),.Y(g28082),.A(I36687));
  NOT NOT1_11366(.VSS(VSS),.VDD(VDD),.Y(I36690),.A(g27319));
  NOT NOT1_11367(.VSS(VSS),.VDD(VDD),.Y(g28083),.A(I36690));
  NOT NOT1_11368(.VSS(VSS),.VDD(VDD),.Y(I36693),.A(g27320));
  NOT NOT1_11369(.VSS(VSS),.VDD(VDD),.Y(g28084),.A(I36693));
  NOT NOT1_11370(.VSS(VSS),.VDD(VDD),.Y(I36696),.A(g27321));
  NOT NOT1_11371(.VSS(VSS),.VDD(VDD),.Y(g28085),.A(I36696));
  NOT NOT1_11372(.VSS(VSS),.VDD(VDD),.Y(I36702),.A(g27322));
  NOT NOT1_11373(.VSS(VSS),.VDD(VDD),.Y(g28089),.A(I36702));
  NOT NOT1_11374(.VSS(VSS),.VDD(VDD),.Y(I36705),.A(g27323));
  NOT NOT1_11375(.VSS(VSS),.VDD(VDD),.Y(g28090),.A(I36705));
  NOT NOT1_11376(.VSS(VSS),.VDD(VDD),.Y(I36708),.A(g27324));
  NOT NOT1_11377(.VSS(VSS),.VDD(VDD),.Y(g28091),.A(I36708));
  NOT NOT1_11378(.VSS(VSS),.VDD(VDD),.Y(I36711),.A(g27325));
  NOT NOT1_11379(.VSS(VSS),.VDD(VDD),.Y(g28092),.A(I36711));
  NOT NOT1_11380(.VSS(VSS),.VDD(VDD),.Y(I36714),.A(g27326));
  NOT NOT1_11381(.VSS(VSS),.VDD(VDD),.Y(g28093),.A(I36714));
  NOT NOT1_11382(.VSS(VSS),.VDD(VDD),.Y(I36718),.A(g27327));
  NOT NOT1_11383(.VSS(VSS),.VDD(VDD),.Y(g28095),.A(I36718));
  NOT NOT1_11384(.VSS(VSS),.VDD(VDD),.Y(I36721),.A(g27328));
  NOT NOT1_11385(.VSS(VSS),.VDD(VDD),.Y(g28096),.A(I36721));
  NOT NOT1_11386(.VSS(VSS),.VDD(VDD),.Y(I36724),.A(g27329));
  NOT NOT1_11387(.VSS(VSS),.VDD(VDD),.Y(g28097),.A(I36724));
  NOT NOT1_11388(.VSS(VSS),.VDD(VDD),.Y(I36728),.A(g27330));
  NOT NOT1_11389(.VSS(VSS),.VDD(VDD),.Y(g28099),.A(I36728));
  NOT NOT1_11390(.VSS(VSS),.VDD(VDD),.Y(I36738),.A(g27331));
  NOT NOT1_11391(.VSS(VSS),.VDD(VDD),.Y(g28101),.A(I36738));
  NOT NOT1_11392(.VSS(VSS),.VDD(VDD),.Y(I36741),.A(g27332));
  NOT NOT1_11393(.VSS(VSS),.VDD(VDD),.Y(g28102),.A(I36741));
  NOT NOT1_11394(.VSS(VSS),.VDD(VDD),.Y(I36744),.A(g27333));
  NOT NOT1_11395(.VSS(VSS),.VDD(VDD),.Y(g28103),.A(I36744));
  NOT NOT1_11396(.VSS(VSS),.VDD(VDD),.Y(I36749),.A(g27334));
  NOT NOT1_11397(.VSS(VSS),.VDD(VDD),.Y(g28106),.A(I36749));
  NOT NOT1_11398(.VSS(VSS),.VDD(VDD),.Y(I36752),.A(g27335));
  NOT NOT1_11399(.VSS(VSS),.VDD(VDD),.Y(g28107),.A(I36752));
  NOT NOT1_11400(.VSS(VSS),.VDD(VDD),.Y(I36755),.A(g27336));
  NOT NOT1_11401(.VSS(VSS),.VDD(VDD),.Y(g28108),.A(I36755));
  NOT NOT1_11402(.VSS(VSS),.VDD(VDD),.Y(I36758),.A(g27337));
  NOT NOT1_11403(.VSS(VSS),.VDD(VDD),.Y(g28109),.A(I36758));
  NOT NOT1_11404(.VSS(VSS),.VDD(VDD),.Y(I36761),.A(g27338));
  NOT NOT1_11405(.VSS(VSS),.VDD(VDD),.Y(g28110),.A(I36761));
  NOT NOT1_11406(.VSS(VSS),.VDD(VDD),.Y(I36766),.A(g27339));
  NOT NOT1_11407(.VSS(VSS),.VDD(VDD),.Y(g28113),.A(I36766));
  NOT NOT1_11408(.VSS(VSS),.VDD(VDD),.Y(I36769),.A(g27340));
  NOT NOT1_11409(.VSS(VSS),.VDD(VDD),.Y(g28114),.A(I36769));
  NOT NOT1_11410(.VSS(VSS),.VDD(VDD),.Y(I36772),.A(g27341));
  NOT NOT1_11411(.VSS(VSS),.VDD(VDD),.Y(g28115),.A(I36772));
  NOT NOT1_11412(.VSS(VSS),.VDD(VDD),.Y(I36776),.A(g27342));
  NOT NOT1_11413(.VSS(VSS),.VDD(VDD),.Y(g28117),.A(I36776));
  NOT NOT1_11414(.VSS(VSS),.VDD(VDD),.Y(I36786),.A(g27343));
  NOT NOT1_11415(.VSS(VSS),.VDD(VDD),.Y(g28119),.A(I36786));
  NOT NOT1_11416(.VSS(VSS),.VDD(VDD),.Y(I36789),.A(g27344));
  NOT NOT1_11417(.VSS(VSS),.VDD(VDD),.Y(g28120),.A(I36789));
  NOT NOT1_11418(.VSS(VSS),.VDD(VDD),.Y(I36792),.A(g27345));
  NOT NOT1_11419(.VSS(VSS),.VDD(VDD),.Y(g28121),.A(I36792));
  NOT NOT1_11420(.VSS(VSS),.VDD(VDD),.Y(I36797),.A(g27346));
  NOT NOT1_11421(.VSS(VSS),.VDD(VDD),.Y(g28124),.A(I36797));
  NOT NOT1_11422(.VSS(VSS),.VDD(VDD),.Y(I36800),.A(g27347));
  NOT NOT1_11423(.VSS(VSS),.VDD(VDD),.Y(g28125),.A(I36800));
  NOT NOT1_11424(.VSS(VSS),.VDD(VDD),.Y(I36803),.A(g27348));
  NOT NOT1_11425(.VSS(VSS),.VDD(VDD),.Y(g28126),.A(I36803));
  NOT NOT1_11426(.VSS(VSS),.VDD(VDD),.Y(g28128),.A(g27528));
  NOT NOT1_11427(.VSS(VSS),.VDD(VDD),.Y(I36808),.A(g27354));
  NOT NOT1_11428(.VSS(VSS),.VDD(VDD),.Y(g28132),.A(I36808));
  NOT NOT1_11429(.VSS(VSS),.VDD(VDD),.Y(g28133),.A(g27550));
  NOT NOT1_11430(.VSS(VSS),.VDD(VDD),.Y(g28137),.A(g27566));
  NOT NOT1_11431(.VSS(VSS),.VDD(VDD),.Y(g28141),.A(g27576));
  NOT NOT1_11432(.VSS(VSS),.VDD(VDD),.Y(g28149),.A(g27667));
  NOT NOT1_11433(.VSS(VSS),.VDD(VDD),.Y(g28150),.A(g27387));
  NOT NOT1_11434(.VSS(VSS),.VDD(VDD),.Y(g28151),.A(g27381));
  NOT NOT1_11435(.VSS(VSS),.VDD(VDD),.Y(g28152),.A(g27391));
  NOT NOT1_11436(.VSS(VSS),.VDD(VDD),.Y(g28153),.A(g27397));
  NOT NOT1_11437(.VSS(VSS),.VDD(VDD),.Y(g28154),.A(g27401));
  NOT NOT1_11438(.VSS(VSS),.VDD(VDD),.Y(g28155),.A(g27404));
  NOT NOT1_11439(.VSS(VSS),.VDD(VDD),.Y(g28156),.A(g27410));
  NOT NOT1_11440(.VSS(VSS),.VDD(VDD),.Y(g28158),.A(g27416));
  NOT NOT1_11441(.VSS(VSS),.VDD(VDD),.Y(g28159),.A(g27419));
  NOT NOT1_11442(.VSS(VSS),.VDD(VDD),.Y(g28160),.A(g27422));
  NOT NOT1_11443(.VSS(VSS),.VDD(VDD),.Y(g28161),.A(g27428));
  NOT NOT1_11444(.VSS(VSS),.VDD(VDD),.Y(g28162),.A(g27432));
  NOT NOT1_11445(.VSS(VSS),.VDD(VDD),.Y(g28163),.A(g27437));
  NOT NOT1_11446(.VSS(VSS),.VDD(VDD),.Y(g28164),.A(g27440));
  NOT NOT1_11447(.VSS(VSS),.VDD(VDD),.Y(g28165),.A(g27443));
  NOT NOT1_11448(.VSS(VSS),.VDD(VDD),.Y(g28166),.A(g27451));
  NOT NOT1_11449(.VSS(VSS),.VDD(VDD),.Y(g28167),.A(g27456));
  NOT NOT1_11450(.VSS(VSS),.VDD(VDD),.Y(g28168),.A(g27459));
  NOT NOT1_11451(.VSS(VSS),.VDD(VDD),.Y(g28169),.A(g27467));
  NOT NOT1_11452(.VSS(VSS),.VDD(VDD),.Y(g28170),.A(g27472));
  NOT NOT1_11453(.VSS(VSS),.VDD(VDD),.Y(g28172),.A(g27475));
  NOT NOT1_11454(.VSS(VSS),.VDD(VDD),.Y(g28173),.A(g27486));
  NOT NOT1_11455(.VSS(VSS),.VDD(VDD),.Y(g28174),.A(g27489));
  NOT NOT1_11456(.VSS(VSS),.VDD(VDD),.Y(g28175),.A(g27498));
  NOT NOT1_11457(.VSS(VSS),.VDD(VDD),.Y(g28177),.A(g27510));
  NOT NOT1_11458(.VSS(VSS),.VDD(VDD),.Y(g28178),.A(g27518));
  NOT NOT1_11459(.VSS(VSS),.VDD(VDD),.Y(I36848),.A(g27383));
  NOT NOT1_11460(.VSS(VSS),.VDD(VDD),.Y(g28179),.A(I36848));
  NOT NOT1_11461(.VSS(VSS),.VDD(VDD),.Y(g28186),.A(g27535));
  NOT NOT1_11462(.VSS(VSS),.VDD(VDD),.Y(g28187),.A(g27543));
  NOT NOT1_11463(.VSS(VSS),.VDD(VDD),.Y(g28190),.A(g27555));
  NOT NOT1_11464(.VSS(VSS),.VDD(VDD),.Y(I36860),.A(g27386));
  NOT NOT1_11465(.VSS(VSS),.VDD(VDD),.Y(g28194),.A(I36860));
  NOT NOT1_11466(.VSS(VSS),.VDD(VDD),.Y(I36864),.A(g27384));
  NOT NOT1_11467(.VSS(VSS),.VDD(VDD),.Y(g28200),.A(I36864));
  NOT NOT1_11468(.VSS(VSS),.VDD(VDD),.Y(I36867),.A(g27786));
  NOT NOT1_11469(.VSS(VSS),.VDD(VDD),.Y(g28206),.A(I36867));
  NOT NOT1_11470(.VSS(VSS),.VDD(VDD),.Y(I36870),.A(g27955));
  NOT NOT1_11471(.VSS(VSS),.VDD(VDD),.Y(g28207),.A(I36870));
  NOT NOT1_11472(.VSS(VSS),.VDD(VDD),.Y(I36873),.A(g27971));
  NOT NOT1_11473(.VSS(VSS),.VDD(VDD),.Y(g28208),.A(I36873));
  NOT NOT1_11474(.VSS(VSS),.VDD(VDD),.Y(I36876),.A(g27986));
  NOT NOT1_11475(.VSS(VSS),.VDD(VDD),.Y(g28209),.A(I36876));
  NOT NOT1_11476(.VSS(VSS),.VDD(VDD),.Y(I36879),.A(g27972));
  NOT NOT1_11477(.VSS(VSS),.VDD(VDD),.Y(g28210),.A(I36879));
  NOT NOT1_11478(.VSS(VSS),.VDD(VDD),.Y(I36882),.A(g27987));
  NOT NOT1_11479(.VSS(VSS),.VDD(VDD),.Y(g28211),.A(I36882));
  NOT NOT1_11480(.VSS(VSS),.VDD(VDD),.Y(I36885),.A(g28003));
  NOT NOT1_11481(.VSS(VSS),.VDD(VDD),.Y(g28212),.A(I36885));
  NOT NOT1_11482(.VSS(VSS),.VDD(VDD),.Y(I36888),.A(g27988));
  NOT NOT1_11483(.VSS(VSS),.VDD(VDD),.Y(g28213),.A(I36888));
  NOT NOT1_11484(.VSS(VSS),.VDD(VDD),.Y(I36891),.A(g28004));
  NOT NOT1_11485(.VSS(VSS),.VDD(VDD),.Y(g28214),.A(I36891));
  NOT NOT1_11486(.VSS(VSS),.VDD(VDD),.Y(I36894),.A(g28022));
  NOT NOT1_11487(.VSS(VSS),.VDD(VDD),.Y(g28215),.A(I36894));
  NOT NOT1_11488(.VSS(VSS),.VDD(VDD),.Y(I36897),.A(g28005));
  NOT NOT1_11489(.VSS(VSS),.VDD(VDD),.Y(g28216),.A(I36897));
  NOT NOT1_11490(.VSS(VSS),.VDD(VDD),.Y(I36900),.A(g28023));
  NOT NOT1_11491(.VSS(VSS),.VDD(VDD),.Y(g28217),.A(I36900));
  NOT NOT1_11492(.VSS(VSS),.VDD(VDD),.Y(I36903),.A(g28045));
  NOT NOT1_11493(.VSS(VSS),.VDD(VDD),.Y(g28218),.A(I36903));
  NOT NOT1_11494(.VSS(VSS),.VDD(VDD),.Y(I36906),.A(g27989));
  NOT NOT1_11495(.VSS(VSS),.VDD(VDD),.Y(g28219),.A(I36906));
  NOT NOT1_11496(.VSS(VSS),.VDD(VDD),.Y(I36909),.A(g28006));
  NOT NOT1_11497(.VSS(VSS),.VDD(VDD),.Y(g28220),.A(I36909));
  NOT NOT1_11498(.VSS(VSS),.VDD(VDD),.Y(I36912),.A(g28024));
  NOT NOT1_11499(.VSS(VSS),.VDD(VDD),.Y(g28221),.A(I36912));
  NOT NOT1_11500(.VSS(VSS),.VDD(VDD),.Y(I36915),.A(g28007));
  NOT NOT1_11501(.VSS(VSS),.VDD(VDD),.Y(g28222),.A(I36915));
  NOT NOT1_11502(.VSS(VSS),.VDD(VDD),.Y(I36918),.A(g28025));
  NOT NOT1_11503(.VSS(VSS),.VDD(VDD),.Y(g28223),.A(I36918));
  NOT NOT1_11504(.VSS(VSS),.VDD(VDD),.Y(I36921),.A(g28047));
  NOT NOT1_11505(.VSS(VSS),.VDD(VDD),.Y(g28224),.A(I36921));
  NOT NOT1_11506(.VSS(VSS),.VDD(VDD),.Y(I36924),.A(g28026));
  NOT NOT1_11507(.VSS(VSS),.VDD(VDD),.Y(g28225),.A(I36924));
  NOT NOT1_11508(.VSS(VSS),.VDD(VDD),.Y(I36927),.A(g28048));
  NOT NOT1_11509(.VSS(VSS),.VDD(VDD),.Y(g28226),.A(I36927));
  NOT NOT1_11510(.VSS(VSS),.VDD(VDD),.Y(I36930),.A(g28071));
  NOT NOT1_11511(.VSS(VSS),.VDD(VDD),.Y(g28227),.A(I36930));
  NOT NOT1_11512(.VSS(VSS),.VDD(VDD),.Y(I36933),.A(g28049));
  NOT NOT1_11513(.VSS(VSS),.VDD(VDD),.Y(g28228),.A(I36933));
  NOT NOT1_11514(.VSS(VSS),.VDD(VDD),.Y(I36936),.A(g28072));
  NOT NOT1_11515(.VSS(VSS),.VDD(VDD),.Y(g28229),.A(I36936));
  NOT NOT1_11516(.VSS(VSS),.VDD(VDD),.Y(I36939),.A(g28095));
  NOT NOT1_11517(.VSS(VSS),.VDD(VDD),.Y(g28230),.A(I36939));
  NOT NOT1_11518(.VSS(VSS),.VDD(VDD),.Y(I36942),.A(g27905));
  NOT NOT1_11519(.VSS(VSS),.VDD(VDD),.Y(g28231),.A(I36942));
  NOT NOT1_11520(.VSS(VSS),.VDD(VDD),.Y(I36945),.A(g27793));
  NOT NOT1_11521(.VSS(VSS),.VDD(VDD),.Y(g28232),.A(I36945));
  NOT NOT1_11522(.VSS(VSS),.VDD(VDD),.Y(I36948),.A(g27976));
  NOT NOT1_11523(.VSS(VSS),.VDD(VDD),.Y(g28233),.A(I36948));
  NOT NOT1_11524(.VSS(VSS),.VDD(VDD),.Y(I36951),.A(g27992));
  NOT NOT1_11525(.VSS(VSS),.VDD(VDD),.Y(g28234),.A(I36951));
  NOT NOT1_11526(.VSS(VSS),.VDD(VDD),.Y(I36954),.A(g28010));
  NOT NOT1_11527(.VSS(VSS),.VDD(VDD),.Y(g28235),.A(I36954));
  NOT NOT1_11528(.VSS(VSS),.VDD(VDD),.Y(I36957),.A(g27993));
  NOT NOT1_11529(.VSS(VSS),.VDD(VDD),.Y(g28236),.A(I36957));
  NOT NOT1_11530(.VSS(VSS),.VDD(VDD),.Y(I36960),.A(g28011));
  NOT NOT1_11531(.VSS(VSS),.VDD(VDD),.Y(g28237),.A(I36960));
  NOT NOT1_11532(.VSS(VSS),.VDD(VDD),.Y(I36963),.A(g28030));
  NOT NOT1_11533(.VSS(VSS),.VDD(VDD),.Y(g28238),.A(I36963));
  NOT NOT1_11534(.VSS(VSS),.VDD(VDD),.Y(I36966),.A(g28012));
  NOT NOT1_11535(.VSS(VSS),.VDD(VDD),.Y(g28239),.A(I36966));
  NOT NOT1_11536(.VSS(VSS),.VDD(VDD),.Y(I36969),.A(g28031));
  NOT NOT1_11537(.VSS(VSS),.VDD(VDD),.Y(g28240),.A(I36969));
  NOT NOT1_11538(.VSS(VSS),.VDD(VDD),.Y(I36972),.A(g28052));
  NOT NOT1_11539(.VSS(VSS),.VDD(VDD),.Y(g28241),.A(I36972));
  NOT NOT1_11540(.VSS(VSS),.VDD(VDD),.Y(I36975),.A(g28032));
  NOT NOT1_11541(.VSS(VSS),.VDD(VDD),.Y(g28242),.A(I36975));
  NOT NOT1_11542(.VSS(VSS),.VDD(VDD),.Y(I36978),.A(g28053));
  NOT NOT1_11543(.VSS(VSS),.VDD(VDD),.Y(g28243),.A(I36978));
  NOT NOT1_11544(.VSS(VSS),.VDD(VDD),.Y(I36981),.A(g28074));
  NOT NOT1_11545(.VSS(VSS),.VDD(VDD),.Y(g28244),.A(I36981));
  NOT NOT1_11546(.VSS(VSS),.VDD(VDD),.Y(I36984),.A(g28013));
  NOT NOT1_11547(.VSS(VSS),.VDD(VDD),.Y(g28245),.A(I36984));
  NOT NOT1_11548(.VSS(VSS),.VDD(VDD),.Y(I36987),.A(g28033));
  NOT NOT1_11549(.VSS(VSS),.VDD(VDD),.Y(g28246),.A(I36987));
  NOT NOT1_11550(.VSS(VSS),.VDD(VDD),.Y(I36990),.A(g28054));
  NOT NOT1_11551(.VSS(VSS),.VDD(VDD),.Y(g28247),.A(I36990));
  NOT NOT1_11552(.VSS(VSS),.VDD(VDD),.Y(I36993),.A(g28034));
  NOT NOT1_11553(.VSS(VSS),.VDD(VDD),.Y(g28248),.A(I36993));
  NOT NOT1_11554(.VSS(VSS),.VDD(VDD),.Y(I36996),.A(g28055));
  NOT NOT1_11555(.VSS(VSS),.VDD(VDD),.Y(g28249),.A(I36996));
  NOT NOT1_11556(.VSS(VSS),.VDD(VDD),.Y(I36999),.A(g28076));
  NOT NOT1_11557(.VSS(VSS),.VDD(VDD),.Y(g28250),.A(I36999));
  NOT NOT1_11558(.VSS(VSS),.VDD(VDD),.Y(I37002),.A(g28056));
  NOT NOT1_11559(.VSS(VSS),.VDD(VDD),.Y(g28251),.A(I37002));
  NOT NOT1_11560(.VSS(VSS),.VDD(VDD),.Y(I37005),.A(g28077));
  NOT NOT1_11561(.VSS(VSS),.VDD(VDD),.Y(g28252),.A(I37005));
  NOT NOT1_11562(.VSS(VSS),.VDD(VDD),.Y(I37008),.A(g28096));
  NOT NOT1_11563(.VSS(VSS),.VDD(VDD),.Y(g28253),.A(I37008));
  NOT NOT1_11564(.VSS(VSS),.VDD(VDD),.Y(I37011),.A(g28078));
  NOT NOT1_11565(.VSS(VSS),.VDD(VDD),.Y(g28254),.A(I37011));
  NOT NOT1_11566(.VSS(VSS),.VDD(VDD),.Y(I37014),.A(g28097));
  NOT NOT1_11567(.VSS(VSS),.VDD(VDD),.Y(g28255),.A(I37014));
  NOT NOT1_11568(.VSS(VSS),.VDD(VDD),.Y(I37017),.A(g28113));
  NOT NOT1_11569(.VSS(VSS),.VDD(VDD),.Y(g28256),.A(I37017));
  NOT NOT1_11570(.VSS(VSS),.VDD(VDD),.Y(I37020),.A(g27910));
  NOT NOT1_11571(.VSS(VSS),.VDD(VDD),.Y(g28257),.A(I37020));
  NOT NOT1_11572(.VSS(VSS),.VDD(VDD),.Y(I37023),.A(g27799));
  NOT NOT1_11573(.VSS(VSS),.VDD(VDD),.Y(g28258),.A(I37023));
  NOT NOT1_11574(.VSS(VSS),.VDD(VDD),.Y(I37026),.A(g27998));
  NOT NOT1_11575(.VSS(VSS),.VDD(VDD),.Y(g28259),.A(I37026));
  NOT NOT1_11576(.VSS(VSS),.VDD(VDD),.Y(I37029),.A(g28016));
  NOT NOT1_11577(.VSS(VSS),.VDD(VDD),.Y(g28260),.A(I37029));
  NOT NOT1_11578(.VSS(VSS),.VDD(VDD),.Y(I37032),.A(g28037));
  NOT NOT1_11579(.VSS(VSS),.VDD(VDD),.Y(g28261),.A(I37032));
  NOT NOT1_11580(.VSS(VSS),.VDD(VDD),.Y(I37035),.A(g28017));
  NOT NOT1_11581(.VSS(VSS),.VDD(VDD),.Y(g28262),.A(I37035));
  NOT NOT1_11582(.VSS(VSS),.VDD(VDD),.Y(I37038),.A(g28038));
  NOT NOT1_11583(.VSS(VSS),.VDD(VDD),.Y(g28263),.A(I37038));
  NOT NOT1_11584(.VSS(VSS),.VDD(VDD),.Y(I37041),.A(g28060));
  NOT NOT1_11585(.VSS(VSS),.VDD(VDD),.Y(g28264),.A(I37041));
  NOT NOT1_11586(.VSS(VSS),.VDD(VDD),.Y(I37044),.A(g28039));
  NOT NOT1_11587(.VSS(VSS),.VDD(VDD),.Y(g28265),.A(I37044));
  NOT NOT1_11588(.VSS(VSS),.VDD(VDD),.Y(I37047),.A(g28061));
  NOT NOT1_11589(.VSS(VSS),.VDD(VDD),.Y(g28266),.A(I37047));
  NOT NOT1_11590(.VSS(VSS),.VDD(VDD),.Y(I37050),.A(g28081));
  NOT NOT1_11591(.VSS(VSS),.VDD(VDD),.Y(g28267),.A(I37050));
  NOT NOT1_11592(.VSS(VSS),.VDD(VDD),.Y(I37053),.A(g28062));
  NOT NOT1_11593(.VSS(VSS),.VDD(VDD),.Y(g28268),.A(I37053));
  NOT NOT1_11594(.VSS(VSS),.VDD(VDD),.Y(I37056),.A(g28082));
  NOT NOT1_11595(.VSS(VSS),.VDD(VDD),.Y(g28269),.A(I37056));
  NOT NOT1_11596(.VSS(VSS),.VDD(VDD),.Y(I37059),.A(g28099));
  NOT NOT1_11597(.VSS(VSS),.VDD(VDD),.Y(g28270),.A(I37059));
  NOT NOT1_11598(.VSS(VSS),.VDD(VDD),.Y(I37062),.A(g28040));
  NOT NOT1_11599(.VSS(VSS),.VDD(VDD),.Y(g28271),.A(I37062));
  NOT NOT1_11600(.VSS(VSS),.VDD(VDD),.Y(I37065),.A(g28063));
  NOT NOT1_11601(.VSS(VSS),.VDD(VDD),.Y(g28272),.A(I37065));
  NOT NOT1_11602(.VSS(VSS),.VDD(VDD),.Y(I37068),.A(g28083));
  NOT NOT1_11603(.VSS(VSS),.VDD(VDD),.Y(g28273),.A(I37068));
  NOT NOT1_11604(.VSS(VSS),.VDD(VDD),.Y(I37071),.A(g28064));
  NOT NOT1_11605(.VSS(VSS),.VDD(VDD),.Y(g28274),.A(I37071));
  NOT NOT1_11606(.VSS(VSS),.VDD(VDD),.Y(I37074),.A(g28084));
  NOT NOT1_11607(.VSS(VSS),.VDD(VDD),.Y(g28275),.A(I37074));
  NOT NOT1_11608(.VSS(VSS),.VDD(VDD),.Y(I37077),.A(g28101));
  NOT NOT1_11609(.VSS(VSS),.VDD(VDD),.Y(g28276),.A(I37077));
  NOT NOT1_11610(.VSS(VSS),.VDD(VDD),.Y(I37080),.A(g28085));
  NOT NOT1_11611(.VSS(VSS),.VDD(VDD),.Y(g28277),.A(I37080));
  NOT NOT1_11612(.VSS(VSS),.VDD(VDD),.Y(I37083),.A(g28102));
  NOT NOT1_11613(.VSS(VSS),.VDD(VDD),.Y(g28278),.A(I37083));
  NOT NOT1_11614(.VSS(VSS),.VDD(VDD),.Y(I37086),.A(g28114));
  NOT NOT1_11615(.VSS(VSS),.VDD(VDD),.Y(g28279),.A(I37086));
  NOT NOT1_11616(.VSS(VSS),.VDD(VDD),.Y(I37089),.A(g28103));
  NOT NOT1_11617(.VSS(VSS),.VDD(VDD),.Y(g28280),.A(I37089));
  NOT NOT1_11618(.VSS(VSS),.VDD(VDD),.Y(I37092),.A(g28115));
  NOT NOT1_11619(.VSS(VSS),.VDD(VDD),.Y(g28281),.A(I37092));
  NOT NOT1_11620(.VSS(VSS),.VDD(VDD),.Y(I37095),.A(g28124));
  NOT NOT1_11621(.VSS(VSS),.VDD(VDD),.Y(g28282),.A(I37095));
  NOT NOT1_11622(.VSS(VSS),.VDD(VDD),.Y(I37098),.A(g27918));
  NOT NOT1_11623(.VSS(VSS),.VDD(VDD),.Y(g28283),.A(I37098));
  NOT NOT1_11624(.VSS(VSS),.VDD(VDD),.Y(I37101),.A(g27805));
  NOT NOT1_11625(.VSS(VSS),.VDD(VDD),.Y(g28284),.A(I37101));
  NOT NOT1_11626(.VSS(VSS),.VDD(VDD),.Y(I37104),.A(g28021));
  NOT NOT1_11627(.VSS(VSS),.VDD(VDD),.Y(g28285),.A(I37104));
  NOT NOT1_11628(.VSS(VSS),.VDD(VDD),.Y(I37107),.A(g28043));
  NOT NOT1_11629(.VSS(VSS),.VDD(VDD),.Y(g28286),.A(I37107));
  NOT NOT1_11630(.VSS(VSS),.VDD(VDD),.Y(I37110),.A(g28067));
  NOT NOT1_11631(.VSS(VSS),.VDD(VDD),.Y(g28287),.A(I37110));
  NOT NOT1_11632(.VSS(VSS),.VDD(VDD),.Y(I37113),.A(g28044));
  NOT NOT1_11633(.VSS(VSS),.VDD(VDD),.Y(g28288),.A(I37113));
  NOT NOT1_11634(.VSS(VSS),.VDD(VDD),.Y(I37116),.A(g28068));
  NOT NOT1_11635(.VSS(VSS),.VDD(VDD),.Y(g28289),.A(I37116));
  NOT NOT1_11636(.VSS(VSS),.VDD(VDD),.Y(I37119),.A(g28089));
  NOT NOT1_11637(.VSS(VSS),.VDD(VDD),.Y(g28290),.A(I37119));
  NOT NOT1_11638(.VSS(VSS),.VDD(VDD),.Y(I37122),.A(g28069));
  NOT NOT1_11639(.VSS(VSS),.VDD(VDD),.Y(g28291),.A(I37122));
  NOT NOT1_11640(.VSS(VSS),.VDD(VDD),.Y(I37125),.A(g28090));
  NOT NOT1_11641(.VSS(VSS),.VDD(VDD),.Y(g28292),.A(I37125));
  NOT NOT1_11642(.VSS(VSS),.VDD(VDD),.Y(I37128),.A(g28106));
  NOT NOT1_11643(.VSS(VSS),.VDD(VDD),.Y(g28293),.A(I37128));
  NOT NOT1_11644(.VSS(VSS),.VDD(VDD),.Y(I37131),.A(g28091));
  NOT NOT1_11645(.VSS(VSS),.VDD(VDD),.Y(g28294),.A(I37131));
  NOT NOT1_11646(.VSS(VSS),.VDD(VDD),.Y(I37134),.A(g28107));
  NOT NOT1_11647(.VSS(VSS),.VDD(VDD),.Y(g28295),.A(I37134));
  NOT NOT1_11648(.VSS(VSS),.VDD(VDD),.Y(I37137),.A(g28117));
  NOT NOT1_11649(.VSS(VSS),.VDD(VDD),.Y(g28296),.A(I37137));
  NOT NOT1_11650(.VSS(VSS),.VDD(VDD),.Y(I37140),.A(g28070));
  NOT NOT1_11651(.VSS(VSS),.VDD(VDD),.Y(g28297),.A(I37140));
  NOT NOT1_11652(.VSS(VSS),.VDD(VDD),.Y(I37143),.A(g28092));
  NOT NOT1_11653(.VSS(VSS),.VDD(VDD),.Y(g28298),.A(I37143));
  NOT NOT1_11654(.VSS(VSS),.VDD(VDD),.Y(I37146),.A(g28108));
  NOT NOT1_11655(.VSS(VSS),.VDD(VDD),.Y(g28299),.A(I37146));
  NOT NOT1_11656(.VSS(VSS),.VDD(VDD),.Y(I37149),.A(g28093));
  NOT NOT1_11657(.VSS(VSS),.VDD(VDD),.Y(g28300),.A(I37149));
  NOT NOT1_11658(.VSS(VSS),.VDD(VDD),.Y(I37152),.A(g28109));
  NOT NOT1_11659(.VSS(VSS),.VDD(VDD),.Y(g28301),.A(I37152));
  NOT NOT1_11660(.VSS(VSS),.VDD(VDD),.Y(I37155),.A(g28119));
  NOT NOT1_11661(.VSS(VSS),.VDD(VDD),.Y(g28302),.A(I37155));
  NOT NOT1_11662(.VSS(VSS),.VDD(VDD),.Y(I37158),.A(g28110));
  NOT NOT1_11663(.VSS(VSS),.VDD(VDD),.Y(g28303),.A(I37158));
  NOT NOT1_11664(.VSS(VSS),.VDD(VDD),.Y(I37161),.A(g28120));
  NOT NOT1_11665(.VSS(VSS),.VDD(VDD),.Y(g28304),.A(I37161));
  NOT NOT1_11666(.VSS(VSS),.VDD(VDD),.Y(I37164),.A(g28125));
  NOT NOT1_11667(.VSS(VSS),.VDD(VDD),.Y(g28305),.A(I37164));
  NOT NOT1_11668(.VSS(VSS),.VDD(VDD),.Y(I37167),.A(g28121));
  NOT NOT1_11669(.VSS(VSS),.VDD(VDD),.Y(g28306),.A(I37167));
  NOT NOT1_11670(.VSS(VSS),.VDD(VDD),.Y(I37170),.A(g28126));
  NOT NOT1_11671(.VSS(VSS),.VDD(VDD),.Y(g28307),.A(I37170));
  NOT NOT1_11672(.VSS(VSS),.VDD(VDD),.Y(I37173),.A(g28132));
  NOT NOT1_11673(.VSS(VSS),.VDD(VDD),.Y(g28308),.A(I37173));
  NOT NOT1_11674(.VSS(VSS),.VDD(VDD),.Y(I37176),.A(g27927));
  NOT NOT1_11675(.VSS(VSS),.VDD(VDD),.Y(g28309),.A(I37176));
  NOT NOT1_11676(.VSS(VSS),.VDD(VDD),.Y(I37179),.A(g27784));
  NOT NOT1_11677(.VSS(VSS),.VDD(VDD),.Y(g28310),.A(I37179));
  NOT NOT1_11678(.VSS(VSS),.VDD(VDD),.Y(I37182),.A(g27791));
  NOT NOT1_11679(.VSS(VSS),.VDD(VDD),.Y(g28311),.A(I37182));
  NOT NOT1_11680(.VSS(VSS),.VDD(VDD),.Y(I37185),.A(g27797));
  NOT NOT1_11681(.VSS(VSS),.VDD(VDD),.Y(g28312),.A(I37185));
  NOT NOT1_11682(.VSS(VSS),.VDD(VDD),.Y(I37188),.A(g27785));
  NOT NOT1_11683(.VSS(VSS),.VDD(VDD),.Y(g28313),.A(I37188));
  NOT NOT1_11684(.VSS(VSS),.VDD(VDD),.Y(I37191),.A(g27792));
  NOT NOT1_11685(.VSS(VSS),.VDD(VDD),.Y(g28314),.A(I37191));
  NOT NOT1_11686(.VSS(VSS),.VDD(VDD),.Y(I37194),.A(g27800));
  NOT NOT1_11687(.VSS(VSS),.VDD(VDD),.Y(g28315),.A(I37194));
  NOT NOT1_11688(.VSS(VSS),.VDD(VDD),.Y(I37197),.A(g27903));
  NOT NOT1_11689(.VSS(VSS),.VDD(VDD),.Y(g28316),.A(I37197));
  NOT NOT1_11690(.VSS(VSS),.VDD(VDD),.Y(I37200),.A(g27907));
  NOT NOT1_11691(.VSS(VSS),.VDD(VDD),.Y(g28317),.A(I37200));
  NOT NOT1_11692(.VSS(VSS),.VDD(VDD),.Y(I37203),.A(g27912));
  NOT NOT1_11693(.VSS(VSS),.VDD(VDD),.Y(g28318),.A(I37203));
  NOT NOT1_11694(.VSS(VSS),.VDD(VDD),.Y(I37228),.A(g28194));
  NOT NOT1_11695(.VSS(VSS),.VDD(VDD),.Y(g28341),.A(I37228));
  NOT NOT1_11696(.VSS(VSS),.VDD(VDD),.Y(I37232),.A(g28200));
  NOT NOT1_11697(.VSS(VSS),.VDD(VDD),.Y(g28343),.A(I37232));
  NOT NOT1_11698(.VSS(VSS),.VDD(VDD),.Y(I37238),.A(g28179));
  NOT NOT1_11699(.VSS(VSS),.VDD(VDD),.Y(g28347),.A(I37238));
  NOT NOT1_11700(.VSS(VSS),.VDD(VDD),.Y(I37252),.A(g28200));
  NOT NOT1_11701(.VSS(VSS),.VDD(VDD),.Y(g28359),.A(I37252));
  NOT NOT1_11702(.VSS(VSS),.VDD(VDD),.Y(I37260),.A(g28179));
  NOT NOT1_11703(.VSS(VSS),.VDD(VDD),.Y(g28365),.A(I37260));
  NOT NOT1_11704(.VSS(VSS),.VDD(VDD),.Y(I37266),.A(g28200));
  NOT NOT1_11705(.VSS(VSS),.VDD(VDD),.Y(g28369),.A(I37266));
  NOT NOT1_11706(.VSS(VSS),.VDD(VDD),.Y(I37269),.A(g28145));
  NOT NOT1_11707(.VSS(VSS),.VDD(VDD),.Y(g28370),.A(I37269));
  NOT NOT1_11708(.VSS(VSS),.VDD(VDD),.Y(I37273),.A(g28179));
  NOT NOT1_11709(.VSS(VSS),.VDD(VDD),.Y(g28372),.A(I37273));
  NOT NOT1_11710(.VSS(VSS),.VDD(VDD),.Y(I37277),.A(g28146));
  NOT NOT1_11711(.VSS(VSS),.VDD(VDD),.Y(g28374),.A(I37277));
  NOT NOT1_11712(.VSS(VSS),.VDD(VDD),.Y(I37280),.A(g28179));
  NOT NOT1_11713(.VSS(VSS),.VDD(VDD),.Y(g28375),.A(I37280));
  NOT NOT1_11714(.VSS(VSS),.VDD(VDD),.Y(I37284),.A(g28147));
  NOT NOT1_11715(.VSS(VSS),.VDD(VDD),.Y(g28377),.A(I37284));
  NOT NOT1_11716(.VSS(VSS),.VDD(VDD),.Y(I37291),.A(g28148));
  NOT NOT1_11717(.VSS(VSS),.VDD(VDD),.Y(g28382),.A(I37291));
  NOT NOT1_11718(.VSS(VSS),.VDD(VDD),.Y(I37319),.A(g28149));
  NOT NOT1_11719(.VSS(VSS),.VDD(VDD),.Y(g28390),.A(I37319));
  NOT NOT1_11720(.VSS(VSS),.VDD(VDD),.Y(I37330),.A(g28194));
  NOT NOT1_11721(.VSS(VSS),.VDD(VDD),.Y(g28393),.A(I37330));
  NOT NOT1_11722(.VSS(VSS),.VDD(VDD),.Y(I37334),.A(g28194));
  NOT NOT1_11723(.VSS(VSS),.VDD(VDD),.Y(g28395),.A(I37334));
  NOT NOT1_11724(.VSS(VSS),.VDD(VDD),.Y(g28419),.A(g28151));
  NOT NOT1_11725(.VSS(VSS),.VDD(VDD),.Y(I37379),.A(g28199));
  NOT NOT1_11726(.VSS(VSS),.VDD(VDD),.Y(g28432),.A(I37379));
  NOT NOT1_11727(.VSS(VSS),.VDD(VDD),.Y(I37386),.A(g28194));
  NOT NOT1_11728(.VSS(VSS),.VDD(VDD),.Y(g28437),.A(I37386));
  NOT NOT1_11729(.VSS(VSS),.VDD(VDD),.Y(I37394),.A(g27718));
  NOT NOT1_11730(.VSS(VSS),.VDD(VDD),.Y(g28443),.A(I37394));
  NOT NOT1_11731(.VSS(VSS),.VDD(VDD),.Y(I37400),.A(g28200));
  NOT NOT1_11732(.VSS(VSS),.VDD(VDD),.Y(g28447),.A(I37400));
  NOT NOT1_11733(.VSS(VSS),.VDD(VDD),.Y(I37410),.A(g27722));
  NOT NOT1_11734(.VSS(VSS),.VDD(VDD),.Y(g28455),.A(I37410));
  NOT NOT1_11735(.VSS(VSS),.VDD(VDD),.Y(I37415),.A(g28179));
  NOT NOT1_11736(.VSS(VSS),.VDD(VDD),.Y(g28458),.A(I37415));
  NOT NOT1_11737(.VSS(VSS),.VDD(VDD),.Y(I37426),.A(g27724));
  NOT NOT1_11738(.VSS(VSS),.VDD(VDD),.Y(g28467),.A(I37426));
  NOT NOT1_11739(.VSS(VSS),.VDD(VDD),.Y(g28483),.A(g27776));
  NOT NOT1_11740(.VSS(VSS),.VDD(VDD),.Y(g28491),.A(g27780));
  NOT NOT1_11741(.VSS(VSS),.VDD(VDD),.Y(g28496),.A(g27787));
  NOT NOT1_11742(.VSS(VSS),.VDD(VDD),.Y(I37459),.A(g27759));
  NOT NOT1_11743(.VSS(VSS),.VDD(VDD),.Y(g28498),.A(I37459));
  NOT NOT1_11744(.VSS(VSS),.VDD(VDD),.Y(g28500),.A(g27794));
  NOT NOT1_11745(.VSS(VSS),.VDD(VDD),.Y(I37467),.A(g27760));
  NOT NOT1_11746(.VSS(VSS),.VDD(VDD),.Y(g28524),.A(I37467));
  NOT NOT1_11747(.VSS(VSS),.VDD(VDD),.Y(I37471),.A(g27761));
  NOT NOT1_11748(.VSS(VSS),.VDD(VDD),.Y(g28526),.A(I37471));
  NOT NOT1_11749(.VSS(VSS),.VDD(VDD),.Y(I37474),.A(g27762));
  NOT NOT1_11750(.VSS(VSS),.VDD(VDD),.Y(g28527),.A(I37474));
  NOT NOT1_11751(.VSS(VSS),.VDD(VDD),.Y(I37481),.A(g27763));
  NOT NOT1_11752(.VSS(VSS),.VDD(VDD),.Y(g28552),.A(I37481));
  NOT NOT1_11753(.VSS(VSS),.VDD(VDD),.Y(I37484),.A(g27764));
  NOT NOT1_11754(.VSS(VSS),.VDD(VDD),.Y(g28553),.A(I37484));
  NOT NOT1_11755(.VSS(VSS),.VDD(VDD),.Y(g28554),.A(g27806));
  NOT NOT1_11756(.VSS(VSS),.VDD(VDD),.Y(I37488),.A(g27765));
  NOT NOT1_11757(.VSS(VSS),.VDD(VDD),.Y(g28555),.A(I37488));
  NOT NOT1_11758(.VSS(VSS),.VDD(VDD),.Y(I37494),.A(g27766));
  NOT NOT1_11759(.VSS(VSS),.VDD(VDD),.Y(g28579),.A(I37494));
  NOT NOT1_11760(.VSS(VSS),.VDD(VDD),.Y(I37497),.A(g27767));
  NOT NOT1_11761(.VSS(VSS),.VDD(VDD),.Y(g28580),.A(I37497));
  NOT NOT1_11762(.VSS(VSS),.VDD(VDD),.Y(g28581),.A(g27817));
  NOT NOT1_11763(.VSS(VSS),.VDD(VDD),.Y(g28582),.A(g27820));
  NOT NOT1_11764(.VSS(VSS),.VDD(VDD),.Y(I37502),.A(g27768));
  NOT NOT1_11765(.VSS(VSS),.VDD(VDD),.Y(g28583),.A(I37502));
  NOT NOT1_11766(.VSS(VSS),.VDD(VDD),.Y(I37508),.A(g27769));
  NOT NOT1_11767(.VSS(VSS),.VDD(VDD),.Y(g28607),.A(I37508));
  NOT NOT1_11768(.VSS(VSS),.VDD(VDD),.Y(g28608),.A(g27831));
  NOT NOT1_11769(.VSS(VSS),.VDD(VDD),.Y(g28609),.A(g27839));
  NOT NOT1_11770(.VSS(VSS),.VDD(VDD),.Y(g28610),.A(g27843));
  NOT NOT1_11771(.VSS(VSS),.VDD(VDD),.Y(I37514),.A(g27771));
  NOT NOT1_11772(.VSS(VSS),.VDD(VDD),.Y(g28611),.A(I37514));
  NOT NOT1_11773(.VSS(VSS),.VDD(VDD),.Y(g28612),.A(g28046));
  NOT NOT1_11774(.VSS(VSS),.VDD(VDD),.Y(g28616),.A(g27847));
  NOT NOT1_11775(.VSS(VSS),.VDD(VDD),.Y(g28617),.A(g27858));
  NOT NOT1_11776(.VSS(VSS),.VDD(VDD),.Y(g28618),.A(g27861));
  NOT NOT1_11777(.VSS(VSS),.VDD(VDD),.Y(g28619),.A(g28075));
  NOT NOT1_11778(.VSS(VSS),.VDD(VDD),.Y(g28623),.A(g27872));
  NOT NOT1_11779(.VSS(VSS),.VDD(VDD),.Y(g28624),.A(g27879));
  NOT NOT1_11780(.VSS(VSS),.VDD(VDD),.Y(g28625),.A(g28100));
  NOT NOT1_11781(.VSS(VSS),.VDD(VDD),.Y(g28629),.A(g27889));
  NOT NOT1_11782(.VSS(VSS),.VDD(VDD),.Y(g28630),.A(g28118));
  NOT NOT1_11783(.VSS(VSS),.VDD(VDD),.Y(g28638),.A(g28200));
  NOT NOT1_11784(.VSS(VSS),.VDD(VDD),.Y(g28639),.A(g27919));
  NOT NOT1_11785(.VSS(VSS),.VDD(VDD),.Y(g28640),.A(g27928));
  NOT NOT1_11786(.VSS(VSS),.VDD(VDD),.Y(g28641),.A(g27932));
  NOT NOT1_11787(.VSS(VSS),.VDD(VDD),.Y(g28642),.A(g27939));
  NOT NOT1_11788(.VSS(VSS),.VDD(VDD),.Y(g28643),.A(g27942));
  NOT NOT1_11789(.VSS(VSS),.VDD(VDD),.Y(g28644),.A(g27946));
  NOT NOT1_11790(.VSS(VSS),.VDD(VDD),.Y(g28645),.A(g27952));
  NOT NOT1_11791(.VSS(VSS),.VDD(VDD),.Y(g28646),.A(g27956));
  NOT NOT1_11792(.VSS(VSS),.VDD(VDD),.Y(g28647),.A(g27959));
  NOT NOT1_11793(.VSS(VSS),.VDD(VDD),.Y(g28648),.A(g27965));
  NOT NOT1_11794(.VSS(VSS),.VDD(VDD),.Y(g28649),.A(g27973));
  NOT NOT1_11795(.VSS(VSS),.VDD(VDD),.Y(g28650),.A(g27977));
  NOT NOT1_11796(.VSS(VSS),.VDD(VDD),.Y(g28651),.A(g27981));
  NOT NOT1_11797(.VSS(VSS),.VDD(VDD),.Y(g28652),.A(g27994));
  NOT NOT1_11798(.VSS(VSS),.VDD(VDD),.Y(g28653),.A(g27999));
  NOT NOT1_11799(.VSS(VSS),.VDD(VDD),.Y(g28655),.A(g28018));
  NOT NOT1_11800(.VSS(VSS),.VDD(VDD),.Y(I37566),.A(g28370));
  NOT NOT1_11801(.VSS(VSS),.VDD(VDD),.Y(g28673),.A(I37566));
  NOT NOT1_11802(.VSS(VSS),.VDD(VDD),.Y(I37569),.A(g28498));
  NOT NOT1_11803(.VSS(VSS),.VDD(VDD),.Y(g28674),.A(I37569));
  NOT NOT1_11804(.VSS(VSS),.VDD(VDD),.Y(I37572),.A(g28524));
  NOT NOT1_11805(.VSS(VSS),.VDD(VDD),.Y(g28675),.A(I37572));
  NOT NOT1_11806(.VSS(VSS),.VDD(VDD),.Y(I37575),.A(g28527));
  NOT NOT1_11807(.VSS(VSS),.VDD(VDD),.Y(g28676),.A(I37575));
  NOT NOT1_11808(.VSS(VSS),.VDD(VDD),.Y(I37578),.A(g28432));
  NOT NOT1_11809(.VSS(VSS),.VDD(VDD),.Y(g28677),.A(I37578));
  NOT NOT1_11810(.VSS(VSS),.VDD(VDD),.Y(I37581),.A(g28374));
  NOT NOT1_11811(.VSS(VSS),.VDD(VDD),.Y(g28678),.A(I37581));
  NOT NOT1_11812(.VSS(VSS),.VDD(VDD),.Y(I37584),.A(g28526));
  NOT NOT1_11813(.VSS(VSS),.VDD(VDD),.Y(g28679),.A(I37584));
  NOT NOT1_11814(.VSS(VSS),.VDD(VDD),.Y(I37587),.A(g28552));
  NOT NOT1_11815(.VSS(VSS),.VDD(VDD),.Y(g28680),.A(I37587));
  NOT NOT1_11816(.VSS(VSS),.VDD(VDD),.Y(I37590),.A(g28555));
  NOT NOT1_11817(.VSS(VSS),.VDD(VDD),.Y(g28681),.A(I37590));
  NOT NOT1_11818(.VSS(VSS),.VDD(VDD),.Y(I37593),.A(g28443));
  NOT NOT1_11819(.VSS(VSS),.VDD(VDD),.Y(g28682),.A(I37593));
  NOT NOT1_11820(.VSS(VSS),.VDD(VDD),.Y(I37596),.A(g28377));
  NOT NOT1_11821(.VSS(VSS),.VDD(VDD),.Y(g28683),.A(I37596));
  NOT NOT1_11822(.VSS(VSS),.VDD(VDD),.Y(I37599),.A(g28553));
  NOT NOT1_11823(.VSS(VSS),.VDD(VDD),.Y(g28684),.A(I37599));
  NOT NOT1_11824(.VSS(VSS),.VDD(VDD),.Y(I37602),.A(g28579));
  NOT NOT1_11825(.VSS(VSS),.VDD(VDD),.Y(g28685),.A(I37602));
  NOT NOT1_11826(.VSS(VSS),.VDD(VDD),.Y(I37605),.A(g28583));
  NOT NOT1_11827(.VSS(VSS),.VDD(VDD),.Y(g28686),.A(I37605));
  NOT NOT1_11828(.VSS(VSS),.VDD(VDD),.Y(I37608),.A(g28455));
  NOT NOT1_11829(.VSS(VSS),.VDD(VDD),.Y(g28687),.A(I37608));
  NOT NOT1_11830(.VSS(VSS),.VDD(VDD),.Y(I37611),.A(g28382));
  NOT NOT1_11831(.VSS(VSS),.VDD(VDD),.Y(g28688),.A(I37611));
  NOT NOT1_11832(.VSS(VSS),.VDD(VDD),.Y(I37614),.A(g28580));
  NOT NOT1_11833(.VSS(VSS),.VDD(VDD),.Y(g28689),.A(I37614));
  NOT NOT1_11834(.VSS(VSS),.VDD(VDD),.Y(I37617),.A(g28607));
  NOT NOT1_11835(.VSS(VSS),.VDD(VDD),.Y(g28690),.A(I37617));
  NOT NOT1_11836(.VSS(VSS),.VDD(VDD),.Y(I37620),.A(g28611));
  NOT NOT1_11837(.VSS(VSS),.VDD(VDD),.Y(g28691),.A(I37620));
  NOT NOT1_11838(.VSS(VSS),.VDD(VDD),.Y(I37623),.A(g28467));
  NOT NOT1_11839(.VSS(VSS),.VDD(VDD),.Y(g28692),.A(I37623));
  NOT NOT1_11840(.VSS(VSS),.VDD(VDD),.Y(I37626),.A(g28393));
  NOT NOT1_11841(.VSS(VSS),.VDD(VDD),.Y(g28693),.A(I37626));
  NOT NOT1_11842(.VSS(VSS),.VDD(VDD),.Y(I37629),.A(g28369));
  NOT NOT1_11843(.VSS(VSS),.VDD(VDD),.Y(g28694),.A(I37629));
  NOT NOT1_11844(.VSS(VSS),.VDD(VDD),.Y(I37632),.A(g28372));
  NOT NOT1_11845(.VSS(VSS),.VDD(VDD),.Y(g28695),.A(I37632));
  NOT NOT1_11846(.VSS(VSS),.VDD(VDD),.Y(I37635),.A(g28390));
  NOT NOT1_11847(.VSS(VSS),.VDD(VDD),.Y(g28696),.A(I37635));
  NOT NOT1_11848(.VSS(VSS),.VDD(VDD),.Y(I37638),.A(g28395));
  NOT NOT1_11849(.VSS(VSS),.VDD(VDD),.Y(g28697),.A(I37638));
  NOT NOT1_11850(.VSS(VSS),.VDD(VDD),.Y(I37641),.A(g28375));
  NOT NOT1_11851(.VSS(VSS),.VDD(VDD),.Y(g28698),.A(I37641));
  NOT NOT1_11852(.VSS(VSS),.VDD(VDD),.Y(I37644),.A(g28341));
  NOT NOT1_11853(.VSS(VSS),.VDD(VDD),.Y(g28699),.A(I37644));
  NOT NOT1_11854(.VSS(VSS),.VDD(VDD),.Y(I37647),.A(g28343));
  NOT NOT1_11855(.VSS(VSS),.VDD(VDD),.Y(g28700),.A(I37647));
  NOT NOT1_11856(.VSS(VSS),.VDD(VDD),.Y(I37650),.A(g28347));
  NOT NOT1_11857(.VSS(VSS),.VDD(VDD),.Y(g28701),.A(I37650));
  NOT NOT1_11858(.VSS(VSS),.VDD(VDD),.Y(I37653),.A(g28359));
  NOT NOT1_11859(.VSS(VSS),.VDD(VDD),.Y(g28702),.A(I37653));
  NOT NOT1_11860(.VSS(VSS),.VDD(VDD),.Y(I37656),.A(g28365));
  NOT NOT1_11861(.VSS(VSS),.VDD(VDD),.Y(g28703),.A(I37656));
  NOT NOT1_11862(.VSS(VSS),.VDD(VDD),.Y(I37659),.A(g28437));
  NOT NOT1_11863(.VSS(VSS),.VDD(VDD),.Y(g28704),.A(I37659));
  NOT NOT1_11864(.VSS(VSS),.VDD(VDD),.Y(I37662),.A(g28447));
  NOT NOT1_11865(.VSS(VSS),.VDD(VDD),.Y(g28705),.A(I37662));
  NOT NOT1_11866(.VSS(VSS),.VDD(VDD),.Y(I37665),.A(g28458));
  NOT NOT1_11867(.VSS(VSS),.VDD(VDD),.Y(g28706),.A(I37665));
  NOT NOT1_11868(.VSS(VSS),.VDD(VDD),.Y(g28720),.A(g28495));
  NOT NOT1_11869(.VSS(VSS),.VDD(VDD),.Y(g28721),.A(g28490));
  NOT NOT1_11870(.VSS(VSS),.VDD(VDD),.Y(g28723),.A(g28528));
  NOT NOT1_11871(.VSS(VSS),.VDD(VDD),.Y(g28725),.A(g28499));
  NOT NOT1_11872(.VSS(VSS),.VDD(VDD),.Y(g28727),.A(g28489));
  NOT NOT1_11873(.VSS(VSS),.VDD(VDD),.Y(g28730),.A(g28470));
  NOT NOT1_11874(.VSS(VSS),.VDD(VDD),.Y(g28734),.A(g28525));
  NOT NOT1_11875(.VSS(VSS),.VDD(VDD),.Y(g28740),.A(g28488));
  NOT NOT1_11876(.VSS(VSS),.VDD(VDD),.Y(I37702),.A(g28512));
  NOT NOT1_11877(.VSS(VSS),.VDD(VDD),.Y(g28741),.A(I37702));
  NOT NOT1_11878(.VSS(VSS),.VDD(VDD),.Y(I37712),.A(g28512));
  NOT NOT1_11879(.VSS(VSS),.VDD(VDD),.Y(g28751),.A(I37712));
  NOT NOT1_11880(.VSS(VSS),.VDD(VDD),.Y(I37716),.A(g28540));
  NOT NOT1_11881(.VSS(VSS),.VDD(VDD),.Y(g28755),.A(I37716));
  NOT NOT1_11882(.VSS(VSS),.VDD(VDD),.Y(I37725),.A(g28540));
  NOT NOT1_11883(.VSS(VSS),.VDD(VDD),.Y(g28764),.A(I37725));
  NOT NOT1_11884(.VSS(VSS),.VDD(VDD),.Y(I37729),.A(g28567));
  NOT NOT1_11885(.VSS(VSS),.VDD(VDD),.Y(g28768),.A(I37729));
  NOT NOT1_11886(.VSS(VSS),.VDD(VDD),.Y(I37736),.A(g28567));
  NOT NOT1_11887(.VSS(VSS),.VDD(VDD),.Y(g28775),.A(I37736));
  NOT NOT1_11888(.VSS(VSS),.VDD(VDD),.Y(I37740),.A(g28595));
  NOT NOT1_11889(.VSS(VSS),.VDD(VDD),.Y(g28779),.A(I37740));
  NOT NOT1_11890(.VSS(VSS),.VDD(VDD),.Y(I37746),.A(g28595));
  NOT NOT1_11891(.VSS(VSS),.VDD(VDD),.Y(g28785),.A(I37746));
  NOT NOT1_11892(.VSS(VSS),.VDD(VDD),.Y(I37752),.A(g28512));
  NOT NOT1_11893(.VSS(VSS),.VDD(VDD),.Y(g28791),.A(I37752));
  NOT NOT1_11894(.VSS(VSS),.VDD(VDD),.Y(I37757),.A(g28512));
  NOT NOT1_11895(.VSS(VSS),.VDD(VDD),.Y(g28796),.A(I37757));
  NOT NOT1_11896(.VSS(VSS),.VDD(VDD),.Y(I37760),.A(g28540));
  NOT NOT1_11897(.VSS(VSS),.VDD(VDD),.Y(g28799),.A(I37760));
  NOT NOT1_11898(.VSS(VSS),.VDD(VDD),.Y(I37765),.A(g28512));
  NOT NOT1_11899(.VSS(VSS),.VDD(VDD),.Y(g28804),.A(I37765));
  NOT NOT1_11900(.VSS(VSS),.VDD(VDD),.Y(I37768),.A(g28540));
  NOT NOT1_11901(.VSS(VSS),.VDD(VDD),.Y(g28807),.A(I37768));
  NOT NOT1_11902(.VSS(VSS),.VDD(VDD),.Y(I37771),.A(g28567));
  NOT NOT1_11903(.VSS(VSS),.VDD(VDD),.Y(g28810),.A(I37771));
  NOT NOT1_11904(.VSS(VSS),.VDD(VDD),.Y(I37775),.A(g28540));
  NOT NOT1_11905(.VSS(VSS),.VDD(VDD),.Y(g28814),.A(I37775));
  NOT NOT1_11906(.VSS(VSS),.VDD(VDD),.Y(I37778),.A(g28567));
  NOT NOT1_11907(.VSS(VSS),.VDD(VDD),.Y(g28817),.A(I37778));
  NOT NOT1_11908(.VSS(VSS),.VDD(VDD),.Y(I37781),.A(g28595));
  NOT NOT1_11909(.VSS(VSS),.VDD(VDD),.Y(g28820),.A(I37781));
  NOT NOT1_11910(.VSS(VSS),.VDD(VDD),.Y(I37784),.A(g28567));
  NOT NOT1_11911(.VSS(VSS),.VDD(VDD),.Y(g28823),.A(I37784));
  NOT NOT1_11912(.VSS(VSS),.VDD(VDD),.Y(I37787),.A(g28595));
  NOT NOT1_11913(.VSS(VSS),.VDD(VDD),.Y(g28826),.A(I37787));
  NOT NOT1_11914(.VSS(VSS),.VDD(VDD),.Y(I37790),.A(g28595));
  NOT NOT1_11915(.VSS(VSS),.VDD(VDD),.Y(g28829),.A(I37790));
  NOT NOT1_11916(.VSS(VSS),.VDD(VDD),.Y(I37793),.A(g28638));
  NOT NOT1_11917(.VSS(VSS),.VDD(VDD),.Y(g28832),.A(I37793));
  NOT NOT1_11918(.VSS(VSS),.VDD(VDD),.Y(I37796),.A(g28634));
  NOT NOT1_11919(.VSS(VSS),.VDD(VDD),.Y(g28833),.A(I37796));
  NOT NOT1_11920(.VSS(VSS),.VDD(VDD),.Y(I37800),.A(g28635));
  NOT NOT1_11921(.VSS(VSS),.VDD(VDD),.Y(g28835),.A(I37800));
  NOT NOT1_11922(.VSS(VSS),.VDD(VDD),.Y(I37804),.A(g28636));
  NOT NOT1_11923(.VSS(VSS),.VDD(VDD),.Y(g28837),.A(I37804));
  NOT NOT1_11924(.VSS(VSS),.VDD(VDD),.Y(I37808),.A(g28637));
  NOT NOT1_11925(.VSS(VSS),.VDD(VDD),.Y(g28839),.A(I37808));
  NOT NOT1_11926(.VSS(VSS),.VDD(VDD),.Y(g28855),.A(g28409));
  NOT NOT1_11927(.VSS(VSS),.VDD(VDD),.Y(g28859),.A(g28413));
  NOT NOT1_11928(.VSS(VSS),.VDD(VDD),.Y(g28863),.A(g28417));
  NOT NOT1_11929(.VSS(VSS),.VDD(VDD),.Y(g28867),.A(g28418));
  NOT NOT1_11930(.VSS(VSS),.VDD(VDD),.Y(I37842),.A(g28501));
  NOT NOT1_11931(.VSS(VSS),.VDD(VDD),.Y(g28871),.A(I37842));
  NOT NOT1_11932(.VSS(VSS),.VDD(VDD),.Y(I37846),.A(g28501));
  NOT NOT1_11933(.VSS(VSS),.VDD(VDD),.Y(g28877),.A(I37846));
  NOT NOT1_11934(.VSS(VSS),.VDD(VDD),.Y(I37851),.A(g28668));
  NOT NOT1_11935(.VSS(VSS),.VDD(VDD),.Y(g28882),.A(I37851));
  NOT NOT1_11936(.VSS(VSS),.VDD(VDD),.Y(I37854),.A(g28529));
  NOT NOT1_11937(.VSS(VSS),.VDD(VDD),.Y(g28883),.A(I37854));
  NOT NOT1_11938(.VSS(VSS),.VDD(VDD),.Y(I37858),.A(g28501));
  NOT NOT1_11939(.VSS(VSS),.VDD(VDD),.Y(g28889),.A(I37858));
  NOT NOT1_11940(.VSS(VSS),.VDD(VDD),.Y(I37863),.A(g28529));
  NOT NOT1_11941(.VSS(VSS),.VDD(VDD),.Y(g28894),.A(I37863));
  NOT NOT1_11942(.VSS(VSS),.VDD(VDD),.Y(I37868),.A(g28321));
  NOT NOT1_11943(.VSS(VSS),.VDD(VDD),.Y(g28899),.A(I37868));
  NOT NOT1_11944(.VSS(VSS),.VDD(VDD),.Y(I37871),.A(g28556));
  NOT NOT1_11945(.VSS(VSS),.VDD(VDD),.Y(g28900),.A(I37871));
  NOT NOT1_11946(.VSS(VSS),.VDD(VDD),.Y(I37875),.A(g28501));
  NOT NOT1_11947(.VSS(VSS),.VDD(VDD),.Y(g28906),.A(I37875));
  NOT NOT1_11948(.VSS(VSS),.VDD(VDD),.Y(I37880),.A(g28529));
  NOT NOT1_11949(.VSS(VSS),.VDD(VDD),.Y(g28911),.A(I37880));
  NOT NOT1_11950(.VSS(VSS),.VDD(VDD),.Y(I37885),.A(g28556));
  NOT NOT1_11951(.VSS(VSS),.VDD(VDD),.Y(g28916),.A(I37885));
  NOT NOT1_11952(.VSS(VSS),.VDD(VDD),.Y(I37891),.A(g28325));
  NOT NOT1_11953(.VSS(VSS),.VDD(VDD),.Y(g28924),.A(I37891));
  NOT NOT1_11954(.VSS(VSS),.VDD(VDD),.Y(I37894),.A(g28584));
  NOT NOT1_11955(.VSS(VSS),.VDD(VDD),.Y(g28925),.A(I37894));
  NOT NOT1_11956(.VSS(VSS),.VDD(VDD),.Y(I37897),.A(g28501));
  NOT NOT1_11957(.VSS(VSS),.VDD(VDD),.Y(g28928),.A(I37897));
  NOT NOT1_11958(.VSS(VSS),.VDD(VDD),.Y(I37901),.A(g28529));
  NOT NOT1_11959(.VSS(VSS),.VDD(VDD),.Y(g28932),.A(I37901));
  NOT NOT1_11960(.VSS(VSS),.VDD(VDD),.Y(I37906),.A(g28556));
  NOT NOT1_11961(.VSS(VSS),.VDD(VDD),.Y(g28937),.A(I37906));
  NOT NOT1_11962(.VSS(VSS),.VDD(VDD),.Y(I37912),.A(g28584));
  NOT NOT1_11963(.VSS(VSS),.VDD(VDD),.Y(g28945),.A(I37912));
  NOT NOT1_11964(.VSS(VSS),.VDD(VDD),.Y(I37917),.A(g28328));
  NOT NOT1_11965(.VSS(VSS),.VDD(VDD),.Y(g28950),.A(I37917));
  NOT NOT1_11966(.VSS(VSS),.VDD(VDD),.Y(I37920),.A(g28501));
  NOT NOT1_11967(.VSS(VSS),.VDD(VDD),.Y(g28951),.A(I37920));
  NOT NOT1_11968(.VSS(VSS),.VDD(VDD),.Y(I37924),.A(g28529));
  NOT NOT1_11969(.VSS(VSS),.VDD(VDD),.Y(g28955),.A(I37924));
  NOT NOT1_11970(.VSS(VSS),.VDD(VDD),.Y(I37928),.A(g28556));
  NOT NOT1_11971(.VSS(VSS),.VDD(VDD),.Y(g28959),.A(I37928));
  NOT NOT1_11972(.VSS(VSS),.VDD(VDD),.Y(I37934),.A(g28584));
  NOT NOT1_11973(.VSS(VSS),.VDD(VDD),.Y(g28967),.A(I37934));
  NOT NOT1_11974(.VSS(VSS),.VDD(VDD),.Y(I37939),.A(g28501));
  NOT NOT1_11975(.VSS(VSS),.VDD(VDD),.Y(g28972),.A(I37939));
  NOT NOT1_11976(.VSS(VSS),.VDD(VDD),.Y(I37942),.A(g28501));
  NOT NOT1_11977(.VSS(VSS),.VDD(VDD),.Y(g28975),.A(I37942));
  NOT NOT1_11978(.VSS(VSS),.VDD(VDD),.Y(I37946),.A(g28529));
  NOT NOT1_11979(.VSS(VSS),.VDD(VDD),.Y(g28979),.A(I37946));
  NOT NOT1_11980(.VSS(VSS),.VDD(VDD),.Y(I37950),.A(g28556));
  NOT NOT1_11981(.VSS(VSS),.VDD(VDD),.Y(g28983),.A(I37950));
  NOT NOT1_11982(.VSS(VSS),.VDD(VDD),.Y(I37956),.A(g28584));
  NOT NOT1_11983(.VSS(VSS),.VDD(VDD),.Y(g28993),.A(I37956));
  NOT NOT1_11984(.VSS(VSS),.VDD(VDD),.Y(I37961),.A(g28501));
  NOT NOT1_11985(.VSS(VSS),.VDD(VDD),.Y(g28998),.A(I37961));
  NOT NOT1_11986(.VSS(VSS),.VDD(VDD),.Y(I37965),.A(g28529));
  NOT NOT1_11987(.VSS(VSS),.VDD(VDD),.Y(g29002),.A(I37965));
  NOT NOT1_11988(.VSS(VSS),.VDD(VDD),.Y(I37968),.A(g28529));
  NOT NOT1_11989(.VSS(VSS),.VDD(VDD),.Y(g29005),.A(I37968));
  NOT NOT1_11990(.VSS(VSS),.VDD(VDD),.Y(I37973),.A(g28556));
  NOT NOT1_11991(.VSS(VSS),.VDD(VDD),.Y(g29010),.A(I37973));
  NOT NOT1_11992(.VSS(VSS),.VDD(VDD),.Y(I37978),.A(g28584));
  NOT NOT1_11993(.VSS(VSS),.VDD(VDD),.Y(g29019),.A(I37978));
  NOT NOT1_11994(.VSS(VSS),.VDD(VDD),.Y(I37982),.A(g28501));
  NOT NOT1_11995(.VSS(VSS),.VDD(VDD),.Y(g29023),.A(I37982));
  NOT NOT1_11996(.VSS(VSS),.VDD(VDD),.Y(I37986),.A(g28529));
  NOT NOT1_11997(.VSS(VSS),.VDD(VDD),.Y(g29027),.A(I37986));
  NOT NOT1_11998(.VSS(VSS),.VDD(VDD),.Y(I37991),.A(g28556));
  NOT NOT1_11999(.VSS(VSS),.VDD(VDD),.Y(g29032),.A(I37991));
  NOT NOT1_12000(.VSS(VSS),.VDD(VDD),.Y(I37994),.A(g28556));
  NOT NOT1_12001(.VSS(VSS),.VDD(VDD),.Y(g29035),.A(I37994));
  NOT NOT1_12002(.VSS(VSS),.VDD(VDD),.Y(I37999),.A(g28584));
  NOT NOT1_12003(.VSS(VSS),.VDD(VDD),.Y(g29042),.A(I37999));
  NOT NOT1_12004(.VSS(VSS),.VDD(VDD),.Y(I38003),.A(g28529));
  NOT NOT1_12005(.VSS(VSS),.VDD(VDD),.Y(g29046),.A(I38003));
  NOT NOT1_12006(.VSS(VSS),.VDD(VDD),.Y(I38007),.A(g28556));
  NOT NOT1_12007(.VSS(VSS),.VDD(VDD),.Y(g29050),.A(I38007));
  NOT NOT1_12008(.VSS(VSS),.VDD(VDD),.Y(I38011),.A(g28584));
  NOT NOT1_12009(.VSS(VSS),.VDD(VDD),.Y(g29054),.A(I38011));
  NOT NOT1_12010(.VSS(VSS),.VDD(VDD),.Y(I38014),.A(g28584));
  NOT NOT1_12011(.VSS(VSS),.VDD(VDD),.Y(g29057),.A(I38014));
  NOT NOT1_12012(.VSS(VSS),.VDD(VDD),.Y(I38018),.A(g28342));
  NOT NOT1_12013(.VSS(VSS),.VDD(VDD),.Y(g29061),.A(I38018));
  NOT NOT1_12014(.VSS(VSS),.VDD(VDD),.Y(I38024),.A(g28556));
  NOT NOT1_12015(.VSS(VSS),.VDD(VDD),.Y(g29065),.A(I38024));
  NOT NOT1_12016(.VSS(VSS),.VDD(VDD),.Y(I38028),.A(g28584));
  NOT NOT1_12017(.VSS(VSS),.VDD(VDD),.Y(g29069),.A(I38028));
  NOT NOT1_12018(.VSS(VSS),.VDD(VDD),.Y(I38032),.A(g28344));
  NOT NOT1_12019(.VSS(VSS),.VDD(VDD),.Y(g29073),.A(I38032));
  NOT NOT1_12020(.VSS(VSS),.VDD(VDD),.Y(I38035),.A(g28345));
  NOT NOT1_12021(.VSS(VSS),.VDD(VDD),.Y(g29074),.A(I38035));
  NOT NOT1_12022(.VSS(VSS),.VDD(VDD),.Y(I38038),.A(g28346));
  NOT NOT1_12023(.VSS(VSS),.VDD(VDD),.Y(g29075),.A(I38038));
  NOT NOT1_12024(.VSS(VSS),.VDD(VDD),.Y(I38042),.A(g28584));
  NOT NOT1_12025(.VSS(VSS),.VDD(VDD),.Y(g29077),.A(I38042));
  NOT NOT1_12026(.VSS(VSS),.VDD(VDD),.Y(I38046),.A(g28348));
  NOT NOT1_12027(.VSS(VSS),.VDD(VDD),.Y(g29081),.A(I38046));
  NOT NOT1_12028(.VSS(VSS),.VDD(VDD),.Y(I38049),.A(g28349));
  NOT NOT1_12029(.VSS(VSS),.VDD(VDD),.Y(g29082),.A(I38049));
  NOT NOT1_12030(.VSS(VSS),.VDD(VDD),.Y(I38053),.A(g28350));
  NOT NOT1_12031(.VSS(VSS),.VDD(VDD),.Y(g29084),.A(I38053));
  NOT NOT1_12032(.VSS(VSS),.VDD(VDD),.Y(I38056),.A(g28351));
  NOT NOT1_12033(.VSS(VSS),.VDD(VDD),.Y(g29085),.A(I38056));
  NOT NOT1_12034(.VSS(VSS),.VDD(VDD),.Y(I38059),.A(g28352));
  NOT NOT1_12035(.VSS(VSS),.VDD(VDD),.Y(g29086),.A(I38059));
  NOT NOT1_12036(.VSS(VSS),.VDD(VDD),.Y(I38064),.A(g28353));
  NOT NOT1_12037(.VSS(VSS),.VDD(VDD),.Y(g29089),.A(I38064));
  NOT NOT1_12038(.VSS(VSS),.VDD(VDD),.Y(I38068),.A(g28354));
  NOT NOT1_12039(.VSS(VSS),.VDD(VDD),.Y(g29091),.A(I38068));
  NOT NOT1_12040(.VSS(VSS),.VDD(VDD),.Y(I38071),.A(g28355));
  NOT NOT1_12041(.VSS(VSS),.VDD(VDD),.Y(g29092),.A(I38071));
  NOT NOT1_12042(.VSS(VSS),.VDD(VDD),.Y(I38074),.A(g28356));
  NOT NOT1_12043(.VSS(VSS),.VDD(VDD),.Y(g29093),.A(I38074));
  NOT NOT1_12044(.VSS(VSS),.VDD(VDD),.Y(I38077),.A(g28357));
  NOT NOT1_12045(.VSS(VSS),.VDD(VDD),.Y(g29094),.A(I38077));
  NOT NOT1_12046(.VSS(VSS),.VDD(VDD),.Y(I38080),.A(g28358));
  NOT NOT1_12047(.VSS(VSS),.VDD(VDD),.Y(g29095),.A(I38080));
  NOT NOT1_12048(.VSS(VSS),.VDD(VDD),.Y(I38085),.A(g28360));
  NOT NOT1_12049(.VSS(VSS),.VDD(VDD),.Y(g29098),.A(I38085));
  NOT NOT1_12050(.VSS(VSS),.VDD(VDD),.Y(I38088),.A(g28361));
  NOT NOT1_12051(.VSS(VSS),.VDD(VDD),.Y(g29099),.A(I38088));
  NOT NOT1_12052(.VSS(VSS),.VDD(VDD),.Y(I38091),.A(g28362));
  NOT NOT1_12053(.VSS(VSS),.VDD(VDD),.Y(g29100),.A(I38091));
  NOT NOT1_12054(.VSS(VSS),.VDD(VDD),.Y(I38094),.A(g28363));
  NOT NOT1_12055(.VSS(VSS),.VDD(VDD),.Y(g29101),.A(I38094));
  NOT NOT1_12056(.VSS(VSS),.VDD(VDD),.Y(I38097),.A(g28364));
  NOT NOT1_12057(.VSS(VSS),.VDD(VDD),.Y(g29102),.A(I38097));
  NOT NOT1_12058(.VSS(VSS),.VDD(VDD),.Y(I38101),.A(g28366));
  NOT NOT1_12059(.VSS(VSS),.VDD(VDD),.Y(g29104),.A(I38101));
  NOT NOT1_12060(.VSS(VSS),.VDD(VDD),.Y(I38104),.A(g28367));
  NOT NOT1_12061(.VSS(VSS),.VDD(VDD),.Y(g29105),.A(I38104));
  NOT NOT1_12062(.VSS(VSS),.VDD(VDD),.Y(I38107),.A(g28368));
  NOT NOT1_12063(.VSS(VSS),.VDD(VDD),.Y(g29106),.A(I38107));
  NOT NOT1_12064(.VSS(VSS),.VDD(VDD),.Y(I38111),.A(g28371));
  NOT NOT1_12065(.VSS(VSS),.VDD(VDD),.Y(g29108),.A(I38111));
  NOT NOT1_12066(.VSS(VSS),.VDD(VDD),.Y(I38119),.A(g28420));
  NOT NOT1_12067(.VSS(VSS),.VDD(VDD),.Y(g29117),.A(I38119));
  NOT NOT1_12068(.VSS(VSS),.VDD(VDD),.Y(I38122),.A(g28421));
  NOT NOT1_12069(.VSS(VSS),.VDD(VDD),.Y(g29118),.A(I38122));
  NOT NOT1_12070(.VSS(VSS),.VDD(VDD),.Y(I38125),.A(g28425));
  NOT NOT1_12071(.VSS(VSS),.VDD(VDD),.Y(g29119),.A(I38125));
  NOT NOT1_12072(.VSS(VSS),.VDD(VDD),.Y(I38128),.A(g28419));
  NOT NOT1_12073(.VSS(VSS),.VDD(VDD),.Y(g29120),.A(I38128));
  NOT NOT1_12074(.VSS(VSS),.VDD(VDD),.Y(I38136),.A(g28833));
  NOT NOT1_12075(.VSS(VSS),.VDD(VDD),.Y(g29131),.A(I38136));
  NOT NOT1_12076(.VSS(VSS),.VDD(VDD),.Y(I38139),.A(g29061));
  NOT NOT1_12077(.VSS(VSS),.VDD(VDD),.Y(g29132),.A(I38139));
  NOT NOT1_12078(.VSS(VSS),.VDD(VDD),.Y(I38142),.A(g29073));
  NOT NOT1_12079(.VSS(VSS),.VDD(VDD),.Y(g29133),.A(I38142));
  NOT NOT1_12080(.VSS(VSS),.VDD(VDD),.Y(I38145),.A(g29081));
  NOT NOT1_12081(.VSS(VSS),.VDD(VDD),.Y(g29134),.A(I38145));
  NOT NOT1_12082(.VSS(VSS),.VDD(VDD),.Y(I38148),.A(g29074));
  NOT NOT1_12083(.VSS(VSS),.VDD(VDD),.Y(g29135),.A(I38148));
  NOT NOT1_12084(.VSS(VSS),.VDD(VDD),.Y(I38151),.A(g29082));
  NOT NOT1_12085(.VSS(VSS),.VDD(VDD),.Y(g29136),.A(I38151));
  NOT NOT1_12086(.VSS(VSS),.VDD(VDD),.Y(I38154),.A(g29089));
  NOT NOT1_12087(.VSS(VSS),.VDD(VDD),.Y(g29137),.A(I38154));
  NOT NOT1_12088(.VSS(VSS),.VDD(VDD),.Y(I38157),.A(g28882));
  NOT NOT1_12089(.VSS(VSS),.VDD(VDD),.Y(g29138),.A(I38157));
  NOT NOT1_12090(.VSS(VSS),.VDD(VDD),.Y(I38160),.A(g28835));
  NOT NOT1_12091(.VSS(VSS),.VDD(VDD),.Y(g29139),.A(I38160));
  NOT NOT1_12092(.VSS(VSS),.VDD(VDD),.Y(I38163),.A(g29075));
  NOT NOT1_12093(.VSS(VSS),.VDD(VDD),.Y(g29140),.A(I38163));
  NOT NOT1_12094(.VSS(VSS),.VDD(VDD),.Y(I38166),.A(g29084));
  NOT NOT1_12095(.VSS(VSS),.VDD(VDD),.Y(g29141),.A(I38166));
  NOT NOT1_12096(.VSS(VSS),.VDD(VDD),.Y(I38169),.A(g29091));
  NOT NOT1_12097(.VSS(VSS),.VDD(VDD),.Y(g29142),.A(I38169));
  NOT NOT1_12098(.VSS(VSS),.VDD(VDD),.Y(I38172),.A(g29085));
  NOT NOT1_12099(.VSS(VSS),.VDD(VDD),.Y(g29143),.A(I38172));
  NOT NOT1_12100(.VSS(VSS),.VDD(VDD),.Y(I38175),.A(g29092));
  NOT NOT1_12101(.VSS(VSS),.VDD(VDD),.Y(g29144),.A(I38175));
  NOT NOT1_12102(.VSS(VSS),.VDD(VDD),.Y(I38178),.A(g29098));
  NOT NOT1_12103(.VSS(VSS),.VDD(VDD),.Y(g29145),.A(I38178));
  NOT NOT1_12104(.VSS(VSS),.VDD(VDD),.Y(I38181),.A(g28899));
  NOT NOT1_12105(.VSS(VSS),.VDD(VDD),.Y(g29146),.A(I38181));
  NOT NOT1_12106(.VSS(VSS),.VDD(VDD),.Y(I38184),.A(g28837));
  NOT NOT1_12107(.VSS(VSS),.VDD(VDD),.Y(g29147),.A(I38184));
  NOT NOT1_12108(.VSS(VSS),.VDD(VDD),.Y(I38187),.A(g29086));
  NOT NOT1_12109(.VSS(VSS),.VDD(VDD),.Y(g29148),.A(I38187));
  NOT NOT1_12110(.VSS(VSS),.VDD(VDD),.Y(I38190),.A(g29093));
  NOT NOT1_12111(.VSS(VSS),.VDD(VDD),.Y(g29149),.A(I38190));
  NOT NOT1_12112(.VSS(VSS),.VDD(VDD),.Y(I38193),.A(g29099));
  NOT NOT1_12113(.VSS(VSS),.VDD(VDD),.Y(g29150),.A(I38193));
  NOT NOT1_12114(.VSS(VSS),.VDD(VDD),.Y(I38196),.A(g29094));
  NOT NOT1_12115(.VSS(VSS),.VDD(VDD),.Y(g29151),.A(I38196));
  NOT NOT1_12116(.VSS(VSS),.VDD(VDD),.Y(I38199),.A(g29100));
  NOT NOT1_12117(.VSS(VSS),.VDD(VDD),.Y(g29152),.A(I38199));
  NOT NOT1_12118(.VSS(VSS),.VDD(VDD),.Y(I38202),.A(g29104));
  NOT NOT1_12119(.VSS(VSS),.VDD(VDD),.Y(g29153),.A(I38202));
  NOT NOT1_12120(.VSS(VSS),.VDD(VDD),.Y(I38205),.A(g28924));
  NOT NOT1_12121(.VSS(VSS),.VDD(VDD),.Y(g29154),.A(I38205));
  NOT NOT1_12122(.VSS(VSS),.VDD(VDD),.Y(I38208),.A(g28839));
  NOT NOT1_12123(.VSS(VSS),.VDD(VDD),.Y(g29155),.A(I38208));
  NOT NOT1_12124(.VSS(VSS),.VDD(VDD),.Y(I38211),.A(g29095));
  NOT NOT1_12125(.VSS(VSS),.VDD(VDD),.Y(g29156),.A(I38211));
  NOT NOT1_12126(.VSS(VSS),.VDD(VDD),.Y(I38214),.A(g29101));
  NOT NOT1_12127(.VSS(VSS),.VDD(VDD),.Y(g29157),.A(I38214));
  NOT NOT1_12128(.VSS(VSS),.VDD(VDD),.Y(I38217),.A(g29105));
  NOT NOT1_12129(.VSS(VSS),.VDD(VDD),.Y(g29158),.A(I38217));
  NOT NOT1_12130(.VSS(VSS),.VDD(VDD),.Y(I38220),.A(g29102));
  NOT NOT1_12131(.VSS(VSS),.VDD(VDD),.Y(g29159),.A(I38220));
  NOT NOT1_12132(.VSS(VSS),.VDD(VDD),.Y(I38223),.A(g29106));
  NOT NOT1_12133(.VSS(VSS),.VDD(VDD),.Y(g29160),.A(I38223));
  NOT NOT1_12134(.VSS(VSS),.VDD(VDD),.Y(I38226),.A(g29108));
  NOT NOT1_12135(.VSS(VSS),.VDD(VDD),.Y(g29161),.A(I38226));
  NOT NOT1_12136(.VSS(VSS),.VDD(VDD),.Y(I38229),.A(g28950));
  NOT NOT1_12137(.VSS(VSS),.VDD(VDD),.Y(g29162),.A(I38229));
  NOT NOT1_12138(.VSS(VSS),.VDD(VDD),.Y(I38232),.A(g29117));
  NOT NOT1_12139(.VSS(VSS),.VDD(VDD),.Y(g29163),.A(I38232));
  NOT NOT1_12140(.VSS(VSS),.VDD(VDD),.Y(I38235),.A(g29118));
  NOT NOT1_12141(.VSS(VSS),.VDD(VDD),.Y(g29164),.A(I38235));
  NOT NOT1_12142(.VSS(VSS),.VDD(VDD),.Y(I38238),.A(g29119));
  NOT NOT1_12143(.VSS(VSS),.VDD(VDD),.Y(g29165),.A(I38238));
  NOT NOT1_12144(.VSS(VSS),.VDD(VDD),.Y(I38241),.A(g28832));
  NOT NOT1_12145(.VSS(VSS),.VDD(VDD),.Y(g29166),.A(I38241));
  NOT NOT1_12146(.VSS(VSS),.VDD(VDD),.Y(I38245),.A(g28920));
  NOT NOT1_12147(.VSS(VSS),.VDD(VDD),.Y(g29168),.A(I38245));
  NOT NOT1_12148(.VSS(VSS),.VDD(VDD),.Y(I38250),.A(g28941));
  NOT NOT1_12149(.VSS(VSS),.VDD(VDD),.Y(g29171),.A(I38250));
  NOT NOT1_12150(.VSS(VSS),.VDD(VDD),.Y(I38258),.A(g28963));
  NOT NOT1_12151(.VSS(VSS),.VDD(VDD),.Y(g29177),.A(I38258));
  NOT NOT1_12152(.VSS(VSS),.VDD(VDD),.Y(I38272),.A(g29013));
  NOT NOT1_12153(.VSS(VSS),.VDD(VDD),.Y(g29189),.A(I38272));
  NOT NOT1_12154(.VSS(VSS),.VDD(VDD),.Y(I38275),.A(g28987));
  NOT NOT1_12155(.VSS(VSS),.VDD(VDD),.Y(g29190),.A(I38275));
  NOT NOT1_12156(.VSS(VSS),.VDD(VDD),.Y(I38278),.A(g28963));
  NOT NOT1_12157(.VSS(VSS),.VDD(VDD),.Y(g29191),.A(I38278));
  NOT NOT1_12158(.VSS(VSS),.VDD(VDD),.Y(g29192),.A(g28954));
  NOT NOT1_12159(.VSS(VSS),.VDD(VDD),.Y(I38282),.A(g28941));
  NOT NOT1_12160(.VSS(VSS),.VDD(VDD),.Y(g29193),.A(I38282));
  NOT NOT1_12161(.VSS(VSS),.VDD(VDD),.Y(I38321),.A(g29113));
  NOT NOT1_12162(.VSS(VSS),.VDD(VDD),.Y(g29230),.A(I38321));
  NOT NOT1_12163(.VSS(VSS),.VDD(VDD),.Y(I38330),.A(g29120));
  NOT NOT1_12164(.VSS(VSS),.VDD(VDD),.Y(g29237),.A(I38330));
  NOT NOT1_12165(.VSS(VSS),.VDD(VDD),.Y(I38339),.A(g29120));
  NOT NOT1_12166(.VSS(VSS),.VDD(VDD),.Y(g29244),.A(I38339));
  NOT NOT1_12167(.VSS(VSS),.VDD(VDD),.Y(I38342),.A(g28886));
  NOT NOT1_12168(.VSS(VSS),.VDD(VDD),.Y(g29245),.A(I38342));
  NOT NOT1_12169(.VSS(VSS),.VDD(VDD),.Y(I38345),.A(g29109));
  NOT NOT1_12170(.VSS(VSS),.VDD(VDD),.Y(g29246),.A(I38345));
  NOT NOT1_12171(.VSS(VSS),.VDD(VDD),.Y(I38348),.A(g28874));
  NOT NOT1_12172(.VSS(VSS),.VDD(VDD),.Y(g29247),.A(I38348));
  NOT NOT1_12173(.VSS(VSS),.VDD(VDD),.Y(I38352),.A(g29110));
  NOT NOT1_12174(.VSS(VSS),.VDD(VDD),.Y(g29249),.A(I38352));
  NOT NOT1_12175(.VSS(VSS),.VDD(VDD),.Y(I38355),.A(g29039));
  NOT NOT1_12176(.VSS(VSS),.VDD(VDD),.Y(g29250),.A(I38355));
  NOT NOT1_12177(.VSS(VSS),.VDD(VDD),.Y(I38360),.A(g29111));
  NOT NOT1_12178(.VSS(VSS),.VDD(VDD),.Y(g29253),.A(I38360));
  NOT NOT1_12179(.VSS(VSS),.VDD(VDD),.Y(I38363),.A(g29016));
  NOT NOT1_12180(.VSS(VSS),.VDD(VDD),.Y(g29254),.A(I38363));
  NOT NOT1_12181(.VSS(VSS),.VDD(VDD),.Y(I38369),.A(g29112));
  NOT NOT1_12182(.VSS(VSS),.VDD(VDD),.Y(g29258),.A(I38369));
  NOT NOT1_12183(.VSS(VSS),.VDD(VDD),.Y(g29266),.A(g28741));
  NOT NOT1_12184(.VSS(VSS),.VDD(VDD),.Y(I38386),.A(g28734));
  NOT NOT1_12185(.VSS(VSS),.VDD(VDD),.Y(g29267),.A(I38386));
  NOT NOT1_12186(.VSS(VSS),.VDD(VDD),.Y(g29268),.A(g28751));
  NOT NOT1_12187(.VSS(VSS),.VDD(VDD),.Y(g29269),.A(g28755));
  NOT NOT1_12188(.VSS(VSS),.VDD(VDD),.Y(I38391),.A(g28730));
  NOT NOT1_12189(.VSS(VSS),.VDD(VDD),.Y(g29270),.A(I38391));
  NOT NOT1_12190(.VSS(VSS),.VDD(VDD),.Y(g29271),.A(g28764));
  NOT NOT1_12191(.VSS(VSS),.VDD(VDD),.Y(g29272),.A(g28768));
  NOT NOT1_12192(.VSS(VSS),.VDD(VDD),.Y(I38396),.A(g28727));
  NOT NOT1_12193(.VSS(VSS),.VDD(VDD),.Y(g29273),.A(I38396));
  NOT NOT1_12194(.VSS(VSS),.VDD(VDD),.Y(g29274),.A(g28775));
  NOT NOT1_12195(.VSS(VSS),.VDD(VDD),.Y(g29275),.A(g28779));
  NOT NOT1_12196(.VSS(VSS),.VDD(VDD),.Y(I38401),.A(g28725));
  NOT NOT1_12197(.VSS(VSS),.VDD(VDD),.Y(g29276),.A(I38401));
  NOT NOT1_12198(.VSS(VSS),.VDD(VDD),.Y(g29277),.A(g28785));
  NOT NOT1_12199(.VSS(VSS),.VDD(VDD),.Y(I38405),.A(g28723));
  NOT NOT1_12200(.VSS(VSS),.VDD(VDD),.Y(g29278),.A(I38405));
  NOT NOT1_12201(.VSS(VSS),.VDD(VDD),.Y(I38408),.A(g28721));
  NOT NOT1_12202(.VSS(VSS),.VDD(VDD),.Y(g29279),.A(I38408));
  NOT NOT1_12203(.VSS(VSS),.VDD(VDD),.Y(g29280),.A(g28791));
  NOT NOT1_12204(.VSS(VSS),.VDD(VDD),.Y(I38412),.A(g28720));
  NOT NOT1_12205(.VSS(VSS),.VDD(VDD),.Y(g29281),.A(I38412));
  NOT NOT1_12206(.VSS(VSS),.VDD(VDD),.Y(g29282),.A(g28796));
  NOT NOT1_12207(.VSS(VSS),.VDD(VDD),.Y(g29283),.A(g28799));
  NOT NOT1_12208(.VSS(VSS),.VDD(VDD),.Y(g29285),.A(g28804));
  NOT NOT1_12209(.VSS(VSS),.VDD(VDD),.Y(g29286),.A(g28807));
  NOT NOT1_12210(.VSS(VSS),.VDD(VDD),.Y(g29287),.A(g28810));
  NOT NOT1_12211(.VSS(VSS),.VDD(VDD),.Y(I38421),.A(g28740));
  NOT NOT1_12212(.VSS(VSS),.VDD(VDD),.Y(g29288),.A(I38421));
  NOT NOT1_12213(.VSS(VSS),.VDD(VDD),.Y(g29290),.A(g28814));
  NOT NOT1_12214(.VSS(VSS),.VDD(VDD),.Y(g29291),.A(g28817));
  NOT NOT1_12215(.VSS(VSS),.VDD(VDD),.Y(g29292),.A(g28820));
  NOT NOT1_12216(.VSS(VSS),.VDD(VDD),.Y(I38428),.A(g28732));
  NOT NOT1_12217(.VSS(VSS),.VDD(VDD),.Y(g29293),.A(I38428));
  NOT NOT1_12218(.VSS(VSS),.VDD(VDD),.Y(g29295),.A(g28823));
  NOT NOT1_12219(.VSS(VSS),.VDD(VDD),.Y(g29296),.A(g28826));
  NOT NOT1_12220(.VSS(VSS),.VDD(VDD),.Y(I38434),.A(g28735));
  NOT NOT1_12221(.VSS(VSS),.VDD(VDD),.Y(g29297),.A(I38434));
  NOT NOT1_12222(.VSS(VSS),.VDD(VDD),.Y(I38437),.A(g28736));
  NOT NOT1_12223(.VSS(VSS),.VDD(VDD),.Y(g29298),.A(I38437));
  NOT NOT1_12224(.VSS(VSS),.VDD(VDD),.Y(I38440),.A(g28738));
  NOT NOT1_12225(.VSS(VSS),.VDD(VDD),.Y(g29299),.A(I38440));
  NOT NOT1_12226(.VSS(VSS),.VDD(VDD),.Y(g29301),.A(g28829));
  NOT NOT1_12227(.VSS(VSS),.VDD(VDD),.Y(I38447),.A(g28744));
  NOT NOT1_12228(.VSS(VSS),.VDD(VDD),.Y(g29304),.A(I38447));
  NOT NOT1_12229(.VSS(VSS),.VDD(VDD),.Y(I38450),.A(g28745));
  NOT NOT1_12230(.VSS(VSS),.VDD(VDD),.Y(g29305),.A(I38450));
  NOT NOT1_12231(.VSS(VSS),.VDD(VDD),.Y(I38453),.A(g28746));
  NOT NOT1_12232(.VSS(VSS),.VDD(VDD),.Y(g29306),.A(I38453));
  NOT NOT1_12233(.VSS(VSS),.VDD(VDD),.Y(I38456),.A(g28747));
  NOT NOT1_12234(.VSS(VSS),.VDD(VDD),.Y(g29307),.A(I38456));
  NOT NOT1_12235(.VSS(VSS),.VDD(VDD),.Y(I38459),.A(g28749));
  NOT NOT1_12236(.VSS(VSS),.VDD(VDD),.Y(g29308),.A(I38459));
  NOT NOT1_12237(.VSS(VSS),.VDD(VDD),.Y(I38462),.A(g29120));
  NOT NOT1_12238(.VSS(VSS),.VDD(VDD),.Y(g29309),.A(I38462));
  NOT NOT1_12239(.VSS(VSS),.VDD(VDD),.Y(I38466),.A(g28754));
  NOT NOT1_12240(.VSS(VSS),.VDD(VDD),.Y(g29311),.A(I38466));
  NOT NOT1_12241(.VSS(VSS),.VDD(VDD),.Y(I38471),.A(g28758));
  NOT NOT1_12242(.VSS(VSS),.VDD(VDD),.Y(g29314),.A(I38471));
  NOT NOT1_12243(.VSS(VSS),.VDD(VDD),.Y(I38474),.A(g28759));
  NOT NOT1_12244(.VSS(VSS),.VDD(VDD),.Y(g29315),.A(I38474));
  NOT NOT1_12245(.VSS(VSS),.VDD(VDD),.Y(I38477),.A(g28760));
  NOT NOT1_12246(.VSS(VSS),.VDD(VDD),.Y(g29316),.A(I38477));
  NOT NOT1_12247(.VSS(VSS),.VDD(VDD),.Y(I38480),.A(g28761));
  NOT NOT1_12248(.VSS(VSS),.VDD(VDD),.Y(g29317),.A(I38480));
  NOT NOT1_12249(.VSS(VSS),.VDD(VDD),.Y(I38483),.A(g28990));
  NOT NOT1_12250(.VSS(VSS),.VDD(VDD),.Y(g29318),.A(I38483));
  NOT NOT1_12251(.VSS(VSS),.VDD(VDD),.Y(I38486),.A(g28763));
  NOT NOT1_12252(.VSS(VSS),.VDD(VDD),.Y(g29319),.A(I38486));
  NOT NOT1_12253(.VSS(VSS),.VDD(VDD),.Y(I38491),.A(g28767));
  NOT NOT1_12254(.VSS(VSS),.VDD(VDD),.Y(g29322),.A(I38491));
  NOT NOT1_12255(.VSS(VSS),.VDD(VDD),.Y(I38496),.A(g28771));
  NOT NOT1_12256(.VSS(VSS),.VDD(VDD),.Y(g29325),.A(I38496));
  NOT NOT1_12257(.VSS(VSS),.VDD(VDD),.Y(I38499),.A(g28772));
  NOT NOT1_12258(.VSS(VSS),.VDD(VDD),.Y(g29326),.A(I38499));
  NOT NOT1_12259(.VSS(VSS),.VDD(VDD),.Y(I38502),.A(g28773));
  NOT NOT1_12260(.VSS(VSS),.VDD(VDD),.Y(g29327),.A(I38502));
  NOT NOT1_12261(.VSS(VSS),.VDD(VDD),.Y(I38505),.A(g28774));
  NOT NOT1_12262(.VSS(VSS),.VDD(VDD),.Y(g29328),.A(I38505));
  NOT NOT1_12263(.VSS(VSS),.VDD(VDD),.Y(I38510),.A(g28778));
  NOT NOT1_12264(.VSS(VSS),.VDD(VDD),.Y(g29331),.A(I38510));
  NOT NOT1_12265(.VSS(VSS),.VDD(VDD),.Y(I38515),.A(g28782));
  NOT NOT1_12266(.VSS(VSS),.VDD(VDD),.Y(g29334),.A(I38515));
  NOT NOT1_12267(.VSS(VSS),.VDD(VDD),.Y(I38518),.A(g28783));
  NOT NOT1_12268(.VSS(VSS),.VDD(VDD),.Y(g29335),.A(I38518));
  NOT NOT1_12269(.VSS(VSS),.VDD(VDD),.Y(I38524),.A(g28788));
  NOT NOT1_12270(.VSS(VSS),.VDD(VDD),.Y(g29339),.A(I38524));
  NOT NOT1_12271(.VSS(VSS),.VDD(VDD),.Y(I38536),.A(g28920));
  NOT NOT1_12272(.VSS(VSS),.VDD(VDD),.Y(g29349),.A(I38536));
  NOT NOT1_12273(.VSS(VSS),.VDD(VDD),.Y(I38539),.A(g29113));
  NOT NOT1_12274(.VSS(VSS),.VDD(VDD),.Y(g29350),.A(I38539));
  NOT NOT1_12275(.VSS(VSS),.VDD(VDD),.Y(g29356),.A(g29120));
  NOT NOT1_12276(.VSS(VSS),.VDD(VDD),.Y(g29358),.A(g29120));
  NOT NOT1_12277(.VSS(VSS),.VDD(VDD),.Y(I38548),.A(g28903));
  NOT NOT1_12278(.VSS(VSS),.VDD(VDD),.Y(g29359),.A(I38548));
  NOT NOT1_12279(.VSS(VSS),.VDD(VDD),.Y(g29360),.A(g28871));
  NOT NOT1_12280(.VSS(VSS),.VDD(VDD),.Y(g29361),.A(g28877));
  NOT NOT1_12281(.VSS(VSS),.VDD(VDD),.Y(g29362),.A(g28883));
  NOT NOT1_12282(.VSS(VSS),.VDD(VDD),.Y(g29363),.A(g28889));
  NOT NOT1_12283(.VSS(VSS),.VDD(VDD),.Y(g29364),.A(g28894));
  NOT NOT1_12284(.VSS(VSS),.VDD(VDD),.Y(g29365),.A(g28900));
  NOT NOT1_12285(.VSS(VSS),.VDD(VDD),.Y(g29366),.A(g28906));
  NOT NOT1_12286(.VSS(VSS),.VDD(VDD),.Y(g29367),.A(g28911));
  NOT NOT1_12287(.VSS(VSS),.VDD(VDD),.Y(g29368),.A(g28916));
  NOT NOT1_12288(.VSS(VSS),.VDD(VDD),.Y(g29369),.A(g28925));
  NOT NOT1_12289(.VSS(VSS),.VDD(VDD),.Y(g29370),.A(g28928));
  NOT NOT1_12290(.VSS(VSS),.VDD(VDD),.Y(g29371),.A(g28932));
  NOT NOT1_12291(.VSS(VSS),.VDD(VDD),.Y(g29372),.A(g28937));
  NOT NOT1_12292(.VSS(VSS),.VDD(VDD),.Y(g29373),.A(g28945));
  NOT NOT1_12293(.VSS(VSS),.VDD(VDD),.Y(g29374),.A(g28951));
  NOT NOT1_12294(.VSS(VSS),.VDD(VDD),.Y(g29375),.A(g28955));
  NOT NOT1_12295(.VSS(VSS),.VDD(VDD),.Y(g29376),.A(g28959));
  NOT NOT1_12296(.VSS(VSS),.VDD(VDD),.Y(g29377),.A(g28967));
  NOT NOT1_12297(.VSS(VSS),.VDD(VDD),.Y(g29378),.A(g28972));
  NOT NOT1_12298(.VSS(VSS),.VDD(VDD),.Y(g29379),.A(g28975));
  NOT NOT1_12299(.VSS(VSS),.VDD(VDD),.Y(g29380),.A(g28979));
  NOT NOT1_12300(.VSS(VSS),.VDD(VDD),.Y(g29381),.A(g28983));
  NOT NOT1_12301(.VSS(VSS),.VDD(VDD),.Y(g29382),.A(g28993));
  NOT NOT1_12302(.VSS(VSS),.VDD(VDD),.Y(g29383),.A(g28998));
  NOT NOT1_12303(.VSS(VSS),.VDD(VDD),.Y(g29384),.A(g29002));
  NOT NOT1_12304(.VSS(VSS),.VDD(VDD),.Y(g29385),.A(g29005));
  NOT NOT1_12305(.VSS(VSS),.VDD(VDD),.Y(g29386),.A(g29010));
  NOT NOT1_12306(.VSS(VSS),.VDD(VDD),.Y(g29387),.A(g29019));
  NOT NOT1_12307(.VSS(VSS),.VDD(VDD),.Y(g29388),.A(g29023));
  NOT NOT1_12308(.VSS(VSS),.VDD(VDD),.Y(g29389),.A(g29027));
  NOT NOT1_12309(.VSS(VSS),.VDD(VDD),.Y(g29390),.A(g29032));
  NOT NOT1_12310(.VSS(VSS),.VDD(VDD),.Y(g29391),.A(g29035));
  NOT NOT1_12311(.VSS(VSS),.VDD(VDD),.Y(g29392),.A(g29042));
  NOT NOT1_12312(.VSS(VSS),.VDD(VDD),.Y(g29393),.A(g29046));
  NOT NOT1_12313(.VSS(VSS),.VDD(VDD),.Y(g29394),.A(g29050));
  NOT NOT1_12314(.VSS(VSS),.VDD(VDD),.Y(g29395),.A(g29054));
  NOT NOT1_12315(.VSS(VSS),.VDD(VDD),.Y(g29396),.A(g29057));
  NOT NOT1_12316(.VSS(VSS),.VDD(VDD),.Y(g29397),.A(g29065));
  NOT NOT1_12317(.VSS(VSS),.VDD(VDD),.Y(g29398),.A(g29069));
  NOT NOT1_12318(.VSS(VSS),.VDD(VDD),.Y(I38591),.A(g28987));
  NOT NOT1_12319(.VSS(VSS),.VDD(VDD),.Y(g29400),.A(I38591));
  NOT NOT1_12320(.VSS(VSS),.VDD(VDD),.Y(I38594),.A(g28990));
  NOT NOT1_12321(.VSS(VSS),.VDD(VDD),.Y(g29401),.A(I38594));
  NOT NOT1_12322(.VSS(VSS),.VDD(VDD),.Y(g29402),.A(g29077));
  NOT NOT1_12323(.VSS(VSS),.VDD(VDD),.Y(I38599),.A(g29013));
  NOT NOT1_12324(.VSS(VSS),.VDD(VDD),.Y(g29404),.A(I38599));
  NOT NOT1_12325(.VSS(VSS),.VDD(VDD),.Y(I38602),.A(g29016));
  NOT NOT1_12326(.VSS(VSS),.VDD(VDD),.Y(g29405),.A(I38602));
  NOT NOT1_12327(.VSS(VSS),.VDD(VDD),.Y(I38606),.A(g29039));
  NOT NOT1_12328(.VSS(VSS),.VDD(VDD),.Y(g29407),.A(I38606));
  NOT NOT1_12329(.VSS(VSS),.VDD(VDD),.Y(I38609),.A(g28874));
  NOT NOT1_12330(.VSS(VSS),.VDD(VDD),.Y(g29408),.A(I38609));
  NOT NOT1_12331(.VSS(VSS),.VDD(VDD),.Y(I38613),.A(g28886));
  NOT NOT1_12332(.VSS(VSS),.VDD(VDD),.Y(g29410),.A(I38613));
  NOT NOT1_12333(.VSS(VSS),.VDD(VDD),.Y(I38617),.A(g28903));
  NOT NOT1_12334(.VSS(VSS),.VDD(VDD),.Y(g29412),.A(I38617));
  NOT NOT1_12335(.VSS(VSS),.VDD(VDD),.Y(I38620),.A(g29246));
  NOT NOT1_12336(.VSS(VSS),.VDD(VDD),.Y(g29413),.A(I38620));
  NOT NOT1_12337(.VSS(VSS),.VDD(VDD),.Y(I38623),.A(g29293));
  NOT NOT1_12338(.VSS(VSS),.VDD(VDD),.Y(g29414),.A(I38623));
  NOT NOT1_12339(.VSS(VSS),.VDD(VDD),.Y(I38626),.A(g29297));
  NOT NOT1_12340(.VSS(VSS),.VDD(VDD),.Y(g29415),.A(I38626));
  NOT NOT1_12341(.VSS(VSS),.VDD(VDD),.Y(I38629),.A(g29304));
  NOT NOT1_12342(.VSS(VSS),.VDD(VDD),.Y(g29416),.A(I38629));
  NOT NOT1_12343(.VSS(VSS),.VDD(VDD),.Y(I38632),.A(g29298));
  NOT NOT1_12344(.VSS(VSS),.VDD(VDD),.Y(g29417),.A(I38632));
  NOT NOT1_12345(.VSS(VSS),.VDD(VDD),.Y(I38635),.A(g29305));
  NOT NOT1_12346(.VSS(VSS),.VDD(VDD),.Y(g29418),.A(I38635));
  NOT NOT1_12347(.VSS(VSS),.VDD(VDD),.Y(I38638),.A(g29311));
  NOT NOT1_12348(.VSS(VSS),.VDD(VDD),.Y(g29419),.A(I38638));
  NOT NOT1_12349(.VSS(VSS),.VDD(VDD),.Y(I38641),.A(g29249));
  NOT NOT1_12350(.VSS(VSS),.VDD(VDD),.Y(g29420),.A(I38641));
  NOT NOT1_12351(.VSS(VSS),.VDD(VDD),.Y(I38644),.A(g29299));
  NOT NOT1_12352(.VSS(VSS),.VDD(VDD),.Y(g29421),.A(I38644));
  NOT NOT1_12353(.VSS(VSS),.VDD(VDD),.Y(I38647),.A(g29306));
  NOT NOT1_12354(.VSS(VSS),.VDD(VDD),.Y(g29422),.A(I38647));
  NOT NOT1_12355(.VSS(VSS),.VDD(VDD),.Y(I38650),.A(g29314));
  NOT NOT1_12356(.VSS(VSS),.VDD(VDD),.Y(g29423),.A(I38650));
  NOT NOT1_12357(.VSS(VSS),.VDD(VDD),.Y(I38653),.A(g29307));
  NOT NOT1_12358(.VSS(VSS),.VDD(VDD),.Y(g29424),.A(I38653));
  NOT NOT1_12359(.VSS(VSS),.VDD(VDD),.Y(I38656),.A(g29315));
  NOT NOT1_12360(.VSS(VSS),.VDD(VDD),.Y(g29425),.A(I38656));
  NOT NOT1_12361(.VSS(VSS),.VDD(VDD),.Y(I38659),.A(g29322));
  NOT NOT1_12362(.VSS(VSS),.VDD(VDD),.Y(g29426),.A(I38659));
  NOT NOT1_12363(.VSS(VSS),.VDD(VDD),.Y(I38662),.A(g29253));
  NOT NOT1_12364(.VSS(VSS),.VDD(VDD),.Y(g29427),.A(I38662));
  NOT NOT1_12365(.VSS(VSS),.VDD(VDD),.Y(I38665),.A(g29412));
  NOT NOT1_12366(.VSS(VSS),.VDD(VDD),.Y(g29428),.A(I38665));
  NOT NOT1_12367(.VSS(VSS),.VDD(VDD),.Y(I38668),.A(g29168));
  NOT NOT1_12368(.VSS(VSS),.VDD(VDD),.Y(g29429),.A(I38668));
  NOT NOT1_12369(.VSS(VSS),.VDD(VDD),.Y(I38671),.A(g29171));
  NOT NOT1_12370(.VSS(VSS),.VDD(VDD),.Y(g29430),.A(I38671));
  NOT NOT1_12371(.VSS(VSS),.VDD(VDD),.Y(I38674),.A(g29177));
  NOT NOT1_12372(.VSS(VSS),.VDD(VDD),.Y(g29431),.A(I38674));
  NOT NOT1_12373(.VSS(VSS),.VDD(VDD),.Y(I38677),.A(g29400));
  NOT NOT1_12374(.VSS(VSS),.VDD(VDD),.Y(g29432),.A(I38677));
  NOT NOT1_12375(.VSS(VSS),.VDD(VDD),.Y(I38680),.A(g29404));
  NOT NOT1_12376(.VSS(VSS),.VDD(VDD),.Y(g29433),.A(I38680));
  NOT NOT1_12377(.VSS(VSS),.VDD(VDD),.Y(I38683),.A(g29308));
  NOT NOT1_12378(.VSS(VSS),.VDD(VDD),.Y(g29434),.A(I38683));
  NOT NOT1_12379(.VSS(VSS),.VDD(VDD),.Y(I38686),.A(g29316));
  NOT NOT1_12380(.VSS(VSS),.VDD(VDD),.Y(g29435),.A(I38686));
  NOT NOT1_12381(.VSS(VSS),.VDD(VDD),.Y(I38689),.A(g29325));
  NOT NOT1_12382(.VSS(VSS),.VDD(VDD),.Y(g29436),.A(I38689));
  NOT NOT1_12383(.VSS(VSS),.VDD(VDD),.Y(I38692),.A(g29317));
  NOT NOT1_12384(.VSS(VSS),.VDD(VDD),.Y(g29437),.A(I38692));
  NOT NOT1_12385(.VSS(VSS),.VDD(VDD),.Y(I38695),.A(g29326));
  NOT NOT1_12386(.VSS(VSS),.VDD(VDD),.Y(g29438),.A(I38695));
  NOT NOT1_12387(.VSS(VSS),.VDD(VDD),.Y(I38698),.A(g29331));
  NOT NOT1_12388(.VSS(VSS),.VDD(VDD),.Y(g29439),.A(I38698));
  NOT NOT1_12389(.VSS(VSS),.VDD(VDD),.Y(I38701),.A(g29401));
  NOT NOT1_12390(.VSS(VSS),.VDD(VDD),.Y(g29440),.A(I38701));
  NOT NOT1_12391(.VSS(VSS),.VDD(VDD),.Y(I38704),.A(g29405));
  NOT NOT1_12392(.VSS(VSS),.VDD(VDD),.Y(g29441),.A(I38704));
  NOT NOT1_12393(.VSS(VSS),.VDD(VDD),.Y(I38707),.A(g29407));
  NOT NOT1_12394(.VSS(VSS),.VDD(VDD),.Y(g29442),.A(I38707));
  NOT NOT1_12395(.VSS(VSS),.VDD(VDD),.Y(I38710),.A(g29408));
  NOT NOT1_12396(.VSS(VSS),.VDD(VDD),.Y(g29443),.A(I38710));
  NOT NOT1_12397(.VSS(VSS),.VDD(VDD),.Y(I38713),.A(g29410));
  NOT NOT1_12398(.VSS(VSS),.VDD(VDD),.Y(g29444),.A(I38713));
  NOT NOT1_12399(.VSS(VSS),.VDD(VDD),.Y(I38716),.A(g29230));
  NOT NOT1_12400(.VSS(VSS),.VDD(VDD),.Y(g29445),.A(I38716));
  NOT NOT1_12401(.VSS(VSS),.VDD(VDD),.Y(I38719),.A(g29258));
  NOT NOT1_12402(.VSS(VSS),.VDD(VDD),.Y(g29446),.A(I38719));
  NOT NOT1_12403(.VSS(VSS),.VDD(VDD),.Y(I38722),.A(g29319));
  NOT NOT1_12404(.VSS(VSS),.VDD(VDD),.Y(g29447),.A(I38722));
  NOT NOT1_12405(.VSS(VSS),.VDD(VDD),.Y(I38725),.A(g29327));
  NOT NOT1_12406(.VSS(VSS),.VDD(VDD),.Y(g29448),.A(I38725));
  NOT NOT1_12407(.VSS(VSS),.VDD(VDD),.Y(I38728),.A(g29334));
  NOT NOT1_12408(.VSS(VSS),.VDD(VDD),.Y(g29449),.A(I38728));
  NOT NOT1_12409(.VSS(VSS),.VDD(VDD),.Y(I38731),.A(g29328));
  NOT NOT1_12410(.VSS(VSS),.VDD(VDD),.Y(g29450),.A(I38731));
  NOT NOT1_12411(.VSS(VSS),.VDD(VDD),.Y(I38734),.A(g29335));
  NOT NOT1_12412(.VSS(VSS),.VDD(VDD),.Y(g29451),.A(I38734));
  NOT NOT1_12413(.VSS(VSS),.VDD(VDD),.Y(I38737),.A(g29339));
  NOT NOT1_12414(.VSS(VSS),.VDD(VDD),.Y(g29452),.A(I38737));
  NOT NOT1_12415(.VSS(VSS),.VDD(VDD),.Y(I38740),.A(g29288));
  NOT NOT1_12416(.VSS(VSS),.VDD(VDD),.Y(g29453),.A(I38740));
  NOT NOT1_12417(.VSS(VSS),.VDD(VDD),.Y(I38743),.A(g29267));
  NOT NOT1_12418(.VSS(VSS),.VDD(VDD),.Y(g29454),.A(I38743));
  NOT NOT1_12419(.VSS(VSS),.VDD(VDD),.Y(I38746),.A(g29270));
  NOT NOT1_12420(.VSS(VSS),.VDD(VDD),.Y(g29455),.A(I38746));
  NOT NOT1_12421(.VSS(VSS),.VDD(VDD),.Y(I38749),.A(g29273));
  NOT NOT1_12422(.VSS(VSS),.VDD(VDD),.Y(g29456),.A(I38749));
  NOT NOT1_12423(.VSS(VSS),.VDD(VDD),.Y(I38752),.A(g29276));
  NOT NOT1_12424(.VSS(VSS),.VDD(VDD),.Y(g29457),.A(I38752));
  NOT NOT1_12425(.VSS(VSS),.VDD(VDD),.Y(I38755),.A(g29278));
  NOT NOT1_12426(.VSS(VSS),.VDD(VDD),.Y(g29458),.A(I38755));
  NOT NOT1_12427(.VSS(VSS),.VDD(VDD),.Y(I38758),.A(g29279));
  NOT NOT1_12428(.VSS(VSS),.VDD(VDD),.Y(g29459),.A(I38758));
  NOT NOT1_12429(.VSS(VSS),.VDD(VDD),.Y(I38761),.A(g29281));
  NOT NOT1_12430(.VSS(VSS),.VDD(VDD),.Y(g29460),.A(I38761));
  NOT NOT1_12431(.VSS(VSS),.VDD(VDD),.Y(I38764),.A(g29237));
  NOT NOT1_12432(.VSS(VSS),.VDD(VDD),.Y(g29461),.A(I38764));
  NOT NOT1_12433(.VSS(VSS),.VDD(VDD),.Y(I38767),.A(g29244));
  NOT NOT1_12434(.VSS(VSS),.VDD(VDD),.Y(g29462),.A(I38767));
  NOT NOT1_12435(.VSS(VSS),.VDD(VDD),.Y(I38770),.A(g29309));
  NOT NOT1_12436(.VSS(VSS),.VDD(VDD),.Y(g29463),.A(I38770));
  NOT NOT1_12437(.VSS(VSS),.VDD(VDD),.Y(g29491),.A(g29350));
  NOT NOT1_12438(.VSS(VSS),.VDD(VDD),.Y(I38801),.A(g29358));
  NOT NOT1_12439(.VSS(VSS),.VDD(VDD),.Y(g29495),.A(I38801));
  NOT NOT1_12440(.VSS(VSS),.VDD(VDD),.Y(I38804),.A(g29353));
  NOT NOT1_12441(.VSS(VSS),.VDD(VDD),.Y(g29496),.A(I38804));
  NOT NOT1_12442(.VSS(VSS),.VDD(VDD),.Y(I38807),.A(g29356));
  NOT NOT1_12443(.VSS(VSS),.VDD(VDD),.Y(g29497),.A(I38807));
  NOT NOT1_12444(.VSS(VSS),.VDD(VDD),.Y(I38817),.A(g29354));
  NOT NOT1_12445(.VSS(VSS),.VDD(VDD),.Y(g29499),.A(I38817));
  NOT NOT1_12446(.VSS(VSS),.VDD(VDD),.Y(I38827),.A(g29355));
  NOT NOT1_12447(.VSS(VSS),.VDD(VDD),.Y(g29501),.A(I38827));
  NOT NOT1_12448(.VSS(VSS),.VDD(VDD),.Y(I38838),.A(g29357));
  NOT NOT1_12449(.VSS(VSS),.VDD(VDD),.Y(g29504),.A(I38838));
  NOT NOT1_12450(.VSS(VSS),.VDD(VDD),.Y(I38848),.A(g29167));
  NOT NOT1_12451(.VSS(VSS),.VDD(VDD),.Y(g29506),.A(I38848));
  NOT NOT1_12452(.VSS(VSS),.VDD(VDD),.Y(I38851),.A(g29169));
  NOT NOT1_12453(.VSS(VSS),.VDD(VDD),.Y(g29507),.A(I38851));
  NOT NOT1_12454(.VSS(VSS),.VDD(VDD),.Y(I38854),.A(g29170));
  NOT NOT1_12455(.VSS(VSS),.VDD(VDD),.Y(g29508),.A(I38854));
  NOT NOT1_12456(.VSS(VSS),.VDD(VDD),.Y(I38857),.A(g29172));
  NOT NOT1_12457(.VSS(VSS),.VDD(VDD),.Y(g29509),.A(I38857));
  NOT NOT1_12458(.VSS(VSS),.VDD(VDD),.Y(I38860),.A(g29173));
  NOT NOT1_12459(.VSS(VSS),.VDD(VDD),.Y(g29510),.A(I38860));
  NOT NOT1_12460(.VSS(VSS),.VDD(VDD),.Y(I38863),.A(g29178));
  NOT NOT1_12461(.VSS(VSS),.VDD(VDD),.Y(g29511),.A(I38863));
  NOT NOT1_12462(.VSS(VSS),.VDD(VDD),.Y(I38866),.A(g29179));
  NOT NOT1_12463(.VSS(VSS),.VDD(VDD),.Y(g29512),.A(I38866));
  NOT NOT1_12464(.VSS(VSS),.VDD(VDD),.Y(I38869),.A(g29181));
  NOT NOT1_12465(.VSS(VSS),.VDD(VDD),.Y(g29513),.A(I38869));
  NOT NOT1_12466(.VSS(VSS),.VDD(VDD),.Y(I38872),.A(g29182));
  NOT NOT1_12467(.VSS(VSS),.VDD(VDD),.Y(g29514),.A(I38872));
  NOT NOT1_12468(.VSS(VSS),.VDD(VDD),.Y(I38875),.A(g29184));
  NOT NOT1_12469(.VSS(VSS),.VDD(VDD),.Y(g29515),.A(I38875));
  NOT NOT1_12470(.VSS(VSS),.VDD(VDD),.Y(I38878),.A(g29185));
  NOT NOT1_12471(.VSS(VSS),.VDD(VDD),.Y(g29516),.A(I38878));
  NOT NOT1_12472(.VSS(VSS),.VDD(VDD),.Y(I38881),.A(g29187));
  NOT NOT1_12473(.VSS(VSS),.VDD(VDD),.Y(g29517),.A(I38881));
  NOT NOT1_12474(.VSS(VSS),.VDD(VDD),.Y(I38885),.A(g29192));
  NOT NOT1_12475(.VSS(VSS),.VDD(VDD),.Y(g29519),.A(I38885));
  NOT NOT1_12476(.VSS(VSS),.VDD(VDD),.Y(I38898),.A(g29194));
  NOT NOT1_12477(.VSS(VSS),.VDD(VDD),.Y(g29530),.A(I38898));
  NOT NOT1_12478(.VSS(VSS),.VDD(VDD),.Y(I38905),.A(g29197));
  NOT NOT1_12479(.VSS(VSS),.VDD(VDD),.Y(g29535),.A(I38905));
  NOT NOT1_12480(.VSS(VSS),.VDD(VDD),.Y(I38909),.A(g29198));
  NOT NOT1_12481(.VSS(VSS),.VDD(VDD),.Y(g29537),.A(I38909));
  NOT NOT1_12482(.VSS(VSS),.VDD(VDD),.Y(I38916),.A(g29201));
  NOT NOT1_12483(.VSS(VSS),.VDD(VDD),.Y(g29542),.A(I38916));
  NOT NOT1_12484(.VSS(VSS),.VDD(VDD),.Y(I38920),.A(g29204));
  NOT NOT1_12485(.VSS(VSS),.VDD(VDD),.Y(g29544),.A(I38920));
  NOT NOT1_12486(.VSS(VSS),.VDD(VDD),.Y(I38924),.A(g29205));
  NOT NOT1_12487(.VSS(VSS),.VDD(VDD),.Y(g29546),.A(I38924));
  NOT NOT1_12488(.VSS(VSS),.VDD(VDD),.Y(I38931),.A(g29209));
  NOT NOT1_12489(.VSS(VSS),.VDD(VDD),.Y(g29551),.A(I38931));
  NOT NOT1_12490(.VSS(VSS),.VDD(VDD),.Y(I38936),.A(g29212));
  NOT NOT1_12491(.VSS(VSS),.VDD(VDD),.Y(g29554),.A(I38936));
  NOT NOT1_12492(.VSS(VSS),.VDD(VDD),.Y(I38940),.A(g29213));
  NOT NOT1_12493(.VSS(VSS),.VDD(VDD),.Y(g29556),.A(I38940));
  NOT NOT1_12494(.VSS(VSS),.VDD(VDD),.Y(I38947),.A(g29218));
  NOT NOT1_12495(.VSS(VSS),.VDD(VDD),.Y(g29561),.A(I38947));
  NOT NOT1_12496(.VSS(VSS),.VDD(VDD),.Y(I38951),.A(g29221));
  NOT NOT1_12497(.VSS(VSS),.VDD(VDD),.Y(g29563),.A(I38951));
  NOT NOT1_12498(.VSS(VSS),.VDD(VDD),.Y(I38958),.A(g29226));
  NOT NOT1_12499(.VSS(VSS),.VDD(VDD),.Y(g29568),.A(I38958));
  NOT NOT1_12500(.VSS(VSS),.VDD(VDD),.Y(I38975),.A(g29348));
  NOT NOT1_12501(.VSS(VSS),.VDD(VDD),.Y(g29583),.A(I38975));
  NOT NOT1_12502(.VSS(VSS),.VDD(VDD),.Y(I38999),.A(g29496));
  NOT NOT1_12503(.VSS(VSS),.VDD(VDD),.Y(g29627),.A(I38999));
  NOT NOT1_12504(.VSS(VSS),.VDD(VDD),.Y(I39002),.A(g29506));
  NOT NOT1_12505(.VSS(VSS),.VDD(VDD),.Y(g29628),.A(I39002));
  NOT NOT1_12506(.VSS(VSS),.VDD(VDD),.Y(I39005),.A(g29507));
  NOT NOT1_12507(.VSS(VSS),.VDD(VDD),.Y(g29629),.A(I39005));
  NOT NOT1_12508(.VSS(VSS),.VDD(VDD),.Y(I39008),.A(g29509));
  NOT NOT1_12509(.VSS(VSS),.VDD(VDD),.Y(g29630),.A(I39008));
  NOT NOT1_12510(.VSS(VSS),.VDD(VDD),.Y(I39011),.A(g29530));
  NOT NOT1_12511(.VSS(VSS),.VDD(VDD),.Y(g29631),.A(I39011));
  NOT NOT1_12512(.VSS(VSS),.VDD(VDD),.Y(I39014),.A(g29535));
  NOT NOT1_12513(.VSS(VSS),.VDD(VDD),.Y(g29632),.A(I39014));
  NOT NOT1_12514(.VSS(VSS),.VDD(VDD),.Y(I39017),.A(g29542));
  NOT NOT1_12515(.VSS(VSS),.VDD(VDD),.Y(g29633),.A(I39017));
  NOT NOT1_12516(.VSS(VSS),.VDD(VDD),.Y(I39020),.A(g29499));
  NOT NOT1_12517(.VSS(VSS),.VDD(VDD),.Y(g29634),.A(I39020));
  NOT NOT1_12518(.VSS(VSS),.VDD(VDD),.Y(I39023),.A(g29508));
  NOT NOT1_12519(.VSS(VSS),.VDD(VDD),.Y(g29635),.A(I39023));
  NOT NOT1_12520(.VSS(VSS),.VDD(VDD),.Y(I39026),.A(g29510));
  NOT NOT1_12521(.VSS(VSS),.VDD(VDD),.Y(g29636),.A(I39026));
  NOT NOT1_12522(.VSS(VSS),.VDD(VDD),.Y(I39029),.A(g29512));
  NOT NOT1_12523(.VSS(VSS),.VDD(VDD),.Y(g29637),.A(I39029));
  NOT NOT1_12524(.VSS(VSS),.VDD(VDD),.Y(I39032),.A(g29537));
  NOT NOT1_12525(.VSS(VSS),.VDD(VDD),.Y(g29638),.A(I39032));
  NOT NOT1_12526(.VSS(VSS),.VDD(VDD),.Y(I39035),.A(g29544));
  NOT NOT1_12527(.VSS(VSS),.VDD(VDD),.Y(g29639),.A(I39035));
  NOT NOT1_12528(.VSS(VSS),.VDD(VDD),.Y(I39038),.A(g29551));
  NOT NOT1_12529(.VSS(VSS),.VDD(VDD),.Y(g29640),.A(I39038));
  NOT NOT1_12530(.VSS(VSS),.VDD(VDD),.Y(I39041),.A(g29501));
  NOT NOT1_12531(.VSS(VSS),.VDD(VDD),.Y(g29641),.A(I39041));
  NOT NOT1_12532(.VSS(VSS),.VDD(VDD),.Y(I39044),.A(g29511));
  NOT NOT1_12533(.VSS(VSS),.VDD(VDD),.Y(g29642),.A(I39044));
  NOT NOT1_12534(.VSS(VSS),.VDD(VDD),.Y(I39047),.A(g29513));
  NOT NOT1_12535(.VSS(VSS),.VDD(VDD),.Y(g29643),.A(I39047));
  NOT NOT1_12536(.VSS(VSS),.VDD(VDD),.Y(I39050),.A(g29515));
  NOT NOT1_12537(.VSS(VSS),.VDD(VDD),.Y(g29644),.A(I39050));
  NOT NOT1_12538(.VSS(VSS),.VDD(VDD),.Y(I39053),.A(g29546));
  NOT NOT1_12539(.VSS(VSS),.VDD(VDD),.Y(g29645),.A(I39053));
  NOT NOT1_12540(.VSS(VSS),.VDD(VDD),.Y(I39056),.A(g29554));
  NOT NOT1_12541(.VSS(VSS),.VDD(VDD),.Y(g29646),.A(I39056));
  NOT NOT1_12542(.VSS(VSS),.VDD(VDD),.Y(I39059),.A(g29561));
  NOT NOT1_12543(.VSS(VSS),.VDD(VDD),.Y(g29647),.A(I39059));
  NOT NOT1_12544(.VSS(VSS),.VDD(VDD),.Y(I39062),.A(g29504));
  NOT NOT1_12545(.VSS(VSS),.VDD(VDD),.Y(g29648),.A(I39062));
  NOT NOT1_12546(.VSS(VSS),.VDD(VDD),.Y(I39065),.A(g29514));
  NOT NOT1_12547(.VSS(VSS),.VDD(VDD),.Y(g29649),.A(I39065));
  NOT NOT1_12548(.VSS(VSS),.VDD(VDD),.Y(I39068),.A(g29516));
  NOT NOT1_12549(.VSS(VSS),.VDD(VDD),.Y(g29650),.A(I39068));
  NOT NOT1_12550(.VSS(VSS),.VDD(VDD),.Y(I39071),.A(g29517));
  NOT NOT1_12551(.VSS(VSS),.VDD(VDD),.Y(g29651),.A(I39071));
  NOT NOT1_12552(.VSS(VSS),.VDD(VDD),.Y(I39074),.A(g29556));
  NOT NOT1_12553(.VSS(VSS),.VDD(VDD),.Y(g29652),.A(I39074));
  NOT NOT1_12554(.VSS(VSS),.VDD(VDD),.Y(I39077),.A(g29563));
  NOT NOT1_12555(.VSS(VSS),.VDD(VDD),.Y(g29653),.A(I39077));
  NOT NOT1_12556(.VSS(VSS),.VDD(VDD),.Y(I39080),.A(g29568));
  NOT NOT1_12557(.VSS(VSS),.VDD(VDD),.Y(g29654),.A(I39080));
  NOT NOT1_12558(.VSS(VSS),.VDD(VDD),.Y(I39083),.A(g29519));
  NOT NOT1_12559(.VSS(VSS),.VDD(VDD),.Y(g29655),.A(I39083));
  NOT NOT1_12560(.VSS(VSS),.VDD(VDD),.Y(I39086),.A(g29497));
  NOT NOT1_12561(.VSS(VSS),.VDD(VDD),.Y(g29656),.A(I39086));
  NOT NOT1_12562(.VSS(VSS),.VDD(VDD),.Y(I39089),.A(g29495));
  NOT NOT1_12563(.VSS(VSS),.VDD(VDD),.Y(g29657),.A(I39089));
  NOT NOT1_12564(.VSS(VSS),.VDD(VDD),.Y(g29658),.A(g29574));
  NOT NOT1_12565(.VSS(VSS),.VDD(VDD),.Y(g29659),.A(g29571));
  NOT NOT1_12566(.VSS(VSS),.VDD(VDD),.Y(g29660),.A(g29578));
  NOT NOT1_12567(.VSS(VSS),.VDD(VDD),.Y(g29661),.A(g29576));
  NOT NOT1_12568(.VSS(VSS),.VDD(VDD),.Y(g29662),.A(g29570));
  NOT NOT1_12569(.VSS(VSS),.VDD(VDD),.Y(g29664),.A(g29552));
  NOT NOT1_12570(.VSS(VSS),.VDD(VDD),.Y(g29666),.A(g29577));
  NOT NOT1_12571(.VSS(VSS),.VDD(VDD),.Y(g29668),.A(g29569));
  NOT NOT1_12572(.VSS(VSS),.VDD(VDD),.Y(g29673),.A(g29583));
  NOT NOT1_12573(.VSS(VSS),.VDD(VDD),.Y(I39121),.A(g29579));
  NOT NOT1_12574(.VSS(VSS),.VDD(VDD),.Y(g29689),.A(I39121));
  NOT NOT1_12575(.VSS(VSS),.VDD(VDD),.Y(I39124),.A(g29606));
  NOT NOT1_12576(.VSS(VSS),.VDD(VDD),.Y(g29690),.A(I39124));
  NOT NOT1_12577(.VSS(VSS),.VDD(VDD),.Y(I39127),.A(g29608));
  NOT NOT1_12578(.VSS(VSS),.VDD(VDD),.Y(g29691),.A(I39127));
  NOT NOT1_12579(.VSS(VSS),.VDD(VDD),.Y(I39130),.A(g29580));
  NOT NOT1_12580(.VSS(VSS),.VDD(VDD),.Y(g29692),.A(I39130));
  NOT NOT1_12581(.VSS(VSS),.VDD(VDD),.Y(I39133),.A(g29609));
  NOT NOT1_12582(.VSS(VSS),.VDD(VDD),.Y(g29693),.A(I39133));
  NOT NOT1_12583(.VSS(VSS),.VDD(VDD),.Y(I39136),.A(g29611));
  NOT NOT1_12584(.VSS(VSS),.VDD(VDD),.Y(g29694),.A(I39136));
  NOT NOT1_12585(.VSS(VSS),.VDD(VDD),.Y(I39139),.A(g29612));
  NOT NOT1_12586(.VSS(VSS),.VDD(VDD),.Y(g29695),.A(I39139));
  NOT NOT1_12587(.VSS(VSS),.VDD(VDD),.Y(I39142),.A(g29581));
  NOT NOT1_12588(.VSS(VSS),.VDD(VDD),.Y(g29696),.A(I39142));
  NOT NOT1_12589(.VSS(VSS),.VDD(VDD),.Y(I39145),.A(g29613));
  NOT NOT1_12590(.VSS(VSS),.VDD(VDD),.Y(g29697),.A(I39145));
  NOT NOT1_12591(.VSS(VSS),.VDD(VDD),.Y(I39148),.A(g29616));
  NOT NOT1_12592(.VSS(VSS),.VDD(VDD),.Y(g29698),.A(I39148));
  NOT NOT1_12593(.VSS(VSS),.VDD(VDD),.Y(I39151),.A(g29617));
  NOT NOT1_12594(.VSS(VSS),.VDD(VDD),.Y(g29699),.A(I39151));
  NOT NOT1_12595(.VSS(VSS),.VDD(VDD),.Y(I39154),.A(g29582));
  NOT NOT1_12596(.VSS(VSS),.VDD(VDD),.Y(g29700),.A(I39154));
  NOT NOT1_12597(.VSS(VSS),.VDD(VDD),.Y(I39157),.A(g29618));
  NOT NOT1_12598(.VSS(VSS),.VDD(VDD),.Y(g29701),.A(I39157));
  NOT NOT1_12599(.VSS(VSS),.VDD(VDD),.Y(I39160),.A(g29620));
  NOT NOT1_12600(.VSS(VSS),.VDD(VDD),.Y(g29702),.A(I39160));
  NOT NOT1_12601(.VSS(VSS),.VDD(VDD),.Y(I39164),.A(g29621));
  NOT NOT1_12602(.VSS(VSS),.VDD(VDD),.Y(g29704),.A(I39164));
  NOT NOT1_12603(.VSS(VSS),.VDD(VDD),.Y(I39168),.A(g29623));
  NOT NOT1_12604(.VSS(VSS),.VDD(VDD),.Y(g29708),.A(I39168));
  NOT NOT1_12605(.VSS(VSS),.VDD(VDD),.Y(g29716),.A(g29498));
  NOT NOT1_12606(.VSS(VSS),.VDD(VDD),.Y(g29724),.A(g29500));
  NOT NOT1_12607(.VSS(VSS),.VDD(VDD),.Y(g29726),.A(g29503));
  NOT NOT1_12608(.VSS(VSS),.VDD(VDD),.Y(g29739),.A(g29505));
  NOT NOT1_12609(.VSS(VSS),.VDD(VDD),.Y(I39234),.A(g29689));
  NOT NOT1_12610(.VSS(VSS),.VDD(VDD),.Y(g29794),.A(I39234));
  NOT NOT1_12611(.VSS(VSS),.VDD(VDD),.Y(I39237),.A(g29690));
  NOT NOT1_12612(.VSS(VSS),.VDD(VDD),.Y(g29795),.A(I39237));
  NOT NOT1_12613(.VSS(VSS),.VDD(VDD),.Y(I39240),.A(g29691));
  NOT NOT1_12614(.VSS(VSS),.VDD(VDD),.Y(g29796),.A(I39240));
  NOT NOT1_12615(.VSS(VSS),.VDD(VDD),.Y(I39243),.A(g29694));
  NOT NOT1_12616(.VSS(VSS),.VDD(VDD),.Y(g29797),.A(I39243));
  NOT NOT1_12617(.VSS(VSS),.VDD(VDD),.Y(I39246),.A(g29692));
  NOT NOT1_12618(.VSS(VSS),.VDD(VDD),.Y(g29798),.A(I39246));
  NOT NOT1_12619(.VSS(VSS),.VDD(VDD),.Y(I39249),.A(g29693));
  NOT NOT1_12620(.VSS(VSS),.VDD(VDD),.Y(g29799),.A(I39249));
  NOT NOT1_12621(.VSS(VSS),.VDD(VDD),.Y(I39252),.A(g29695));
  NOT NOT1_12622(.VSS(VSS),.VDD(VDD),.Y(g29800),.A(I39252));
  NOT NOT1_12623(.VSS(VSS),.VDD(VDD),.Y(I39255),.A(g29698));
  NOT NOT1_12624(.VSS(VSS),.VDD(VDD),.Y(g29801),.A(I39255));
  NOT NOT1_12625(.VSS(VSS),.VDD(VDD),.Y(I39258),.A(g29696));
  NOT NOT1_12626(.VSS(VSS),.VDD(VDD),.Y(g29802),.A(I39258));
  NOT NOT1_12627(.VSS(VSS),.VDD(VDD),.Y(I39261),.A(g29697));
  NOT NOT1_12628(.VSS(VSS),.VDD(VDD),.Y(g29803),.A(I39261));
  NOT NOT1_12629(.VSS(VSS),.VDD(VDD),.Y(I39264),.A(g29699));
  NOT NOT1_12630(.VSS(VSS),.VDD(VDD),.Y(g29804),.A(I39264));
  NOT NOT1_12631(.VSS(VSS),.VDD(VDD),.Y(I39267),.A(g29702));
  NOT NOT1_12632(.VSS(VSS),.VDD(VDD),.Y(g29805),.A(I39267));
  NOT NOT1_12633(.VSS(VSS),.VDD(VDD),.Y(I39270),.A(g29700));
  NOT NOT1_12634(.VSS(VSS),.VDD(VDD),.Y(g29806),.A(I39270));
  NOT NOT1_12635(.VSS(VSS),.VDD(VDD),.Y(I39273),.A(g29701));
  NOT NOT1_12636(.VSS(VSS),.VDD(VDD),.Y(g29807),.A(I39273));
  NOT NOT1_12637(.VSS(VSS),.VDD(VDD),.Y(I39276),.A(g29704));
  NOT NOT1_12638(.VSS(VSS),.VDD(VDD),.Y(g29808),.A(I39276));
  NOT NOT1_12639(.VSS(VSS),.VDD(VDD),.Y(I39279),.A(g29708));
  NOT NOT1_12640(.VSS(VSS),.VDD(VDD),.Y(g29809),.A(I39279));
  NOT NOT1_12641(.VSS(VSS),.VDD(VDD),.Y(g29823),.A(g29663));
  NOT NOT1_12642(.VSS(VSS),.VDD(VDD),.Y(g29829),.A(g29665));
  NOT NOT1_12643(.VSS(VSS),.VDD(VDD),.Y(g29835),.A(g29667));
  NOT NOT1_12644(.VSS(VSS),.VDD(VDD),.Y(g29840),.A(g29669));
  NOT NOT1_12645(.VSS(VSS),.VDD(VDD),.Y(g29844),.A(g29670));
  NOT NOT1_12646(.VSS(VSS),.VDD(VDD),.Y(g29848),.A(g29761));
  NOT NOT1_12647(.VSS(VSS),.VDD(VDD),.Y(g29849),.A(g29671));
  NOT NOT1_12648(.VSS(VSS),.VDD(VDD),.Y(g29853),.A(g29672));
  NOT NOT1_12649(.VSS(VSS),.VDD(VDD),.Y(g29857),.A(g29676));
  NOT NOT1_12650(.VSS(VSS),.VDD(VDD),.Y(g29861),.A(g29677));
  NOT NOT1_12651(.VSS(VSS),.VDD(VDD),.Y(g29865),.A(g29678));
  NOT NOT1_12652(.VSS(VSS),.VDD(VDD),.Y(g29869),.A(g29679));
  NOT NOT1_12653(.VSS(VSS),.VDD(VDD),.Y(g29873),.A(g29680));
  NOT NOT1_12654(.VSS(VSS),.VDD(VDD),.Y(g29877),.A(g29681));
  NOT NOT1_12655(.VSS(VSS),.VDD(VDD),.Y(g29881),.A(g29682));
  NOT NOT1_12656(.VSS(VSS),.VDD(VDD),.Y(g29885),.A(g29683));
  NOT NOT1_12657(.VSS(VSS),.VDD(VDD),.Y(g29889),.A(g29684));
  NOT NOT1_12658(.VSS(VSS),.VDD(VDD),.Y(g29893),.A(g29685));
  NOT NOT1_12659(.VSS(VSS),.VDD(VDD),.Y(g29897),.A(g29686));
  NOT NOT1_12660(.VSS(VSS),.VDD(VDD),.Y(g29901),.A(g29687));
  NOT NOT1_12661(.VSS(VSS),.VDD(VDD),.Y(g29905),.A(g29688));
  NOT NOT1_12662(.VSS(VSS),.VDD(VDD),.Y(I39398),.A(g29664));
  NOT NOT1_12663(.VSS(VSS),.VDD(VDD),.Y(g29932),.A(I39398));
  NOT NOT1_12664(.VSS(VSS),.VDD(VDD),.Y(I39401),.A(g29662));
  NOT NOT1_12665(.VSS(VSS),.VDD(VDD),.Y(g29933),.A(I39401));
  NOT NOT1_12666(.VSS(VSS),.VDD(VDD),.Y(I39404),.A(g29661));
  NOT NOT1_12667(.VSS(VSS),.VDD(VDD),.Y(g29934),.A(I39404));
  NOT NOT1_12668(.VSS(VSS),.VDD(VDD),.Y(I39407),.A(g29660));
  NOT NOT1_12669(.VSS(VSS),.VDD(VDD),.Y(g29935),.A(I39407));
  NOT NOT1_12670(.VSS(VSS),.VDD(VDD),.Y(I39411),.A(g29659));
  NOT NOT1_12671(.VSS(VSS),.VDD(VDD),.Y(g29937),.A(I39411));
  NOT NOT1_12672(.VSS(VSS),.VDD(VDD),.Y(I39414),.A(g29658));
  NOT NOT1_12673(.VSS(VSS),.VDD(VDD),.Y(g29938),.A(I39414));
  NOT NOT1_12674(.VSS(VSS),.VDD(VDD),.Y(I39418),.A(g29668));
  NOT NOT1_12675(.VSS(VSS),.VDD(VDD),.Y(g29940),.A(I39418));
  NOT NOT1_12676(.VSS(VSS),.VDD(VDD),.Y(I39423),.A(g29666));
  NOT NOT1_12677(.VSS(VSS),.VDD(VDD),.Y(g29943),.A(I39423));
  NOT NOT1_12678(.VSS(VSS),.VDD(VDD),.Y(I39454),.A(g29940));
  NOT NOT1_12679(.VSS(VSS),.VDD(VDD),.Y(g29972),.A(I39454));
  NOT NOT1_12680(.VSS(VSS),.VDD(VDD),.Y(I39457),.A(g29943));
  NOT NOT1_12681(.VSS(VSS),.VDD(VDD),.Y(g29973),.A(I39457));
  NOT NOT1_12682(.VSS(VSS),.VDD(VDD),.Y(I39460),.A(g29932));
  NOT NOT1_12683(.VSS(VSS),.VDD(VDD),.Y(g29974),.A(I39460));
  NOT NOT1_12684(.VSS(VSS),.VDD(VDD),.Y(I39463),.A(g29933));
  NOT NOT1_12685(.VSS(VSS),.VDD(VDD),.Y(g29975),.A(I39463));
  NOT NOT1_12686(.VSS(VSS),.VDD(VDD),.Y(I39466),.A(g29934));
  NOT NOT1_12687(.VSS(VSS),.VDD(VDD),.Y(g29976),.A(I39466));
  NOT NOT1_12688(.VSS(VSS),.VDD(VDD),.Y(I39469),.A(g29935));
  NOT NOT1_12689(.VSS(VSS),.VDD(VDD),.Y(g29977),.A(I39469));
  NOT NOT1_12690(.VSS(VSS),.VDD(VDD),.Y(I39472),.A(g29937));
  NOT NOT1_12691(.VSS(VSS),.VDD(VDD),.Y(g29978),.A(I39472));
  NOT NOT1_12692(.VSS(VSS),.VDD(VDD),.Y(I39475),.A(g29938));
  NOT NOT1_12693(.VSS(VSS),.VDD(VDD),.Y(g29979),.A(I39475));
  NOT NOT1_12694(.VSS(VSS),.VDD(VDD),.Y(g30036),.A(g29912));
  NOT NOT1_12695(.VSS(VSS),.VDD(VDD),.Y(g30040),.A(g29914));
  NOT NOT1_12696(.VSS(VSS),.VDD(VDD),.Y(g30044),.A(g29916));
  NOT NOT1_12697(.VSS(VSS),.VDD(VDD),.Y(g30048),.A(g29920));
  NOT NOT1_12698(.VSS(VSS),.VDD(VDD),.Y(I39550),.A(g29848));
  NOT NOT1_12699(.VSS(VSS),.VDD(VDD),.Y(g30052),.A(I39550));
  NOT NOT1_12700(.VSS(VSS),.VDD(VDD),.Y(I39573),.A(g29936));
  NOT NOT1_12701(.VSS(VSS),.VDD(VDD),.Y(g30076),.A(I39573));
  NOT NOT1_12702(.VSS(VSS),.VDD(VDD),.Y(I39577),.A(g29939));
  NOT NOT1_12703(.VSS(VSS),.VDD(VDD),.Y(g30078),.A(I39577));
  NOT NOT1_12704(.VSS(VSS),.VDD(VDD),.Y(I39585),.A(g29941));
  NOT NOT1_12705(.VSS(VSS),.VDD(VDD),.Y(g30084),.A(I39585));
  NOT NOT1_12706(.VSS(VSS),.VDD(VDD),.Y(I39622),.A(g30052));
  NOT NOT1_12707(.VSS(VSS),.VDD(VDD),.Y(g30119),.A(I39622));
  NOT NOT1_12708(.VSS(VSS),.VDD(VDD),.Y(I39625),.A(g30076));
  NOT NOT1_12709(.VSS(VSS),.VDD(VDD),.Y(g30120),.A(I39625));
  NOT NOT1_12710(.VSS(VSS),.VDD(VDD),.Y(I39628),.A(g30078));
  NOT NOT1_12711(.VSS(VSS),.VDD(VDD),.Y(g30121),.A(I39628));
  NOT NOT1_12712(.VSS(VSS),.VDD(VDD),.Y(I39631),.A(g30084));
  NOT NOT1_12713(.VSS(VSS),.VDD(VDD),.Y(g30122),.A(I39631));
  NOT NOT1_12714(.VSS(VSS),.VDD(VDD),.Y(I39635),.A(g30055));
  NOT NOT1_12715(.VSS(VSS),.VDD(VDD),.Y(g30124),.A(I39635));
  NOT NOT1_12716(.VSS(VSS),.VDD(VDD),.Y(I39638),.A(g30056));
  NOT NOT1_12717(.VSS(VSS),.VDD(VDD),.Y(g30125),.A(I39638));
  NOT NOT1_12718(.VSS(VSS),.VDD(VDD),.Y(I39641),.A(g30057));
  NOT NOT1_12719(.VSS(VSS),.VDD(VDD),.Y(g30126),.A(I39641));
  NOT NOT1_12720(.VSS(VSS),.VDD(VDD),.Y(I39647),.A(g30058));
  NOT NOT1_12721(.VSS(VSS),.VDD(VDD),.Y(g30130),.A(I39647));
  NOT NOT1_12722(.VSS(VSS),.VDD(VDD),.Y(g30134),.A(g30010));
  NOT NOT1_12723(.VSS(VSS),.VDD(VDD),.Y(g30139),.A(g30011));
  NOT NOT1_12724(.VSS(VSS),.VDD(VDD),.Y(g30143),.A(g30012));
  NOT NOT1_12725(.VSS(VSS),.VDD(VDD),.Y(g30147),.A(g30013));
  NOT NOT1_12726(.VSS(VSS),.VDD(VDD),.Y(g30151),.A(g30014));
  NOT NOT1_12727(.VSS(VSS),.VDD(VDD),.Y(g30155),.A(g30015));
  NOT NOT1_12728(.VSS(VSS),.VDD(VDD),.Y(g30159),.A(g30016));
  NOT NOT1_12729(.VSS(VSS),.VDD(VDD),.Y(g30163),.A(g30017));
  NOT NOT1_12730(.VSS(VSS),.VDD(VDD),.Y(g30167),.A(g30018));
  NOT NOT1_12731(.VSS(VSS),.VDD(VDD),.Y(g30171),.A(g30019));
  NOT NOT1_12732(.VSS(VSS),.VDD(VDD),.Y(g30175),.A(g30020));
  NOT NOT1_12733(.VSS(VSS),.VDD(VDD),.Y(g30179),.A(g30021));
  NOT NOT1_12734(.VSS(VSS),.VDD(VDD),.Y(g30183),.A(g30022));
  NOT NOT1_12735(.VSS(VSS),.VDD(VDD),.Y(g30187),.A(g30023));
  NOT NOT1_12736(.VSS(VSS),.VDD(VDD),.Y(g30191),.A(g30024));
  NOT NOT1_12737(.VSS(VSS),.VDD(VDD),.Y(g30195),.A(g30025));
  NOT NOT1_12738(.VSS(VSS),.VDD(VDD),.Y(g30199),.A(g30026));
  NOT NOT1_12739(.VSS(VSS),.VDD(VDD),.Y(g30203),.A(g30027));
  NOT NOT1_12740(.VSS(VSS),.VDD(VDD),.Y(g30207),.A(g30028));
  NOT NOT1_12741(.VSS(VSS),.VDD(VDD),.Y(g30211),.A(g30029));
  NOT NOT1_12742(.VSS(VSS),.VDD(VDD),.Y(I39674),.A(g30072));
  NOT NOT1_12743(.VSS(VSS),.VDD(VDD),.Y(g30215),.A(I39674));
  NOT NOT1_12744(.VSS(VSS),.VDD(VDD),.Y(g30229),.A(g30030));
  NOT NOT1_12745(.VSS(VSS),.VDD(VDD),.Y(g30233),.A(g30031));
  NOT NOT1_12746(.VSS(VSS),.VDD(VDD),.Y(g30237),.A(g30032));
  NOT NOT1_12747(.VSS(VSS),.VDD(VDD),.Y(g30241),.A(g30033));
  NOT NOT1_12748(.VSS(VSS),.VDD(VDD),.Y(I39761),.A(g30072));
  NOT NOT1_12749(.VSS(VSS),.VDD(VDD),.Y(g30306),.A(I39761));
  NOT NOT1_12750(.VSS(VSS),.VDD(VDD),.Y(I39764),.A(g30060));
  NOT NOT1_12751(.VSS(VSS),.VDD(VDD),.Y(g30307),.A(I39764));
  NOT NOT1_12752(.VSS(VSS),.VDD(VDD),.Y(I39767),.A(g30061));
  NOT NOT1_12753(.VSS(VSS),.VDD(VDD),.Y(g30308),.A(I39767));
  NOT NOT1_12754(.VSS(VSS),.VDD(VDD),.Y(I39770),.A(g30063));
  NOT NOT1_12755(.VSS(VSS),.VDD(VDD),.Y(g30309),.A(I39770));
  NOT NOT1_12756(.VSS(VSS),.VDD(VDD),.Y(I39773),.A(g30064));
  NOT NOT1_12757(.VSS(VSS),.VDD(VDD),.Y(g30310),.A(I39773));
  NOT NOT1_12758(.VSS(VSS),.VDD(VDD),.Y(I39776),.A(g30066));
  NOT NOT1_12759(.VSS(VSS),.VDD(VDD),.Y(g30311),.A(I39776));
  NOT NOT1_12760(.VSS(VSS),.VDD(VDD),.Y(I39779),.A(g30053));
  NOT NOT1_12761(.VSS(VSS),.VDD(VDD),.Y(g30312),.A(I39779));
  NOT NOT1_12762(.VSS(VSS),.VDD(VDD),.Y(I39782),.A(g30054));
  NOT NOT1_12763(.VSS(VSS),.VDD(VDD),.Y(g30313),.A(I39782));
  NOT NOT1_12764(.VSS(VSS),.VDD(VDD),.Y(I39785),.A(g30124));
  NOT NOT1_12765(.VSS(VSS),.VDD(VDD),.Y(g30314),.A(I39785));
  NOT NOT1_12766(.VSS(VSS),.VDD(VDD),.Y(I39788),.A(g30125));
  NOT NOT1_12767(.VSS(VSS),.VDD(VDD),.Y(g30315),.A(I39788));
  NOT NOT1_12768(.VSS(VSS),.VDD(VDD),.Y(I39791),.A(g30126));
  NOT NOT1_12769(.VSS(VSS),.VDD(VDD),.Y(g30316),.A(I39791));
  NOT NOT1_12770(.VSS(VSS),.VDD(VDD),.Y(I39794),.A(g30130));
  NOT NOT1_12771(.VSS(VSS),.VDD(VDD),.Y(g30317),.A(I39794));
  NOT NOT1_12772(.VSS(VSS),.VDD(VDD),.Y(I39797),.A(g30307));
  NOT NOT1_12773(.VSS(VSS),.VDD(VDD),.Y(g30318),.A(I39797));
  NOT NOT1_12774(.VSS(VSS),.VDD(VDD),.Y(I39800),.A(g30309));
  NOT NOT1_12775(.VSS(VSS),.VDD(VDD),.Y(g30319),.A(I39800));
  NOT NOT1_12776(.VSS(VSS),.VDD(VDD),.Y(I39803),.A(g30308));
  NOT NOT1_12777(.VSS(VSS),.VDD(VDD),.Y(g30320),.A(I39803));
  NOT NOT1_12778(.VSS(VSS),.VDD(VDD),.Y(I39806),.A(g30310));
  NOT NOT1_12779(.VSS(VSS),.VDD(VDD),.Y(g30321),.A(I39806));
  NOT NOT1_12780(.VSS(VSS),.VDD(VDD),.Y(I39809),.A(g30311));
  NOT NOT1_12781(.VSS(VSS),.VDD(VDD),.Y(g30322),.A(I39809));
  NOT NOT1_12782(.VSS(VSS),.VDD(VDD),.Y(I39812),.A(g30312));
  NOT NOT1_12783(.VSS(VSS),.VDD(VDD),.Y(g30323),.A(I39812));
  NOT NOT1_12784(.VSS(VSS),.VDD(VDD),.Y(I39815),.A(g30313));
  NOT NOT1_12785(.VSS(VSS),.VDD(VDD),.Y(g30324),.A(I39815));
  NOT NOT1_12786(.VSS(VSS),.VDD(VDD),.Y(I39818),.A(g30215));
  NOT NOT1_12787(.VSS(VSS),.VDD(VDD),.Y(g30325),.A(I39818));
  NOT NOT1_12788(.VSS(VSS),.VDD(VDD),.Y(I39821),.A(g30267));
  NOT NOT1_12789(.VSS(VSS),.VDD(VDD),.Y(g30326),.A(I39821));
  NOT NOT1_12790(.VSS(VSS),.VDD(VDD),.Y(I39825),.A(g30268));
  NOT NOT1_12791(.VSS(VSS),.VDD(VDD),.Y(g30328),.A(I39825));
  NOT NOT1_12792(.VSS(VSS),.VDD(VDD),.Y(I39828),.A(g30269));
  NOT NOT1_12793(.VSS(VSS),.VDD(VDD),.Y(g30329),.A(I39828));
  NOT NOT1_12794(.VSS(VSS),.VDD(VDD),.Y(I39832),.A(g30270));
  NOT NOT1_12795(.VSS(VSS),.VDD(VDD),.Y(g30331),.A(I39832));
  NOT NOT1_12796(.VSS(VSS),.VDD(VDD),.Y(I39835),.A(g30271));
  NOT NOT1_12797(.VSS(VSS),.VDD(VDD),.Y(g30332),.A(I39835));
  NOT NOT1_12798(.VSS(VSS),.VDD(VDD),.Y(I39840),.A(g30272));
  NOT NOT1_12799(.VSS(VSS),.VDD(VDD),.Y(g30335),.A(I39840));
  NOT NOT1_12800(.VSS(VSS),.VDD(VDD),.Y(I39843),.A(g30273));
  NOT NOT1_12801(.VSS(VSS),.VDD(VDD),.Y(g30336),.A(I39843));
  NOT NOT1_12802(.VSS(VSS),.VDD(VDD),.Y(I39848),.A(g30274));
  NOT NOT1_12803(.VSS(VSS),.VDD(VDD),.Y(g30339),.A(I39848));
  NOT NOT1_12804(.VSS(VSS),.VDD(VDD),.Y(I39853),.A(g30275));
  NOT NOT1_12805(.VSS(VSS),.VDD(VDD),.Y(g30342),.A(I39853));
  NOT NOT1_12806(.VSS(VSS),.VDD(VDD),.Y(I39856),.A(g30276));
  NOT NOT1_12807(.VSS(VSS),.VDD(VDD),.Y(g30343),.A(I39856));
  NOT NOT1_12808(.VSS(VSS),.VDD(VDD),.Y(I39859),.A(g30277));
  NOT NOT1_12809(.VSS(VSS),.VDD(VDD),.Y(g30344),.A(I39859));
  NOT NOT1_12810(.VSS(VSS),.VDD(VDD),.Y(I39863),.A(g30278));
  NOT NOT1_12811(.VSS(VSS),.VDD(VDD),.Y(g30346),.A(I39863));
  NOT NOT1_12812(.VSS(VSS),.VDD(VDD),.Y(I39866),.A(g30279));
  NOT NOT1_12813(.VSS(VSS),.VDD(VDD),.Y(g30347),.A(I39866));
  NOT NOT1_12814(.VSS(VSS),.VDD(VDD),.Y(I39870),.A(g30280));
  NOT NOT1_12815(.VSS(VSS),.VDD(VDD),.Y(g30349),.A(I39870));
  NOT NOT1_12816(.VSS(VSS),.VDD(VDD),.Y(I39873),.A(g30281));
  NOT NOT1_12817(.VSS(VSS),.VDD(VDD),.Y(g30350),.A(I39873));
  NOT NOT1_12818(.VSS(VSS),.VDD(VDD),.Y(I39878),.A(g30282));
  NOT NOT1_12819(.VSS(VSS),.VDD(VDD),.Y(g30353),.A(I39878));
  NOT NOT1_12820(.VSS(VSS),.VDD(VDD),.Y(I39881),.A(g30283));
  NOT NOT1_12821(.VSS(VSS),.VDD(VDD),.Y(g30354),.A(I39881));
  NOT NOT1_12822(.VSS(VSS),.VDD(VDD),.Y(I39886),.A(g30284));
  NOT NOT1_12823(.VSS(VSS),.VDD(VDD),.Y(g30357),.A(I39886));
  NOT NOT1_12824(.VSS(VSS),.VDD(VDD),.Y(I39889),.A(g30285));
  NOT NOT1_12825(.VSS(VSS),.VDD(VDD),.Y(g30358),.A(I39889));
  NOT NOT1_12826(.VSS(VSS),.VDD(VDD),.Y(I39892),.A(g30286));
  NOT NOT1_12827(.VSS(VSS),.VDD(VDD),.Y(g30359),.A(I39892));
  NOT NOT1_12828(.VSS(VSS),.VDD(VDD),.Y(I39895),.A(g30287));
  NOT NOT1_12829(.VSS(VSS),.VDD(VDD),.Y(g30360),.A(I39895));
  NOT NOT1_12830(.VSS(VSS),.VDD(VDD),.Y(I39899),.A(g30288));
  NOT NOT1_12831(.VSS(VSS),.VDD(VDD),.Y(g30362),.A(I39899));
  NOT NOT1_12832(.VSS(VSS),.VDD(VDD),.Y(I39902),.A(g30289));
  NOT NOT1_12833(.VSS(VSS),.VDD(VDD),.Y(g30363),.A(I39902));
  NOT NOT1_12834(.VSS(VSS),.VDD(VDD),.Y(I39906),.A(g30290));
  NOT NOT1_12835(.VSS(VSS),.VDD(VDD),.Y(g30365),.A(I39906));
  NOT NOT1_12836(.VSS(VSS),.VDD(VDD),.Y(I39909),.A(g30291));
  NOT NOT1_12837(.VSS(VSS),.VDD(VDD),.Y(g30366),.A(I39909));
  NOT NOT1_12838(.VSS(VSS),.VDD(VDD),.Y(I39913),.A(g30292));
  NOT NOT1_12839(.VSS(VSS),.VDD(VDD),.Y(g30368),.A(I39913));
  NOT NOT1_12840(.VSS(VSS),.VDD(VDD),.Y(I39916),.A(g30293));
  NOT NOT1_12841(.VSS(VSS),.VDD(VDD),.Y(g30369),.A(I39916));
  NOT NOT1_12842(.VSS(VSS),.VDD(VDD),.Y(I39919),.A(g30294));
  NOT NOT1_12843(.VSS(VSS),.VDD(VDD),.Y(g30370),.A(I39919));
  NOT NOT1_12844(.VSS(VSS),.VDD(VDD),.Y(I39922),.A(g30295));
  NOT NOT1_12845(.VSS(VSS),.VDD(VDD),.Y(g30371),.A(I39922));
  NOT NOT1_12846(.VSS(VSS),.VDD(VDD),.Y(I39926),.A(g30296));
  NOT NOT1_12847(.VSS(VSS),.VDD(VDD),.Y(g30373),.A(I39926));
  NOT NOT1_12848(.VSS(VSS),.VDD(VDD),.Y(I39930),.A(g30297));
  NOT NOT1_12849(.VSS(VSS),.VDD(VDD),.Y(g30375),.A(I39930));
  NOT NOT1_12850(.VSS(VSS),.VDD(VDD),.Y(I39933),.A(g30298));
  NOT NOT1_12851(.VSS(VSS),.VDD(VDD),.Y(g30376),.A(I39933));
  NOT NOT1_12852(.VSS(VSS),.VDD(VDD),.Y(I39936),.A(g30299));
  NOT NOT1_12853(.VSS(VSS),.VDD(VDD),.Y(g30377),.A(I39936));
  NOT NOT1_12854(.VSS(VSS),.VDD(VDD),.Y(I39939),.A(g30300));
  NOT NOT1_12855(.VSS(VSS),.VDD(VDD),.Y(g30378),.A(I39939));
  NOT NOT1_12856(.VSS(VSS),.VDD(VDD),.Y(I39942),.A(g30301));
  NOT NOT1_12857(.VSS(VSS),.VDD(VDD),.Y(g30379),.A(I39942));
  NOT NOT1_12858(.VSS(VSS),.VDD(VDD),.Y(I39945),.A(g30302));
  NOT NOT1_12859(.VSS(VSS),.VDD(VDD),.Y(g30380),.A(I39945));
  NOT NOT1_12860(.VSS(VSS),.VDD(VDD),.Y(I39948),.A(g30303));
  NOT NOT1_12861(.VSS(VSS),.VDD(VDD),.Y(g30381),.A(I39948));
  NOT NOT1_12862(.VSS(VSS),.VDD(VDD),.Y(I39951),.A(g30304));
  NOT NOT1_12863(.VSS(VSS),.VDD(VDD),.Y(g30382),.A(I39951));
  NOT NOT1_12864(.VSS(VSS),.VDD(VDD),.Y(g30383),.A(g30306));
  NOT NOT1_12865(.VSS(VSS),.VDD(VDD),.Y(I39976),.A(g30245));
  NOT NOT1_12866(.VSS(VSS),.VDD(VDD),.Y(g30408),.A(I39976));
  NOT NOT1_12867(.VSS(VSS),.VDD(VDD),.Y(I39982),.A(g30305));
  NOT NOT1_12868(.VSS(VSS),.VDD(VDD),.Y(g30412),.A(I39982));
  NOT NOT1_12869(.VSS(VSS),.VDD(VDD),.Y(I39985),.A(g30246));
  NOT NOT1_12870(.VSS(VSS),.VDD(VDD),.Y(g30435),.A(I39985));
  NOT NOT1_12871(.VSS(VSS),.VDD(VDD),.Y(I39991),.A(g30247));
  NOT NOT1_12872(.VSS(VSS),.VDD(VDD),.Y(g30439),.A(I39991));
  NOT NOT1_12873(.VSS(VSS),.VDD(VDD),.Y(I39997),.A(g30248));
  NOT NOT1_12874(.VSS(VSS),.VDD(VDD),.Y(g30443),.A(I39997));
  NOT NOT1_12875(.VSS(VSS),.VDD(VDD),.Y(I40002),.A(g30249));
  NOT NOT1_12876(.VSS(VSS),.VDD(VDD),.Y(g30446),.A(I40002));
  NOT NOT1_12877(.VSS(VSS),.VDD(VDD),.Y(I40008),.A(g30250));
  NOT NOT1_12878(.VSS(VSS),.VDD(VDD),.Y(g30450),.A(I40008));
  NOT NOT1_12879(.VSS(VSS),.VDD(VDD),.Y(I40016),.A(g30251));
  NOT NOT1_12880(.VSS(VSS),.VDD(VDD),.Y(g30456),.A(I40016));
  NOT NOT1_12881(.VSS(VSS),.VDD(VDD),.Y(I40021),.A(g30252));
  NOT NOT1_12882(.VSS(VSS),.VDD(VDD),.Y(g30459),.A(I40021));
  NOT NOT1_12883(.VSS(VSS),.VDD(VDD),.Y(I40027),.A(g30253));
  NOT NOT1_12884(.VSS(VSS),.VDD(VDD),.Y(g30463),.A(I40027));
  NOT NOT1_12885(.VSS(VSS),.VDD(VDD),.Y(I40032),.A(g30254));
  NOT NOT1_12886(.VSS(VSS),.VDD(VDD),.Y(g30466),.A(I40032));
  NOT NOT1_12887(.VSS(VSS),.VDD(VDD),.Y(I40039),.A(g30255));
  NOT NOT1_12888(.VSS(VSS),.VDD(VDD),.Y(g30471),.A(I40039));
  NOT NOT1_12889(.VSS(VSS),.VDD(VDD),.Y(I40044),.A(g30256));
  NOT NOT1_12890(.VSS(VSS),.VDD(VDD),.Y(g30474),.A(I40044));
  NOT NOT1_12891(.VSS(VSS),.VDD(VDD),.Y(I40051),.A(g30257));
  NOT NOT1_12892(.VSS(VSS),.VDD(VDD),.Y(g30479),.A(I40051));
  NOT NOT1_12893(.VSS(VSS),.VDD(VDD),.Y(I40054),.A(g30258));
  NOT NOT1_12894(.VSS(VSS),.VDD(VDD),.Y(g30480),.A(I40054));
  NOT NOT1_12895(.VSS(VSS),.VDD(VDD),.Y(I40059),.A(g30259));
  NOT NOT1_12896(.VSS(VSS),.VDD(VDD),.Y(g30483),.A(I40059));
  NOT NOT1_12897(.VSS(VSS),.VDD(VDD),.Y(I40066),.A(g30260));
  NOT NOT1_12898(.VSS(VSS),.VDD(VDD),.Y(g30488),.A(I40066));
  NOT NOT1_12899(.VSS(VSS),.VDD(VDD),.Y(I40071),.A(g30261));
  NOT NOT1_12900(.VSS(VSS),.VDD(VDD),.Y(g30491),.A(I40071));
  NOT NOT1_12901(.VSS(VSS),.VDD(VDD),.Y(I40075),.A(g30262));
  NOT NOT1_12902(.VSS(VSS),.VDD(VDD),.Y(g30493),.A(I40075));
  NOT NOT1_12903(.VSS(VSS),.VDD(VDD),.Y(I40078),.A(g30263));
  NOT NOT1_12904(.VSS(VSS),.VDD(VDD),.Y(g30494),.A(I40078));
  NOT NOT1_12905(.VSS(VSS),.VDD(VDD),.Y(I40083),.A(g30264));
  NOT NOT1_12906(.VSS(VSS),.VDD(VDD),.Y(g30497),.A(I40083));
  NOT NOT1_12907(.VSS(VSS),.VDD(VDD),.Y(I40086),.A(g30265));
  NOT NOT1_12908(.VSS(VSS),.VDD(VDD),.Y(g30498),.A(I40086));
  NOT NOT1_12909(.VSS(VSS),.VDD(VDD),.Y(I40091),.A(g30266));
  NOT NOT1_12910(.VSS(VSS),.VDD(VDD),.Y(g30501),.A(I40091));
  NOT NOT1_12911(.VSS(VSS),.VDD(VDD),.Y(I40098),.A(g30491));
  NOT NOT1_12912(.VSS(VSS),.VDD(VDD),.Y(g30506),.A(I40098));
  NOT NOT1_12913(.VSS(VSS),.VDD(VDD),.Y(I40101),.A(g30326));
  NOT NOT1_12914(.VSS(VSS),.VDD(VDD),.Y(g30507),.A(I40101));
  NOT NOT1_12915(.VSS(VSS),.VDD(VDD),.Y(I40104),.A(g30342));
  NOT NOT1_12916(.VSS(VSS),.VDD(VDD),.Y(g30508),.A(I40104));
  NOT NOT1_12917(.VSS(VSS),.VDD(VDD),.Y(I40107),.A(g30343));
  NOT NOT1_12918(.VSS(VSS),.VDD(VDD),.Y(g30509),.A(I40107));
  NOT NOT1_12919(.VSS(VSS),.VDD(VDD),.Y(I40110),.A(g30357));
  NOT NOT1_12920(.VSS(VSS),.VDD(VDD),.Y(g30510),.A(I40110));
  NOT NOT1_12921(.VSS(VSS),.VDD(VDD),.Y(I40113),.A(g30368));
  NOT NOT1_12922(.VSS(VSS),.VDD(VDD),.Y(g30511),.A(I40113));
  NOT NOT1_12923(.VSS(VSS),.VDD(VDD),.Y(I40116),.A(g30408));
  NOT NOT1_12924(.VSS(VSS),.VDD(VDD),.Y(g30512),.A(I40116));
  NOT NOT1_12925(.VSS(VSS),.VDD(VDD),.Y(I40119),.A(g30435));
  NOT NOT1_12926(.VSS(VSS),.VDD(VDD),.Y(g30513),.A(I40119));
  NOT NOT1_12927(.VSS(VSS),.VDD(VDD),.Y(I40122),.A(g30443));
  NOT NOT1_12928(.VSS(VSS),.VDD(VDD),.Y(g30514),.A(I40122));
  NOT NOT1_12929(.VSS(VSS),.VDD(VDD),.Y(I40125),.A(g30466));
  NOT NOT1_12930(.VSS(VSS),.VDD(VDD),.Y(g30515),.A(I40125));
  NOT NOT1_12931(.VSS(VSS),.VDD(VDD),.Y(I40128),.A(g30479));
  NOT NOT1_12932(.VSS(VSS),.VDD(VDD),.Y(g30516),.A(I40128));
  NOT NOT1_12933(.VSS(VSS),.VDD(VDD),.Y(I40131),.A(g30493));
  NOT NOT1_12934(.VSS(VSS),.VDD(VDD),.Y(g30517),.A(I40131));
  NOT NOT1_12935(.VSS(VSS),.VDD(VDD),.Y(I40134),.A(g30480));
  NOT NOT1_12936(.VSS(VSS),.VDD(VDD),.Y(g30518),.A(I40134));
  NOT NOT1_12937(.VSS(VSS),.VDD(VDD),.Y(I40137),.A(g30494));
  NOT NOT1_12938(.VSS(VSS),.VDD(VDD),.Y(g30519),.A(I40137));
  NOT NOT1_12939(.VSS(VSS),.VDD(VDD),.Y(I40140),.A(g30328));
  NOT NOT1_12940(.VSS(VSS),.VDD(VDD),.Y(g30520),.A(I40140));
  NOT NOT1_12941(.VSS(VSS),.VDD(VDD),.Y(I40143),.A(g30329));
  NOT NOT1_12942(.VSS(VSS),.VDD(VDD),.Y(g30521),.A(I40143));
  NOT NOT1_12943(.VSS(VSS),.VDD(VDD),.Y(I40146),.A(g30344));
  NOT NOT1_12944(.VSS(VSS),.VDD(VDD),.Y(g30522),.A(I40146));
  NOT NOT1_12945(.VSS(VSS),.VDD(VDD),.Y(I40149),.A(g30358));
  NOT NOT1_12946(.VSS(VSS),.VDD(VDD),.Y(g30523),.A(I40149));
  NOT NOT1_12947(.VSS(VSS),.VDD(VDD),.Y(I40152),.A(g30359));
  NOT NOT1_12948(.VSS(VSS),.VDD(VDD),.Y(g30524),.A(I40152));
  NOT NOT1_12949(.VSS(VSS),.VDD(VDD),.Y(I40155),.A(g30369));
  NOT NOT1_12950(.VSS(VSS),.VDD(VDD),.Y(g30525),.A(I40155));
  NOT NOT1_12951(.VSS(VSS),.VDD(VDD),.Y(I40158),.A(g30376));
  NOT NOT1_12952(.VSS(VSS),.VDD(VDD),.Y(g30526),.A(I40158));
  NOT NOT1_12953(.VSS(VSS),.VDD(VDD),.Y(I40161),.A(g30439));
  NOT NOT1_12954(.VSS(VSS),.VDD(VDD),.Y(g30527),.A(I40161));
  NOT NOT1_12955(.VSS(VSS),.VDD(VDD),.Y(I40164),.A(g30446));
  NOT NOT1_12956(.VSS(VSS),.VDD(VDD),.Y(g30528),.A(I40164));
  NOT NOT1_12957(.VSS(VSS),.VDD(VDD),.Y(I40167),.A(g30456));
  NOT NOT1_12958(.VSS(VSS),.VDD(VDD),.Y(g30529),.A(I40167));
  NOT NOT1_12959(.VSS(VSS),.VDD(VDD),.Y(I40170),.A(g30483));
  NOT NOT1_12960(.VSS(VSS),.VDD(VDD),.Y(g30530),.A(I40170));
  NOT NOT1_12961(.VSS(VSS),.VDD(VDD),.Y(I40173),.A(g30497));
  NOT NOT1_12962(.VSS(VSS),.VDD(VDD),.Y(g30531),.A(I40173));
  NOT NOT1_12963(.VSS(VSS),.VDD(VDD),.Y(I40176),.A(g30331));
  NOT NOT1_12964(.VSS(VSS),.VDD(VDD),.Y(g30532),.A(I40176));
  NOT NOT1_12965(.VSS(VSS),.VDD(VDD),.Y(I40179),.A(g30498));
  NOT NOT1_12966(.VSS(VSS),.VDD(VDD),.Y(g30533),.A(I40179));
  NOT NOT1_12967(.VSS(VSS),.VDD(VDD),.Y(I40182),.A(g30332));
  NOT NOT1_12968(.VSS(VSS),.VDD(VDD),.Y(g30534),.A(I40182));
  NOT NOT1_12969(.VSS(VSS),.VDD(VDD),.Y(I40185),.A(g30346));
  NOT NOT1_12970(.VSS(VSS),.VDD(VDD),.Y(g30535),.A(I40185));
  NOT NOT1_12971(.VSS(VSS),.VDD(VDD),.Y(I40188),.A(g30347));
  NOT NOT1_12972(.VSS(VSS),.VDD(VDD),.Y(g30536),.A(I40188));
  NOT NOT1_12973(.VSS(VSS),.VDD(VDD),.Y(I40191),.A(g30360));
  NOT NOT1_12974(.VSS(VSS),.VDD(VDD),.Y(g30537),.A(I40191));
  NOT NOT1_12975(.VSS(VSS),.VDD(VDD),.Y(I40194),.A(g30370));
  NOT NOT1_12976(.VSS(VSS),.VDD(VDD),.Y(g30538),.A(I40194));
  NOT NOT1_12977(.VSS(VSS),.VDD(VDD),.Y(I40197),.A(g30371));
  NOT NOT1_12978(.VSS(VSS),.VDD(VDD),.Y(g30539),.A(I40197));
  NOT NOT1_12979(.VSS(VSS),.VDD(VDD),.Y(I40200),.A(g30377));
  NOT NOT1_12980(.VSS(VSS),.VDD(VDD),.Y(g30540),.A(I40200));
  NOT NOT1_12981(.VSS(VSS),.VDD(VDD),.Y(I40203),.A(g30380));
  NOT NOT1_12982(.VSS(VSS),.VDD(VDD),.Y(g30541),.A(I40203));
  NOT NOT1_12983(.VSS(VSS),.VDD(VDD),.Y(I40206),.A(g30450));
  NOT NOT1_12984(.VSS(VSS),.VDD(VDD),.Y(g30542),.A(I40206));
  NOT NOT1_12985(.VSS(VSS),.VDD(VDD),.Y(I40209),.A(g30459));
  NOT NOT1_12986(.VSS(VSS),.VDD(VDD),.Y(g30543),.A(I40209));
  NOT NOT1_12987(.VSS(VSS),.VDD(VDD),.Y(I40212),.A(g30471));
  NOT NOT1_12988(.VSS(VSS),.VDD(VDD),.Y(g30544),.A(I40212));
  NOT NOT1_12989(.VSS(VSS),.VDD(VDD),.Y(I40215),.A(g30501));
  NOT NOT1_12990(.VSS(VSS),.VDD(VDD),.Y(g30545),.A(I40215));
  NOT NOT1_12991(.VSS(VSS),.VDD(VDD),.Y(I40218),.A(g30335));
  NOT NOT1_12992(.VSS(VSS),.VDD(VDD),.Y(g30546),.A(I40218));
  NOT NOT1_12993(.VSS(VSS),.VDD(VDD),.Y(I40221),.A(g30349));
  NOT NOT1_12994(.VSS(VSS),.VDD(VDD),.Y(g30547),.A(I40221));
  NOT NOT1_12995(.VSS(VSS),.VDD(VDD),.Y(I40224),.A(g30336));
  NOT NOT1_12996(.VSS(VSS),.VDD(VDD),.Y(g30548),.A(I40224));
  NOT NOT1_12997(.VSS(VSS),.VDD(VDD),.Y(I40227),.A(g30350));
  NOT NOT1_12998(.VSS(VSS),.VDD(VDD),.Y(g30549),.A(I40227));
  NOT NOT1_12999(.VSS(VSS),.VDD(VDD),.Y(I40230),.A(g30362));
  NOT NOT1_13000(.VSS(VSS),.VDD(VDD),.Y(g30550),.A(I40230));
  NOT NOT1_13001(.VSS(VSS),.VDD(VDD),.Y(I40233),.A(g30363));
  NOT NOT1_13002(.VSS(VSS),.VDD(VDD),.Y(g30551),.A(I40233));
  NOT NOT1_13003(.VSS(VSS),.VDD(VDD),.Y(I40236),.A(g30373));
  NOT NOT1_13004(.VSS(VSS),.VDD(VDD),.Y(g30552),.A(I40236));
  NOT NOT1_13005(.VSS(VSS),.VDD(VDD),.Y(I40239),.A(g30378));
  NOT NOT1_13006(.VSS(VSS),.VDD(VDD),.Y(g30553),.A(I40239));
  NOT NOT1_13007(.VSS(VSS),.VDD(VDD),.Y(I40242),.A(g30379));
  NOT NOT1_13008(.VSS(VSS),.VDD(VDD),.Y(g30554),.A(I40242));
  NOT NOT1_13009(.VSS(VSS),.VDD(VDD),.Y(I40245),.A(g30381));
  NOT NOT1_13010(.VSS(VSS),.VDD(VDD),.Y(g30555),.A(I40245));
  NOT NOT1_13011(.VSS(VSS),.VDD(VDD),.Y(I40248),.A(g30382));
  NOT NOT1_13012(.VSS(VSS),.VDD(VDD),.Y(g30556),.A(I40248));
  NOT NOT1_13013(.VSS(VSS),.VDD(VDD),.Y(I40251),.A(g30463));
  NOT NOT1_13014(.VSS(VSS),.VDD(VDD),.Y(g30557),.A(I40251));
  NOT NOT1_13015(.VSS(VSS),.VDD(VDD),.Y(I40254),.A(g30474));
  NOT NOT1_13016(.VSS(VSS),.VDD(VDD),.Y(g30558),.A(I40254));
  NOT NOT1_13017(.VSS(VSS),.VDD(VDD),.Y(I40257),.A(g30488));
  NOT NOT1_13018(.VSS(VSS),.VDD(VDD),.Y(g30559),.A(I40257));
  NOT NOT1_13019(.VSS(VSS),.VDD(VDD),.Y(I40260),.A(g30339));
  NOT NOT1_13020(.VSS(VSS),.VDD(VDD),.Y(g30560),.A(I40260));
  NOT NOT1_13021(.VSS(VSS),.VDD(VDD),.Y(I40263),.A(g30353));
  NOT NOT1_13022(.VSS(VSS),.VDD(VDD),.Y(g30561),.A(I40263));
  NOT NOT1_13023(.VSS(VSS),.VDD(VDD),.Y(I40266),.A(g30365));
  NOT NOT1_13024(.VSS(VSS),.VDD(VDD),.Y(g30562),.A(I40266));
  NOT NOT1_13025(.VSS(VSS),.VDD(VDD),.Y(I40269),.A(g30354));
  NOT NOT1_13026(.VSS(VSS),.VDD(VDD),.Y(g30563),.A(I40269));
  NOT NOT1_13027(.VSS(VSS),.VDD(VDD),.Y(I40272),.A(g30366));
  NOT NOT1_13028(.VSS(VSS),.VDD(VDD),.Y(g30564),.A(I40272));
  NOT NOT1_13029(.VSS(VSS),.VDD(VDD),.Y(I40275),.A(g30375));
  NOT NOT1_13030(.VSS(VSS),.VDD(VDD),.Y(g30565),.A(I40275));
  NOT NOT1_13031(.VSS(VSS),.VDD(VDD),.Y(g30567),.A(g30403));
  NOT NOT1_13032(.VSS(VSS),.VDD(VDD),.Y(g30568),.A(g30402));
  NOT NOT1_13033(.VSS(VSS),.VDD(VDD),.Y(g30569),.A(g30406));
  NOT NOT1_13034(.VSS(VSS),.VDD(VDD),.Y(g30570),.A(g30404));
  NOT NOT1_13035(.VSS(VSS),.VDD(VDD),.Y(g30571),.A(g30401));
  NOT NOT1_13036(.VSS(VSS),.VDD(VDD),.Y(g30572),.A(g30399));
  NOT NOT1_13037(.VSS(VSS),.VDD(VDD),.Y(g30573),.A(g30405));
  NOT NOT1_13038(.VSS(VSS),.VDD(VDD),.Y(g30574),.A(g30400));
  NOT NOT1_13039(.VSS(VSS),.VDD(VDD),.Y(g30575),.A(g30412));
  NOT NOT1_13040(.VSS(VSS),.VDD(VDD),.Y(I40288),.A(g30455));
  NOT NOT1_13041(.VSS(VSS),.VDD(VDD),.Y(g30578),.A(I40288));
  NOT NOT1_13042(.VSS(VSS),.VDD(VDD),.Y(I40291),.A(g30468));
  NOT NOT1_13043(.VSS(VSS),.VDD(VDD),.Y(g30579),.A(I40291));
  NOT NOT1_13044(.VSS(VSS),.VDD(VDD),.Y(I40294),.A(g30470));
  NOT NOT1_13045(.VSS(VSS),.VDD(VDD),.Y(g30580),.A(I40294));
  NOT NOT1_13046(.VSS(VSS),.VDD(VDD),.Y(I40297),.A(g30482));
  NOT NOT1_13047(.VSS(VSS),.VDD(VDD),.Y(g30581),.A(I40297));
  NOT NOT1_13048(.VSS(VSS),.VDD(VDD),.Y(I40300),.A(g30485));
  NOT NOT1_13049(.VSS(VSS),.VDD(VDD),.Y(g30582),.A(I40300));
  NOT NOT1_13050(.VSS(VSS),.VDD(VDD),.Y(I40303),.A(g30487));
  NOT NOT1_13051(.VSS(VSS),.VDD(VDD),.Y(g30583),.A(I40303));
  NOT NOT1_13052(.VSS(VSS),.VDD(VDD),.Y(I40307),.A(g30500));
  NOT NOT1_13053(.VSS(VSS),.VDD(VDD),.Y(g30585),.A(I40307));
  NOT NOT1_13054(.VSS(VSS),.VDD(VDD),.Y(I40310),.A(g30503));
  NOT NOT1_13055(.VSS(VSS),.VDD(VDD),.Y(g30586),.A(I40310));
  NOT NOT1_13056(.VSS(VSS),.VDD(VDD),.Y(I40313),.A(g30505));
  NOT NOT1_13057(.VSS(VSS),.VDD(VDD),.Y(g30587),.A(I40313));
  NOT NOT1_13058(.VSS(VSS),.VDD(VDD),.Y(I40317),.A(g30338));
  NOT NOT1_13059(.VSS(VSS),.VDD(VDD),.Y(g30591),.A(I40317));
  NOT NOT1_13060(.VSS(VSS),.VDD(VDD),.Y(I40320),.A(g30341));
  NOT NOT1_13061(.VSS(VSS),.VDD(VDD),.Y(g30592),.A(I40320));
  NOT NOT1_13062(.VSS(VSS),.VDD(VDD),.Y(I40326),.A(g30356));
  NOT NOT1_13063(.VSS(VSS),.VDD(VDD),.Y(g30600),.A(I40326));
  NOT NOT1_13064(.VSS(VSS),.VDD(VDD),.Y(I40420),.A(g30578));
  NOT NOT1_13065(.VSS(VSS),.VDD(VDD),.Y(g30710),.A(I40420));
  NOT NOT1_13066(.VSS(VSS),.VDD(VDD),.Y(I40423),.A(g30579));
  NOT NOT1_13067(.VSS(VSS),.VDD(VDD),.Y(g30711),.A(I40423));
  NOT NOT1_13068(.VSS(VSS),.VDD(VDD),.Y(I40426),.A(g30581));
  NOT NOT1_13069(.VSS(VSS),.VDD(VDD),.Y(g30712),.A(I40426));
  NOT NOT1_13070(.VSS(VSS),.VDD(VDD),.Y(I40429),.A(g30580));
  NOT NOT1_13071(.VSS(VSS),.VDD(VDD),.Y(g30713),.A(I40429));
  NOT NOT1_13072(.VSS(VSS),.VDD(VDD),.Y(I40432),.A(g30582));
  NOT NOT1_13073(.VSS(VSS),.VDD(VDD),.Y(g30714),.A(I40432));
  NOT NOT1_13074(.VSS(VSS),.VDD(VDD),.Y(I40435),.A(g30585));
  NOT NOT1_13075(.VSS(VSS),.VDD(VDD),.Y(g30715),.A(I40435));
  NOT NOT1_13076(.VSS(VSS),.VDD(VDD),.Y(I40438),.A(g30583));
  NOT NOT1_13077(.VSS(VSS),.VDD(VDD),.Y(g30716),.A(I40438));
  NOT NOT1_13078(.VSS(VSS),.VDD(VDD),.Y(I40441),.A(g30586));
  NOT NOT1_13079(.VSS(VSS),.VDD(VDD),.Y(g30717),.A(I40441));
  NOT NOT1_13080(.VSS(VSS),.VDD(VDD),.Y(I40444),.A(g30591));
  NOT NOT1_13081(.VSS(VSS),.VDD(VDD),.Y(g30718),.A(I40444));
  NOT NOT1_13082(.VSS(VSS),.VDD(VDD),.Y(I40447),.A(g30587));
  NOT NOT1_13083(.VSS(VSS),.VDD(VDD),.Y(g30719),.A(I40447));
  NOT NOT1_13084(.VSS(VSS),.VDD(VDD),.Y(I40450),.A(g30592));
  NOT NOT1_13085(.VSS(VSS),.VDD(VDD),.Y(g30720),.A(I40450));
  NOT NOT1_13086(.VSS(VSS),.VDD(VDD),.Y(I40453),.A(g30600));
  NOT NOT1_13087(.VSS(VSS),.VDD(VDD),.Y(g30721),.A(I40453));
  NOT NOT1_13088(.VSS(VSS),.VDD(VDD),.Y(I40456),.A(g30668));
  NOT NOT1_13089(.VSS(VSS),.VDD(VDD),.Y(g30722),.A(I40456));
  NOT NOT1_13090(.VSS(VSS),.VDD(VDD),.Y(I40459),.A(g30669));
  NOT NOT1_13091(.VSS(VSS),.VDD(VDD),.Y(g30723),.A(I40459));
  NOT NOT1_13092(.VSS(VSS),.VDD(VDD),.Y(I40462),.A(g30670));
  NOT NOT1_13093(.VSS(VSS),.VDD(VDD),.Y(g30724),.A(I40462));
  NOT NOT1_13094(.VSS(VSS),.VDD(VDD),.Y(I40465),.A(g30671));
  NOT NOT1_13095(.VSS(VSS),.VDD(VDD),.Y(g30725),.A(I40465));
  NOT NOT1_13096(.VSS(VSS),.VDD(VDD),.Y(I40468),.A(g30672));
  NOT NOT1_13097(.VSS(VSS),.VDD(VDD),.Y(g30726),.A(I40468));
  NOT NOT1_13098(.VSS(VSS),.VDD(VDD),.Y(I40471),.A(g30673));
  NOT NOT1_13099(.VSS(VSS),.VDD(VDD),.Y(g30727),.A(I40471));
  NOT NOT1_13100(.VSS(VSS),.VDD(VDD),.Y(I40475),.A(g30674));
  NOT NOT1_13101(.VSS(VSS),.VDD(VDD),.Y(g30729),.A(I40475));
  NOT NOT1_13102(.VSS(VSS),.VDD(VDD),.Y(I40478),.A(g30675));
  NOT NOT1_13103(.VSS(VSS),.VDD(VDD),.Y(g30730),.A(I40478));
  NOT NOT1_13104(.VSS(VSS),.VDD(VDD),.Y(I40481),.A(g30676));
  NOT NOT1_13105(.VSS(VSS),.VDD(VDD),.Y(g30731),.A(I40481));
  NOT NOT1_13106(.VSS(VSS),.VDD(VDD),.Y(I40484),.A(g30677));
  NOT NOT1_13107(.VSS(VSS),.VDD(VDD),.Y(g30732),.A(I40484));
  NOT NOT1_13108(.VSS(VSS),.VDD(VDD),.Y(I40487),.A(g30678));
  NOT NOT1_13109(.VSS(VSS),.VDD(VDD),.Y(g30733),.A(I40487));
  NOT NOT1_13110(.VSS(VSS),.VDD(VDD),.Y(I40490),.A(g30679));
  NOT NOT1_13111(.VSS(VSS),.VDD(VDD),.Y(g30734),.A(I40490));
  NOT NOT1_13112(.VSS(VSS),.VDD(VDD),.Y(I40495),.A(g30680));
  NOT NOT1_13113(.VSS(VSS),.VDD(VDD),.Y(g30737),.A(I40495));
  NOT NOT1_13114(.VSS(VSS),.VDD(VDD),.Y(I40498),.A(g30681));
  NOT NOT1_13115(.VSS(VSS),.VDD(VDD),.Y(g30738),.A(I40498));
  NOT NOT1_13116(.VSS(VSS),.VDD(VDD),.Y(I40501),.A(g30682));
  NOT NOT1_13117(.VSS(VSS),.VDD(VDD),.Y(g30739),.A(I40501));
  NOT NOT1_13118(.VSS(VSS),.VDD(VDD),.Y(I40504),.A(g30683));
  NOT NOT1_13119(.VSS(VSS),.VDD(VDD),.Y(g30740),.A(I40504));
  NOT NOT1_13120(.VSS(VSS),.VDD(VDD),.Y(I40507),.A(g30684));
  NOT NOT1_13121(.VSS(VSS),.VDD(VDD),.Y(g30741),.A(I40507));
  NOT NOT1_13122(.VSS(VSS),.VDD(VDD),.Y(I40510),.A(g30686));
  NOT NOT1_13123(.VSS(VSS),.VDD(VDD),.Y(g30742),.A(I40510));
  NOT NOT1_13124(.VSS(VSS),.VDD(VDD),.Y(I40515),.A(g30687));
  NOT NOT1_13125(.VSS(VSS),.VDD(VDD),.Y(g30745),.A(I40515));
  NOT NOT1_13126(.VSS(VSS),.VDD(VDD),.Y(I40518),.A(g30688));
  NOT NOT1_13127(.VSS(VSS),.VDD(VDD),.Y(g30746),.A(I40518));
  NOT NOT1_13128(.VSS(VSS),.VDD(VDD),.Y(I40521),.A(g30689));
  NOT NOT1_13129(.VSS(VSS),.VDD(VDD),.Y(g30747),.A(I40521));
  NOT NOT1_13130(.VSS(VSS),.VDD(VDD),.Y(I40524),.A(g30690));
  NOT NOT1_13131(.VSS(VSS),.VDD(VDD),.Y(g30748),.A(I40524));
  NOT NOT1_13132(.VSS(VSS),.VDD(VDD),.Y(I40527),.A(g30691));
  NOT NOT1_13133(.VSS(VSS),.VDD(VDD),.Y(g30749),.A(I40527));
  NOT NOT1_13134(.VSS(VSS),.VDD(VDD),.Y(I40531),.A(g30692));
  NOT NOT1_13135(.VSS(VSS),.VDD(VDD),.Y(g30751),.A(I40531));
  NOT NOT1_13136(.VSS(VSS),.VDD(VDD),.Y(I40534),.A(g30693));
  NOT NOT1_13137(.VSS(VSS),.VDD(VDD),.Y(g30752),.A(I40534));
  NOT NOT1_13138(.VSS(VSS),.VDD(VDD),.Y(I40537),.A(g30694));
  NOT NOT1_13139(.VSS(VSS),.VDD(VDD),.Y(g30753),.A(I40537));
  NOT NOT1_13140(.VSS(VSS),.VDD(VDD),.Y(I40542),.A(g30695));
  NOT NOT1_13141(.VSS(VSS),.VDD(VDD),.Y(g30756),.A(I40542));
  NOT NOT1_13142(.VSS(VSS),.VDD(VDD),.Y(g30765),.A(g30685));
  NOT NOT1_13143(.VSS(VSS),.VDD(VDD),.Y(I40555),.A(g30699));
  NOT NOT1_13144(.VSS(VSS),.VDD(VDD),.Y(g30767),.A(I40555));
  NOT NOT1_13145(.VSS(VSS),.VDD(VDD),.Y(I40565),.A(g30700));
  NOT NOT1_13146(.VSS(VSS),.VDD(VDD),.Y(g30769),.A(I40565));
  NOT NOT1_13147(.VSS(VSS),.VDD(VDD),.Y(I40568),.A(g30701));
  NOT NOT1_13148(.VSS(VSS),.VDD(VDD),.Y(g30770),.A(I40568));
  NOT NOT1_13149(.VSS(VSS),.VDD(VDD),.Y(I40578),.A(g30702));
  NOT NOT1_13150(.VSS(VSS),.VDD(VDD),.Y(g30772),.A(I40578));
  NOT NOT1_13151(.VSS(VSS),.VDD(VDD),.Y(I40581),.A(g30703));
  NOT NOT1_13152(.VSS(VSS),.VDD(VDD),.Y(g30773),.A(I40581));
  NOT NOT1_13153(.VSS(VSS),.VDD(VDD),.Y(I40584),.A(g30704));
  NOT NOT1_13154(.VSS(VSS),.VDD(VDD),.Y(g30774),.A(I40584));
  NOT NOT1_13155(.VSS(VSS),.VDD(VDD),.Y(I40594),.A(g30705));
  NOT NOT1_13156(.VSS(VSS),.VDD(VDD),.Y(g30776),.A(I40594));
  NOT NOT1_13157(.VSS(VSS),.VDD(VDD),.Y(I40597),.A(g30706));
  NOT NOT1_13158(.VSS(VSS),.VDD(VDD),.Y(g30777),.A(I40597));
  NOT NOT1_13159(.VSS(VSS),.VDD(VDD),.Y(I40600),.A(g30707));
  NOT NOT1_13160(.VSS(VSS),.VDD(VDD),.Y(g30778),.A(I40600));
  NOT NOT1_13161(.VSS(VSS),.VDD(VDD),.Y(I40611),.A(g30708));
  NOT NOT1_13162(.VSS(VSS),.VDD(VDD),.Y(g30781),.A(I40611));
  NOT NOT1_13163(.VSS(VSS),.VDD(VDD),.Y(I40614),.A(g30709));
  NOT NOT1_13164(.VSS(VSS),.VDD(VDD),.Y(g30782),.A(I40614));
  NOT NOT1_13165(.VSS(VSS),.VDD(VDD),.Y(I40618),.A(g30566));
  NOT NOT1_13166(.VSS(VSS),.VDD(VDD),.Y(g30784),.A(I40618));
  NOT NOT1_13167(.VSS(VSS),.VDD(VDD),.Y(I40634),.A(g30571));
  NOT NOT1_13168(.VSS(VSS),.VDD(VDD),.Y(g30792),.A(I40634));
  NOT NOT1_13169(.VSS(VSS),.VDD(VDD),.Y(I40637),.A(g30570));
  NOT NOT1_13170(.VSS(VSS),.VDD(VDD),.Y(g30793),.A(I40637));
  NOT NOT1_13171(.VSS(VSS),.VDD(VDD),.Y(I40640),.A(g30569));
  NOT NOT1_13172(.VSS(VSS),.VDD(VDD),.Y(g30794),.A(I40640));
  NOT NOT1_13173(.VSS(VSS),.VDD(VDD),.Y(I40643),.A(g30568));
  NOT NOT1_13174(.VSS(VSS),.VDD(VDD),.Y(g30795),.A(I40643));
  NOT NOT1_13175(.VSS(VSS),.VDD(VDD),.Y(I40647),.A(g30567));
  NOT NOT1_13176(.VSS(VSS),.VDD(VDD),.Y(g30797),.A(I40647));
  NOT NOT1_13177(.VSS(VSS),.VDD(VDD),.Y(I40651),.A(g30574));
  NOT NOT1_13178(.VSS(VSS),.VDD(VDD),.Y(g30799),.A(I40651));
  NOT NOT1_13179(.VSS(VSS),.VDD(VDD),.Y(I40654),.A(g30573));
  NOT NOT1_13180(.VSS(VSS),.VDD(VDD),.Y(g30800),.A(I40654));
  NOT NOT1_13181(.VSS(VSS),.VDD(VDD),.Y(I40658),.A(g30572));
  NOT NOT1_13182(.VSS(VSS),.VDD(VDD),.Y(g30802),.A(I40658));
  NOT NOT1_13183(.VSS(VSS),.VDD(VDD),.Y(I40661),.A(g30635));
  NOT NOT1_13184(.VSS(VSS),.VDD(VDD),.Y(g30803),.A(I40661));
  NOT NOT1_13185(.VSS(VSS),.VDD(VDD),.Y(I40664),.A(g30636));
  NOT NOT1_13186(.VSS(VSS),.VDD(VDD),.Y(g30804),.A(I40664));
  NOT NOT1_13187(.VSS(VSS),.VDD(VDD),.Y(I40667),.A(g30637));
  NOT NOT1_13188(.VSS(VSS),.VDD(VDD),.Y(g30805),.A(I40667));
  NOT NOT1_13189(.VSS(VSS),.VDD(VDD),.Y(I40670),.A(g30638));
  NOT NOT1_13190(.VSS(VSS),.VDD(VDD),.Y(g30806),.A(I40670));
  NOT NOT1_13191(.VSS(VSS),.VDD(VDD),.Y(I40673),.A(g30639));
  NOT NOT1_13192(.VSS(VSS),.VDD(VDD),.Y(g30807),.A(I40673));
  NOT NOT1_13193(.VSS(VSS),.VDD(VDD),.Y(I40676),.A(g30640));
  NOT NOT1_13194(.VSS(VSS),.VDD(VDD),.Y(g30808),.A(I40676));
  NOT NOT1_13195(.VSS(VSS),.VDD(VDD),.Y(I40679),.A(g30641));
  NOT NOT1_13196(.VSS(VSS),.VDD(VDD),.Y(g30809),.A(I40679));
  NOT NOT1_13197(.VSS(VSS),.VDD(VDD),.Y(I40682),.A(g30642));
  NOT NOT1_13198(.VSS(VSS),.VDD(VDD),.Y(g30810),.A(I40682));
  NOT NOT1_13199(.VSS(VSS),.VDD(VDD),.Y(I40685),.A(g30643));
  NOT NOT1_13200(.VSS(VSS),.VDD(VDD),.Y(g30811),.A(I40685));
  NOT NOT1_13201(.VSS(VSS),.VDD(VDD),.Y(I40688),.A(g30644));
  NOT NOT1_13202(.VSS(VSS),.VDD(VDD),.Y(g30812),.A(I40688));
  NOT NOT1_13203(.VSS(VSS),.VDD(VDD),.Y(I40691),.A(g30645));
  NOT NOT1_13204(.VSS(VSS),.VDD(VDD),.Y(g30813),.A(I40691));
  NOT NOT1_13205(.VSS(VSS),.VDD(VDD),.Y(I40694),.A(g30646));
  NOT NOT1_13206(.VSS(VSS),.VDD(VDD),.Y(g30814),.A(I40694));
  NOT NOT1_13207(.VSS(VSS),.VDD(VDD),.Y(I40697),.A(g30647));
  NOT NOT1_13208(.VSS(VSS),.VDD(VDD),.Y(g30815),.A(I40697));
  NOT NOT1_13209(.VSS(VSS),.VDD(VDD),.Y(I40700),.A(g30648));
  NOT NOT1_13210(.VSS(VSS),.VDD(VDD),.Y(g30816),.A(I40700));
  NOT NOT1_13211(.VSS(VSS),.VDD(VDD),.Y(I40703),.A(g30649));
  NOT NOT1_13212(.VSS(VSS),.VDD(VDD),.Y(g30817),.A(I40703));
  NOT NOT1_13213(.VSS(VSS),.VDD(VDD),.Y(I40706),.A(g30650));
  NOT NOT1_13214(.VSS(VSS),.VDD(VDD),.Y(g30818),.A(I40706));
  NOT NOT1_13215(.VSS(VSS),.VDD(VDD),.Y(I40709),.A(g30651));
  NOT NOT1_13216(.VSS(VSS),.VDD(VDD),.Y(g30819),.A(I40709));
  NOT NOT1_13217(.VSS(VSS),.VDD(VDD),.Y(I40712),.A(g30652));
  NOT NOT1_13218(.VSS(VSS),.VDD(VDD),.Y(g30820),.A(I40712));
  NOT NOT1_13219(.VSS(VSS),.VDD(VDD),.Y(I40715),.A(g30653));
  NOT NOT1_13220(.VSS(VSS),.VDD(VDD),.Y(g30821),.A(I40715));
  NOT NOT1_13221(.VSS(VSS),.VDD(VDD),.Y(I40718),.A(g30654));
  NOT NOT1_13222(.VSS(VSS),.VDD(VDD),.Y(g30822),.A(I40718));
  NOT NOT1_13223(.VSS(VSS),.VDD(VDD),.Y(I40721),.A(g30655));
  NOT NOT1_13224(.VSS(VSS),.VDD(VDD),.Y(g30823),.A(I40721));
  NOT NOT1_13225(.VSS(VSS),.VDD(VDD),.Y(I40724),.A(g30656));
  NOT NOT1_13226(.VSS(VSS),.VDD(VDD),.Y(g30824),.A(I40724));
  NOT NOT1_13227(.VSS(VSS),.VDD(VDD),.Y(I40727),.A(g30657));
  NOT NOT1_13228(.VSS(VSS),.VDD(VDD),.Y(g30825),.A(I40727));
  NOT NOT1_13229(.VSS(VSS),.VDD(VDD),.Y(I40730),.A(g30658));
  NOT NOT1_13230(.VSS(VSS),.VDD(VDD),.Y(g30826),.A(I40730));
  NOT NOT1_13231(.VSS(VSS),.VDD(VDD),.Y(I40733),.A(g30659));
  NOT NOT1_13232(.VSS(VSS),.VDD(VDD),.Y(g30827),.A(I40733));
  NOT NOT1_13233(.VSS(VSS),.VDD(VDD),.Y(I40736),.A(g30660));
  NOT NOT1_13234(.VSS(VSS),.VDD(VDD),.Y(g30828),.A(I40736));
  NOT NOT1_13235(.VSS(VSS),.VDD(VDD),.Y(I40739),.A(g30661));
  NOT NOT1_13236(.VSS(VSS),.VDD(VDD),.Y(g30829),.A(I40739));
  NOT NOT1_13237(.VSS(VSS),.VDD(VDD),.Y(I40742),.A(g30662));
  NOT NOT1_13238(.VSS(VSS),.VDD(VDD),.Y(g30830),.A(I40742));
  NOT NOT1_13239(.VSS(VSS),.VDD(VDD),.Y(I40745),.A(g30663));
  NOT NOT1_13240(.VSS(VSS),.VDD(VDD),.Y(g30831),.A(I40745));
  NOT NOT1_13241(.VSS(VSS),.VDD(VDD),.Y(I40748),.A(g30664));
  NOT NOT1_13242(.VSS(VSS),.VDD(VDD),.Y(g30832),.A(I40748));
  NOT NOT1_13243(.VSS(VSS),.VDD(VDD),.Y(I40751),.A(g30665));
  NOT NOT1_13244(.VSS(VSS),.VDD(VDD),.Y(g30833),.A(I40751));
  NOT NOT1_13245(.VSS(VSS),.VDD(VDD),.Y(I40754),.A(g30666));
  NOT NOT1_13246(.VSS(VSS),.VDD(VDD),.Y(g30834),.A(I40754));
  NOT NOT1_13247(.VSS(VSS),.VDD(VDD),.Y(I40757),.A(g30667));
  NOT NOT1_13248(.VSS(VSS),.VDD(VDD),.Y(g30835),.A(I40757));
  NOT NOT1_13249(.VSS(VSS),.VDD(VDD),.Y(I40760),.A(g30722));
  NOT NOT1_13250(.VSS(VSS),.VDD(VDD),.Y(g30836),.A(I40760));
  NOT NOT1_13251(.VSS(VSS),.VDD(VDD),.Y(I40763),.A(g30729));
  NOT NOT1_13252(.VSS(VSS),.VDD(VDD),.Y(g30837),.A(I40763));
  NOT NOT1_13253(.VSS(VSS),.VDD(VDD),.Y(I40766),.A(g30737));
  NOT NOT1_13254(.VSS(VSS),.VDD(VDD),.Y(g30838),.A(I40766));
  NOT NOT1_13255(.VSS(VSS),.VDD(VDD),.Y(I40769),.A(g30803));
  NOT NOT1_13256(.VSS(VSS),.VDD(VDD),.Y(g30839),.A(I40769));
  NOT NOT1_13257(.VSS(VSS),.VDD(VDD),.Y(I40772),.A(g30804));
  NOT NOT1_13258(.VSS(VSS),.VDD(VDD),.Y(g30840),.A(I40772));
  NOT NOT1_13259(.VSS(VSS),.VDD(VDD),.Y(I40775),.A(g30807));
  NOT NOT1_13260(.VSS(VSS),.VDD(VDD),.Y(g30841),.A(I40775));
  NOT NOT1_13261(.VSS(VSS),.VDD(VDD),.Y(I40778),.A(g30805));
  NOT NOT1_13262(.VSS(VSS),.VDD(VDD),.Y(g30842),.A(I40778));
  NOT NOT1_13263(.VSS(VSS),.VDD(VDD),.Y(I40781),.A(g30808));
  NOT NOT1_13264(.VSS(VSS),.VDD(VDD),.Y(g30843),.A(I40781));
  NOT NOT1_13265(.VSS(VSS),.VDD(VDD),.Y(I40784),.A(g30813));
  NOT NOT1_13266(.VSS(VSS),.VDD(VDD),.Y(g30844),.A(I40784));
  NOT NOT1_13267(.VSS(VSS),.VDD(VDD),.Y(I40787),.A(g30809));
  NOT NOT1_13268(.VSS(VSS),.VDD(VDD),.Y(g30845),.A(I40787));
  NOT NOT1_13269(.VSS(VSS),.VDD(VDD),.Y(I40790),.A(g30814));
  NOT NOT1_13270(.VSS(VSS),.VDD(VDD),.Y(g30846),.A(I40790));
  NOT NOT1_13271(.VSS(VSS),.VDD(VDD),.Y(I40793),.A(g30821));
  NOT NOT1_13272(.VSS(VSS),.VDD(VDD),.Y(g30847),.A(I40793));
  NOT NOT1_13273(.VSS(VSS),.VDD(VDD),.Y(I40796),.A(g30829));
  NOT NOT1_13274(.VSS(VSS),.VDD(VDD),.Y(g30848),.A(I40796));
  NOT NOT1_13275(.VSS(VSS),.VDD(VDD),.Y(I40799),.A(g30723));
  NOT NOT1_13276(.VSS(VSS),.VDD(VDD),.Y(g30849),.A(I40799));
  NOT NOT1_13277(.VSS(VSS),.VDD(VDD),.Y(I40802),.A(g30730));
  NOT NOT1_13278(.VSS(VSS),.VDD(VDD),.Y(g30850),.A(I40802));
  NOT NOT1_13279(.VSS(VSS),.VDD(VDD),.Y(I40805),.A(g30767));
  NOT NOT1_13280(.VSS(VSS),.VDD(VDD),.Y(g30851),.A(I40805));
  NOT NOT1_13281(.VSS(VSS),.VDD(VDD),.Y(I40808),.A(g30769));
  NOT NOT1_13282(.VSS(VSS),.VDD(VDD),.Y(g30852),.A(I40808));
  NOT NOT1_13283(.VSS(VSS),.VDD(VDD),.Y(I40811),.A(g30772));
  NOT NOT1_13284(.VSS(VSS),.VDD(VDD),.Y(g30853),.A(I40811));
  NOT NOT1_13285(.VSS(VSS),.VDD(VDD),.Y(I40814),.A(g30731));
  NOT NOT1_13286(.VSS(VSS),.VDD(VDD),.Y(g30854),.A(I40814));
  NOT NOT1_13287(.VSS(VSS),.VDD(VDD),.Y(I40817),.A(g30738));
  NOT NOT1_13288(.VSS(VSS),.VDD(VDD),.Y(g30855),.A(I40817));
  NOT NOT1_13289(.VSS(VSS),.VDD(VDD),.Y(I40820),.A(g30745));
  NOT NOT1_13290(.VSS(VSS),.VDD(VDD),.Y(g30856),.A(I40820));
  NOT NOT1_13291(.VSS(VSS),.VDD(VDD),.Y(I40823),.A(g30806));
  NOT NOT1_13292(.VSS(VSS),.VDD(VDD),.Y(g30857),.A(I40823));
  NOT NOT1_13293(.VSS(VSS),.VDD(VDD),.Y(I40826),.A(g30810));
  NOT NOT1_13294(.VSS(VSS),.VDD(VDD),.Y(g30858),.A(I40826));
  NOT NOT1_13295(.VSS(VSS),.VDD(VDD),.Y(I40829),.A(g30815));
  NOT NOT1_13296(.VSS(VSS),.VDD(VDD),.Y(g30859),.A(I40829));
  NOT NOT1_13297(.VSS(VSS),.VDD(VDD),.Y(I40832),.A(g30811));
  NOT NOT1_13298(.VSS(VSS),.VDD(VDD),.Y(g30860),.A(I40832));
  NOT NOT1_13299(.VSS(VSS),.VDD(VDD),.Y(I40835),.A(g30816));
  NOT NOT1_13300(.VSS(VSS),.VDD(VDD),.Y(g30861),.A(I40835));
  NOT NOT1_13301(.VSS(VSS),.VDD(VDD),.Y(I40838),.A(g30822));
  NOT NOT1_13302(.VSS(VSS),.VDD(VDD),.Y(g30862),.A(I40838));
  NOT NOT1_13303(.VSS(VSS),.VDD(VDD),.Y(I40841),.A(g30817));
  NOT NOT1_13304(.VSS(VSS),.VDD(VDD),.Y(g30863),.A(I40841));
  NOT NOT1_13305(.VSS(VSS),.VDD(VDD),.Y(I40844),.A(g30823));
  NOT NOT1_13306(.VSS(VSS),.VDD(VDD),.Y(g30864),.A(I40844));
  NOT NOT1_13307(.VSS(VSS),.VDD(VDD),.Y(I40847),.A(g30830));
  NOT NOT1_13308(.VSS(VSS),.VDD(VDD),.Y(g30865),.A(I40847));
  NOT NOT1_13309(.VSS(VSS),.VDD(VDD),.Y(I40850),.A(g30724));
  NOT NOT1_13310(.VSS(VSS),.VDD(VDD),.Y(g30866),.A(I40850));
  NOT NOT1_13311(.VSS(VSS),.VDD(VDD),.Y(I40853),.A(g30732));
  NOT NOT1_13312(.VSS(VSS),.VDD(VDD),.Y(g30867),.A(I40853));
  NOT NOT1_13313(.VSS(VSS),.VDD(VDD),.Y(I40856),.A(g30739));
  NOT NOT1_13314(.VSS(VSS),.VDD(VDD),.Y(g30868),.A(I40856));
  NOT NOT1_13315(.VSS(VSS),.VDD(VDD),.Y(I40859),.A(g30770));
  NOT NOT1_13316(.VSS(VSS),.VDD(VDD),.Y(g30869),.A(I40859));
  NOT NOT1_13317(.VSS(VSS),.VDD(VDD),.Y(I40862),.A(g30773));
  NOT NOT1_13318(.VSS(VSS),.VDD(VDD),.Y(g30870),.A(I40862));
  NOT NOT1_13319(.VSS(VSS),.VDD(VDD),.Y(I40865),.A(g30776));
  NOT NOT1_13320(.VSS(VSS),.VDD(VDD),.Y(g30871),.A(I40865));
  NOT NOT1_13321(.VSS(VSS),.VDD(VDD),.Y(I40868),.A(g30740));
  NOT NOT1_13322(.VSS(VSS),.VDD(VDD),.Y(g30872),.A(I40868));
  NOT NOT1_13323(.VSS(VSS),.VDD(VDD),.Y(I40871),.A(g30746));
  NOT NOT1_13324(.VSS(VSS),.VDD(VDD),.Y(g30873),.A(I40871));
  NOT NOT1_13325(.VSS(VSS),.VDD(VDD),.Y(I40874),.A(g30751));
  NOT NOT1_13326(.VSS(VSS),.VDD(VDD),.Y(g30874),.A(I40874));
  NOT NOT1_13327(.VSS(VSS),.VDD(VDD),.Y(I40877),.A(g30812));
  NOT NOT1_13328(.VSS(VSS),.VDD(VDD),.Y(g30875),.A(I40877));
  NOT NOT1_13329(.VSS(VSS),.VDD(VDD),.Y(I40880),.A(g30818));
  NOT NOT1_13330(.VSS(VSS),.VDD(VDD),.Y(g30876),.A(I40880));
  NOT NOT1_13331(.VSS(VSS),.VDD(VDD),.Y(I40883),.A(g30824));
  NOT NOT1_13332(.VSS(VSS),.VDD(VDD),.Y(g30877),.A(I40883));
  NOT NOT1_13333(.VSS(VSS),.VDD(VDD),.Y(I40886),.A(g30819));
  NOT NOT1_13334(.VSS(VSS),.VDD(VDD),.Y(g30878),.A(I40886));
  NOT NOT1_13335(.VSS(VSS),.VDD(VDD),.Y(I40889),.A(g30825));
  NOT NOT1_13336(.VSS(VSS),.VDD(VDD),.Y(g30879),.A(I40889));
  NOT NOT1_13337(.VSS(VSS),.VDD(VDD),.Y(I40892),.A(g30831));
  NOT NOT1_13338(.VSS(VSS),.VDD(VDD),.Y(g30880),.A(I40892));
  NOT NOT1_13339(.VSS(VSS),.VDD(VDD),.Y(I40895),.A(g30826));
  NOT NOT1_13340(.VSS(VSS),.VDD(VDD),.Y(g30881),.A(I40895));
  NOT NOT1_13341(.VSS(VSS),.VDD(VDD),.Y(I40898),.A(g30832));
  NOT NOT1_13342(.VSS(VSS),.VDD(VDD),.Y(g30882),.A(I40898));
  NOT NOT1_13343(.VSS(VSS),.VDD(VDD),.Y(I40901),.A(g30725));
  NOT NOT1_13344(.VSS(VSS),.VDD(VDD),.Y(g30883),.A(I40901));
  NOT NOT1_13345(.VSS(VSS),.VDD(VDD),.Y(I40904),.A(g30733));
  NOT NOT1_13346(.VSS(VSS),.VDD(VDD),.Y(g30884),.A(I40904));
  NOT NOT1_13347(.VSS(VSS),.VDD(VDD),.Y(I40907),.A(g30741));
  NOT NOT1_13348(.VSS(VSS),.VDD(VDD),.Y(g30885),.A(I40907));
  NOT NOT1_13349(.VSS(VSS),.VDD(VDD),.Y(I40910),.A(g30747));
  NOT NOT1_13350(.VSS(VSS),.VDD(VDD),.Y(g30886),.A(I40910));
  NOT NOT1_13351(.VSS(VSS),.VDD(VDD),.Y(I40913),.A(g30774));
  NOT NOT1_13352(.VSS(VSS),.VDD(VDD),.Y(g30887),.A(I40913));
  NOT NOT1_13353(.VSS(VSS),.VDD(VDD),.Y(I40916),.A(g30777));
  NOT NOT1_13354(.VSS(VSS),.VDD(VDD),.Y(g30888),.A(I40916));
  NOT NOT1_13355(.VSS(VSS),.VDD(VDD),.Y(I40919),.A(g30781));
  NOT NOT1_13356(.VSS(VSS),.VDD(VDD),.Y(g30889),.A(I40919));
  NOT NOT1_13357(.VSS(VSS),.VDD(VDD),.Y(I40922),.A(g30748));
  NOT NOT1_13358(.VSS(VSS),.VDD(VDD),.Y(g30890),.A(I40922));
  NOT NOT1_13359(.VSS(VSS),.VDD(VDD),.Y(I40925),.A(g30752));
  NOT NOT1_13360(.VSS(VSS),.VDD(VDD),.Y(g30891),.A(I40925));
  NOT NOT1_13361(.VSS(VSS),.VDD(VDD),.Y(I40928),.A(g30756));
  NOT NOT1_13362(.VSS(VSS),.VDD(VDD),.Y(g30892),.A(I40928));
  NOT NOT1_13363(.VSS(VSS),.VDD(VDD),.Y(I40931),.A(g30820));
  NOT NOT1_13364(.VSS(VSS),.VDD(VDD),.Y(g30893),.A(I40931));
  NOT NOT1_13365(.VSS(VSS),.VDD(VDD),.Y(I40934),.A(g30827));
  NOT NOT1_13366(.VSS(VSS),.VDD(VDD),.Y(g30894),.A(I40934));
  NOT NOT1_13367(.VSS(VSS),.VDD(VDD),.Y(I40937),.A(g30833));
  NOT NOT1_13368(.VSS(VSS),.VDD(VDD),.Y(g30895),.A(I40937));
  NOT NOT1_13369(.VSS(VSS),.VDD(VDD),.Y(I40940),.A(g30828));
  NOT NOT1_13370(.VSS(VSS),.VDD(VDD),.Y(g30896),.A(I40940));
  NOT NOT1_13371(.VSS(VSS),.VDD(VDD),.Y(I40943),.A(g30834));
  NOT NOT1_13372(.VSS(VSS),.VDD(VDD),.Y(g30897),.A(I40943));
  NOT NOT1_13373(.VSS(VSS),.VDD(VDD),.Y(I40946),.A(g30726));
  NOT NOT1_13374(.VSS(VSS),.VDD(VDD),.Y(g30898),.A(I40946));
  NOT NOT1_13375(.VSS(VSS),.VDD(VDD),.Y(I40949),.A(g30835));
  NOT NOT1_13376(.VSS(VSS),.VDD(VDD),.Y(g30899),.A(I40949));
  NOT NOT1_13377(.VSS(VSS),.VDD(VDD),.Y(I40952),.A(g30727));
  NOT NOT1_13378(.VSS(VSS),.VDD(VDD),.Y(g30900),.A(I40952));
  NOT NOT1_13379(.VSS(VSS),.VDD(VDD),.Y(I40955),.A(g30734));
  NOT NOT1_13380(.VSS(VSS),.VDD(VDD),.Y(g30901),.A(I40955));
  NOT NOT1_13381(.VSS(VSS),.VDD(VDD),.Y(I40958),.A(g30742));
  NOT NOT1_13382(.VSS(VSS),.VDD(VDD),.Y(g30902),.A(I40958));
  NOT NOT1_13383(.VSS(VSS),.VDD(VDD),.Y(I40961),.A(g30749));
  NOT NOT1_13384(.VSS(VSS),.VDD(VDD),.Y(g30903),.A(I40961));
  NOT NOT1_13385(.VSS(VSS),.VDD(VDD),.Y(I40964),.A(g30753));
  NOT NOT1_13386(.VSS(VSS),.VDD(VDD),.Y(g30904),.A(I40964));
  NOT NOT1_13387(.VSS(VSS),.VDD(VDD),.Y(I40967),.A(g30778));
  NOT NOT1_13388(.VSS(VSS),.VDD(VDD),.Y(g30905),.A(I40967));
  NOT NOT1_13389(.VSS(VSS),.VDD(VDD),.Y(I40970),.A(g30782));
  NOT NOT1_13390(.VSS(VSS),.VDD(VDD),.Y(g30906),.A(I40970));
  NOT NOT1_13391(.VSS(VSS),.VDD(VDD),.Y(I40973),.A(g30784));
  NOT NOT1_13392(.VSS(VSS),.VDD(VDD),.Y(g30907),.A(I40973));
  NOT NOT1_13393(.VSS(VSS),.VDD(VDD),.Y(I40976),.A(g30799));
  NOT NOT1_13394(.VSS(VSS),.VDD(VDD),.Y(g30908),.A(I40976));
  NOT NOT1_13395(.VSS(VSS),.VDD(VDD),.Y(I40979),.A(g30800));
  NOT NOT1_13396(.VSS(VSS),.VDD(VDD),.Y(g30909),.A(I40979));
  NOT NOT1_13397(.VSS(VSS),.VDD(VDD),.Y(I40982),.A(g30802));
  NOT NOT1_13398(.VSS(VSS),.VDD(VDD),.Y(g30910),.A(I40982));
  NOT NOT1_13399(.VSS(VSS),.VDD(VDD),.Y(I40985),.A(g30792));
  NOT NOT1_13400(.VSS(VSS),.VDD(VDD),.Y(g30911),.A(I40985));
  NOT NOT1_13401(.VSS(VSS),.VDD(VDD),.Y(I40988),.A(g30793));
  NOT NOT1_13402(.VSS(VSS),.VDD(VDD),.Y(g30912),.A(I40988));
  NOT NOT1_13403(.VSS(VSS),.VDD(VDD),.Y(I40991),.A(g30794));
  NOT NOT1_13404(.VSS(VSS),.VDD(VDD),.Y(g30913),.A(I40991));
  NOT NOT1_13405(.VSS(VSS),.VDD(VDD),.Y(I40994),.A(g30795));
  NOT NOT1_13406(.VSS(VSS),.VDD(VDD),.Y(g30914),.A(I40994));
  NOT NOT1_13407(.VSS(VSS),.VDD(VDD),.Y(I40997),.A(g30797));
  NOT NOT1_13408(.VSS(VSS),.VDD(VDD),.Y(g30915),.A(I40997));
  NOT NOT1_13409(.VSS(VSS),.VDD(VDD),.Y(I41024),.A(g30765));
  NOT NOT1_13410(.VSS(VSS),.VDD(VDD),.Y(g30928),.A(I41024));
  NOT NOT1_13411(.VSS(VSS),.VDD(VDD),.Y(I41035),.A(g30796));
  NOT NOT1_13412(.VSS(VSS),.VDD(VDD),.Y(g30937),.A(I41035));
  NOT NOT1_13413(.VSS(VSS),.VDD(VDD),.Y(I41038),.A(g30798));
  NOT NOT1_13414(.VSS(VSS),.VDD(VDD),.Y(g30938),.A(I41038));
  NOT NOT1_13415(.VSS(VSS),.VDD(VDD),.Y(I41041),.A(g30801));
  NOT NOT1_13416(.VSS(VSS),.VDD(VDD),.Y(g30939),.A(I41041));
  NOT NOT1_13417(.VSS(VSS),.VDD(VDD),.Y(I41044),.A(g30928));
  NOT NOT1_13418(.VSS(VSS),.VDD(VDD),.Y(g30940),.A(I41044));
  NOT NOT1_13419(.VSS(VSS),.VDD(VDD),.Y(I41047),.A(g30937));
  NOT NOT1_13420(.VSS(VSS),.VDD(VDD),.Y(g30941),.A(I41047));
  NOT NOT1_13421(.VSS(VSS),.VDD(VDD),.Y(I41050),.A(g30938));
  NOT NOT1_13422(.VSS(VSS),.VDD(VDD),.Y(g30942),.A(I41050));
  NOT NOT1_13423(.VSS(VSS),.VDD(VDD),.Y(I41053),.A(g30939));
  NOT NOT1_13424(.VSS(VSS),.VDD(VDD),.Y(g30943),.A(I41053));
  NOT NOT1_13425(.VSS(VSS),.VDD(VDD),.Y(g30962),.A(g30958));
  NOT NOT1_13426(.VSS(VSS),.VDD(VDD),.Y(g30963),.A(g30957));
  NOT NOT1_13427(.VSS(VSS),.VDD(VDD),.Y(g30964),.A(g30961));
  NOT NOT1_13428(.VSS(VSS),.VDD(VDD),.Y(g30965),.A(g30959));
  NOT NOT1_13429(.VSS(VSS),.VDD(VDD),.Y(g30966),.A(g30956));
  NOT NOT1_13430(.VSS(VSS),.VDD(VDD),.Y(g30967),.A(g30954));
  NOT NOT1_13431(.VSS(VSS),.VDD(VDD),.Y(g30968),.A(g30960));
  NOT NOT1_13432(.VSS(VSS),.VDD(VDD),.Y(g30969),.A(g30955));
  NOT NOT1_13433(.VSS(VSS),.VDD(VDD),.Y(g30971),.A(g30970));
  NOT NOT1_13434(.VSS(VSS),.VDD(VDD),.Y(I41090),.A(g30965));
  NOT NOT1_13435(.VSS(VSS),.VDD(VDD),.Y(g30972),.A(I41090));
  NOT NOT1_13436(.VSS(VSS),.VDD(VDD),.Y(I41093),.A(g30964));
  NOT NOT1_13437(.VSS(VSS),.VDD(VDD),.Y(g30973),.A(I41093));
  NOT NOT1_13438(.VSS(VSS),.VDD(VDD),.Y(I41096),.A(g30963));
  NOT NOT1_13439(.VSS(VSS),.VDD(VDD),.Y(g30974),.A(I41096));
  NOT NOT1_13440(.VSS(VSS),.VDD(VDD),.Y(I41099),.A(g30962));
  NOT NOT1_13441(.VSS(VSS),.VDD(VDD),.Y(g30975),.A(I41099));
  NOT NOT1_13442(.VSS(VSS),.VDD(VDD),.Y(I41102),.A(g30969));
  NOT NOT1_13443(.VSS(VSS),.VDD(VDD),.Y(g30976),.A(I41102));
  NOT NOT1_13444(.VSS(VSS),.VDD(VDD),.Y(I41105),.A(g30968));
  NOT NOT1_13445(.VSS(VSS),.VDD(VDD),.Y(g30977),.A(I41105));
  NOT NOT1_13446(.VSS(VSS),.VDD(VDD),.Y(I41108),.A(g30967));
  NOT NOT1_13447(.VSS(VSS),.VDD(VDD),.Y(g30978),.A(I41108));
  NOT NOT1_13448(.VSS(VSS),.VDD(VDD),.Y(I41111),.A(g30966));
  NOT NOT1_13449(.VSS(VSS),.VDD(VDD),.Y(g30979),.A(I41111));
  NOT NOT1_13450(.VSS(VSS),.VDD(VDD),.Y(I41114),.A(g30976));
  NOT NOT1_13451(.VSS(VSS),.VDD(VDD),.Y(g30980),.A(I41114));
  NOT NOT1_13452(.VSS(VSS),.VDD(VDD),.Y(I41117),.A(g30977));
  NOT NOT1_13453(.VSS(VSS),.VDD(VDD),.Y(g30981),.A(I41117));
  NOT NOT1_13454(.VSS(VSS),.VDD(VDD),.Y(I41120),.A(g30978));
  NOT NOT1_13455(.VSS(VSS),.VDD(VDD),.Y(g30982),.A(I41120));
  NOT NOT1_13456(.VSS(VSS),.VDD(VDD),.Y(I41123),.A(g30979));
  NOT NOT1_13457(.VSS(VSS),.VDD(VDD),.Y(g30983),.A(I41123));
  NOT NOT1_13458(.VSS(VSS),.VDD(VDD),.Y(I41126),.A(g30972));
  NOT NOT1_13459(.VSS(VSS),.VDD(VDD),.Y(g30984),.A(I41126));
  NOT NOT1_13460(.VSS(VSS),.VDD(VDD),.Y(I41129),.A(g30973));
  NOT NOT1_13461(.VSS(VSS),.VDD(VDD),.Y(g30985),.A(I41129));
  NOT NOT1_13462(.VSS(VSS),.VDD(VDD),.Y(I41132),.A(g30974));
  NOT NOT1_13463(.VSS(VSS),.VDD(VDD),.Y(g30986),.A(I41132));
  NOT NOT1_13464(.VSS(VSS),.VDD(VDD),.Y(I41135),.A(g30975));
  NOT NOT1_13465(.VSS(VSS),.VDD(VDD),.Y(g30987),.A(I41135));
  NOT NOT1_13466(.VSS(VSS),.VDD(VDD),.Y(I41138),.A(g30971));
  NOT NOT1_13467(.VSS(VSS),.VDD(VDD),.Y(g30988),.A(I41138));
  NOT NOT1_13468(.VSS(VSS),.VDD(VDD),.Y(I41141),.A(g30988));
  NOT NOT1_13469(.VSS(VSS),.VDD(VDD),.Y(g30989),.A(I41141));
//
  AND2 AND2_0(.VSS(VSS),.VDD(VDD),.Y(g5630),.A(g325),.B(g349));
  AND2 AND2_1(.VSS(VSS),.VDD(VDD),.Y(g5649),.A(g331),.B(g351));
  AND2 AND2_2(.VSS(VSS),.VDD(VDD),.Y(g5650),.A(g325),.B(g364));
  AND2 AND2_3(.VSS(VSS),.VDD(VDD),.Y(g5658),.A(g1012),.B(g1036));
  AND2 AND2_4(.VSS(VSS),.VDD(VDD),.Y(g5676),.A(g337),.B(g353));
  AND2 AND2_5(.VSS(VSS),.VDD(VDD),.Y(g5677),.A(g331),.B(g366));
  AND2 AND2_6(.VSS(VSS),.VDD(VDD),.Y(g5678),.A(g325),.B(g379));
  AND2 AND2_7(.VSS(VSS),.VDD(VDD),.Y(g5687),.A(g1018),.B(g1038));
  AND2 AND2_8(.VSS(VSS),.VDD(VDD),.Y(g5688),.A(g1012),.B(g1051));
  AND2 AND2_9(.VSS(VSS),.VDD(VDD),.Y(g5696),.A(g1706),.B(g1730));
  AND2 AND2_10(.VSS(VSS),.VDD(VDD),.Y(g5709),.A(g337),.B(g368));
  AND2 AND2_11(.VSS(VSS),.VDD(VDD),.Y(g5710),.A(g331),.B(g381));
  AND2 AND2_12(.VSS(VSS),.VDD(VDD),.Y(g5711),.A(g325),.B(g394));
  AND2 AND2_13(.VSS(VSS),.VDD(VDD),.Y(g5728),.A(g1024),.B(g1040));
  AND2 AND2_14(.VSS(VSS),.VDD(VDD),.Y(g5729),.A(g1018),.B(g1053));
  AND2 AND2_15(.VSS(VSS),.VDD(VDD),.Y(g5730),.A(g1012),.B(g1066));
  AND2 AND2_16(.VSS(VSS),.VDD(VDD),.Y(g5739),.A(g1712),.B(g1732));
  AND2 AND2_17(.VSS(VSS),.VDD(VDD),.Y(g5740),.A(g1706),.B(g1745));
  AND2 AND2_18(.VSS(VSS),.VDD(VDD),.Y(g5748),.A(g2400),.B(g2424));
  AND2 AND2_19(.VSS(VSS),.VDD(VDD),.Y(g5757),.A(g337),.B(g383));
  AND2 AND2_20(.VSS(VSS),.VDD(VDD),.Y(g5758),.A(g331),.B(g396));
  AND2 AND2_21(.VSS(VSS),.VDD(VDD),.Y(g5767),.A(g1024),.B(g1055));
  AND2 AND2_22(.VSS(VSS),.VDD(VDD),.Y(g5768),.A(g1018),.B(g1068));
  AND2 AND2_23(.VSS(VSS),.VDD(VDD),.Y(g5769),.A(g1012),.B(g1081));
  AND2 AND2_24(.VSS(VSS),.VDD(VDD),.Y(g5786),.A(g1718),.B(g1734));
  AND2 AND2_25(.VSS(VSS),.VDD(VDD),.Y(g5787),.A(g1712),.B(g1747));
  AND2 AND2_26(.VSS(VSS),.VDD(VDD),.Y(g5788),.A(g1706),.B(g1760));
  AND2 AND2_27(.VSS(VSS),.VDD(VDD),.Y(g5797),.A(g2406),.B(g2426));
  AND2 AND2_28(.VSS(VSS),.VDD(VDD),.Y(g5798),.A(g2400),.B(g2439));
  AND2 AND2_29(.VSS(VSS),.VDD(VDD),.Y(g5807),.A(g337),.B(g324));
  AND2 AND2_30(.VSS(VSS),.VDD(VDD),.Y(g5816),.A(g1024),.B(g1070));
  AND2 AND2_31(.VSS(VSS),.VDD(VDD),.Y(g5817),.A(g1018),.B(g1083));
  AND2 AND2_32(.VSS(VSS),.VDD(VDD),.Y(g5826),.A(g1718),.B(g1749));
  AND2 AND2_33(.VSS(VSS),.VDD(VDD),.Y(g5827),.A(g1712),.B(g1762));
  AND2 AND2_34(.VSS(VSS),.VDD(VDD),.Y(g5828),.A(g1706),.B(g1775));
  AND2 AND2_35(.VSS(VSS),.VDD(VDD),.Y(g5845),.A(g2412),.B(g2428));
  AND2 AND2_36(.VSS(VSS),.VDD(VDD),.Y(g5846),.A(g2406),.B(g2441));
  AND2 AND2_37(.VSS(VSS),.VDD(VDD),.Y(g5847),.A(g2400),.B(g2454));
  AND2 AND2_38(.VSS(VSS),.VDD(VDD),.Y(g5863),.A(g1024),.B(g1011));
  AND2 AND2_39(.VSS(VSS),.VDD(VDD),.Y(g5872),.A(g1718),.B(g1764));
  AND2 AND2_40(.VSS(VSS),.VDD(VDD),.Y(g5873),.A(g1712),.B(g1777));
  AND2 AND2_41(.VSS(VSS),.VDD(VDD),.Y(g5882),.A(g2412),.B(g2443));
  AND2 AND2_42(.VSS(VSS),.VDD(VDD),.Y(g5883),.A(g2406),.B(g2456));
  AND2 AND2_43(.VSS(VSS),.VDD(VDD),.Y(g5884),.A(g2400),.B(g2469));
  AND2 AND2_44(.VSS(VSS),.VDD(VDD),.Y(g5910),.A(g1718),.B(g1705));
  AND2 AND2_45(.VSS(VSS),.VDD(VDD),.Y(g5919),.A(g2412),.B(g2458));
  AND2 AND2_46(.VSS(VSS),.VDD(VDD),.Y(g5920),.A(g2406),.B(g2471));
  AND2 AND2_47(.VSS(VSS),.VDD(VDD),.Y(g5949),.A(g2412),.B(g2399));
  AND2 AND2_48(.VSS(VSS),.VDD(VDD),.Y(g8327),.A(g3254),.B(g219));
  AND2 AND2_49(.VSS(VSS),.VDD(VDD),.Y(g8328),.A(g6314),.B(g225));
  AND2 AND2_50(.VSS(VSS),.VDD(VDD),.Y(g8329),.A(g6232),.B(g231));
  AND2 AND2_51(.VSS(VSS),.VDD(VDD),.Y(g8339),.A(g6519),.B(g903));
  AND2 AND2_52(.VSS(VSS),.VDD(VDD),.Y(g8340),.A(g6369),.B(g909));
  AND2 AND2_53(.VSS(VSS),.VDD(VDD),.Y(g8350),.A(g6574),.B(g1594));
  AND2 AND2_54(.VSS(VSS),.VDD(VDD),.Y(g8385),.A(g3254),.B(g228));
  AND2 AND2_55(.VSS(VSS),.VDD(VDD),.Y(g8386),.A(g6314),.B(g234));
  AND2 AND2_56(.VSS(VSS),.VDD(VDD),.Y(g8387),.A(g6232),.B(g240));
  AND2 AND2_57(.VSS(VSS),.VDD(VDD),.Y(g8394),.A(g3410),.B(g906));
  AND2 AND2_58(.VSS(VSS),.VDD(VDD),.Y(g8395),.A(g6519),.B(g912));
  AND2 AND2_59(.VSS(VSS),.VDD(VDD),.Y(g8396),.A(g6369),.B(g918));
  AND2 AND2_60(.VSS(VSS),.VDD(VDD),.Y(g8406),.A(g6783),.B(g1597));
  AND2 AND2_61(.VSS(VSS),.VDD(VDD),.Y(g8407),.A(g6574),.B(g1603));
  AND2 AND2_62(.VSS(VSS),.VDD(VDD),.Y(g8417),.A(g6838),.B(g2288));
  AND2 AND2_63(.VSS(VSS),.VDD(VDD),.Y(g8431),.A(g3254),.B(g237));
  AND2 AND2_64(.VSS(VSS),.VDD(VDD),.Y(g8432),.A(g6314),.B(g243));
  AND2 AND2_65(.VSS(VSS),.VDD(VDD),.Y(g8433),.A(g6232),.B(g249));
  AND2 AND2_66(.VSS(VSS),.VDD(VDD),.Y(g8437),.A(g3410),.B(g915));
  AND2 AND2_67(.VSS(VSS),.VDD(VDD),.Y(g8438),.A(g6519),.B(g921));
  AND2 AND2_68(.VSS(VSS),.VDD(VDD),.Y(g8439),.A(g6369),.B(g927));
  AND2 AND2_69(.VSS(VSS),.VDD(VDD),.Y(g8446),.A(g3566),.B(g1600));
  AND2 AND2_70(.VSS(VSS),.VDD(VDD),.Y(g8447),.A(g6783),.B(g1606));
  AND2 AND2_71(.VSS(VSS),.VDD(VDD),.Y(g8448),.A(g6574),.B(g1612));
  AND2 AND2_72(.VSS(VSS),.VDD(VDD),.Y(g8458),.A(g7085),.B(g2291));
  AND2 AND2_73(.VSS(VSS),.VDD(VDD),.Y(g8459),.A(g6838),.B(g2297));
  AND2 AND2_74(.VSS(VSS),.VDD(VDD),.Y(g8463),.A(g3254),.B(g246));
  AND2 AND2_75(.VSS(VSS),.VDD(VDD),.Y(g8464),.A(g6314),.B(g252));
  AND2 AND2_76(.VSS(VSS),.VDD(VDD),.Y(g8465),.A(g6232),.B(g258));
  AND2 AND2_77(.VSS(VSS),.VDD(VDD),.Y(g8466),.A(g3410),.B(g924));
  AND2 AND2_78(.VSS(VSS),.VDD(VDD),.Y(g8467),.A(g6519),.B(g930));
  AND2 AND2_79(.VSS(VSS),.VDD(VDD),.Y(g8468),.A(g6369),.B(g936));
  AND2 AND2_80(.VSS(VSS),.VDD(VDD),.Y(g8472),.A(g3566),.B(g1609));
  AND2 AND2_81(.VSS(VSS),.VDD(VDD),.Y(g8473),.A(g6783),.B(g1615));
  AND2 AND2_82(.VSS(VSS),.VDD(VDD),.Y(g8474),.A(g6574),.B(g1621));
  AND2 AND2_83(.VSS(VSS),.VDD(VDD),.Y(g8481),.A(g3722),.B(g2294));
  AND2 AND2_84(.VSS(VSS),.VDD(VDD),.Y(g8482),.A(g7085),.B(g2300));
  AND2 AND2_85(.VSS(VSS),.VDD(VDD),.Y(g8483),.A(g6838),.B(g2306));
  AND2 AND2_86(.VSS(VSS),.VDD(VDD),.Y(g8484),.A(g6232),.B(g186));
  AND2 AND2_87(.VSS(VSS),.VDD(VDD),.Y(g8485),.A(g3254),.B(g255));
  AND2 AND2_88(.VSS(VSS),.VDD(VDD),.Y(g8486),.A(g6314),.B(g261));
  AND2 AND2_89(.VSS(VSS),.VDD(VDD),.Y(g8487),.A(g6232),.B(g267));
  AND2 AND2_90(.VSS(VSS),.VDD(VDD),.Y(g8488),.A(g3410),.B(g933));
  AND2 AND2_91(.VSS(VSS),.VDD(VDD),.Y(g8489),.A(g6519),.B(g939));
  AND2 AND2_92(.VSS(VSS),.VDD(VDD),.Y(g8490),.A(g6369),.B(g945));
  AND2 AND2_93(.VSS(VSS),.VDD(VDD),.Y(g8491),.A(g3566),.B(g1618));
  AND2 AND2_94(.VSS(VSS),.VDD(VDD),.Y(g8492),.A(g6783),.B(g1624));
  AND2 AND2_95(.VSS(VSS),.VDD(VDD),.Y(g8493),.A(g6574),.B(g1630));
  AND2 AND2_96(.VSS(VSS),.VDD(VDD),.Y(g8497),.A(g3722),.B(g2303));
  AND2 AND2_97(.VSS(VSS),.VDD(VDD),.Y(g8498),.A(g7085),.B(g2309));
  AND2 AND2_98(.VSS(VSS),.VDD(VDD),.Y(g8499),.A(g6838),.B(g2315));
  AND2 AND2_99(.VSS(VSS),.VDD(VDD),.Y(g8500),.A(g6314),.B(g189));
  AND2 AND2_100(.VSS(VSS),.VDD(VDD),.Y(g8501),.A(g6232),.B(g195));
  AND2 AND2_101(.VSS(VSS),.VDD(VDD),.Y(g8502),.A(g3254),.B(g264));
  AND2 AND2_102(.VSS(VSS),.VDD(VDD),.Y(g8503),.A(g6314),.B(g270));
  AND2 AND2_103(.VSS(VSS),.VDD(VDD),.Y(g8504),.A(g6369),.B(g873));
  AND2 AND2_104(.VSS(VSS),.VDD(VDD),.Y(g8505),.A(g3410),.B(g942));
  AND2 AND2_105(.VSS(VSS),.VDD(VDD),.Y(g8506),.A(g6519),.B(g948));
  AND2 AND2_106(.VSS(VSS),.VDD(VDD),.Y(g8507),.A(g6369),.B(g954));
  AND2 AND2_107(.VSS(VSS),.VDD(VDD),.Y(g8508),.A(g3566),.B(g1627));
  AND2 AND2_108(.VSS(VSS),.VDD(VDD),.Y(g8509),.A(g6783),.B(g1633));
  AND2 AND2_109(.VSS(VSS),.VDD(VDD),.Y(g8510),.A(g6574),.B(g1639));
  AND2 AND2_110(.VSS(VSS),.VDD(VDD),.Y(g8511),.A(g3722),.B(g2312));
  AND2 AND2_111(.VSS(VSS),.VDD(VDD),.Y(g8512),.A(g7085),.B(g2318));
  AND2 AND2_112(.VSS(VSS),.VDD(VDD),.Y(g8513),.A(g6838),.B(g2324));
  AND2 AND2_113(.VSS(VSS),.VDD(VDD),.Y(g8515),.A(g3254),.B(g192));
  AND2 AND2_114(.VSS(VSS),.VDD(VDD),.Y(g8516),.A(g6314),.B(g198));
  AND2 AND2_115(.VSS(VSS),.VDD(VDD),.Y(g8517),.A(g6232),.B(g204));
  AND2 AND2_116(.VSS(VSS),.VDD(VDD),.Y(g8518),.A(g3254),.B(g273));
  AND2 AND2_117(.VSS(VSS),.VDD(VDD),.Y(g8519),.A(g6519),.B(g876));
  AND2 AND2_118(.VSS(VSS),.VDD(VDD),.Y(g8520),.A(g6369),.B(g882));
  AND2 AND2_119(.VSS(VSS),.VDD(VDD),.Y(g8521),.A(g3410),.B(g951));
  AND2 AND2_120(.VSS(VSS),.VDD(VDD),.Y(g8522),.A(g6519),.B(g957));
  AND2 AND2_121(.VSS(VSS),.VDD(VDD),.Y(g8523),.A(g6574),.B(g1567));
  AND2 AND2_122(.VSS(VSS),.VDD(VDD),.Y(g8524),.A(g3566),.B(g1636));
  AND2 AND2_123(.VSS(VSS),.VDD(VDD),.Y(g8525),.A(g6783),.B(g1642));
  AND2 AND2_124(.VSS(VSS),.VDD(VDD),.Y(g8526),.A(g6574),.B(g1648));
  AND2 AND2_125(.VSS(VSS),.VDD(VDD),.Y(g8527),.A(g3722),.B(g2321));
  AND2 AND2_126(.VSS(VSS),.VDD(VDD),.Y(g8528),.A(g7085),.B(g2327));
  AND2 AND2_127(.VSS(VSS),.VDD(VDD),.Y(g8529),.A(g6838),.B(g2333));
  AND2 AND2_128(.VSS(VSS),.VDD(VDD),.Y(g8531),.A(g3254),.B(g201));
  AND2 AND2_129(.VSS(VSS),.VDD(VDD),.Y(g8532),.A(g6314),.B(g207));
  AND2 AND2_130(.VSS(VSS),.VDD(VDD),.Y(g8534),.A(g3410),.B(g879));
  AND2 AND2_131(.VSS(VSS),.VDD(VDD),.Y(g8535),.A(g6519),.B(g885));
  AND2 AND2_132(.VSS(VSS),.VDD(VDD),.Y(g8536),.A(g6369),.B(g891));
  AND2 AND2_133(.VSS(VSS),.VDD(VDD),.Y(g8537),.A(g3410),.B(g960));
  AND2 AND2_134(.VSS(VSS),.VDD(VDD),.Y(g8538),.A(g6783),.B(g1570));
  AND2 AND2_135(.VSS(VSS),.VDD(VDD),.Y(g8539),.A(g6574),.B(g1576));
  AND2 AND2_136(.VSS(VSS),.VDD(VDD),.Y(g8540),.A(g3566),.B(g1645));
  AND2 AND2_137(.VSS(VSS),.VDD(VDD),.Y(g8541),.A(g6783),.B(g1651));
  AND2 AND2_138(.VSS(VSS),.VDD(VDD),.Y(g8542),.A(g6838),.B(g2261));
  AND2 AND2_139(.VSS(VSS),.VDD(VDD),.Y(g8543),.A(g3722),.B(g2330));
  AND2 AND2_140(.VSS(VSS),.VDD(VDD),.Y(g8544),.A(g7085),.B(g2336));
  AND2 AND2_141(.VSS(VSS),.VDD(VDD),.Y(g8545),.A(g6838),.B(g2342));
  AND2 AND2_142(.VSS(VSS),.VDD(VDD),.Y(g8546),.A(g3254),.B(g210));
  AND2 AND2_143(.VSS(VSS),.VDD(VDD),.Y(g8548),.A(g3410),.B(g888));
  AND2 AND2_144(.VSS(VSS),.VDD(VDD),.Y(g8549),.A(g6519),.B(g894));
  AND2 AND2_145(.VSS(VSS),.VDD(VDD),.Y(g8551),.A(g3566),.B(g1573));
  AND2 AND2_146(.VSS(VSS),.VDD(VDD),.Y(g8552),.A(g6783),.B(g1579));
  AND2 AND2_147(.VSS(VSS),.VDD(VDD),.Y(g8553),.A(g6574),.B(g1585));
  AND2 AND2_148(.VSS(VSS),.VDD(VDD),.Y(g8554),.A(g3566),.B(g1654));
  AND2 AND2_149(.VSS(VSS),.VDD(VDD),.Y(g8555),.A(g7085),.B(g2264));
  AND2 AND2_150(.VSS(VSS),.VDD(VDD),.Y(g8556),.A(g6838),.B(g2270));
  AND2 AND2_151(.VSS(VSS),.VDD(VDD),.Y(g8557),.A(g3722),.B(g2339));
  AND2 AND2_152(.VSS(VSS),.VDD(VDD),.Y(g8558),.A(g7085),.B(g2345));
  AND2 AND2_153(.VSS(VSS),.VDD(VDD),.Y(g8559),.A(g3410),.B(g897));
  AND2 AND2_154(.VSS(VSS),.VDD(VDD),.Y(g8561),.A(g3566),.B(g1582));
  AND2 AND2_155(.VSS(VSS),.VDD(VDD),.Y(g8562),.A(g6783),.B(g1588));
  AND2 AND2_156(.VSS(VSS),.VDD(VDD),.Y(g8564),.A(g3722),.B(g2267));
  AND2 AND2_157(.VSS(VSS),.VDD(VDD),.Y(g8565),.A(g7085),.B(g2273));
  AND2 AND2_158(.VSS(VSS),.VDD(VDD),.Y(g8566),.A(g6838),.B(g2279));
  AND2 AND2_159(.VSS(VSS),.VDD(VDD),.Y(g8567),.A(g3722),.B(g2348));
  AND2 AND2_160(.VSS(VSS),.VDD(VDD),.Y(g8570),.A(g3566),.B(g1591));
  AND2 AND2_161(.VSS(VSS),.VDD(VDD),.Y(g8572),.A(g3722),.B(g2276));
  AND2 AND2_162(.VSS(VSS),.VDD(VDD),.Y(g8573),.A(g7085),.B(g2282));
  AND2 AND2_163(.VSS(VSS),.VDD(VDD),.Y(g8576),.A(g3722),.B(g2285));
  AND2 AND2_164(.VSS(VSS),.VDD(VDD),.Y(g8601),.A(g6643),.B(g7153));
  AND2 AND2_165(.VSS(VSS),.VDD(VDD),.Y(g8612),.A(g3338),.B(g6908));
  AND2 AND2_166(.VSS(VSS),.VDD(VDD),.Y(g8613),.A(g6945),.B(g7349));
  AND2 AND2_167(.VSS(VSS),.VDD(VDD),.Y(g8621),.A(g6486),.B(g6672));
  AND2 AND2_168(.VSS(VSS),.VDD(VDD),.Y(g8625),.A(g3494),.B(g7158));
  AND2 AND2_169(.VSS(VSS),.VDD(VDD),.Y(g8626),.A(g7195),.B(g7479));
  AND2 AND2_170(.VSS(VSS),.VDD(VDD),.Y(g8631),.A(g6751),.B(g6974));
  AND2 AND2_171(.VSS(VSS),.VDD(VDD),.Y(g8635),.A(g3650),.B(g7354));
  AND2 AND2_172(.VSS(VSS),.VDD(VDD),.Y(g8636),.A(g7391),.B(g7535));
  AND2 AND2_173(.VSS(VSS),.VDD(VDD),.Y(g8650),.A(g7053),.B(g7224));
  AND2 AND2_174(.VSS(VSS),.VDD(VDD),.Y(g8654),.A(g3806),.B(g7484));
  AND2 AND2_175(.VSS(VSS),.VDD(VDD),.Y(g8666),.A(g7303),.B(g7420));
  AND2 AND2_176(.VSS(VSS),.VDD(VDD),.Y(g8676),.A(g6643),.B(g7838));
  AND2 AND2_177(.VSS(VSS),.VDD(VDD),.Y(g8687),.A(g3338),.B(g7827));
  AND2 AND2_178(.VSS(VSS),.VDD(VDD),.Y(g8688),.A(g6945),.B(g7858));
  AND2 AND2_179(.VSS(VSS),.VDD(VDD),.Y(g8703),.A(g6486),.B(g7819));
  AND2 AND2_180(.VSS(VSS),.VDD(VDD),.Y(g8704),.A(g6643),.B(g7996));
  AND2 AND2_181(.VSS(VSS),.VDD(VDD),.Y(g8705),.A(g3494),.B(g7842));
  AND2 AND2_182(.VSS(VSS),.VDD(VDD),.Y(g8706),.A(g7195),.B(g7888));
  AND2 AND2_183(.VSS(VSS),.VDD(VDD),.Y(g8717),.A(g3338),.B(g7953));
  AND2 AND2_184(.VSS(VSS),.VDD(VDD),.Y(g8722),.A(g6751),.B(g7830));
  AND2 AND2_185(.VSS(VSS),.VDD(VDD),.Y(g8723),.A(g6945),.B(g8071));
  AND2 AND2_186(.VSS(VSS),.VDD(VDD),.Y(g8724),.A(g3650),.B(g7862));
  AND2 AND2_187(.VSS(VSS),.VDD(VDD),.Y(g8725),.A(g7391),.B(g7912));
  AND2 AND2_188(.VSS(VSS),.VDD(VDD),.Y(g8751),.A(g6486),.B(g7906));
  AND2 AND2_189(.VSS(VSS),.VDD(VDD),.Y(g8755),.A(g3494),.B(g8004));
  AND2 AND2_190(.VSS(VSS),.VDD(VDD),.Y(g8760),.A(g7053),.B(g7845));
  AND2 AND2_191(.VSS(VSS),.VDD(VDD),.Y(g8761),.A(g7195),.B(g8156));
  AND2 AND2_192(.VSS(VSS),.VDD(VDD),.Y(g8762),.A(g3806),.B(g7892));
  AND2 AND2_193(.VSS(VSS),.VDD(VDD),.Y(g8774),.A(g6751),.B(g7958));
  AND2 AND2_194(.VSS(VSS),.VDD(VDD),.Y(g8778),.A(g3650),.B(g8079));
  AND2 AND2_195(.VSS(VSS),.VDD(VDD),.Y(g8783),.A(g7303),.B(g7865));
  AND2 AND2_196(.VSS(VSS),.VDD(VDD),.Y(g8784),.A(g7391),.B(g8242));
  AND2 AND2_197(.VSS(VSS),.VDD(VDD),.Y(g8797),.A(g7053),.B(g8009));
  AND2 AND2_198(.VSS(VSS),.VDD(VDD),.Y(g8801),.A(g3806),.B(g8164));
  AND2 AND2_199(.VSS(VSS),.VDD(VDD),.Y(g8816),.A(g7303),.B(g8084));
  AND2 AND2_200(.VSS(VSS),.VDD(VDD),.Y(g8841),.A(g6486),.B(g490));
  AND2 AND2_201(.VSS(VSS),.VDD(VDD),.Y(g8842),.A(g6512),.B(g5508));
  AND2 AND2_202(.VSS(VSS),.VDD(VDD),.Y(g8861),.A(g6643),.B(g493));
  AND2 AND2_203(.VSS(VSS),.VDD(VDD),.Y(g8868),.A(g6751),.B(g1177));
  AND2 AND2_204(.VSS(VSS),.VDD(VDD),.Y(g8869),.A(g6776),.B(g5552));
  AND2 AND2_205(.VSS(VSS),.VDD(VDD),.Y(g8892),.A(g3338),.B(g496));
  AND2 AND2_206(.VSS(VSS),.VDD(VDD),.Y(g8899),.A(g6945),.B(g1180));
  AND2 AND2_207(.VSS(VSS),.VDD(VDD),.Y(g8906),.A(g7053),.B(g1871));
  AND2 AND2_208(.VSS(VSS),.VDD(VDD),.Y(g8907),.A(g7078),.B(g5598));
  AND2 AND2_209(.VSS(VSS),.VDD(VDD),.Y(g8932),.A(g3494),.B(g1183));
  AND2 AND2_210(.VSS(VSS),.VDD(VDD),.Y(g8939),.A(g7195),.B(g1874));
  AND2 AND2_211(.VSS(VSS),.VDD(VDD),.Y(g8946),.A(g7303),.B(g2565));
  AND2 AND2_212(.VSS(VSS),.VDD(VDD),.Y(g8947),.A(g7328),.B(g5615));
  AND2 AND2_213(.VSS(VSS),.VDD(VDD),.Y(g8972),.A(g3650),.B(g1877));
  AND2 AND2_214(.VSS(VSS),.VDD(VDD),.Y(g8979),.A(g7391),.B(g2568));
  AND2 AND2_215(.VSS(VSS),.VDD(VDD),.Y(g9004),.A(g3806),.B(g2571));
  AND2 AND2_216(.VSS(VSS),.VDD(VDD),.Y(g9009),.A(g6486),.B(g565));
  AND2 AND2_217(.VSS(VSS),.VDD(VDD),.Y(g9026),.A(g5438),.B(g7610));
  AND2 AND2_218(.VSS(VSS),.VDD(VDD),.Y(g9033),.A(g6643),.B(g567));
  AND2 AND2_219(.VSS(VSS),.VDD(VDD),.Y(g9034),.A(g6751),.B(g1251));
  AND2 AND2_220(.VSS(VSS),.VDD(VDD),.Y(g9047),.A(g6448),.B(g7616));
  AND2 AND2_221(.VSS(VSS),.VDD(VDD),.Y(g9048),.A(g3338),.B(g489));
  AND2 AND2_222(.VSS(VSS),.VDD(VDD),.Y(g9049),.A(g5473),.B(g7619));
  AND2 AND2_223(.VSS(VSS),.VDD(VDD),.Y(g9056),.A(g6945),.B(g1253));
  AND2 AND2_224(.VSS(VSS),.VDD(VDD),.Y(g9057),.A(g7053),.B(g1945));
  AND2 AND2_225(.VSS(VSS),.VDD(VDD),.Y(g9061),.A(g3306),.B(g7623));
  AND2 AND2_226(.VSS(VSS),.VDD(VDD),.Y(g9062),.A(g5438),.B(g7626));
  AND2 AND2_227(.VSS(VSS),.VDD(VDD),.Y(g9063),.A(g5438),.B(g7629));
  AND2 AND2_228(.VSS(VSS),.VDD(VDD),.Y(g9064),.A(g6713),.B(g7632));
  AND2 AND2_229(.VSS(VSS),.VDD(VDD),.Y(g9065),.A(g3494),.B(g1176));
  AND2 AND2_230(.VSS(VSS),.VDD(VDD),.Y(g9066),.A(g5512),.B(g7635));
  AND2 AND2_231(.VSS(VSS),.VDD(VDD),.Y(g9073),.A(g7195),.B(g1947));
  AND2 AND2_232(.VSS(VSS),.VDD(VDD),.Y(g9074),.A(g7303),.B(g2639));
  AND2 AND2_233(.VSS(VSS),.VDD(VDD),.Y(g9075),.A(g6448),.B(g7643));
  AND2 AND2_234(.VSS(VSS),.VDD(VDD),.Y(g9076),.A(g5438),.B(g7646));
  AND2 AND2_235(.VSS(VSS),.VDD(VDD),.Y(g9077),.A(g6448),.B(g7649));
  AND2 AND2_236(.VSS(VSS),.VDD(VDD),.Y(g9078),.A(g3462),.B(g7652));
  AND2 AND2_237(.VSS(VSS),.VDD(VDD),.Y(g9079),.A(g5473),.B(g7655));
  AND2 AND2_238(.VSS(VSS),.VDD(VDD),.Y(g9080),.A(g5473),.B(g7658));
  AND2 AND2_239(.VSS(VSS),.VDD(VDD),.Y(g9081),.A(g7015),.B(g7661));
  AND2 AND2_240(.VSS(VSS),.VDD(VDD),.Y(g9082),.A(g3650),.B(g1870));
  AND2 AND2_241(.VSS(VSS),.VDD(VDD),.Y(g9083),.A(g5556),.B(g7664));
  AND2 AND2_242(.VSS(VSS),.VDD(VDD),.Y(g9090),.A(g7391),.B(g2641));
  AND2 AND2_243(.VSS(VSS),.VDD(VDD),.Y(g9091),.A(g3306),.B(g7670));
  AND2 AND2_244(.VSS(VSS),.VDD(VDD),.Y(g9092),.A(g6448),.B(g7673));
  AND2 AND2_245(.VSS(VSS),.VDD(VDD),.Y(g9093),.A(g3306),.B(g7676));
  AND2 AND2_246(.VSS(VSS),.VDD(VDD),.Y(g9094),.A(g6713),.B(g7679));
  AND2 AND2_247(.VSS(VSS),.VDD(VDD),.Y(g9095),.A(g5473),.B(g7682));
  AND2 AND2_248(.VSS(VSS),.VDD(VDD),.Y(g9096),.A(g6713),.B(g7685));
  AND2 AND2_249(.VSS(VSS),.VDD(VDD),.Y(g9097),.A(g3618),.B(g7688));
  AND2 AND2_250(.VSS(VSS),.VDD(VDD),.Y(g9098),.A(g5512),.B(g7691));
  AND2 AND2_251(.VSS(VSS),.VDD(VDD),.Y(g9099),.A(g5512),.B(g7694));
  AND2 AND2_252(.VSS(VSS),.VDD(VDD),.Y(g9100),.A(g7265),.B(g7697));
  AND2 AND2_253(.VSS(VSS),.VDD(VDD),.Y(g9101),.A(g3806),.B(g2564));
  AND2 AND2_254(.VSS(VSS),.VDD(VDD),.Y(g9102),.A(g3306),.B(g7703));
  AND2 AND2_255(.VSS(VSS),.VDD(VDD),.Y(g9103),.A(g3462),.B(g7706));
  AND2 AND2_256(.VSS(VSS),.VDD(VDD),.Y(g9104),.A(g6713),.B(g7709));
  AND2 AND2_257(.VSS(VSS),.VDD(VDD),.Y(g9105),.A(g3462),.B(g7712));
  AND2 AND2_258(.VSS(VSS),.VDD(VDD),.Y(g9106),.A(g7015),.B(g7715));
  AND2 AND2_259(.VSS(VSS),.VDD(VDD),.Y(g9107),.A(g5512),.B(g7718));
  AND2 AND2_260(.VSS(VSS),.VDD(VDD),.Y(g9108),.A(g7015),.B(g7721));
  AND2 AND2_261(.VSS(VSS),.VDD(VDD),.Y(g9109),.A(g3774),.B(g7724));
  AND2 AND2_262(.VSS(VSS),.VDD(VDD),.Y(g9110),.A(g5556),.B(g7727));
  AND2 AND2_263(.VSS(VSS),.VDD(VDD),.Y(g9111),.A(g5556),.B(g7730));
  AND2 AND2_264(.VSS(VSS),.VDD(VDD),.Y(g9112),.A(g3462),.B(g7733));
  AND2 AND2_265(.VSS(VSS),.VDD(VDD),.Y(g9113),.A(g3618),.B(g7736));
  AND2 AND2_266(.VSS(VSS),.VDD(VDD),.Y(g9114),.A(g7015),.B(g7739));
  AND2 AND2_267(.VSS(VSS),.VDD(VDD),.Y(g9115),.A(g3618),.B(g7742));
  AND2 AND2_268(.VSS(VSS),.VDD(VDD),.Y(g9116),.A(g7265),.B(g7745));
  AND2 AND2_269(.VSS(VSS),.VDD(VDD),.Y(g9117),.A(g5556),.B(g7748));
  AND2 AND2_270(.VSS(VSS),.VDD(VDD),.Y(g9118),.A(g7265),.B(g7751));
  AND2 AND2_271(.VSS(VSS),.VDD(VDD),.Y(g9119),.A(g5438),.B(g7754));
  AND2 AND2_272(.VSS(VSS),.VDD(VDD),.Y(g9120),.A(g3618),.B(g7757));
  AND2 AND2_273(.VSS(VSS),.VDD(VDD),.Y(g9121),.A(g3774),.B(g7760));
  AND2 AND2_274(.VSS(VSS),.VDD(VDD),.Y(g9122),.A(g7265),.B(g7763));
  AND2 AND2_275(.VSS(VSS),.VDD(VDD),.Y(g9123),.A(g3774),.B(g7766));
  AND2 AND2_276(.VSS(VSS),.VDD(VDD),.Y(g9124),.A(g6448),.B(g7769));
  AND2 AND2_277(.VSS(VSS),.VDD(VDD),.Y(g9125),.A(g5473),.B(g7776));
  AND2 AND2_278(.VSS(VSS),.VDD(VDD),.Y(g9126),.A(g3774),.B(g7779));
  AND2 AND2_279(.VSS(VSS),.VDD(VDD),.Y(g9127),.A(g3306),.B(g7782));
  AND2 AND2_280(.VSS(VSS),.VDD(VDD),.Y(g9131),.A(g6713),.B(g7785));
  AND2 AND2_281(.VSS(VSS),.VDD(VDD),.Y(g9132),.A(g5512),.B(g7792));
  AND2 AND2_282(.VSS(VSS),.VDD(VDD),.Y(g9133),.A(g3462),.B(g7796));
  AND2 AND2_283(.VSS(VSS),.VDD(VDD),.Y(g9137),.A(g7015),.B(g7799));
  AND2 AND2_284(.VSS(VSS),.VDD(VDD),.Y(g9138),.A(g5556),.B(g7806));
  AND2 AND2_285(.VSS(VSS),.VDD(VDD),.Y(g9139),.A(g3618),.B(g7809));
  AND2 AND2_286(.VSS(VSS),.VDD(VDD),.Y(g9143),.A(g7265),.B(g7812));
  AND2 AND2_287(.VSS(VSS),.VDD(VDD),.Y(g9145),.A(g3774),.B(g7823));
  AND2 AND2_288(.VSS(VSS),.VDD(VDD),.Y(g9241),.A(g6232),.B(g7950));
  AND2 AND2_289(.VSS(VSS),.VDD(VDD),.Y(g9301),.A(g6314),.B(g7990));
  AND2 AND2_290(.VSS(VSS),.VDD(VDD),.Y(g9302),.A(g6232),.B(g7993));
  AND2 AND2_291(.VSS(VSS),.VDD(VDD),.Y(g9319),.A(g6369),.B(g8001));
  AND2 AND2_292(.VSS(VSS),.VDD(VDD),.Y(g9364),.A(g3254),.B(g8053));
  AND2 AND2_293(.VSS(VSS),.VDD(VDD),.Y(g9365),.A(g6314),.B(g8056));
  AND2 AND2_294(.VSS(VSS),.VDD(VDD),.Y(g9366),.A(g6232),.B(g8059));
  AND2 AND2_295(.VSS(VSS),.VDD(VDD),.Y(g9367),.A(g6232),.B(g8062));
  AND2 AND2_296(.VSS(VSS),.VDD(VDD),.Y(g9382),.A(g6519),.B(g8065));
  AND2 AND2_297(.VSS(VSS),.VDD(VDD),.Y(g9383),.A(g6369),.B(g8068));
  AND2 AND2_298(.VSS(VSS),.VDD(VDD),.Y(g9400),.A(g6574),.B(g8076));
  AND2 AND2_299(.VSS(VSS),.VDD(VDD),.Y(g9438),.A(g3254),.B(g8123));
  AND2 AND2_300(.VSS(VSS),.VDD(VDD),.Y(g9439),.A(g6314),.B(g8126));
  AND2 AND2_301(.VSS(VSS),.VDD(VDD),.Y(g9440),.A(g6232),.B(g8129));
  AND2 AND2_302(.VSS(VSS),.VDD(VDD),.Y(g9441),.A(g6314),.B(g8132));
  AND2 AND2_303(.VSS(VSS),.VDD(VDD),.Y(g9442),.A(g6232),.B(g8135));
  AND2 AND2_304(.VSS(VSS),.VDD(VDD),.Y(g9461),.A(g3410),.B(g8138));
  AND2 AND2_305(.VSS(VSS),.VDD(VDD),.Y(g9462),.A(g6519),.B(g8141));
  AND2 AND2_306(.VSS(VSS),.VDD(VDD),.Y(g9463),.A(g6369),.B(g8144));
  AND2 AND2_307(.VSS(VSS),.VDD(VDD),.Y(g9464),.A(g6369),.B(g8147));
  AND2 AND2_308(.VSS(VSS),.VDD(VDD),.Y(g9479),.A(g6783),.B(g8150));
  AND2 AND2_309(.VSS(VSS),.VDD(VDD),.Y(g9480),.A(g6574),.B(g8153));
  AND2 AND2_310(.VSS(VSS),.VDD(VDD),.Y(g9497),.A(g6838),.B(g8161));
  AND2 AND2_311(.VSS(VSS),.VDD(VDD),.Y(g9518),.A(g3254),.B(g8191));
  AND2 AND2_312(.VSS(VSS),.VDD(VDD),.Y(g9519),.A(g6314),.B(g8194));
  AND2 AND2_313(.VSS(VSS),.VDD(VDD),.Y(g9520),.A(g6232),.B(g8197));
  AND2 AND2_314(.VSS(VSS),.VDD(VDD),.Y(g9521),.A(g3254),.B(g8200));
  AND2 AND2_315(.VSS(VSS),.VDD(VDD),.Y(g9522),.A(g6314),.B(g8203));
  AND2 AND2_316(.VSS(VSS),.VDD(VDD),.Y(g9523),.A(g6232),.B(g8206));
  AND3 AND3_0(.VSS(VSS),.VDD(VDD),.Y(g9534),.A(g7772),.B(g6135),.C(g538));
  AND2 AND2_317(.VSS(VSS),.VDD(VDD),.Y(g9580),.A(g3410),.B(g8209));
  AND2 AND2_318(.VSS(VSS),.VDD(VDD),.Y(g9581),.A(g6519),.B(g8212));
  AND2 AND2_319(.VSS(VSS),.VDD(VDD),.Y(g9582),.A(g6369),.B(g8215));
  AND2 AND2_320(.VSS(VSS),.VDD(VDD),.Y(g9583),.A(g6519),.B(g8218));
  AND2 AND2_321(.VSS(VSS),.VDD(VDD),.Y(g9584),.A(g6369),.B(g8221));
  AND2 AND2_322(.VSS(VSS),.VDD(VDD),.Y(g9603),.A(g3566),.B(g8224));
  AND2 AND2_323(.VSS(VSS),.VDD(VDD),.Y(g9604),.A(g6783),.B(g8227));
  AND2 AND2_324(.VSS(VSS),.VDD(VDD),.Y(g9605),.A(g6574),.B(g8230));
  AND2 AND2_325(.VSS(VSS),.VDD(VDD),.Y(g9606),.A(g6574),.B(g8233));
  AND2 AND2_326(.VSS(VSS),.VDD(VDD),.Y(g9621),.A(g7085),.B(g8236));
  AND2 AND2_327(.VSS(VSS),.VDD(VDD),.Y(g9622),.A(g6838),.B(g8239));
  AND2 AND2_328(.VSS(VSS),.VDD(VDD),.Y(g9630),.A(g3254),.B(g3922));
  AND2 AND2_329(.VSS(VSS),.VDD(VDD),.Y(g9631),.A(g6314),.B(g3925));
  AND2 AND2_330(.VSS(VSS),.VDD(VDD),.Y(g9632),.A(g6232),.B(g3928));
  AND2 AND2_331(.VSS(VSS),.VDD(VDD),.Y(g9633),.A(g3254),.B(g3931));
  AND2 AND2_332(.VSS(VSS),.VDD(VDD),.Y(g9634),.A(g6314),.B(g3934));
  AND2 AND2_333(.VSS(VSS),.VDD(VDD),.Y(g9635),.A(g6232),.B(g3937));
  AND4 AND4_0(.VSS(VSS),.VDD(VDD),.Y(I16735),.A(g5856),.B(g4338),.C(g4339),.D(g5141));
  AND4 AND4_1(.VSS(VSS),.VDD(VDD),.Y(I16736),.A(g5713),.B(g5958),.C(g4735),.D(g4736));
  AND2 AND2_334(.VSS(VSS),.VDD(VDD),.Y(g9636),.A(I16735),.B(I16736));
  AND2 AND2_335(.VSS(VSS),.VDD(VDD),.Y(g9639),.A(g5438),.B(g408));
  AND2 AND2_336(.VSS(VSS),.VDD(VDD),.Y(g9647),.A(g6678),.B(g3942));
  AND2 AND2_337(.VSS(VSS),.VDD(VDD),.Y(g9648),.A(g6678),.B(g3945));
  AND2 AND2_338(.VSS(VSS),.VDD(VDD),.Y(g9660),.A(g3410),.B(g3948));
  AND2 AND2_339(.VSS(VSS),.VDD(VDD),.Y(g9661),.A(g6519),.B(g3951));
  AND2 AND2_340(.VSS(VSS),.VDD(VDD),.Y(g9662),.A(g6369),.B(g3954));
  AND2 AND2_341(.VSS(VSS),.VDD(VDD),.Y(g9663),.A(g3410),.B(g3957));
  AND2 AND2_342(.VSS(VSS),.VDD(VDD),.Y(g9664),.A(g6519),.B(g3960));
  AND2 AND2_343(.VSS(VSS),.VDD(VDD),.Y(g9665),.A(g6369),.B(g3963));
  AND3 AND3_1(.VSS(VSS),.VDD(VDD),.Y(g9676),.A(g7788),.B(g6145),.C(g1224));
  AND2 AND2_344(.VSS(VSS),.VDD(VDD),.Y(g9722),.A(g3566),.B(g3966));
  AND2 AND2_345(.VSS(VSS),.VDD(VDD),.Y(g9723),.A(g6783),.B(g3969));
  AND2 AND2_346(.VSS(VSS),.VDD(VDD),.Y(g9724),.A(g6574),.B(g3972));
  AND2 AND2_347(.VSS(VSS),.VDD(VDD),.Y(g9725),.A(g6783),.B(g3975));
  AND2 AND2_348(.VSS(VSS),.VDD(VDD),.Y(g9726),.A(g6574),.B(g3978));
  AND2 AND2_349(.VSS(VSS),.VDD(VDD),.Y(g9745),.A(g3722),.B(g3981));
  AND2 AND2_350(.VSS(VSS),.VDD(VDD),.Y(g9746),.A(g7085),.B(g3984));
  AND2 AND2_351(.VSS(VSS),.VDD(VDD),.Y(g9747),.A(g6838),.B(g3987));
  AND2 AND2_352(.VSS(VSS),.VDD(VDD),.Y(g9748),.A(g6838),.B(g3990));
  AND2 AND2_353(.VSS(VSS),.VDD(VDD),.Y(g9759),.A(g3254),.B(g4000));
  AND2 AND2_354(.VSS(VSS),.VDD(VDD),.Y(g9760),.A(g6314),.B(g4003));
  AND2 AND2_355(.VSS(VSS),.VDD(VDD),.Y(g9761),.A(g6232),.B(g4006));
  AND2 AND2_356(.VSS(VSS),.VDD(VDD),.Y(g9762),.A(g3254),.B(g4009));
  AND2 AND2_357(.VSS(VSS),.VDD(VDD),.Y(g9763),.A(g6314),.B(g4012));
  AND2 AND2_358(.VSS(VSS),.VDD(VDD),.Y(g9764),.A(g6448),.B(g411));
  AND2 AND2_359(.VSS(VSS),.VDD(VDD),.Y(g9765),.A(g5438),.B(g417));
  AND2 AND2_360(.VSS(VSS),.VDD(VDD),.Y(g9766),.A(g5438),.B(g4017));
  AND2 AND2_361(.VSS(VSS),.VDD(VDD),.Y(g9773),.A(g6912),.B(g4020));
  AND2 AND2_362(.VSS(VSS),.VDD(VDD),.Y(g9774),.A(g6678),.B(g4023));
  AND2 AND2_363(.VSS(VSS),.VDD(VDD),.Y(g9775),.A(g6912),.B(g4026));
  AND2 AND2_364(.VSS(VSS),.VDD(VDD),.Y(g9776),.A(g3410),.B(g4029));
  AND2 AND2_365(.VSS(VSS),.VDD(VDD),.Y(g9777),.A(g6519),.B(g4032));
  AND2 AND2_366(.VSS(VSS),.VDD(VDD),.Y(g9778),.A(g6369),.B(g4035));
  AND2 AND2_367(.VSS(VSS),.VDD(VDD),.Y(g9779),.A(g3410),.B(g4038));
  AND2 AND2_368(.VSS(VSS),.VDD(VDD),.Y(g9780),.A(g6519),.B(g4041));
  AND2 AND2_369(.VSS(VSS),.VDD(VDD),.Y(g9781),.A(g6369),.B(g4044));
  AND4 AND4_2(.VSS(VSS),.VDD(VDD),.Y(I16826),.A(g5903),.B(g4507),.C(g4508),.D(g5234));
  AND4 AND4_3(.VSS(VSS),.VDD(VDD),.Y(I16827),.A(g5771),.B(g5987),.C(g4911),.D(g4912));
  AND2 AND2_370(.VSS(VSS),.VDD(VDD),.Y(g9782),.A(I16826),.B(I16827));
  AND2 AND2_371(.VSS(VSS),.VDD(VDD),.Y(g9785),.A(g5473),.B(g1095));
  AND2 AND2_372(.VSS(VSS),.VDD(VDD),.Y(g9793),.A(g6980),.B(g4049));
  AND2 AND2_373(.VSS(VSS),.VDD(VDD),.Y(g9794),.A(g6980),.B(g4052));
  AND2 AND2_374(.VSS(VSS),.VDD(VDD),.Y(g9806),.A(g3566),.B(g4055));
  AND2 AND2_375(.VSS(VSS),.VDD(VDD),.Y(g9807),.A(g6783),.B(g4058));
  AND2 AND2_376(.VSS(VSS),.VDD(VDD),.Y(g9808),.A(g6574),.B(g4061));
  AND2 AND2_377(.VSS(VSS),.VDD(VDD),.Y(g9809),.A(g3566),.B(g4064));
  AND2 AND2_378(.VSS(VSS),.VDD(VDD),.Y(g9810),.A(g6783),.B(g4067));
  AND2 AND2_379(.VSS(VSS),.VDD(VDD),.Y(g9811),.A(g6574),.B(g4070));
  AND3 AND3_2(.VSS(VSS),.VDD(VDD),.Y(g9822),.A(g7802),.B(g6166),.C(g1918));
  AND2 AND2_380(.VSS(VSS),.VDD(VDD),.Y(g9868),.A(g3722),.B(g4073));
  AND2 AND2_381(.VSS(VSS),.VDD(VDD),.Y(g9869),.A(g7085),.B(g4076));
  AND2 AND2_382(.VSS(VSS),.VDD(VDD),.Y(g9870),.A(g6838),.B(g4079));
  AND2 AND2_383(.VSS(VSS),.VDD(VDD),.Y(g9871),.A(g7085),.B(g4082));
  AND2 AND2_384(.VSS(VSS),.VDD(VDD),.Y(g9872),.A(g6838),.B(g4085));
  AND2 AND2_385(.VSS(VSS),.VDD(VDD),.Y(g9887),.A(g6232),.B(g4095));
  AND2 AND2_386(.VSS(VSS),.VDD(VDD),.Y(g9888),.A(g3254),.B(g4098));
  AND2 AND2_387(.VSS(VSS),.VDD(VDD),.Y(g9889),.A(g6314),.B(g4101));
  AND2 AND2_388(.VSS(VSS),.VDD(VDD),.Y(g9890),.A(g6232),.B(g4104));
  AND2 AND2_389(.VSS(VSS),.VDD(VDD),.Y(g9891),.A(g3254),.B(g4107));
  AND2 AND2_390(.VSS(VSS),.VDD(VDD),.Y(g9892),.A(g3306),.B(g414));
  AND2 AND2_391(.VSS(VSS),.VDD(VDD),.Y(g9893),.A(g6448),.B(g420));
  AND2 AND2_392(.VSS(VSS),.VDD(VDD),.Y(g9894),.A(g6448),.B(g4112));
  AND2 AND2_393(.VSS(VSS),.VDD(VDD),.Y(g9901),.A(g3366),.B(g4115));
  AND2 AND2_394(.VSS(VSS),.VDD(VDD),.Y(g9902),.A(g6912),.B(g4118));
  AND2 AND2_395(.VSS(VSS),.VDD(VDD),.Y(g9903),.A(g6678),.B(g4121));
  AND2 AND2_396(.VSS(VSS),.VDD(VDD),.Y(g9904),.A(g3366),.B(g4124));
  AND2 AND2_397(.VSS(VSS),.VDD(VDD),.Y(g9905),.A(g3410),.B(g4127));
  AND2 AND2_398(.VSS(VSS),.VDD(VDD),.Y(g9906),.A(g6519),.B(g4130));
  AND2 AND2_399(.VSS(VSS),.VDD(VDD),.Y(g9907),.A(g6369),.B(g4133));
  AND2 AND2_400(.VSS(VSS),.VDD(VDD),.Y(g9908),.A(g3410),.B(g4136));
  AND2 AND2_401(.VSS(VSS),.VDD(VDD),.Y(g9909),.A(g6519),.B(g4139));
  AND2 AND2_402(.VSS(VSS),.VDD(VDD),.Y(g9910),.A(g6713),.B(g1098));
  AND2 AND2_403(.VSS(VSS),.VDD(VDD),.Y(g9911),.A(g5473),.B(g1104));
  AND2 AND2_404(.VSS(VSS),.VDD(VDD),.Y(g9912),.A(g5473),.B(g4144));
  AND2 AND2_405(.VSS(VSS),.VDD(VDD),.Y(g9919),.A(g7162),.B(g4147));
  AND2 AND2_406(.VSS(VSS),.VDD(VDD),.Y(g9920),.A(g6980),.B(g4150));
  AND2 AND2_407(.VSS(VSS),.VDD(VDD),.Y(g9921),.A(g7162),.B(g4153));
  AND2 AND2_408(.VSS(VSS),.VDD(VDD),.Y(g9922),.A(g3566),.B(g4156));
  AND2 AND2_409(.VSS(VSS),.VDD(VDD),.Y(g9923),.A(g6783),.B(g4159));
  AND2 AND2_410(.VSS(VSS),.VDD(VDD),.Y(g9924),.A(g6574),.B(g4162));
  AND2 AND2_411(.VSS(VSS),.VDD(VDD),.Y(g9925),.A(g3566),.B(g4165));
  AND2 AND2_412(.VSS(VSS),.VDD(VDD),.Y(g9926),.A(g6783),.B(g4168));
  AND2 AND2_413(.VSS(VSS),.VDD(VDD),.Y(g9927),.A(g6574),.B(g4171));
  AND4 AND4_4(.VSS(VSS),.VDD(VDD),.Y(I16930),.A(g5942),.B(g4683),.C(g4684),.D(g5297));
  AND4 AND4_5(.VSS(VSS),.VDD(VDD),.Y(I16931),.A(g5830),.B(g6024),.C(g5070),.D(g5071));
  AND2 AND2_414(.VSS(VSS),.VDD(VDD),.Y(g9928),.A(I16930),.B(I16931));
  AND2 AND2_415(.VSS(VSS),.VDD(VDD),.Y(g9931),.A(g5512),.B(g1789));
  AND2 AND2_416(.VSS(VSS),.VDD(VDD),.Y(g9939),.A(g7230),.B(g4176));
  AND2 AND2_417(.VSS(VSS),.VDD(VDD),.Y(g9940),.A(g7230),.B(g4179));
  AND2 AND2_418(.VSS(VSS),.VDD(VDD),.Y(g9952),.A(g3722),.B(g4182));
  AND2 AND2_419(.VSS(VSS),.VDD(VDD),.Y(g9953),.A(g7085),.B(g4185));
  AND2 AND2_420(.VSS(VSS),.VDD(VDD),.Y(g9954),.A(g6838),.B(g4188));
  AND2 AND2_421(.VSS(VSS),.VDD(VDD),.Y(g9955),.A(g3722),.B(g4191));
  AND2 AND2_422(.VSS(VSS),.VDD(VDD),.Y(g9956),.A(g7085),.B(g4194));
  AND2 AND2_423(.VSS(VSS),.VDD(VDD),.Y(g9957),.A(g6838),.B(g4197));
  AND3 AND3_3(.VSS(VSS),.VDD(VDD),.Y(g9968),.A(g7815),.B(g6193),.C(g2612));
  AND2 AND2_424(.VSS(VSS),.VDD(VDD),.Y(g10007),.A(g6314),.B(g4205));
  AND2 AND2_425(.VSS(VSS),.VDD(VDD),.Y(g10008),.A(g6232),.B(g4208));
  AND2 AND2_426(.VSS(VSS),.VDD(VDD),.Y(g10009),.A(g3254),.B(g4211));
  AND2 AND2_427(.VSS(VSS),.VDD(VDD),.Y(g10010),.A(g6314),.B(g4214));
  AND2 AND2_428(.VSS(VSS),.VDD(VDD),.Y(g10011),.A(g5438),.B(g4217));
  AND2 AND2_429(.VSS(VSS),.VDD(VDD),.Y(g10012),.A(g3306),.B(g423));
  AND2 AND2_430(.VSS(VSS),.VDD(VDD),.Y(g10013),.A(g3306),.B(g4221));
  AND2 AND2_431(.VSS(VSS),.VDD(VDD),.Y(g10014),.A(g5438),.B(g429));
  AND2 AND2_432(.VSS(VSS),.VDD(VDD),.Y(g10024),.A(g3398),.B(g6912));
  AND2 AND2_433(.VSS(VSS),.VDD(VDD),.Y(g10035),.A(g3366),.B(g4225));
  AND2 AND2_434(.VSS(VSS),.VDD(VDD),.Y(g10036),.A(g6912),.B(g4228));
  AND2 AND2_435(.VSS(VSS),.VDD(VDD),.Y(g10037),.A(g6678),.B(g4231));
  AND2 AND2_436(.VSS(VSS),.VDD(VDD),.Y(g10041),.A(g6369),.B(g4234));
  AND2 AND2_437(.VSS(VSS),.VDD(VDD),.Y(g10042),.A(g3410),.B(g4237));
  AND2 AND2_438(.VSS(VSS),.VDD(VDD),.Y(g10043),.A(g6519),.B(g4240));
  AND2 AND2_439(.VSS(VSS),.VDD(VDD),.Y(g10044),.A(g6369),.B(g4243));
  AND2 AND2_440(.VSS(VSS),.VDD(VDD),.Y(g10045),.A(g3410),.B(g4246));
  AND2 AND2_441(.VSS(VSS),.VDD(VDD),.Y(g10046),.A(g3462),.B(g1101));
  AND2 AND2_442(.VSS(VSS),.VDD(VDD),.Y(g10047),.A(g6713),.B(g1107));
  AND2 AND2_443(.VSS(VSS),.VDD(VDD),.Y(g10048),.A(g6713),.B(g4251));
  AND2 AND2_444(.VSS(VSS),.VDD(VDD),.Y(g10055),.A(g3522),.B(g4254));
  AND2 AND2_445(.VSS(VSS),.VDD(VDD),.Y(g10056),.A(g7162),.B(g4257));
  AND2 AND2_446(.VSS(VSS),.VDD(VDD),.Y(g10057),.A(g6980),.B(g4260));
  AND2 AND2_447(.VSS(VSS),.VDD(VDD),.Y(g10058),.A(g3522),.B(g4263));
  AND2 AND2_448(.VSS(VSS),.VDD(VDD),.Y(g10059),.A(g3566),.B(g4266));
  AND2 AND2_449(.VSS(VSS),.VDD(VDD),.Y(g10060),.A(g6783),.B(g4269));
  AND2 AND2_450(.VSS(VSS),.VDD(VDD),.Y(g10061),.A(g6574),.B(g4272));
  AND2 AND2_451(.VSS(VSS),.VDD(VDD),.Y(g10062),.A(g3566),.B(g4275));
  AND2 AND2_452(.VSS(VSS),.VDD(VDD),.Y(g10063),.A(g6783),.B(g4278));
  AND2 AND2_453(.VSS(VSS),.VDD(VDD),.Y(g10064),.A(g7015),.B(g1792));
  AND2 AND2_454(.VSS(VSS),.VDD(VDD),.Y(g10065),.A(g5512),.B(g1798));
  AND2 AND2_455(.VSS(VSS),.VDD(VDD),.Y(g10066),.A(g5512),.B(g4283));
  AND2 AND2_456(.VSS(VSS),.VDD(VDD),.Y(g10073),.A(g7358),.B(g4286));
  AND2 AND2_457(.VSS(VSS),.VDD(VDD),.Y(g10074),.A(g7230),.B(g4289));
  AND2 AND2_458(.VSS(VSS),.VDD(VDD),.Y(g10075),.A(g7358),.B(g4292));
  AND2 AND2_459(.VSS(VSS),.VDD(VDD),.Y(g10076),.A(g3722),.B(g4295));
  AND2 AND2_460(.VSS(VSS),.VDD(VDD),.Y(g10077),.A(g7085),.B(g4298));
  AND2 AND2_461(.VSS(VSS),.VDD(VDD),.Y(g10078),.A(g6838),.B(g4301));
  AND2 AND2_462(.VSS(VSS),.VDD(VDD),.Y(g10079),.A(g3722),.B(g4304));
  AND2 AND2_463(.VSS(VSS),.VDD(VDD),.Y(g10080),.A(g7085),.B(g4307));
  AND2 AND2_464(.VSS(VSS),.VDD(VDD),.Y(g10081),.A(g6838),.B(g4310));
  AND4 AND4_6(.VSS(VSS),.VDD(VDD),.Y(I17042),.A(g5976),.B(g4860),.C(g4861),.D(g5334));
  AND4 AND4_7(.VSS(VSS),.VDD(VDD),.Y(I17043),.A(g5886),.B(g6040),.C(g5199),.D(g5200));
  AND2 AND2_465(.VSS(VSS),.VDD(VDD),.Y(g10082),.A(I17042),.B(I17043));
  AND2 AND2_466(.VSS(VSS),.VDD(VDD),.Y(g10085),.A(g5556),.B(g2483));
  AND2 AND2_467(.VSS(VSS),.VDD(VDD),.Y(g10093),.A(g7426),.B(g4315));
  AND2 AND2_468(.VSS(VSS),.VDD(VDD),.Y(g10094),.A(g7426),.B(g4318));
  AND2 AND2_469(.VSS(VSS),.VDD(VDD),.Y(g10101),.A(g3254),.B(g4329));
  AND2 AND2_470(.VSS(VSS),.VDD(VDD),.Y(g10102),.A(g6314),.B(g4332));
  AND2 AND2_471(.VSS(VSS),.VDD(VDD),.Y(g10103),.A(g3254),.B(g4335));
  AND2 AND2_472(.VSS(VSS),.VDD(VDD),.Y(g10104),.A(g6448),.B(g4340));
  AND2 AND2_473(.VSS(VSS),.VDD(VDD),.Y(g10105),.A(g5438),.B(g4343));
  AND2 AND2_474(.VSS(VSS),.VDD(VDD),.Y(g10106),.A(g6448),.B(g432));
  AND2 AND2_475(.VSS(VSS),.VDD(VDD),.Y(g10107),.A(g5438),.B(g438));
  AND2 AND2_476(.VSS(VSS),.VDD(VDD),.Y(g10108),.A(g6486),.B(g569));
  AND2 AND2_477(.VSS(VSS),.VDD(VDD),.Y(g10112),.A(g3366),.B(g4348));
  AND2 AND2_478(.VSS(VSS),.VDD(VDD),.Y(g10113),.A(g6912),.B(g4351));
  AND2 AND2_479(.VSS(VSS),.VDD(VDD),.Y(g10114),.A(g6678),.B(g4354));
  AND2 AND2_480(.VSS(VSS),.VDD(VDD),.Y(g10115),.A(g6678),.B(g4357));
  AND2 AND2_481(.VSS(VSS),.VDD(VDD),.Y(g10116),.A(g6519),.B(g4360));
  AND2 AND2_482(.VSS(VSS),.VDD(VDD),.Y(g10117),.A(g6369),.B(g4363));
  AND2 AND2_483(.VSS(VSS),.VDD(VDD),.Y(g10118),.A(g3410),.B(g4366));
  AND2 AND2_484(.VSS(VSS),.VDD(VDD),.Y(g10119),.A(g6519),.B(g4369));
  AND2 AND2_485(.VSS(VSS),.VDD(VDD),.Y(g10120),.A(g5473),.B(g4372));
  AND2 AND2_486(.VSS(VSS),.VDD(VDD),.Y(g10121),.A(g3462),.B(g1110));
  AND2 AND2_487(.VSS(VSS),.VDD(VDD),.Y(g10122),.A(g3462),.B(g4376));
  AND2 AND2_488(.VSS(VSS),.VDD(VDD),.Y(g10123),.A(g5473),.B(g1116));
  AND2 AND2_489(.VSS(VSS),.VDD(VDD),.Y(g10133),.A(g3554),.B(g7162));
  AND2 AND2_490(.VSS(VSS),.VDD(VDD),.Y(g10144),.A(g3522),.B(g4380));
  AND2 AND2_491(.VSS(VSS),.VDD(VDD),.Y(g10145),.A(g7162),.B(g4383));
  AND2 AND2_492(.VSS(VSS),.VDD(VDD),.Y(g10146),.A(g6980),.B(g4386));
  AND2 AND2_493(.VSS(VSS),.VDD(VDD),.Y(g10150),.A(g6574),.B(g4389));
  AND2 AND2_494(.VSS(VSS),.VDD(VDD),.Y(g10151),.A(g3566),.B(g4392));
  AND2 AND2_495(.VSS(VSS),.VDD(VDD),.Y(g10152),.A(g6783),.B(g4395));
  AND2 AND2_496(.VSS(VSS),.VDD(VDD),.Y(g10153),.A(g6574),.B(g4398));
  AND2 AND2_497(.VSS(VSS),.VDD(VDD),.Y(g10154),.A(g3566),.B(g4401));
  AND2 AND2_498(.VSS(VSS),.VDD(VDD),.Y(g10155),.A(g3618),.B(g1795));
  AND2 AND2_499(.VSS(VSS),.VDD(VDD),.Y(g10156),.A(g7015),.B(g1801));
  AND2 AND2_500(.VSS(VSS),.VDD(VDD),.Y(g10157),.A(g7015),.B(g4406));
  AND2 AND2_501(.VSS(VSS),.VDD(VDD),.Y(g10164),.A(g3678),.B(g4409));
  AND2 AND2_502(.VSS(VSS),.VDD(VDD),.Y(g10165),.A(g7358),.B(g4412));
  AND2 AND2_503(.VSS(VSS),.VDD(VDD),.Y(g10166),.A(g7230),.B(g4415));
  AND2 AND2_504(.VSS(VSS),.VDD(VDD),.Y(g10167),.A(g3678),.B(g4418));
  AND2 AND2_505(.VSS(VSS),.VDD(VDD),.Y(g10168),.A(g3722),.B(g4421));
  AND2 AND2_506(.VSS(VSS),.VDD(VDD),.Y(g10169),.A(g7085),.B(g4424));
  AND2 AND2_507(.VSS(VSS),.VDD(VDD),.Y(g10170),.A(g6838),.B(g4427));
  AND2 AND2_508(.VSS(VSS),.VDD(VDD),.Y(g10171),.A(g3722),.B(g4430));
  AND2 AND2_509(.VSS(VSS),.VDD(VDD),.Y(g10172),.A(g7085),.B(g4433));
  AND2 AND2_510(.VSS(VSS),.VDD(VDD),.Y(g10173),.A(g7265),.B(g2486));
  AND2 AND2_511(.VSS(VSS),.VDD(VDD),.Y(g10174),.A(g5556),.B(g2492));
  AND2 AND2_512(.VSS(VSS),.VDD(VDD),.Y(g10175),.A(g5556),.B(g4438));
  AND2 AND2_513(.VSS(VSS),.VDD(VDD),.Y(g10182),.A(g7488),.B(g4441));
  AND2 AND2_514(.VSS(VSS),.VDD(VDD),.Y(g10183),.A(g7426),.B(g4444));
  AND2 AND2_515(.VSS(VSS),.VDD(VDD),.Y(g10184),.A(g7488),.B(g4447));
  AND4 AND4_8(.VSS(VSS),.VDD(VDD),.Y(I17156),.A(g6898),.B(g2998),.C(g6901),.D(g3002));
  AND4 AND4_9(.VSS(VSS),.VDD(VDD),.Y(g10186),.A(g3013),.B(g7466),.C(g3024),.D(I17156));
  AND2 AND2_516(.VSS(VSS),.VDD(VDD),.Y(g10192),.A(g3254),.B(g4453));
  AND2 AND2_517(.VSS(VSS),.VDD(VDD),.Y(g10193),.A(g3306),.B(g4465));
  AND2 AND2_518(.VSS(VSS),.VDD(VDD),.Y(g10194),.A(g6448),.B(g4468));
  AND2 AND2_519(.VSS(VSS),.VDD(VDD),.Y(g10195),.A(g5438),.B(g4471));
  AND2 AND2_520(.VSS(VSS),.VDD(VDD),.Y(g10196),.A(g3306),.B(g435));
  AND2 AND2_521(.VSS(VSS),.VDD(VDD),.Y(g10197),.A(g6448),.B(g441));
  AND2 AND2_522(.VSS(VSS),.VDD(VDD),.Y(g10198),.A(g6643),.B(g571));
  AND2 AND2_523(.VSS(VSS),.VDD(VDD),.Y(g10199),.A(g6486),.B(g4476));
  AND2 AND2_524(.VSS(VSS),.VDD(VDD),.Y(g10200),.A(g6486),.B(g587));
  AND2 AND2_525(.VSS(VSS),.VDD(VDD),.Y(g10201),.A(g3366),.B(g4480));
  AND2 AND2_526(.VSS(VSS),.VDD(VDD),.Y(g10202),.A(g6912),.B(g4483));
  AND2 AND2_527(.VSS(VSS),.VDD(VDD),.Y(g10203),.A(g6678),.B(g4486));
  AND2 AND2_528(.VSS(VSS),.VDD(VDD),.Y(g10204),.A(g6912),.B(g4489));
  AND2 AND2_529(.VSS(VSS),.VDD(VDD),.Y(g10205),.A(g6678),.B(g4492));
  AND2 AND2_530(.VSS(VSS),.VDD(VDD),.Y(g10206),.A(g3410),.B(g4498));
  AND2 AND2_531(.VSS(VSS),.VDD(VDD),.Y(g10207),.A(g6519),.B(g4501));
  AND2 AND2_532(.VSS(VSS),.VDD(VDD),.Y(g10208),.A(g3410),.B(g4504));
  AND2 AND2_533(.VSS(VSS),.VDD(VDD),.Y(g10209),.A(g6713),.B(g4509));
  AND2 AND2_534(.VSS(VSS),.VDD(VDD),.Y(g10210),.A(g5473),.B(g4512));
  AND2 AND2_535(.VSS(VSS),.VDD(VDD),.Y(g10211),.A(g6713),.B(g1119));
  AND2 AND2_536(.VSS(VSS),.VDD(VDD),.Y(g10212),.A(g5473),.B(g1125));
  AND2 AND2_537(.VSS(VSS),.VDD(VDD),.Y(g10213),.A(g6751),.B(g1255));
  AND2 AND2_538(.VSS(VSS),.VDD(VDD),.Y(g10217),.A(g3522),.B(g4517));
  AND2 AND2_539(.VSS(VSS),.VDD(VDD),.Y(g10218),.A(g7162),.B(g4520));
  AND2 AND2_540(.VSS(VSS),.VDD(VDD),.Y(g10219),.A(g6980),.B(g4523));
  AND2 AND2_541(.VSS(VSS),.VDD(VDD),.Y(g10220),.A(g6980),.B(g4526));
  AND2 AND2_542(.VSS(VSS),.VDD(VDD),.Y(g10221),.A(g6783),.B(g4529));
  AND2 AND2_543(.VSS(VSS),.VDD(VDD),.Y(g10222),.A(g6574),.B(g4532));
  AND2 AND2_544(.VSS(VSS),.VDD(VDD),.Y(g10223),.A(g3566),.B(g4535));
  AND2 AND2_545(.VSS(VSS),.VDD(VDD),.Y(g10224),.A(g6783),.B(g4538));
  AND2 AND2_546(.VSS(VSS),.VDD(VDD),.Y(g10225),.A(g5512),.B(g4541));
  AND2 AND2_547(.VSS(VSS),.VDD(VDD),.Y(g10226),.A(g3618),.B(g1804));
  AND2 AND2_548(.VSS(VSS),.VDD(VDD),.Y(g10227),.A(g3618),.B(g4545));
  AND2 AND2_549(.VSS(VSS),.VDD(VDD),.Y(g10228),.A(g5512),.B(g1810));
  AND2 AND2_550(.VSS(VSS),.VDD(VDD),.Y(g10238),.A(g3710),.B(g7358));
  AND2 AND2_551(.VSS(VSS),.VDD(VDD),.Y(g10249),.A(g3678),.B(g4549));
  AND2 AND2_552(.VSS(VSS),.VDD(VDD),.Y(g10250),.A(g7358),.B(g4552));
  AND2 AND2_553(.VSS(VSS),.VDD(VDD),.Y(g10251),.A(g7230),.B(g4555));
  AND2 AND2_554(.VSS(VSS),.VDD(VDD),.Y(g10255),.A(g6838),.B(g4558));
  AND2 AND2_555(.VSS(VSS),.VDD(VDD),.Y(g10256),.A(g3722),.B(g4561));
  AND2 AND2_556(.VSS(VSS),.VDD(VDD),.Y(g10257),.A(g7085),.B(g4564));
  AND2 AND2_557(.VSS(VSS),.VDD(VDD),.Y(g10258),.A(g6838),.B(g4567));
  AND2 AND2_558(.VSS(VSS),.VDD(VDD),.Y(g10259),.A(g3722),.B(g4570));
  AND2 AND2_559(.VSS(VSS),.VDD(VDD),.Y(g10260),.A(g3774),.B(g2489));
  AND2 AND2_560(.VSS(VSS),.VDD(VDD),.Y(g10261),.A(g7265),.B(g2495));
  AND2 AND2_561(.VSS(VSS),.VDD(VDD),.Y(g10262),.A(g7265),.B(g4575));
  AND2 AND2_562(.VSS(VSS),.VDD(VDD),.Y(g10269),.A(g3834),.B(g4578));
  AND2 AND2_563(.VSS(VSS),.VDD(VDD),.Y(g10270),.A(g7488),.B(g4581));
  AND2 AND2_564(.VSS(VSS),.VDD(VDD),.Y(g10271),.A(g7426),.B(g4584));
  AND2 AND2_565(.VSS(VSS),.VDD(VDD),.Y(g10272),.A(g3834),.B(g4587));
  AND2 AND2_566(.VSS(VSS),.VDD(VDD),.Y(g10279),.A(g3306),.B(g4592));
  AND2 AND2_567(.VSS(VSS),.VDD(VDD),.Y(g10280),.A(g6448),.B(g4595));
  AND2 AND2_568(.VSS(VSS),.VDD(VDD),.Y(g10281),.A(g5438),.B(g4598));
  AND2 AND2_569(.VSS(VSS),.VDD(VDD),.Y(g10282),.A(g3306),.B(g444));
  AND2 AND2_570(.VSS(VSS),.VDD(VDD),.Y(g10283),.A(g3338),.B(g573));
  AND2 AND2_571(.VSS(VSS),.VDD(VDD),.Y(g10284),.A(g6643),.B(g4603));
  AND2 AND2_572(.VSS(VSS),.VDD(VDD),.Y(g10285),.A(g6486),.B(g4606));
  AND2 AND2_573(.VSS(VSS),.VDD(VDD),.Y(g10286),.A(g6643),.B(g590));
  AND2 AND2_574(.VSS(VSS),.VDD(VDD),.Y(g10287),.A(g6486),.B(g596));
  AND2 AND2_575(.VSS(VSS),.VDD(VDD),.Y(g10288),.A(g3366),.B(g4611));
  AND2 AND2_576(.VSS(VSS),.VDD(VDD),.Y(g10289),.A(g6912),.B(g4614));
  AND2 AND2_577(.VSS(VSS),.VDD(VDD),.Y(g10290),.A(g6678),.B(g4617));
  AND2 AND2_578(.VSS(VSS),.VDD(VDD),.Y(g10291),.A(g3366),.B(g4620));
  AND2 AND2_579(.VSS(VSS),.VDD(VDD),.Y(g10292),.A(g6912),.B(g4623));
  AND2 AND2_580(.VSS(VSS),.VDD(VDD),.Y(g10293),.A(g6678),.B(g4626));
  AND2 AND2_581(.VSS(VSS),.VDD(VDD),.Y(g10294),.A(g3410),.B(g4629));
  AND2 AND2_582(.VSS(VSS),.VDD(VDD),.Y(g10295),.A(g3462),.B(g4641));
  AND2 AND2_583(.VSS(VSS),.VDD(VDD),.Y(g10296),.A(g6713),.B(g4644));
  AND2 AND2_584(.VSS(VSS),.VDD(VDD),.Y(g10297),.A(g5473),.B(g4647));
  AND2 AND2_585(.VSS(VSS),.VDD(VDD),.Y(g10298),.A(g3462),.B(g1122));
  AND2 AND2_586(.VSS(VSS),.VDD(VDD),.Y(g10299),.A(g6713),.B(g1128));
  AND2 AND2_587(.VSS(VSS),.VDD(VDD),.Y(g10300),.A(g6945),.B(g1257));
  AND2 AND2_588(.VSS(VSS),.VDD(VDD),.Y(g10301),.A(g6751),.B(g4652));
  AND2 AND2_589(.VSS(VSS),.VDD(VDD),.Y(g10302),.A(g6751),.B(g1273));
  AND2 AND2_590(.VSS(VSS),.VDD(VDD),.Y(g10303),.A(g3522),.B(g4656));
  AND2 AND2_591(.VSS(VSS),.VDD(VDD),.Y(g10304),.A(g7162),.B(g4659));
  AND2 AND2_592(.VSS(VSS),.VDD(VDD),.Y(g10305),.A(g6980),.B(g4662));
  AND2 AND2_593(.VSS(VSS),.VDD(VDD),.Y(g10306),.A(g7162),.B(g4665));
  AND2 AND2_594(.VSS(VSS),.VDD(VDD),.Y(g10307),.A(g6980),.B(g4668));
  AND2 AND2_595(.VSS(VSS),.VDD(VDD),.Y(g10308),.A(g3566),.B(g4674));
  AND2 AND2_596(.VSS(VSS),.VDD(VDD),.Y(g10309),.A(g6783),.B(g4677));
  AND2 AND2_597(.VSS(VSS),.VDD(VDD),.Y(g10310),.A(g3566),.B(g4680));
  AND2 AND2_598(.VSS(VSS),.VDD(VDD),.Y(g10311),.A(g7015),.B(g4685));
  AND2 AND2_599(.VSS(VSS),.VDD(VDD),.Y(g10312),.A(g5512),.B(g4688));
  AND2 AND2_600(.VSS(VSS),.VDD(VDD),.Y(g10313),.A(g7015),.B(g1813));
  AND2 AND2_601(.VSS(VSS),.VDD(VDD),.Y(g10314),.A(g5512),.B(g1819));
  AND2 AND2_602(.VSS(VSS),.VDD(VDD),.Y(g10315),.A(g7053),.B(g1949));
  AND2 AND2_603(.VSS(VSS),.VDD(VDD),.Y(g10319),.A(g3678),.B(g4693));
  AND2 AND2_604(.VSS(VSS),.VDD(VDD),.Y(g10320),.A(g7358),.B(g4696));
  AND2 AND2_605(.VSS(VSS),.VDD(VDD),.Y(g10321),.A(g7230),.B(g4699));
  AND2 AND2_606(.VSS(VSS),.VDD(VDD),.Y(g10322),.A(g7230),.B(g4702));
  AND2 AND2_607(.VSS(VSS),.VDD(VDD),.Y(g10323),.A(g7085),.B(g4705));
  AND2 AND2_608(.VSS(VSS),.VDD(VDD),.Y(g10324),.A(g6838),.B(g4708));
  AND2 AND2_609(.VSS(VSS),.VDD(VDD),.Y(g10325),.A(g3722),.B(g4711));
  AND2 AND2_610(.VSS(VSS),.VDD(VDD),.Y(g10326),.A(g7085),.B(g4714));
  AND2 AND2_611(.VSS(VSS),.VDD(VDD),.Y(g10327),.A(g5556),.B(g4717));
  AND2 AND2_612(.VSS(VSS),.VDD(VDD),.Y(g10328),.A(g3774),.B(g2498));
  AND2 AND2_613(.VSS(VSS),.VDD(VDD),.Y(g10329),.A(g3774),.B(g4721));
  AND2 AND2_614(.VSS(VSS),.VDD(VDD),.Y(g10330),.A(g5556),.B(g2504));
  AND2 AND2_615(.VSS(VSS),.VDD(VDD),.Y(g10340),.A(g3866),.B(g7488));
  AND2 AND2_616(.VSS(VSS),.VDD(VDD),.Y(g10351),.A(g3834),.B(g4725));
  AND2 AND2_617(.VSS(VSS),.VDD(VDD),.Y(g10352),.A(g7488),.B(g4728));
  AND2 AND2_618(.VSS(VSS),.VDD(VDD),.Y(g10353),.A(g7426),.B(g4731));
  AND2 AND2_619(.VSS(VSS),.VDD(VDD),.Y(g10360),.A(g3306),.B(g4737));
  AND2 AND2_620(.VSS(VSS),.VDD(VDD),.Y(g10361),.A(g6448),.B(g4740));
  AND2 AND2_621(.VSS(VSS),.VDD(VDD),.Y(g10362),.A(g3338),.B(g4743));
  AND2 AND2_622(.VSS(VSS),.VDD(VDD),.Y(g10363),.A(g6643),.B(g4746));
  AND2 AND2_623(.VSS(VSS),.VDD(VDD),.Y(g10364),.A(g6486),.B(g4749));
  AND2 AND2_624(.VSS(VSS),.VDD(VDD),.Y(g10365),.A(g3338),.B(g593));
  AND2 AND2_625(.VSS(VSS),.VDD(VDD),.Y(g10366),.A(g6643),.B(g599));
  AND2 AND2_626(.VSS(VSS),.VDD(VDD),.Y(g10367),.A(g3366),.B(g4754));
  AND2 AND2_627(.VSS(VSS),.VDD(VDD),.Y(g10368),.A(g6912),.B(g4757));
  AND2 AND2_628(.VSS(VSS),.VDD(VDD),.Y(g10369),.A(g6678),.B(g4760));
  AND2 AND2_629(.VSS(VSS),.VDD(VDD),.Y(g10370),.A(g3366),.B(g4763));
  AND2 AND2_630(.VSS(VSS),.VDD(VDD),.Y(g10371),.A(g6912),.B(g4766));
  AND2 AND2_631(.VSS(VSS),.VDD(VDD),.Y(g10372),.A(g3462),.B(g4769));
  AND2 AND2_632(.VSS(VSS),.VDD(VDD),.Y(g10373),.A(g6713),.B(g4772));
  AND2 AND2_633(.VSS(VSS),.VDD(VDD),.Y(g10374),.A(g5473),.B(g4775));
  AND2 AND2_634(.VSS(VSS),.VDD(VDD),.Y(g10375),.A(g3462),.B(g1131));
  AND2 AND2_635(.VSS(VSS),.VDD(VDD),.Y(g10376),.A(g3494),.B(g1259));
  AND2 AND2_636(.VSS(VSS),.VDD(VDD),.Y(g10377),.A(g6945),.B(g4780));
  AND2 AND2_637(.VSS(VSS),.VDD(VDD),.Y(g10378),.A(g6751),.B(g4783));
  AND2 AND2_638(.VSS(VSS),.VDD(VDD),.Y(g10379),.A(g6945),.B(g1276));
  AND2 AND2_639(.VSS(VSS),.VDD(VDD),.Y(g10380),.A(g6751),.B(g1282));
  AND2 AND2_640(.VSS(VSS),.VDD(VDD),.Y(g10381),.A(g3522),.B(g4788));
  AND2 AND2_641(.VSS(VSS),.VDD(VDD),.Y(g10382),.A(g7162),.B(g4791));
  AND2 AND2_642(.VSS(VSS),.VDD(VDD),.Y(g10383),.A(g6980),.B(g4794));
  AND2 AND2_643(.VSS(VSS),.VDD(VDD),.Y(g10384),.A(g3522),.B(g4797));
  AND2 AND2_644(.VSS(VSS),.VDD(VDD),.Y(g10385),.A(g7162),.B(g4800));
  AND2 AND2_645(.VSS(VSS),.VDD(VDD),.Y(g10386),.A(g6980),.B(g4803));
  AND2 AND2_646(.VSS(VSS),.VDD(VDD),.Y(g10387),.A(g3566),.B(g4806));
  AND2 AND2_647(.VSS(VSS),.VDD(VDD),.Y(g10388),.A(g3618),.B(g4818));
  AND2 AND2_648(.VSS(VSS),.VDD(VDD),.Y(g10389),.A(g7015),.B(g4821));
  AND2 AND2_649(.VSS(VSS),.VDD(VDD),.Y(g10390),.A(g5512),.B(g4824));
  AND2 AND2_650(.VSS(VSS),.VDD(VDD),.Y(g10391),.A(g3618),.B(g1816));
  AND2 AND2_651(.VSS(VSS),.VDD(VDD),.Y(g10392),.A(g7015),.B(g1822));
  AND2 AND2_652(.VSS(VSS),.VDD(VDD),.Y(g10393),.A(g7195),.B(g1951));
  AND2 AND2_653(.VSS(VSS),.VDD(VDD),.Y(g10394),.A(g7053),.B(g4829));
  AND2 AND2_654(.VSS(VSS),.VDD(VDD),.Y(g10395),.A(g7053),.B(g1967));
  AND2 AND2_655(.VSS(VSS),.VDD(VDD),.Y(g10396),.A(g3678),.B(g4833));
  AND2 AND2_656(.VSS(VSS),.VDD(VDD),.Y(g10397),.A(g7358),.B(g4836));
  AND2 AND2_657(.VSS(VSS),.VDD(VDD),.Y(g10398),.A(g7230),.B(g4839));
  AND2 AND2_658(.VSS(VSS),.VDD(VDD),.Y(g10399),.A(g7358),.B(g4842));
  AND2 AND2_659(.VSS(VSS),.VDD(VDD),.Y(g10400),.A(g7230),.B(g4845));
  AND2 AND2_660(.VSS(VSS),.VDD(VDD),.Y(g10401),.A(g3722),.B(g4851));
  AND2 AND2_661(.VSS(VSS),.VDD(VDD),.Y(g10402),.A(g7085),.B(g4854));
  AND2 AND2_662(.VSS(VSS),.VDD(VDD),.Y(g10403),.A(g3722),.B(g4857));
  AND2 AND2_663(.VSS(VSS),.VDD(VDD),.Y(g10404),.A(g7265),.B(g4862));
  AND2 AND2_664(.VSS(VSS),.VDD(VDD),.Y(g10405),.A(g5556),.B(g4865));
  AND2 AND2_665(.VSS(VSS),.VDD(VDD),.Y(g10406),.A(g7265),.B(g2507));
  AND2 AND2_666(.VSS(VSS),.VDD(VDD),.Y(g10407),.A(g5556),.B(g2513));
  AND2 AND2_667(.VSS(VSS),.VDD(VDD),.Y(g10408),.A(g7303),.B(g2643));
  AND2 AND2_668(.VSS(VSS),.VDD(VDD),.Y(g10412),.A(g3834),.B(g4870));
  AND2 AND2_669(.VSS(VSS),.VDD(VDD),.Y(g10413),.A(g7488),.B(g4873));
  AND2 AND2_670(.VSS(VSS),.VDD(VDD),.Y(g10414),.A(g7426),.B(g4876));
  AND2 AND2_671(.VSS(VSS),.VDD(VDD),.Y(g10415),.A(g7426),.B(g4879));
  AND2 AND2_672(.VSS(VSS),.VDD(VDD),.Y(g10422),.A(g3306),.B(g4882));
  AND2 AND2_673(.VSS(VSS),.VDD(VDD),.Y(g10423),.A(g5438),.B(g4885));
  AND2 AND2_674(.VSS(VSS),.VDD(VDD),.Y(g10430),.A(g3338),.B(g4888));
  AND2 AND2_675(.VSS(VSS),.VDD(VDD),.Y(g10431),.A(g6643),.B(g4891));
  AND2 AND2_676(.VSS(VSS),.VDD(VDD),.Y(g10432),.A(g6486),.B(g4894));
  AND2 AND2_677(.VSS(VSS),.VDD(VDD),.Y(g10433),.A(g3338),.B(g602));
  AND2 AND2_678(.VSS(VSS),.VDD(VDD),.Y(g10434),.A(g6486),.B(g605));
  AND2 AND2_679(.VSS(VSS),.VDD(VDD),.Y(g10435),.A(g3366),.B(g4899));
  AND2 AND2_680(.VSS(VSS),.VDD(VDD),.Y(g10436),.A(g6912),.B(g4902));
  AND2 AND2_681(.VSS(VSS),.VDD(VDD),.Y(g10437),.A(g6678),.B(g4905));
  AND2 AND2_682(.VSS(VSS),.VDD(VDD),.Y(g10438),.A(g3366),.B(g4908));
  AND2 AND2_683(.VSS(VSS),.VDD(VDD),.Y(g10439),.A(g3462),.B(g4913));
  AND2 AND2_684(.VSS(VSS),.VDD(VDD),.Y(g10440),.A(g6713),.B(g4916));
  AND2 AND2_685(.VSS(VSS),.VDD(VDD),.Y(g10441),.A(g3494),.B(g4919));
  AND2 AND2_686(.VSS(VSS),.VDD(VDD),.Y(g10442),.A(g6945),.B(g4922));
  AND2 AND2_687(.VSS(VSS),.VDD(VDD),.Y(g10443),.A(g6751),.B(g4925));
  AND2 AND2_688(.VSS(VSS),.VDD(VDD),.Y(g10444),.A(g3494),.B(g1279));
  AND2 AND2_689(.VSS(VSS),.VDD(VDD),.Y(g10445),.A(g6945),.B(g1285));
  AND2 AND2_690(.VSS(VSS),.VDD(VDD),.Y(g10446),.A(g3522),.B(g4930));
  AND2 AND2_691(.VSS(VSS),.VDD(VDD),.Y(g10447),.A(g7162),.B(g4933));
  AND2 AND2_692(.VSS(VSS),.VDD(VDD),.Y(g10448),.A(g6980),.B(g4936));
  AND2 AND2_693(.VSS(VSS),.VDD(VDD),.Y(g10449),.A(g3522),.B(g4939));
  AND2 AND2_694(.VSS(VSS),.VDD(VDD),.Y(g10450),.A(g7162),.B(g4942));
  AND2 AND2_695(.VSS(VSS),.VDD(VDD),.Y(g10451),.A(g3618),.B(g4945));
  AND2 AND2_696(.VSS(VSS),.VDD(VDD),.Y(g10452),.A(g7015),.B(g4948));
  AND2 AND2_697(.VSS(VSS),.VDD(VDD),.Y(g10453),.A(g5512),.B(g4951));
  AND2 AND2_698(.VSS(VSS),.VDD(VDD),.Y(g10454),.A(g3618),.B(g1825));
  AND2 AND2_699(.VSS(VSS),.VDD(VDD),.Y(g10455),.A(g3650),.B(g1953));
  AND2 AND2_700(.VSS(VSS),.VDD(VDD),.Y(g10456),.A(g7195),.B(g4956));
  AND2 AND2_701(.VSS(VSS),.VDD(VDD),.Y(g10457),.A(g7053),.B(g4959));
  AND2 AND2_702(.VSS(VSS),.VDD(VDD),.Y(g10458),.A(g7195),.B(g1970));
  AND2 AND2_703(.VSS(VSS),.VDD(VDD),.Y(g10459),.A(g7053),.B(g1976));
  AND2 AND2_704(.VSS(VSS),.VDD(VDD),.Y(g10460),.A(g3678),.B(g4964));
  AND2 AND2_705(.VSS(VSS),.VDD(VDD),.Y(g10461),.A(g7358),.B(g4967));
  AND2 AND2_706(.VSS(VSS),.VDD(VDD),.Y(g10462),.A(g7230),.B(g4970));
  AND2 AND2_707(.VSS(VSS),.VDD(VDD),.Y(g10463),.A(g3678),.B(g4973));
  AND2 AND2_708(.VSS(VSS),.VDD(VDD),.Y(g10464),.A(g7358),.B(g4976));
  AND2 AND2_709(.VSS(VSS),.VDD(VDD),.Y(g10465),.A(g7230),.B(g4979));
  AND2 AND2_710(.VSS(VSS),.VDD(VDD),.Y(g10466),.A(g3722),.B(g4982));
  AND2 AND2_711(.VSS(VSS),.VDD(VDD),.Y(g10467),.A(g3774),.B(g4994));
  AND2 AND2_712(.VSS(VSS),.VDD(VDD),.Y(g10468),.A(g7265),.B(g4997));
  AND2 AND2_713(.VSS(VSS),.VDD(VDD),.Y(g10469),.A(g5556),.B(g5000));
  AND2 AND2_714(.VSS(VSS),.VDD(VDD),.Y(g10470),.A(g3774),.B(g2510));
  AND2 AND2_715(.VSS(VSS),.VDD(VDD),.Y(g10471),.A(g7265),.B(g2516));
  AND2 AND2_716(.VSS(VSS),.VDD(VDD),.Y(g10472),.A(g7391),.B(g2645));
  AND2 AND2_717(.VSS(VSS),.VDD(VDD),.Y(g10473),.A(g7303),.B(g5005));
  AND2 AND2_718(.VSS(VSS),.VDD(VDD),.Y(g10474),.A(g7303),.B(g2661));
  AND2 AND2_719(.VSS(VSS),.VDD(VDD),.Y(g10475),.A(g3834),.B(g5009));
  AND2 AND2_720(.VSS(VSS),.VDD(VDD),.Y(g10476),.A(g7488),.B(g5012));
  AND2 AND2_721(.VSS(VSS),.VDD(VDD),.Y(g10477),.A(g7426),.B(g5015));
  AND2 AND2_722(.VSS(VSS),.VDD(VDD),.Y(g10478),.A(g7488),.B(g5018));
  AND2 AND2_723(.VSS(VSS),.VDD(VDD),.Y(g10479),.A(g7426),.B(g5021));
  AND3 AND3_4(.VSS(VSS),.VDD(VDD),.Y(I17429),.A(g6901),.B(g7338),.C(g7146));
  AND3 AND3_5(.VSS(VSS),.VDD(VDD),.Y(g10480),.A(g7466),.B(g7342),.C(I17429));
  AND2 AND2_724(.VSS(VSS),.VDD(VDD),.Y(g10485),.A(g6448),.B(g5024));
  AND2 AND2_725(.VSS(VSS),.VDD(VDD),.Y(g10492),.A(g3338),.B(g5027));
  AND2 AND2_726(.VSS(VSS),.VDD(VDD),.Y(g10493),.A(g6643),.B(g5030));
  AND2 AND2_727(.VSS(VSS),.VDD(VDD),.Y(g10494),.A(g6643),.B(g608));
  AND2 AND2_728(.VSS(VSS),.VDD(VDD),.Y(g10495),.A(g6486),.B(g614));
  AND2 AND2_729(.VSS(VSS),.VDD(VDD),.Y(g10496),.A(g3366),.B(g5035));
  AND2 AND2_730(.VSS(VSS),.VDD(VDD),.Y(g10497),.A(g6912),.B(g5038));
  AND2 AND2_731(.VSS(VSS),.VDD(VDD),.Y(g10498),.A(g3462),.B(g5041));
  AND2 AND2_732(.VSS(VSS),.VDD(VDD),.Y(g10499),.A(g5473),.B(g5044));
  AND2 AND2_733(.VSS(VSS),.VDD(VDD),.Y(g10506),.A(g3494),.B(g5047));
  AND2 AND2_734(.VSS(VSS),.VDD(VDD),.Y(g10507),.A(g6945),.B(g5050));
  AND2 AND2_735(.VSS(VSS),.VDD(VDD),.Y(g10508),.A(g6751),.B(g5053));
  AND2 AND2_736(.VSS(VSS),.VDD(VDD),.Y(g10509),.A(g3494),.B(g1288));
  AND2 AND2_737(.VSS(VSS),.VDD(VDD),.Y(g10510),.A(g6751),.B(g1291));
  AND2 AND2_738(.VSS(VSS),.VDD(VDD),.Y(g10511),.A(g3522),.B(g5058));
  AND2 AND2_739(.VSS(VSS),.VDD(VDD),.Y(g10512),.A(g7162),.B(g5061));
  AND2 AND2_740(.VSS(VSS),.VDD(VDD),.Y(g10513),.A(g6980),.B(g5064));
  AND2 AND2_741(.VSS(VSS),.VDD(VDD),.Y(g10514),.A(g3522),.B(g5067));
  AND2 AND2_742(.VSS(VSS),.VDD(VDD),.Y(g10515),.A(g3618),.B(g5072));
  AND2 AND2_743(.VSS(VSS),.VDD(VDD),.Y(g10516),.A(g7015),.B(g5075));
  AND2 AND2_744(.VSS(VSS),.VDD(VDD),.Y(g10517),.A(g3650),.B(g5078));
  AND2 AND2_745(.VSS(VSS),.VDD(VDD),.Y(g10518),.A(g7195),.B(g5081));
  AND2 AND2_746(.VSS(VSS),.VDD(VDD),.Y(g10519),.A(g7053),.B(g5084));
  AND2 AND2_747(.VSS(VSS),.VDD(VDD),.Y(g10520),.A(g3650),.B(g1973));
  AND2 AND2_748(.VSS(VSS),.VDD(VDD),.Y(g10521),.A(g7195),.B(g1979));
  AND2 AND2_749(.VSS(VSS),.VDD(VDD),.Y(g10522),.A(g3678),.B(g5089));
  AND2 AND2_750(.VSS(VSS),.VDD(VDD),.Y(g10523),.A(g7358),.B(g5092));
  AND2 AND2_751(.VSS(VSS),.VDD(VDD),.Y(g10524),.A(g7230),.B(g5095));
  AND2 AND2_752(.VSS(VSS),.VDD(VDD),.Y(g10525),.A(g3678),.B(g5098));
  AND2 AND2_753(.VSS(VSS),.VDD(VDD),.Y(g10526),.A(g7358),.B(g5101));
  AND2 AND2_754(.VSS(VSS),.VDD(VDD),.Y(g10527),.A(g3774),.B(g5104));
  AND2 AND2_755(.VSS(VSS),.VDD(VDD),.Y(g10528),.A(g7265),.B(g5107));
  AND2 AND2_756(.VSS(VSS),.VDD(VDD),.Y(g10529),.A(g5556),.B(g5110));
  AND2 AND2_757(.VSS(VSS),.VDD(VDD),.Y(g10530),.A(g3774),.B(g2519));
  AND2 AND2_758(.VSS(VSS),.VDD(VDD),.Y(g10531),.A(g3806),.B(g2647));
  AND2 AND2_759(.VSS(VSS),.VDD(VDD),.Y(g10532),.A(g7391),.B(g5115));
  AND2 AND2_760(.VSS(VSS),.VDD(VDD),.Y(g10533),.A(g7303),.B(g5118));
  AND2 AND2_761(.VSS(VSS),.VDD(VDD),.Y(g10534),.A(g7391),.B(g2664));
  AND2 AND2_762(.VSS(VSS),.VDD(VDD),.Y(g10535),.A(g7303),.B(g2670));
  AND2 AND2_763(.VSS(VSS),.VDD(VDD),.Y(g10536),.A(g3834),.B(g5123));
  AND2 AND2_764(.VSS(VSS),.VDD(VDD),.Y(g10537),.A(g7488),.B(g5126));
  AND2 AND2_765(.VSS(VSS),.VDD(VDD),.Y(g10538),.A(g7426),.B(g5129));
  AND2 AND2_766(.VSS(VSS),.VDD(VDD),.Y(g10539),.A(g3834),.B(g5132));
  AND2 AND2_767(.VSS(VSS),.VDD(VDD),.Y(g10540),.A(g7488),.B(g5135));
  AND2 AND2_768(.VSS(VSS),.VDD(VDD),.Y(g10541),.A(g7426),.B(g5138));
  AND2 AND2_769(.VSS(VSS),.VDD(VDD),.Y(g10548),.A(g3306),.B(g5142));
  AND2 AND2_770(.VSS(VSS),.VDD(VDD),.Y(g10555),.A(g3338),.B(g5145));
  AND2 AND2_771(.VSS(VSS),.VDD(VDD),.Y(g10556),.A(g3338),.B(g611));
  AND2 AND2_772(.VSS(VSS),.VDD(VDD),.Y(g10557),.A(g6643),.B(g617));
  AND2 AND2_773(.VSS(VSS),.VDD(VDD),.Y(g10558),.A(g3366),.B(g5150));
  AND2 AND2_774(.VSS(VSS),.VDD(VDD),.Y(g10559),.A(g6713),.B(g5153));
  AND2 AND2_775(.VSS(VSS),.VDD(VDD),.Y(g10566),.A(g3494),.B(g5156));
  AND2 AND2_776(.VSS(VSS),.VDD(VDD),.Y(g10567),.A(g6945),.B(g5159));
  AND2 AND2_777(.VSS(VSS),.VDD(VDD),.Y(g10568),.A(g6945),.B(g1294));
  AND2 AND2_778(.VSS(VSS),.VDD(VDD),.Y(g10569),.A(g6751),.B(g1300));
  AND2 AND2_779(.VSS(VSS),.VDD(VDD),.Y(g10570),.A(g3522),.B(g5164));
  AND2 AND2_780(.VSS(VSS),.VDD(VDD),.Y(g10571),.A(g7162),.B(g5167));
  AND2 AND2_781(.VSS(VSS),.VDD(VDD),.Y(g10572),.A(g3618),.B(g5170));
  AND2 AND2_782(.VSS(VSS),.VDD(VDD),.Y(g10573),.A(g5512),.B(g5173));
  AND2 AND2_783(.VSS(VSS),.VDD(VDD),.Y(g10580),.A(g3650),.B(g5176));
  AND2 AND2_784(.VSS(VSS),.VDD(VDD),.Y(g10581),.A(g7195),.B(g5179));
  AND2 AND2_785(.VSS(VSS),.VDD(VDD),.Y(g10582),.A(g7053),.B(g5182));
  AND2 AND2_786(.VSS(VSS),.VDD(VDD),.Y(g10583),.A(g3650),.B(g1982));
  AND2 AND2_787(.VSS(VSS),.VDD(VDD),.Y(g10584),.A(g7053),.B(g1985));
  AND2 AND2_788(.VSS(VSS),.VDD(VDD),.Y(g10585),.A(g3678),.B(g5187));
  AND2 AND2_789(.VSS(VSS),.VDD(VDD),.Y(g10586),.A(g7358),.B(g5190));
  AND2 AND2_790(.VSS(VSS),.VDD(VDD),.Y(g10587),.A(g7230),.B(g5193));
  AND2 AND2_791(.VSS(VSS),.VDD(VDD),.Y(g10588),.A(g3678),.B(g5196));
  AND2 AND2_792(.VSS(VSS),.VDD(VDD),.Y(g10589),.A(g3774),.B(g5201));
  AND2 AND2_793(.VSS(VSS),.VDD(VDD),.Y(g10590),.A(g7265),.B(g5204));
  AND2 AND2_794(.VSS(VSS),.VDD(VDD),.Y(g10591),.A(g3806),.B(g5207));
  AND2 AND2_795(.VSS(VSS),.VDD(VDD),.Y(g10592),.A(g7391),.B(g5210));
  AND2 AND2_796(.VSS(VSS),.VDD(VDD),.Y(g10593),.A(g7303),.B(g5213));
  AND2 AND2_797(.VSS(VSS),.VDD(VDD),.Y(g10594),.A(g3806),.B(g2667));
  AND2 AND2_798(.VSS(VSS),.VDD(VDD),.Y(g10595),.A(g7391),.B(g2673));
  AND2 AND2_799(.VSS(VSS),.VDD(VDD),.Y(g10596),.A(g3834),.B(g5218));
  AND2 AND2_800(.VSS(VSS),.VDD(VDD),.Y(g10597),.A(g7488),.B(g5221));
  AND2 AND2_801(.VSS(VSS),.VDD(VDD),.Y(g10598),.A(g7426),.B(g5224));
  AND2 AND2_802(.VSS(VSS),.VDD(VDD),.Y(g10599),.A(g3834),.B(g5227));
  AND2 AND2_803(.VSS(VSS),.VDD(VDD),.Y(g10600),.A(g7488),.B(g5230));
  AND2 AND2_804(.VSS(VSS),.VDD(VDD),.Y(g10604),.A(g3338),.B(g620));
  AND2 AND2_805(.VSS(VSS),.VDD(VDD),.Y(g10605),.A(g3462),.B(g5235));
  AND2 AND2_806(.VSS(VSS),.VDD(VDD),.Y(g10612),.A(g3494),.B(g5238));
  AND2 AND2_807(.VSS(VSS),.VDD(VDD),.Y(g10613),.A(g3494),.B(g1297));
  AND2 AND2_808(.VSS(VSS),.VDD(VDD),.Y(g10614),.A(g6945),.B(g1303));
  AND2 AND2_809(.VSS(VSS),.VDD(VDD),.Y(g10615),.A(g3522),.B(g5243));
  AND2 AND2_810(.VSS(VSS),.VDD(VDD),.Y(g10616),.A(g7015),.B(g5246));
  AND2 AND2_811(.VSS(VSS),.VDD(VDD),.Y(g10623),.A(g3650),.B(g5249));
  AND2 AND2_812(.VSS(VSS),.VDD(VDD),.Y(g10624),.A(g7195),.B(g5252));
  AND2 AND2_813(.VSS(VSS),.VDD(VDD),.Y(g10625),.A(g7195),.B(g1988));
  AND2 AND2_814(.VSS(VSS),.VDD(VDD),.Y(g10626),.A(g7053),.B(g1994));
  AND2 AND2_815(.VSS(VSS),.VDD(VDD),.Y(g10627),.A(g3678),.B(g5257));
  AND2 AND2_816(.VSS(VSS),.VDD(VDD),.Y(g10628),.A(g7358),.B(g5260));
  AND2 AND2_817(.VSS(VSS),.VDD(VDD),.Y(g10629),.A(g3774),.B(g5263));
  AND2 AND2_818(.VSS(VSS),.VDD(VDD),.Y(g10630),.A(g5556),.B(g5266));
  AND2 AND2_819(.VSS(VSS),.VDD(VDD),.Y(g10637),.A(g3806),.B(g5269));
  AND2 AND2_820(.VSS(VSS),.VDD(VDD),.Y(g10638),.A(g7391),.B(g5272));
  AND2 AND2_821(.VSS(VSS),.VDD(VDD),.Y(g10639),.A(g7303),.B(g5275));
  AND2 AND2_822(.VSS(VSS),.VDD(VDD),.Y(g10640),.A(g3806),.B(g2676));
  AND2 AND2_823(.VSS(VSS),.VDD(VDD),.Y(g10641),.A(g7303),.B(g2679));
  AND2 AND2_824(.VSS(VSS),.VDD(VDD),.Y(g10642),.A(g3834),.B(g5280));
  AND2 AND2_825(.VSS(VSS),.VDD(VDD),.Y(g10643),.A(g7488),.B(g5283));
  AND2 AND2_826(.VSS(VSS),.VDD(VDD),.Y(g10644),.A(g7426),.B(g5286));
  AND2 AND2_827(.VSS(VSS),.VDD(VDD),.Y(g10645),.A(g3834),.B(g5289));
  AND2 AND2_828(.VSS(VSS),.VDD(VDD),.Y(g10650),.A(g6678),.B(g5293));
  AND2 AND2_829(.VSS(VSS),.VDD(VDD),.Y(g10651),.A(g3494),.B(g1306));
  AND2 AND2_830(.VSS(VSS),.VDD(VDD),.Y(g10652),.A(g3618),.B(g5298));
  AND2 AND2_831(.VSS(VSS),.VDD(VDD),.Y(g10659),.A(g3650),.B(g5301));
  AND2 AND2_832(.VSS(VSS),.VDD(VDD),.Y(g10660),.A(g3650),.B(g1991));
  AND2 AND2_833(.VSS(VSS),.VDD(VDD),.Y(g10661),.A(g7195),.B(g1997));
  AND2 AND2_834(.VSS(VSS),.VDD(VDD),.Y(g10662),.A(g3678),.B(g5306));
  AND2 AND2_835(.VSS(VSS),.VDD(VDD),.Y(g10663),.A(g7265),.B(g5309));
  AND2 AND2_836(.VSS(VSS),.VDD(VDD),.Y(g10670),.A(g3806),.B(g5312));
  AND2 AND2_837(.VSS(VSS),.VDD(VDD),.Y(g10671),.A(g7391),.B(g5315));
  AND2 AND2_838(.VSS(VSS),.VDD(VDD),.Y(g10672),.A(g7391),.B(g2682));
  AND2 AND2_839(.VSS(VSS),.VDD(VDD),.Y(g10673),.A(g7303),.B(g2688));
  AND2 AND2_840(.VSS(VSS),.VDD(VDD),.Y(g10674),.A(g3834),.B(g5320));
  AND2 AND2_841(.VSS(VSS),.VDD(VDD),.Y(g10675),.A(g7488),.B(g5323));
  AND2 AND2_842(.VSS(VSS),.VDD(VDD),.Y(g10678),.A(g6912),.B(g5327));
  AND2 AND2_843(.VSS(VSS),.VDD(VDD),.Y(g10680),.A(g6980),.B(g5330));
  AND2 AND2_844(.VSS(VSS),.VDD(VDD),.Y(g10681),.A(g3650),.B(g2000));
  AND2 AND2_845(.VSS(VSS),.VDD(VDD),.Y(g10682),.A(g3774),.B(g5335));
  AND2 AND2_846(.VSS(VSS),.VDD(VDD),.Y(g10689),.A(g3806),.B(g5338));
  AND2 AND2_847(.VSS(VSS),.VDD(VDD),.Y(g10690),.A(g3806),.B(g2685));
  AND2 AND2_848(.VSS(VSS),.VDD(VDD),.Y(g10691),.A(g7391),.B(g2691));
  AND2 AND2_849(.VSS(VSS),.VDD(VDD),.Y(g10692),.A(g3834),.B(g5343));
  AND4 AND4_10(.VSS(VSS),.VDD(VDD),.Y(g10693),.A(g7462),.B(g7522),.C(g2924),.D(g7545));
  AND2 AND2_850(.VSS(VSS),.VDD(VDD),.Y(g10704),.A(g3366),.B(g5352));
  AND2 AND2_851(.VSS(VSS),.VDD(VDD),.Y(g10707),.A(g7162),.B(g5355));
  AND2 AND2_852(.VSS(VSS),.VDD(VDD),.Y(g10709),.A(g7230),.B(g5358));
  AND2 AND2_853(.VSS(VSS),.VDD(VDD),.Y(g10710),.A(g3806),.B(g2694));
  AND3 AND3_6(.VSS(VSS),.VDD(VDD),.Y(I17599),.A(g7566),.B(g7583),.C(g7587));
  AND3 AND3_7(.VSS(VSS),.VDD(VDD),.Y(g10711),.A(g7595),.B(g7600),.C(I17599));
  AND2 AND2_854(.VSS(VSS),.VDD(VDD),.Y(g10724),.A(g3522),.B(g5369));
  AND2 AND2_855(.VSS(VSS),.VDD(VDD),.Y(g10727),.A(g7358),.B(g5372));
  AND2 AND2_856(.VSS(VSS),.VDD(VDD),.Y(g10729),.A(g7426),.B(g5375));
  AND2 AND2_857(.VSS(VSS),.VDD(VDD),.Y(g10745),.A(g3678),.B(g5382));
  AND2 AND2_858(.VSS(VSS),.VDD(VDD),.Y(g10748),.A(g7488),.B(g5385));
  AND2 AND2_859(.VSS(VSS),.VDD(VDD),.Y(g10764),.A(g3834),.B(g5391));
  AND2 AND2_860(.VSS(VSS),.VDD(VDD),.Y(g11347),.A(g6232),.B(g213));
  AND2 AND2_861(.VSS(VSS),.VDD(VDD),.Y(g11420),.A(g6314),.B(g216));
  AND2 AND2_862(.VSS(VSS),.VDD(VDD),.Y(g11421),.A(g6232),.B(g222));
  AND2 AND2_863(.VSS(VSS),.VDD(VDD),.Y(g11431),.A(g6369),.B(g900));
  AND2 AND2_864(.VSS(VSS),.VDD(VDD),.Y(g11607),.A(g5871),.B(g8360));
  AND2 AND2_865(.VSS(VSS),.VDD(VDD),.Y(g11612),.A(g5881),.B(g8378));
  AND2 AND2_866(.VSS(VSS),.VDD(VDD),.Y(g11637),.A(g5918),.B(g8427));
  AND2 AND2_867(.VSS(VSS),.VDD(VDD),.Y(g11771),.A(g554),.B(g8622));
  AND2 AND2_868(.VSS(VSS),.VDD(VDD),.Y(g11788),.A(g1240),.B(g8632));
  AND2 AND2_869(.VSS(VSS),.VDD(VDD),.Y(g11805),.A(g6173),.B(g8643));
  AND2 AND2_870(.VSS(VSS),.VDD(VDD),.Y(g11814),.A(g1934),.B(g8651));
  AND2 AND2_871(.VSS(VSS),.VDD(VDD),.Y(g11816),.A(g7869),.B(g8655));
  AND2 AND2_872(.VSS(VSS),.VDD(VDD),.Y(g11838),.A(g6205),.B(g8659));
  AND2 AND2_873(.VSS(VSS),.VDD(VDD),.Y(g11847),.A(g2628),.B(g8667));
  AND2 AND2_874(.VSS(VSS),.VDD(VDD),.Y(g11851),.A(g7849),.B(g8670));
  AND2 AND2_875(.VSS(VSS),.VDD(VDD),.Y(g11880),.A(g6294),.B(g8678));
  AND2 AND2_876(.VSS(VSS),.VDD(VDD),.Y(g11885),.A(g7834),.B(g8684));
  AND2 AND2_877(.VSS(VSS),.VDD(VDD),.Y(g11922),.A(g6431),.B(g8690));
  AND2 AND2_878(.VSS(VSS),.VDD(VDD),.Y(g11926),.A(g8169),.B(g8696));
  AND2 AND2_879(.VSS(VSS),.VDD(VDD),.Y(g11966),.A(g8090),.B(g8708));
  AND2 AND2_880(.VSS(VSS),.VDD(VDD),.Y(g11967),.A(g7967),.B(g8711));
  AND2 AND2_881(.VSS(VSS),.VDD(VDD),.Y(g12012),.A(g8015),.B(g8745));
  AND2 AND2_882(.VSS(VSS),.VDD(VDD),.Y(g12069),.A(g7964),.B(g8763));
  AND2 AND2_883(.VSS(VSS),.VDD(VDD),.Y(g12070),.A(g8018),.B(g8766));
  AND2 AND2_884(.VSS(VSS),.VDD(VDD),.Y(g12128),.A(g7916),.B(g8785));
  AND2 AND2_885(.VSS(VSS),.VDD(VDD),.Y(g12129),.A(g7872),.B(g8788));
  AND2 AND2_886(.VSS(VSS),.VDD(VDD),.Y(g12186),.A(g8093),.B(g8805));
  AND2 AND2_887(.VSS(VSS),.VDD(VDD),.Y(g12273),.A(g8172),.B(g8829));
  AND2 AND2_888(.VSS(VSS),.VDD(VDD),.Y(g12274),.A(g7900),.B(g8832));
  AND2 AND2_889(.VSS(VSS),.VDD(VDD),.Y(g12307),.A(g7919),.B(g8853));
  AND2 AND2_890(.VSS(VSS),.VDD(VDD),.Y(g12330),.A(g8246),.B(g8879));
  AND2 AND2_891(.VSS(VSS),.VDD(VDD),.Y(g12331),.A(g7927),.B(g8882));
  AND2 AND2_892(.VSS(VSS),.VDD(VDD),.Y(g12353),.A(g7852),.B(g8915));
  AND2 AND2_893(.VSS(VSS),.VDD(VDD),.Y(g12376),.A(g7974),.B(g8949));
  AND2 AND2_894(.VSS(VSS),.VDD(VDD),.Y(g12419),.A(g8028),.B(g9006));
  AND2 AND2_895(.VSS(VSS),.VDD(VDD),.Y(g12429),.A(g8101),.B(g9044));
  AND2 AND2_896(.VSS(VSS),.VDD(VDD),.Y(g12477),.A(g7822),.B(g9128));
  AND2 AND2_897(.VSS(VSS),.VDD(VDD),.Y(g12494),.A(g7833),.B(g9134));
  AND2 AND2_898(.VSS(VSS),.VDD(VDD),.Y(g12514),.A(g7848),.B(g9140));
  AND2 AND2_899(.VSS(VSS),.VDD(VDD),.Y(g12531),.A(g7868),.B(g9146));
  AND2 AND2_900(.VSS(VSS),.VDD(VDD),.Y(g12650),.A(g6149),.B(g9290));
  AND4 AND4_11(.VSS(VSS),.VDD(VDD),.Y(I19937),.A(g9507),.B(g9427),.C(g9356),.D(g9293));
  AND4 AND4_12(.VSS(VSS),.VDD(VDD),.Y(I19938),.A(g9232),.B(g9187),.C(g9161),.D(g9150));
  AND2 AND2_901(.VSS(VSS),.VDD(VDD),.Y(g12876),.A(I19937),.B(I19938));
  AND2 AND2_902(.VSS(VSS),.VDD(VDD),.Y(g12908),.A(g7899),.B(g10004));
  AND4 AND4_13(.VSS(VSS),.VDD(VDD),.Y(I19971),.A(g9649),.B(g9569),.C(g9453),.D(g9374));
  AND4 AND4_14(.VSS(VSS),.VDD(VDD),.Y(I19972),.A(g9310),.B(g9248),.C(g9203),.D(g9174));
  AND2 AND2_903(.VSS(VSS),.VDD(VDD),.Y(g12916),.A(I19971),.B(I19972));
  AND2 AND2_904(.VSS(VSS),.VDD(VDD),.Y(g12938),.A(g8179),.B(g10096));
  AND4 AND4_15(.VSS(VSS),.VDD(VDD),.Y(I19996),.A(g9795),.B(g9711),.C(g9595),.D(g9471));
  AND4 AND4_16(.VSS(VSS),.VDD(VDD),.Y(I19997),.A(g9391),.B(g9326),.C(g9264),.D(g9216));
  AND2 AND2_905(.VSS(VSS),.VDD(VDD),.Y(g12945),.A(I19996),.B(I19997));
  AND2 AND2_906(.VSS(VSS),.VDD(VDD),.Y(g12966),.A(g7926),.B(g10189));
  AND4 AND4_17(.VSS(VSS),.VDD(VDD),.Y(I20021),.A(g9941),.B(g9857),.C(g9737),.D(g9613));
  AND4 AND4_18(.VSS(VSS),.VDD(VDD),.Y(I20022),.A(g9488),.B(g9407),.C(g9342),.D(g9277));
  AND2 AND2_907(.VSS(VSS),.VDD(VDD),.Y(g12974),.A(I20021),.B(I20022));
  AND2 AND2_908(.VSS(VSS),.VDD(VDD),.Y(g12989),.A(g8254),.B(g10273));
  AND2 AND2_909(.VSS(VSS),.VDD(VDD),.Y(g12990),.A(g8180),.B(g10276));
  AND2 AND2_910(.VSS(VSS),.VDD(VDD),.Y(g13000),.A(g7973),.B(g10357));
  AND2 AND2_911(.VSS(VSS),.VDD(VDD),.Y(g13004),.A(g10186),.B(g8317));
  AND2 AND2_912(.VSS(VSS),.VDD(VDD),.Y(g13009),.A(g3995),.B(g10416));
  AND2 AND2_913(.VSS(VSS),.VDD(VDD),.Y(g13010),.A(g8255),.B(g10419));
  AND2 AND2_914(.VSS(VSS),.VDD(VDD),.Y(g13023),.A(g8027),.B(g10482));
  AND2 AND2_915(.VSS(VSS),.VDD(VDD),.Y(g13031),.A(g7879),.B(g10542));
  AND2 AND2_916(.VSS(VSS),.VDD(VDD),.Y(g13032),.A(g3996),.B(g10545));
  AND2 AND2_917(.VSS(VSS),.VDD(VDD),.Y(g13042),.A(g8100),.B(g10601));
  AND3 AND3_8(.VSS(VSS),.VDD(VDD),.Y(I20100),.A(g10186),.B(g3018),.C(g3028));
  AND3 AND3_9(.VSS(VSS),.VDD(VDD),.Y(g13055),.A(g7471),.B(g7570),.C(I20100));
  AND2 AND2_918(.VSS(VSS),.VDD(VDD),.Y(g13056),.A(g4092),.B(g10646));
  AND4 AND4_19(.VSS(VSS),.VDD(VDD),.Y(I20131),.A(g8313),.B(g7542),.C(g2888),.D(g7566));
  AND4 AND4_20(.VSS(VSS),.VDD(VDD),.Y(I20132),.A(g2892),.B(g2903),.C(g7595),.D(g2908));
  AND2 AND2_919(.VSS(VSS),.VDD(VDD),.Y(g13082),.A(I20131),.B(I20132));
  AND4 AND4_21(.VSS(VSS),.VDD(VDD),.Y(g13110),.A(g10693),.B(g2883),.C(g7562),.D(g10711));
  AND2 AND2_920(.VSS(VSS),.VDD(VDD),.Y(g13247),.A(g298),.B(g11032));
  AND2 AND2_921(.VSS(VSS),.VDD(VDD),.Y(g13266),.A(g5628),.B(g11088));
  AND2 AND2_922(.VSS(VSS),.VDD(VDD),.Y(g13270),.A(g985),.B(g11102));
  AND2 AND2_923(.VSS(VSS),.VDD(VDD),.Y(g13289),.A(g5647),.B(g11141));
  AND2 AND2_924(.VSS(VSS),.VDD(VDD),.Y(g13291),.A(g5656),.B(g11154));
  AND2 AND2_925(.VSS(VSS),.VDD(VDD),.Y(g13295),.A(g1679),.B(g11170));
  AND2 AND2_926(.VSS(VSS),.VDD(VDD),.Y(g13316),.A(g5675),.B(g11210));
  AND2 AND2_927(.VSS(VSS),.VDD(VDD),.Y(g13320),.A(g5685),.B(g11225));
  AND2 AND2_928(.VSS(VSS),.VDD(VDD),.Y(g13322),.A(g5694),.B(g11240));
  AND2 AND2_929(.VSS(VSS),.VDD(VDD),.Y(g13326),.A(g2373),.B(g11256));
  AND2 AND2_930(.VSS(VSS),.VDD(VDD),.Y(g13335),.A(g5708),.B(g11278));
  AND2 AND2_931(.VSS(VSS),.VDD(VDD),.Y(g13340),.A(g5727),.B(g11294));
  AND2 AND2_932(.VSS(VSS),.VDD(VDD),.Y(g13343),.A(g5737),.B(g11309));
  AND2 AND2_933(.VSS(VSS),.VDD(VDD),.Y(g13345),.A(g5746),.B(g11324));
  AND2 AND2_934(.VSS(VSS),.VDD(VDD),.Y(g13355),.A(g5756),.B(g11355));
  AND2 AND2_935(.VSS(VSS),.VDD(VDD),.Y(g13360),.A(g5766),.B(g11373));
  AND2 AND2_936(.VSS(VSS),.VDD(VDD),.Y(g13365),.A(g5785),.B(g11389));
  AND2 AND2_937(.VSS(VSS),.VDD(VDD),.Y(g13368),.A(g5795),.B(g11404));
  AND2 AND2_938(.VSS(VSS),.VDD(VDD),.Y(g13385),.A(g5815),.B(g11441));
  AND2 AND2_939(.VSS(VSS),.VDD(VDD),.Y(g13390),.A(g5825),.B(g11459));
  AND2 AND2_940(.VSS(VSS),.VDD(VDD),.Y(g13395),.A(g5844),.B(g11475));
  AND2 AND2_941(.VSS(VSS),.VDD(VDD),.Y(g13477),.A(g6016),.B(g12191));
  AND2 AND2_942(.VSS(VSS),.VDD(VDD),.Y(g13479),.A(g6017),.B(g12196));
  AND2 AND2_943(.VSS(VSS),.VDD(VDD),.Y(g13480),.A(g6018),.B(g12197));
  AND2 AND2_944(.VSS(VSS),.VDD(VDD),.Y(g13481),.A(g5864),.B(g11603));
  AND2 AND2_945(.VSS(VSS),.VDD(VDD),.Y(g13483),.A(g6020),.B(g12209));
  AND2 AND2_946(.VSS(VSS),.VDD(VDD),.Y(g13484),.A(g6021),.B(g12210));
  AND2 AND2_947(.VSS(VSS),.VDD(VDD),.Y(g13485),.A(g6022),.B(g12211));
  AND2 AND2_948(.VSS(VSS),.VDD(VDD),.Y(g13486),.A(g6023),.B(g12212));
  AND2 AND2_949(.VSS(VSS),.VDD(VDD),.Y(g13487),.A(g5874),.B(g11608));
  AND2 AND2_950(.VSS(VSS),.VDD(VDD),.Y(g13488),.A(g6025),.B(g12218));
  AND2 AND2_951(.VSS(VSS),.VDD(VDD),.Y(g13489),.A(g6026),.B(g12219));
  AND2 AND2_952(.VSS(VSS),.VDD(VDD),.Y(g13490),.A(g6027),.B(g12220));
  AND2 AND2_953(.VSS(VSS),.VDD(VDD),.Y(g13491),.A(g6028),.B(g12221));
  AND2 AND2_954(.VSS(VSS),.VDD(VDD),.Y(g13492),.A(g2371),.B(g12222));
  AND2 AND2_955(.VSS(VSS),.VDD(VDD),.Y(g13493),.A(g5887),.B(g11613));
  AND2 AND2_956(.VSS(VSS),.VDD(VDD),.Y(g13496),.A(g6032),.B(g12246));
  AND2 AND2_957(.VSS(VSS),.VDD(VDD),.Y(g13498),.A(g6033),.B(g12251));
  AND2 AND2_958(.VSS(VSS),.VDD(VDD),.Y(g13499),.A(g6034),.B(g12252));
  AND2 AND2_959(.VSS(VSS),.VDD(VDD),.Y(g13500),.A(g5911),.B(g11633));
  AND2 AND2_960(.VSS(VSS),.VDD(VDD),.Y(g13502),.A(g6036),.B(g12264));
  AND2 AND2_961(.VSS(VSS),.VDD(VDD),.Y(g13503),.A(g6037),.B(g12265));
  AND2 AND2_962(.VSS(VSS),.VDD(VDD),.Y(g13504),.A(g6038),.B(g12266));
  AND2 AND2_963(.VSS(VSS),.VDD(VDD),.Y(g13505),.A(g6039),.B(g12267));
  AND2 AND2_964(.VSS(VSS),.VDD(VDD),.Y(g13506),.A(g5921),.B(g11638));
  AND2 AND2_965(.VSS(VSS),.VDD(VDD),.Y(g13513),.A(g6043),.B(g12289));
  AND2 AND2_966(.VSS(VSS),.VDD(VDD),.Y(g13515),.A(g6044),.B(g12294));
  AND2 AND2_967(.VSS(VSS),.VDD(VDD),.Y(g13516),.A(g6045),.B(g12295));
  AND2 AND2_968(.VSS(VSS),.VDD(VDD),.Y(g13517),.A(g5950),.B(g11656));
  AND2 AND2_969(.VSS(VSS),.VDD(VDD),.Y(g13527),.A(g6047),.B(g12325));
  AND2 AND2_970(.VSS(VSS),.VDD(VDD),.Y(g13609),.A(g6141),.B(g12456));
  AND2 AND2_971(.VSS(VSS),.VDD(VDD),.Y(g13619),.A(g6162),.B(g12466));
  AND2 AND2_972(.VSS(VSS),.VDD(VDD),.Y(g13623),.A(g5428),.B(g12472));
  AND2 AND2_973(.VSS(VSS),.VDD(VDD),.Y(g13625),.A(g6173),.B(g12476));
  AND2 AND2_974(.VSS(VSS),.VDD(VDD),.Y(g13631),.A(g6189),.B(g12481));
  AND2 AND2_975(.VSS(VSS),.VDD(VDD),.Y(g13634),.A(g12776),.B(g8617));
  AND2 AND2_976(.VSS(VSS),.VDD(VDD),.Y(g13636),.A(g6205),.B(g12493));
  AND2 AND2_977(.VSS(VSS),.VDD(VDD),.Y(g13642),.A(g6221),.B(g12498));
  AND2 AND2_978(.VSS(VSS),.VDD(VDD),.Y(g13643),.A(g5431),.B(g12502));
  AND2 AND2_979(.VSS(VSS),.VDD(VDD),.Y(g13645),.A(g6281),.B(g12504));
  AND2 AND2_980(.VSS(VSS),.VDD(VDD),.Y(g13646),.A(g7772),.B(g12505));
  AND2 AND2_981(.VSS(VSS),.VDD(VDD),.Y(g13648),.A(g6294),.B(g12513));
  AND2 AND2_982(.VSS(VSS),.VDD(VDD),.Y(g13654),.A(g8093),.B(g11791));
  AND2 AND2_983(.VSS(VSS),.VDD(VDD),.Y(g13655),.A(g7540),.B(g12518));
  AND2 AND2_984(.VSS(VSS),.VDD(VDD),.Y(g13656),.A(g12776),.B(g8640));
  AND2 AND2_985(.VSS(VSS),.VDD(VDD),.Y(g13671),.A(g6418),.B(g12521));
  AND2 AND2_986(.VSS(VSS),.VDD(VDD),.Y(g13672),.A(g7788),.B(g12522));
  AND2 AND2_987(.VSS(VSS),.VDD(VDD),.Y(g13674),.A(g6431),.B(g12530));
  AND2 AND2_988(.VSS(VSS),.VDD(VDD),.Y(g13675),.A(g7561),.B(g12532));
  AND2 AND2_989(.VSS(VSS),.VDD(VDD),.Y(g13676),.A(g5434),.B(g12533));
  AND2 AND2_990(.VSS(VSS),.VDD(VDD),.Y(g13701),.A(g6623),.B(g12536));
  AND2 AND2_991(.VSS(VSS),.VDD(VDD),.Y(g13702),.A(g7802),.B(g12537));
  AND2 AND2_992(.VSS(VSS),.VDD(VDD),.Y(g13703),.A(g8018),.B(g11848));
  AND2 AND2_993(.VSS(VSS),.VDD(VDD),.Y(g13704),.A(g7581),.B(g12542));
  AND2 AND2_994(.VSS(VSS),.VDD(VDD),.Y(g13705),.A(g12776),.B(g8673));
  AND2 AND2_995(.VSS(VSS),.VDD(VDD),.Y(g13738),.A(g6887),.B(g12545));
  AND2 AND2_996(.VSS(VSS),.VDD(VDD),.Y(g13739),.A(g7815),.B(g12546));
  AND2 AND2_997(.VSS(VSS),.VDD(VDD),.Y(g13740),.A(g6636),.B(g12547));
  AND2 AND2_998(.VSS(VSS),.VDD(VDD),.Y(g13755),.A(g7347),.B(g12551));
  AND2 AND2_999(.VSS(VSS),.VDD(VDD),.Y(g13787),.A(g7967),.B(g11923));
  AND2 AND2_1000(.VSS(VSS),.VDD(VDD),.Y(g13788),.A(g6897),.B(g12553));
  AND2 AND2_1001(.VSS(VSS),.VDD(VDD),.Y(g13789),.A(g7140),.B(g12554));
  AND2 AND2_1002(.VSS(VSS),.VDD(VDD),.Y(g13790),.A(g7475),.B(g12558));
  AND2 AND2_1003(.VSS(VSS),.VDD(VDD),.Y(g13796),.A(g7477),.B(g12559));
  AND2 AND2_1004(.VSS(VSS),.VDD(VDD),.Y(g13815),.A(g7139),.B(g12560));
  AND2 AND2_1005(.VSS(VSS),.VDD(VDD),.Y(g13816),.A(g7530),.B(g12596));
  AND2 AND2_1006(.VSS(VSS),.VDD(VDD),.Y(g13818),.A(g7531),.B(g12597));
  AND2 AND2_1007(.VSS(VSS),.VDD(VDD),.Y(g13824),.A(g7533),.B(g12598));
  AND2 AND2_1008(.VSS(VSS),.VDD(VDD),.Y(g13833),.A(g7919),.B(g12009));
  AND2 AND2_1009(.VSS(VSS),.VDD(VDD),.Y(g13834),.A(g7336),.B(g12599));
  AND2 AND2_1010(.VSS(VSS),.VDD(VDD),.Y(g13835),.A(g7461),.B(g12600));
  AND2 AND2_1011(.VSS(VSS),.VDD(VDD),.Y(g13837),.A(g7556),.B(g12642));
  AND2 AND2_1012(.VSS(VSS),.VDD(VDD),.Y(g13839),.A(g7557),.B(g12643));
  AND2 AND2_1013(.VSS(VSS),.VDD(VDD),.Y(g13845),.A(g7559),.B(g12644));
  AND2 AND2_1014(.VSS(VSS),.VDD(VDD),.Y(g13846),.A(g7460),.B(g12645));
  AND2 AND2_1015(.VSS(VSS),.VDD(VDD),.Y(g13847),.A(g7521),.B(g12646));
  AND2 AND2_1016(.VSS(VSS),.VDD(VDD),.Y(g13851),.A(g7579),.B(g12688));
  AND2 AND2_1017(.VSS(VSS),.VDD(VDD),.Y(g13853),.A(g7580),.B(g12689));
  AND2 AND2_1018(.VSS(VSS),.VDD(VDD),.Y(g13854),.A(g5349),.B(g12690));
  AND2 AND2_1019(.VSS(VSS),.VDD(VDD),.Y(g13855),.A(g7541),.B(g12691));
  AND2 AND2_1020(.VSS(VSS),.VDD(VDD),.Y(g13860),.A(g7593),.B(g12742));
  AND2 AND2_1021(.VSS(VSS),.VDD(VDD),.Y(g13862),.A(g5366),.B(g12743));
  AND2 AND2_1022(.VSS(VSS),.VDD(VDD),.Y(g13865),.A(g548),.B(g12748));
  AND2 AND2_1023(.VSS(VSS),.VDD(VDD),.Y(g13870),.A(g7582),.B(g12768));
  AND2 AND2_1024(.VSS(VSS),.VDD(VDD),.Y(g13871),.A(g7898),.B(g12775));
  AND2 AND2_1025(.VSS(VSS),.VDD(VDD),.Y(g13878),.A(g7610),.B(g12782));
  AND2 AND2_1026(.VSS(VSS),.VDD(VDD),.Y(g13880),.A(g1234),.B(g12790));
  AND2 AND2_1027(.VSS(VSS),.VDD(VDD),.Y(g13884),.A(g7594),.B(g12807));
  AND2 AND2_1028(.VSS(VSS),.VDD(VDD),.Y(g13892),.A(g7616),.B(g12815));
  AND2 AND2_1029(.VSS(VSS),.VDD(VDD),.Y(g13900),.A(g7619),.B(g12821));
  AND2 AND2_1030(.VSS(VSS),.VDD(VDD),.Y(g13902),.A(g1928),.B(g12829));
  AND2 AND2_1031(.VSS(VSS),.VDD(VDD),.Y(g13904),.A(g7337),.B(g12843));
  AND2 AND2_1032(.VSS(VSS),.VDD(VDD),.Y(g13905),.A(g7925),.B(g12847));
  AND2 AND2_1033(.VSS(VSS),.VDD(VDD),.Y(g13913),.A(g7623),.B(g12850));
  AND2 AND2_1034(.VSS(VSS),.VDD(VDD),.Y(g13914),.A(g7626),.B(g12851));
  AND2 AND2_1035(.VSS(VSS),.VDD(VDD),.Y(g13933),.A(g7632),.B(g12853));
  AND2 AND2_1036(.VSS(VSS),.VDD(VDD),.Y(g13941),.A(g7635),.B(g12859));
  AND2 AND2_1037(.VSS(VSS),.VDD(VDD),.Y(g13943),.A(g2622),.B(g12867));
  AND2 AND2_1038(.VSS(VSS),.VDD(VDD),.Y(g13944),.A(g7141),.B(g12874));
  AND2 AND2_1039(.VSS(VSS),.VDD(VDD),.Y(g13952),.A(g7643),.B(g12881));
  AND2 AND2_1040(.VSS(VSS),.VDD(VDD),.Y(g13953),.A(g7646),.B(g12882));
  AND2 AND2_1041(.VSS(VSS),.VDD(VDD),.Y(g13969),.A(g7652),.B(g12891));
  AND2 AND2_1042(.VSS(VSS),.VDD(VDD),.Y(g13970),.A(g7655),.B(g12892));
  AND2 AND2_1043(.VSS(VSS),.VDD(VDD),.Y(g13989),.A(g7661),.B(g12894));
  AND2 AND2_1044(.VSS(VSS),.VDD(VDD),.Y(g13997),.A(g7664),.B(g12900));
  AND2 AND2_1045(.VSS(VSS),.VDD(VDD),.Y(g13998),.A(g7972),.B(g12907));
  AND2 AND2_1046(.VSS(VSS),.VDD(VDD),.Y(g14006),.A(g7670),.B(g12914));
  AND2 AND2_1047(.VSS(VSS),.VDD(VDD),.Y(g14007),.A(g7673),.B(g12915));
  AND2 AND2_1048(.VSS(VSS),.VDD(VDD),.Y(g14022),.A(g7679),.B(g12921));
  AND2 AND2_1049(.VSS(VSS),.VDD(VDD),.Y(g14023),.A(g7682),.B(g12922));
  AND2 AND2_1050(.VSS(VSS),.VDD(VDD),.Y(g14039),.A(g7688),.B(g12931));
  AND2 AND2_1051(.VSS(VSS),.VDD(VDD),.Y(g14040),.A(g7691),.B(g12932));
  AND2 AND2_1052(.VSS(VSS),.VDD(VDD),.Y(g14059),.A(g7697),.B(g12934));
  AND2 AND2_1053(.VSS(VSS),.VDD(VDD),.Y(g14067),.A(g7703),.B(g12940));
  AND2 AND2_1054(.VSS(VSS),.VDD(VDD),.Y(g14097),.A(g7706),.B(g12943));
  AND2 AND2_1055(.VSS(VSS),.VDD(VDD),.Y(g14098),.A(g7709),.B(g12944));
  AND2 AND2_1056(.VSS(VSS),.VDD(VDD),.Y(g14113),.A(g7715),.B(g12950));
  AND2 AND2_1057(.VSS(VSS),.VDD(VDD),.Y(g14114),.A(g7718),.B(g12951));
  AND2 AND2_1058(.VSS(VSS),.VDD(VDD),.Y(g14130),.A(g7724),.B(g12960));
  AND2 AND2_1059(.VSS(VSS),.VDD(VDD),.Y(g14131),.A(g7727),.B(g12961));
  AND2 AND2_1060(.VSS(VSS),.VDD(VDD),.Y(g14143),.A(g8026),.B(g12965));
  AND2 AND2_1061(.VSS(VSS),.VDD(VDD),.Y(g14182),.A(g7733),.B(g12969));
  AND2 AND2_1062(.VSS(VSS),.VDD(VDD),.Y(g14212),.A(g7736),.B(g12972));
  AND2 AND2_1063(.VSS(VSS),.VDD(VDD),.Y(g14213),.A(g7739),.B(g12973));
  AND2 AND2_1064(.VSS(VSS),.VDD(VDD),.Y(g14228),.A(g7745),.B(g12979));
  AND2 AND2_1065(.VSS(VSS),.VDD(VDD),.Y(g14229),.A(g7748),.B(g12980));
  AND2 AND2_1066(.VSS(VSS),.VDD(VDD),.Y(g14297),.A(g7757),.B(g12993));
  AND2 AND2_1067(.VSS(VSS),.VDD(VDD),.Y(g14327),.A(g7760),.B(g12996));
  AND2 AND2_1068(.VSS(VSS),.VDD(VDD),.Y(g14328),.A(g7763),.B(g12997));
  AND2 AND2_1069(.VSS(VSS),.VDD(VDD),.Y(g14336),.A(g8099),.B(g12998));
  AND2 AND2_1070(.VSS(VSS),.VDD(VDD),.Y(g14419),.A(g7779),.B(g13003));
  AND2 AND2_1071(.VSS(VSS),.VDD(VDD),.Y(g14690),.A(g7841),.B(g13101));
  AND2 AND2_1072(.VSS(VSS),.VDD(VDD),.Y(g14724),.A(g7861),.B(g13117));
  AND2 AND2_1073(.VSS(VSS),.VDD(VDD),.Y(g14752),.A(g7891),.B(g13130));
  AND2 AND2_1074(.VSS(VSS),.VDD(VDD),.Y(g14767),.A(g13245),.B(g10765));
  AND2 AND2_1075(.VSS(VSS),.VDD(VDD),.Y(g14773),.A(g7915),.B(g13141));
  AND2 AND2_1076(.VSS(VSS),.VDD(VDD),.Y(g14884),.A(g8169),.B(g12548));
  AND2 AND2_1077(.VSS(VSS),.VDD(VDD),.Y(g14894),.A(g3940),.B(g13148));
  AND2 AND2_1078(.VSS(VSS),.VDD(VDD),.Y(g14956),.A(g11059),.B(g13151));
  AND2 AND2_1079(.VSS(VSS),.VDD(VDD),.Y(g14957),.A(g4015),.B(g13152));
  AND2 AND2_1080(.VSS(VSS),.VDD(VDD),.Y(g14958),.A(g4016),.B(g13153));
  AND2 AND2_1081(.VSS(VSS),.VDD(VDD),.Y(g14975),.A(g4047),.B(g13154));
  AND2 AND2_1082(.VSS(VSS),.VDD(VDD),.Y(g15020),.A(g8090),.B(g12561));
  AND2 AND2_1083(.VSS(VSS),.VDD(VDD),.Y(g15030),.A(g4110),.B(g13158));
  AND2 AND2_1084(.VSS(VSS),.VDD(VDD),.Y(g15031),.A(g4111),.B(g13159));
  AND2 AND2_1085(.VSS(VSS),.VDD(VDD),.Y(g15046),.A(g4142),.B(g13161));
  AND2 AND2_1086(.VSS(VSS),.VDD(VDD),.Y(g15047),.A(g4143),.B(g13162));
  AND2 AND2_1087(.VSS(VSS),.VDD(VDD),.Y(g15064),.A(g4174),.B(g13163));
  AND2 AND2_1088(.VSS(VSS),.VDD(VDD),.Y(g15093),.A(g7869),.B(g12601));
  AND2 AND2_1089(.VSS(VSS),.VDD(VDD),.Y(g15094),.A(g7872),.B(g12604));
  AND2 AND2_1090(.VSS(VSS),.VDD(VDD),.Y(g15104),.A(g4220),.B(g13167));
  AND2 AND2_1091(.VSS(VSS),.VDD(VDD),.Y(g15105),.A(g4224),.B(g13168));
  AND2 AND2_1092(.VSS(VSS),.VDD(VDD),.Y(g15126),.A(g4249),.B(g13169));
  AND2 AND2_1093(.VSS(VSS),.VDD(VDD),.Y(g15127),.A(g4250),.B(g13170));
  AND2 AND2_1094(.VSS(VSS),.VDD(VDD),.Y(g15142),.A(g4281),.B(g13172));
  AND2 AND2_1095(.VSS(VSS),.VDD(VDD),.Y(g15143),.A(g4282),.B(g13173));
  AND2 AND2_1096(.VSS(VSS),.VDD(VDD),.Y(g15160),.A(g4313),.B(g13174));
  AND2 AND2_1097(.VSS(VSS),.VDD(VDD),.Y(g15171),.A(g8015),.B(g12647));
  AND2 AND2_1098(.VSS(VSS),.VDD(VDD),.Y(g15172),.A(g4346),.B(g13176));
  AND2 AND2_1099(.VSS(VSS),.VDD(VDD),.Y(g15173),.A(g4347),.B(g13177));
  AND2 AND2_1100(.VSS(VSS),.VDD(VDD),.Y(g15178),.A(g640),.B(g12651));
  AND2 AND2_1101(.VSS(VSS),.VDD(VDD),.Y(g15196),.A(g4375),.B(g13178));
  AND2 AND2_1102(.VSS(VSS),.VDD(VDD),.Y(g15197),.A(g4379),.B(g13179));
  AND2 AND2_1103(.VSS(VSS),.VDD(VDD),.Y(g15218),.A(g4404),.B(g13180));
  AND2 AND2_1104(.VSS(VSS),.VDD(VDD),.Y(g15219),.A(g4405),.B(g13181));
  AND2 AND2_1105(.VSS(VSS),.VDD(VDD),.Y(g15234),.A(g4436),.B(g13183));
  AND2 AND2_1106(.VSS(VSS),.VDD(VDD),.Y(g15235),.A(g4437),.B(g13184));
  AND2 AND2_1107(.VSS(VSS),.VDD(VDD),.Y(g15243),.A(g7849),.B(g12692));
  AND2 AND2_1108(.VSS(VSS),.VDD(VDD),.Y(g15244),.A(g7852),.B(g12695));
  AND2 AND2_1109(.VSS(VSS),.VDD(VDD),.Y(g15245),.A(g4474),.B(g13185));
  AND2 AND2_1110(.VSS(VSS),.VDD(VDD),.Y(g15246),.A(g4475),.B(g13186));
  AND2 AND2_1111(.VSS(VSS),.VDD(VDD),.Y(g15247),.A(g4479),.B(g13187));
  AND2 AND2_1112(.VSS(VSS),.VDD(VDD),.Y(g15257),.A(g4357),.B(g12702));
  AND2 AND2_1113(.VSS(VSS),.VDD(VDD),.Y(g15258),.A(g4515),.B(g13188));
  AND2 AND2_1114(.VSS(VSS),.VDD(VDD),.Y(g15259),.A(g4516),.B(g13189));
  AND2 AND2_1115(.VSS(VSS),.VDD(VDD),.Y(g15264),.A(g1326),.B(g12705));
  AND2 AND2_1116(.VSS(VSS),.VDD(VDD),.Y(g15282),.A(g4544),.B(g13190));
  AND2 AND2_1117(.VSS(VSS),.VDD(VDD),.Y(g15283),.A(g4548),.B(g13191));
  AND2 AND2_1118(.VSS(VSS),.VDD(VDD),.Y(g15304),.A(g4573),.B(g13192));
  AND2 AND2_1119(.VSS(VSS),.VDD(VDD),.Y(g15305),.A(g4574),.B(g13193));
  AND2 AND2_1120(.VSS(VSS),.VDD(VDD),.Y(g15320),.A(g7964),.B(g12744));
  AND2 AND2_1121(.VSS(VSS),.VDD(VDD),.Y(g15321),.A(g4601),.B(g13195));
  AND2 AND2_1122(.VSS(VSS),.VDD(VDD),.Y(g15324),.A(g4609),.B(g13196));
  AND2 AND2_1123(.VSS(VSS),.VDD(VDD),.Y(g15325),.A(g4610),.B(g13197));
  AND2 AND2_1124(.VSS(VSS),.VDD(VDD),.Y(g15335),.A(g4489),.B(g12749));
  AND2 AND2_1125(.VSS(VSS),.VDD(VDD),.Y(g15336),.A(g4492),.B(g12752));
  AND2 AND2_1126(.VSS(VSS),.VDD(VDD),.Y(g15337),.A(g4650),.B(g13198));
  AND2 AND2_1127(.VSS(VSS),.VDD(VDD),.Y(g15338),.A(g4651),.B(g13199));
  AND2 AND2_1128(.VSS(VSS),.VDD(VDD),.Y(g15339),.A(g4655),.B(g13200));
  AND2 AND2_1129(.VSS(VSS),.VDD(VDD),.Y(g15349),.A(g4526),.B(g12759));
  AND2 AND2_1130(.VSS(VSS),.VDD(VDD),.Y(g15350),.A(g4691),.B(g13201));
  AND2 AND2_1131(.VSS(VSS),.VDD(VDD),.Y(g15351),.A(g4692),.B(g13202));
  AND2 AND2_1132(.VSS(VSS),.VDD(VDD),.Y(g15356),.A(g2020),.B(g12762));
  AND2 AND2_1133(.VSS(VSS),.VDD(VDD),.Y(g15374),.A(g4720),.B(g13203));
  AND2 AND2_1134(.VSS(VSS),.VDD(VDD),.Y(g15375),.A(g4724),.B(g13204));
  AND2 AND2_1135(.VSS(VSS),.VDD(VDD),.Y(g15388),.A(g7834),.B(g12769));
  AND2 AND2_1136(.VSS(VSS),.VDD(VDD),.Y(g15389),.A(g8246),.B(g12772));
  AND2 AND2_1137(.VSS(VSS),.VDD(VDD),.Y(g15391),.A(g4752),.B(g13205));
  AND2 AND2_1138(.VSS(VSS),.VDD(VDD),.Y(g15392),.A(g4753),.B(g13206));
  AND2 AND2_1139(.VSS(VSS),.VDD(VDD),.Y(g15402),.A(g4620),.B(g12783));
  AND2 AND2_1140(.VSS(VSS),.VDD(VDD),.Y(g15403),.A(g4623),.B(g12786));
  AND2 AND2_1141(.VSS(VSS),.VDD(VDD),.Y(g15407),.A(g4778),.B(g13207));
  AND2 AND2_1142(.VSS(VSS),.VDD(VDD),.Y(g15410),.A(g4786),.B(g13208));
  AND2 AND2_1143(.VSS(VSS),.VDD(VDD),.Y(g15411),.A(g4787),.B(g13209));
  AND2 AND2_1144(.VSS(VSS),.VDD(VDD),.Y(g15421),.A(g4665),.B(g12791));
  AND2 AND2_1145(.VSS(VSS),.VDD(VDD),.Y(g15422),.A(g4668),.B(g12794));
  AND2 AND2_1146(.VSS(VSS),.VDD(VDD),.Y(g15423),.A(g4827),.B(g13210));
  AND2 AND2_1147(.VSS(VSS),.VDD(VDD),.Y(g15424),.A(g4828),.B(g13211));
  AND2 AND2_1148(.VSS(VSS),.VDD(VDD),.Y(g15425),.A(g4832),.B(g13212));
  AND2 AND2_1149(.VSS(VSS),.VDD(VDD),.Y(g15435),.A(g4702),.B(g12801));
  AND2 AND2_1150(.VSS(VSS),.VDD(VDD),.Y(g15436),.A(g4868),.B(g13213));
  AND2 AND2_1151(.VSS(VSS),.VDD(VDD),.Y(g15437),.A(g4869),.B(g13214));
  AND2 AND2_1152(.VSS(VSS),.VDD(VDD),.Y(g15442),.A(g2714),.B(g12804));
  AND2 AND2_1153(.VSS(VSS),.VDD(VDD),.Y(g15452),.A(g7916),.B(g12808));
  AND2 AND2_1154(.VSS(VSS),.VDD(VDD),.Y(g15453),.A(g6898),.B(g12811));
  AND2 AND2_1155(.VSS(VSS),.VDD(VDD),.Y(g15459),.A(g4897),.B(g13218));
  AND2 AND2_1156(.VSS(VSS),.VDD(VDD),.Y(g15460),.A(g4898),.B(g13219));
  AND2 AND2_1157(.VSS(VSS),.VDD(VDD),.Y(g15470),.A(g4763),.B(g12816));
  AND2 AND2_1158(.VSS(VSS),.VDD(VDD),.Y(g15475),.A(g4928),.B(g13220));
  AND2 AND2_1159(.VSS(VSS),.VDD(VDD),.Y(g15476),.A(g4929),.B(g13221));
  AND2 AND2_1160(.VSS(VSS),.VDD(VDD),.Y(g15486),.A(g4797),.B(g12822));
  AND2 AND2_1161(.VSS(VSS),.VDD(VDD),.Y(g15487),.A(g4800),.B(g12825));
  AND2 AND2_1162(.VSS(VSS),.VDD(VDD),.Y(g15491),.A(g4954),.B(g13222));
  AND2 AND2_1163(.VSS(VSS),.VDD(VDD),.Y(g15494),.A(g4962),.B(g13223));
  AND2 AND2_1164(.VSS(VSS),.VDD(VDD),.Y(g15495),.A(g4963),.B(g13224));
  AND2 AND2_1165(.VSS(VSS),.VDD(VDD),.Y(g15505),.A(g4842),.B(g12830));
  AND2 AND2_1166(.VSS(VSS),.VDD(VDD),.Y(g15506),.A(g4845),.B(g12833));
  AND2 AND2_1167(.VSS(VSS),.VDD(VDD),.Y(g15507),.A(g5003),.B(g13225));
  AND2 AND2_1168(.VSS(VSS),.VDD(VDD),.Y(g15508),.A(g5004),.B(g13226));
  AND2 AND2_1169(.VSS(VSS),.VDD(VDD),.Y(g15509),.A(g5008),.B(g13227));
  AND2 AND2_1170(.VSS(VSS),.VDD(VDD),.Y(g15519),.A(g4879),.B(g12840));
  AND2 AND2_1171(.VSS(VSS),.VDD(VDD),.Y(g15520),.A(g8172),.B(g12844));
  AND2 AND2_1172(.VSS(VSS),.VDD(VDD),.Y(g15526),.A(g5033),.B(g13232));
  AND2 AND2_1173(.VSS(VSS),.VDD(VDD),.Y(g15527),.A(g5034),.B(g13233));
  AND2 AND2_1174(.VSS(VSS),.VDD(VDD),.Y(g15545),.A(g5056),.B(g13237));
  AND2 AND2_1175(.VSS(VSS),.VDD(VDD),.Y(g15546),.A(g5057),.B(g13238));
  AND2 AND2_1176(.VSS(VSS),.VDD(VDD),.Y(g15556),.A(g4939),.B(g12854));
  AND2 AND2_1177(.VSS(VSS),.VDD(VDD),.Y(g15561),.A(g5087),.B(g13239));
  AND2 AND2_1178(.VSS(VSS),.VDD(VDD),.Y(g15562),.A(g5088),.B(g13240));
  AND2 AND2_1179(.VSS(VSS),.VDD(VDD),.Y(g15572),.A(g4973),.B(g12860));
  AND2 AND2_1180(.VSS(VSS),.VDD(VDD),.Y(g15573),.A(g4976),.B(g12863));
  AND2 AND2_1181(.VSS(VSS),.VDD(VDD),.Y(g15577),.A(g5113),.B(g13241));
  AND2 AND2_1182(.VSS(VSS),.VDD(VDD),.Y(g15580),.A(g5121),.B(g13242));
  AND2 AND2_1183(.VSS(VSS),.VDD(VDD),.Y(g15581),.A(g5122),.B(g13243));
  AND2 AND2_1184(.VSS(VSS),.VDD(VDD),.Y(g15591),.A(g5018),.B(g12868));
  AND2 AND2_1185(.VSS(VSS),.VDD(VDD),.Y(g15592),.A(g5021),.B(g12871));
  AND2 AND2_1186(.VSS(VSS),.VDD(VDD),.Y(g15593),.A(g7897),.B(g13244));
  AND2 AND2_1187(.VSS(VSS),.VDD(VDD),.Y(g15594),.A(g5148),.B(g13249));
  AND2 AND2_1188(.VSS(VSS),.VDD(VDD),.Y(g15595),.A(g5149),.B(g13250));
  AND2 AND2_1189(.VSS(VSS),.VDD(VDD),.Y(g15604),.A(g5162),.B(g13255));
  AND2 AND2_1190(.VSS(VSS),.VDD(VDD),.Y(g15605),.A(g5163),.B(g13256));
  AND2 AND2_1191(.VSS(VSS),.VDD(VDD),.Y(g15623),.A(g5185),.B(g13260));
  AND2 AND2_1192(.VSS(VSS),.VDD(VDD),.Y(g15624),.A(g5186),.B(g13261));
  AND2 AND2_1193(.VSS(VSS),.VDD(VDD),.Y(g15634),.A(g5098),.B(g12895));
  AND2 AND2_1194(.VSS(VSS),.VDD(VDD),.Y(g15639),.A(g5216),.B(g13262));
  AND2 AND2_1195(.VSS(VSS),.VDD(VDD),.Y(g15640),.A(g5217),.B(g13263));
  AND2 AND2_1196(.VSS(VSS),.VDD(VDD),.Y(g15650),.A(g5132),.B(g12901));
  AND2 AND2_1197(.VSS(VSS),.VDD(VDD),.Y(g15651),.A(g5135),.B(g12904));
  AND2 AND2_1198(.VSS(VSS),.VDD(VDD),.Y(g15658),.A(g8177),.B(g13264));
  AND2 AND2_1199(.VSS(VSS),.VDD(VDD),.Y(g15666),.A(g5233),.B(g13268));
  AND2 AND2_1200(.VSS(VSS),.VDD(VDD),.Y(g15670),.A(g5241),.B(g13272));
  AND2 AND2_1201(.VSS(VSS),.VDD(VDD),.Y(g15671),.A(g5242),.B(g13273));
  AND2 AND2_1202(.VSS(VSS),.VDD(VDD),.Y(g15680),.A(g5255),.B(g13278));
  AND2 AND2_1203(.VSS(VSS),.VDD(VDD),.Y(g15681),.A(g5256),.B(g13279));
  AND2 AND2_1204(.VSS(VSS),.VDD(VDD),.Y(g15699),.A(g5278),.B(g13283));
  AND2 AND2_1205(.VSS(VSS),.VDD(VDD),.Y(g15700),.A(g5279),.B(g13284));
  AND2 AND2_1206(.VSS(VSS),.VDD(VDD),.Y(g15710),.A(g5227),.B(g12935));
  AND2 AND2_1207(.VSS(VSS),.VDD(VDD),.Y(g15717),.A(g7924),.B(g13285));
  AND2 AND2_1208(.VSS(VSS),.VDD(VDD),.Y(g15725),.A(g5296),.B(g13293));
  AND2 AND2_1209(.VSS(VSS),.VDD(VDD),.Y(g15729),.A(g5304),.B(g13297));
  AND2 AND2_1210(.VSS(VSS),.VDD(VDD),.Y(g15730),.A(g5305),.B(g13298));
  AND2 AND2_1211(.VSS(VSS),.VDD(VDD),.Y(g15739),.A(g5318),.B(g13303));
  AND2 AND2_1212(.VSS(VSS),.VDD(VDD),.Y(g15740),.A(g5319),.B(g13304));
  AND2 AND2_1213(.VSS(VSS),.VDD(VDD),.Y(g15753),.A(g7542),.B(g12962));
  AND2 AND2_1214(.VSS(VSS),.VDD(VDD),.Y(g15754),.A(g7837),.B(g13308));
  AND2 AND2_1215(.VSS(VSS),.VDD(VDD),.Y(g15755),.A(g8178),.B(g13309));
  AND2 AND2_1216(.VSS(VSS),.VDD(VDD),.Y(g15765),.A(g5333),.B(g13324));
  AND2 AND2_1217(.VSS(VSS),.VDD(VDD),.Y(g15769),.A(g5341),.B(g13328));
  AND2 AND2_1218(.VSS(VSS),.VDD(VDD),.Y(g15770),.A(g5342),.B(g13329));
  AND3 AND3_10(.VSS(VSS),.VDD(VDD),.Y(I22028),.A(g13004),.B(g3018),.C(g7549));
  AND3 AND3_11(.VSS(VSS),.VDD(VDD),.Y(g15780),.A(g7471),.B(g3032),.C(I22028));
  AND2 AND2_1219(.VSS(VSS),.VDD(VDD),.Y(g15781),.A(g7971),.B(g13330));
  AND2 AND2_1220(.VSS(VSS),.VDD(VDD),.Y(g15793),.A(g5361),.B(g13347));
  AND2 AND2_1221(.VSS(VSS),.VDD(VDD),.Y(g15801),.A(g7856),.B(g13351));
  AND2 AND2_1222(.VSS(VSS),.VDD(VDD),.Y(g15802),.A(g8253),.B(g13352));
  AND2 AND2_1223(.VSS(VSS),.VDD(VDD),.Y(g15817),.A(g8025),.B(g13373));
  AND2 AND2_1224(.VSS(VSS),.VDD(VDD),.Y(g15828),.A(g7877),.B(g13398));
  AND2 AND2_1225(.VSS(VSS),.VDD(VDD),.Y(g15829),.A(g7857),.B(g13400));
  AND2 AND2_1226(.VSS(VSS),.VDD(VDD),.Y(g15840),.A(g8098),.B(g11620));
  AND2 AND2_1227(.VSS(VSS),.VDD(VDD),.Y(g15852),.A(g7878),.B(g11642));
  AND3 AND3_12(.VSS(VSS),.VDD(VDD),.Y(I22136),.A(g13082),.B(g2912),.C(g7522));
  AND3 AND3_13(.VSS(VSS),.VDD(VDD),.Y(g15902),.A(g7607),.B(g2920),.C(I22136));
  AND2 AND2_1228(.VSS(VSS),.VDD(VDD),.Y(g15998),.A(g5469),.B(g11732));
  AND2 AND2_1229(.VSS(VSS),.VDD(VDD),.Y(g16003),.A(g12013),.B(g10826));
  AND2 AND2_1230(.VSS(VSS),.VDD(VDD),.Y(g16004),.A(g5587),.B(g11734));
  AND2 AND2_1231(.VSS(VSS),.VDD(VDD),.Y(g16008),.A(g5504),.B(g11735));
  AND2 AND2_1232(.VSS(VSS),.VDD(VDD),.Y(g16009),.A(g12071),.B(g10843));
  AND2 AND2_1233(.VSS(VSS),.VDD(VDD),.Y(g16010),.A(g7639),.B(g11736));
  AND2 AND2_1234(.VSS(VSS),.VDD(VDD),.Y(g16015),.A(g12013),.B(g10859));
  AND2 AND2_1235(.VSS(VSS),.VDD(VDD),.Y(g16016),.A(g5601),.B(g11740));
  AND2 AND2_1236(.VSS(VSS),.VDD(VDD),.Y(g16017),.A(g12130),.B(g10862));
  AND2 AND2_1237(.VSS(VSS),.VDD(VDD),.Y(g16018),.A(g6149),.B(g11741));
  AND2 AND2_1238(.VSS(VSS),.VDD(VDD),.Y(g16019),.A(g5507),.B(g11742));
  AND2 AND2_1239(.VSS(VSS),.VDD(VDD),.Y(g16028),.A(g5543),.B(g11745));
  AND2 AND2_1240(.VSS(VSS),.VDD(VDD),.Y(g16029),.A(g12071),.B(g10877));
  AND2 AND2_1241(.VSS(VSS),.VDD(VDD),.Y(g16030),.A(g7667),.B(g11746));
  AND2 AND2_1242(.VSS(VSS),.VDD(VDD),.Y(g16031),.A(g6227),.B(g11747));
  AND2 AND2_1243(.VSS(VSS),.VDD(VDD),.Y(g16032),.A(g12187),.B(g10883));
  AND2 AND2_1244(.VSS(VSS),.VDD(VDD),.Y(g16033),.A(g5546),.B(g11748));
  AND2 AND2_1245(.VSS(VSS),.VDD(VDD),.Y(g16045),.A(g12013),.B(g10892));
  AND2 AND2_1246(.VSS(VSS),.VDD(VDD),.Y(g16046),.A(g5618),.B(g11761));
  AND2 AND2_1247(.VSS(VSS),.VDD(VDD),.Y(g16047),.A(g12130),.B(g10895));
  AND2 AND2_1248(.VSS(VSS),.VDD(VDD),.Y(g16048),.A(g6170),.B(g11762));
  AND2 AND2_1249(.VSS(VSS),.VDD(VDD),.Y(g16049),.A(g6638),.B(g11763));
  AND2 AND2_1250(.VSS(VSS),.VDD(VDD),.Y(g16050),.A(g5590),.B(g11764));
  AND2 AND2_1251(.VSS(VSS),.VDD(VDD),.Y(g16051),.A(g12235),.B(g10901));
  AND2 AND2_1252(.VSS(VSS),.VDD(VDD),.Y(g16052),.A(g5591),.B(g11765));
  AND2 AND2_1253(.VSS(VSS),.VDD(VDD),.Y(g16053),.A(g297),.B(g11770));
  AND2 AND2_1254(.VSS(VSS),.VDD(VDD),.Y(g16066),.A(g12071),.B(g10912));
  AND2 AND2_1255(.VSS(VSS),.VDD(VDD),.Y(g16067),.A(g7700),.B(g11774));
  AND2 AND2_1256(.VSS(VSS),.VDD(VDD),.Y(g16068),.A(g6310),.B(g11775));
  AND2 AND2_1257(.VSS(VSS),.VDD(VDD),.Y(g16069),.A(g5346),.B(g11776));
  AND2 AND2_1258(.VSS(VSS),.VDD(VDD),.Y(g16070),.A(g12187),.B(g10921));
  AND2 AND2_1259(.VSS(VSS),.VDD(VDD),.Y(g16071),.A(g5604),.B(g11777));
  AND2 AND2_1260(.VSS(VSS),.VDD(VDD),.Y(g16072),.A(g12275),.B(g10924));
  AND2 AND2_1261(.VSS(VSS),.VDD(VDD),.Y(g16073),.A(g5605),.B(g11778));
  AND2 AND2_1262(.VSS(VSS),.VDD(VDD),.Y(g16074),.A(g5646),.B(g11782));
  AND2 AND2_1263(.VSS(VSS),.VDD(VDD),.Y(g16081),.A(g3304),.B(g11783));
  AND2 AND2_1264(.VSS(VSS),.VDD(VDD),.Y(g16089),.A(g984),.B(g11787));
  AND2 AND2_1265(.VSS(VSS),.VDD(VDD),.Y(g16100),.A(g12130),.B(g10937));
  AND2 AND2_1266(.VSS(VSS),.VDD(VDD),.Y(g16101),.A(g6197),.B(g11794));
  AND2 AND2_1267(.VSS(VSS),.VDD(VDD),.Y(g16102),.A(g6905),.B(g11795));
  AND2 AND2_1268(.VSS(VSS),.VDD(VDD),.Y(g16103),.A(g5621),.B(g11796));
  AND2 AND2_1269(.VSS(VSS),.VDD(VDD),.Y(g16104),.A(g12235),.B(g10946));
  AND2 AND2_1270(.VSS(VSS),.VDD(VDD),.Y(g16105),.A(g5622),.B(g11797));
  AND2 AND2_1271(.VSS(VSS),.VDD(VDD),.Y(g16106),.A(g12308),.B(g10949));
  AND2 AND2_1272(.VSS(VSS),.VDD(VDD),.Y(g16107),.A(g5666),.B(g11801));
  AND2 AND2_1273(.VSS(VSS),.VDD(VDD),.Y(g16108),.A(g5667),.B(g11802));
  AND2 AND2_1274(.VSS(VSS),.VDD(VDD),.Y(g16109),.A(g8277),.B(g11803));
  AND2 AND2_1275(.VSS(VSS),.VDD(VDD),.Y(g16110),.A(g516),.B(g11804));
  AND2 AND2_1276(.VSS(VSS),.VDD(VDD),.Y(g16111),.A(g5551),.B(g13215));
  AND2 AND2_1277(.VSS(VSS),.VDD(VDD),.Y(g16112),.A(g5684),.B(g11808));
  AND2 AND2_1278(.VSS(VSS),.VDD(VDD),.Y(g16119),.A(g3460),.B(g11809));
  AND2 AND2_1279(.VSS(VSS),.VDD(VDD),.Y(g16127),.A(g1678),.B(g11813));
  AND2 AND2_1280(.VSS(VSS),.VDD(VDD),.Y(g16133),.A(g6444),.B(g11817));
  AND2 AND2_1281(.VSS(VSS),.VDD(VDD),.Y(g16134),.A(g5363),.B(g11818));
  AND2 AND2_1282(.VSS(VSS),.VDD(VDD),.Y(g16135),.A(g12187),.B(g10980));
  AND2 AND2_1283(.VSS(VSS),.VDD(VDD),.Y(g16136),.A(g5640),.B(g11819));
  AND2 AND2_1284(.VSS(VSS),.VDD(VDD),.Y(g16137),.A(g12275),.B(g10983));
  AND2 AND2_1285(.VSS(VSS),.VDD(VDD),.Y(g16138),.A(g5641),.B(g11820));
  AND2 AND2_1286(.VSS(VSS),.VDD(VDD),.Y(g16139),.A(g5704),.B(g11824));
  AND2 AND2_1287(.VSS(VSS),.VDD(VDD),.Y(g16140),.A(g5705),.B(g11825));
  AND2 AND2_1288(.VSS(VSS),.VDD(VDD),.Y(g16141),.A(g5706),.B(g11826));
  AND2 AND2_1289(.VSS(VSS),.VDD(VDD),.Y(g16152),.A(g517),.B(g11829));
  AND2 AND2_1290(.VSS(VSS),.VDD(VDD),.Y(g16153),.A(g5592),.B(g13229));
  AND2 AND2_1291(.VSS(VSS),.VDD(VDD),.Y(g16158),.A(g5718),.B(g11834));
  AND2 AND2_1292(.VSS(VSS),.VDD(VDD),.Y(g16159),.A(g5719),.B(g11835));
  AND2 AND2_1293(.VSS(VSS),.VDD(VDD),.Y(g16160),.A(g8286),.B(g11836));
  AND2 AND2_1294(.VSS(VSS),.VDD(VDD),.Y(g16161),.A(g1202),.B(g11837));
  AND2 AND2_1295(.VSS(VSS),.VDD(VDD),.Y(g16162),.A(g5597),.B(g13234));
  AND2 AND2_1296(.VSS(VSS),.VDD(VDD),.Y(g16163),.A(g5736),.B(g11841));
  AND2 AND2_1297(.VSS(VSS),.VDD(VDD),.Y(g16170),.A(g3616),.B(g11842));
  AND2 AND2_1298(.VSS(VSS),.VDD(VDD),.Y(g16178),.A(g2372),.B(g11846));
  AND2 AND2_1299(.VSS(VSS),.VDD(VDD),.Y(g16182),.A(g7149),.B(g11852));
  AND2 AND2_1300(.VSS(VSS),.VDD(VDD),.Y(g16183),.A(g12235),.B(g11014));
  AND2 AND2_1301(.VSS(VSS),.VDD(VDD),.Y(g16184),.A(g5663),.B(g11853));
  AND2 AND2_1302(.VSS(VSS),.VDD(VDD),.Y(g16185),.A(g12308),.B(g11017));
  AND2 AND2_1303(.VSS(VSS),.VDD(VDD),.Y(g16186),.A(g5753),.B(g11856));
  AND2 AND2_1304(.VSS(VSS),.VDD(VDD),.Y(g16187),.A(g5754),.B(g11857));
  AND2 AND2_1305(.VSS(VSS),.VDD(VDD),.Y(g16188),.A(g5755),.B(g11858));
  AND2 AND2_1306(.VSS(VSS),.VDD(VDD),.Y(g16197),.A(g518),.B(g11862));
  AND2 AND2_1307(.VSS(VSS),.VDD(VDD),.Y(g16198),.A(g5762),.B(g11866));
  AND2 AND2_1308(.VSS(VSS),.VDD(VDD),.Y(g16199),.A(g5763),.B(g11867));
  AND2 AND2_1309(.VSS(VSS),.VDD(VDD),.Y(g16200),.A(g5764),.B(g11868));
  AND2 AND2_1310(.VSS(VSS),.VDD(VDD),.Y(g16211),.A(g1203),.B(g11871));
  AND2 AND2_1311(.VSS(VSS),.VDD(VDD),.Y(g16212),.A(g5609),.B(g13252));
  AND2 AND2_1312(.VSS(VSS),.VDD(VDD),.Y(g16217),.A(g5776),.B(g11876));
  AND2 AND2_1313(.VSS(VSS),.VDD(VDD),.Y(g16218),.A(g5777),.B(g11877));
  AND2 AND2_1314(.VSS(VSS),.VDD(VDD),.Y(g16219),.A(g8295),.B(g11878));
  AND2 AND2_1315(.VSS(VSS),.VDD(VDD),.Y(g16220),.A(g1896),.B(g11879));
  AND2 AND2_1316(.VSS(VSS),.VDD(VDD),.Y(g16221),.A(g5614),.B(g13257));
  AND2 AND2_1317(.VSS(VSS),.VDD(VDD),.Y(g16222),.A(g5794),.B(g11883));
  AND2 AND2_1318(.VSS(VSS),.VDD(VDD),.Y(g16229),.A(g3772),.B(g11884));
  AND2 AND2_1319(.VSS(VSS),.VDD(VDD),.Y(g16237),.A(g5379),.B(g11886));
  AND2 AND2_1320(.VSS(VSS),.VDD(VDD),.Y(g16238),.A(g12275),.B(g11066));
  AND2 AND2_1321(.VSS(VSS),.VDD(VDD),.Y(g16239),.A(g5700),.B(g11887));
  AND2 AND2_1322(.VSS(VSS),.VDD(VDD),.Y(g16240),.A(g5804),.B(g11891));
  AND2 AND2_1323(.VSS(VSS),.VDD(VDD),.Y(g16241),.A(g5805),.B(g11892));
  AND2 AND2_1324(.VSS(VSS),.VDD(VDD),.Y(g16242),.A(g5806),.B(g11893));
  AND2 AND2_1325(.VSS(VSS),.VDD(VDD),.Y(g16250),.A(g519),.B(g11895));
  AND2 AND2_1326(.VSS(VSS),.VDD(VDD),.Y(g16251),.A(g5812),.B(g11898));
  AND2 AND2_1327(.VSS(VSS),.VDD(VDD),.Y(g16252),.A(g5813),.B(g11899));
  AND2 AND2_1328(.VSS(VSS),.VDD(VDD),.Y(g16253),.A(g5814),.B(g11900));
  AND2 AND2_1329(.VSS(VSS),.VDD(VDD),.Y(g16262),.A(g1204),.B(g11904));
  AND2 AND2_1330(.VSS(VSS),.VDD(VDD),.Y(g16263),.A(g5821),.B(g11908));
  AND2 AND2_1331(.VSS(VSS),.VDD(VDD),.Y(g16264),.A(g5822),.B(g11909));
  AND2 AND2_1332(.VSS(VSS),.VDD(VDD),.Y(g16265),.A(g5823),.B(g11910));
  AND2 AND2_1333(.VSS(VSS),.VDD(VDD),.Y(g16276),.A(g1897),.B(g11913));
  AND2 AND2_1334(.VSS(VSS),.VDD(VDD),.Y(g16277),.A(g5634),.B(g13275));
  AND2 AND2_1335(.VSS(VSS),.VDD(VDD),.Y(g16282),.A(g5835),.B(g11918));
  AND2 AND2_1336(.VSS(VSS),.VDD(VDD),.Y(g16283),.A(g5836),.B(g11919));
  AND2 AND2_1337(.VSS(VSS),.VDD(VDD),.Y(g16284),.A(g8304),.B(g11920));
  AND2 AND2_1338(.VSS(VSS),.VDD(VDD),.Y(g16285),.A(g2590),.B(g11921));
  AND2 AND2_1339(.VSS(VSS),.VDD(VDD),.Y(g16286),.A(g5639),.B(g13280));
  AND2 AND2_1340(.VSS(VSS),.VDD(VDD),.Y(g16288),.A(g12308),.B(g11129));
  AND2 AND2_1341(.VSS(VSS),.VDD(VDD),.Y(g16289),.A(g5853),.B(g11929));
  AND2 AND2_1342(.VSS(VSS),.VDD(VDD),.Y(g16290),.A(g5854),.B(g11930));
  AND2 AND2_1343(.VSS(VSS),.VDD(VDD),.Y(g16291),.A(g5855),.B(g11931));
  AND2 AND2_1344(.VSS(VSS),.VDD(VDD),.Y(g16292),.A(g294),.B(g11932));
  AND2 AND2_1345(.VSS(VSS),.VDD(VDD),.Y(g16298),.A(g520),.B(g11936));
  AND2 AND2_1346(.VSS(VSS),.VDD(VDD),.Y(g16299),.A(g5860),.B(g11941));
  AND2 AND2_1347(.VSS(VSS),.VDD(VDD),.Y(g16300),.A(g5861),.B(g11942));
  AND2 AND2_1348(.VSS(VSS),.VDD(VDD),.Y(g16301),.A(g5862),.B(g11943));
  AND2 AND2_1349(.VSS(VSS),.VDD(VDD),.Y(g16309),.A(g1205),.B(g11945));
  AND2 AND2_1350(.VSS(VSS),.VDD(VDD),.Y(g16310),.A(g5868),.B(g11948));
  AND2 AND2_1351(.VSS(VSS),.VDD(VDD),.Y(g16311),.A(g5869),.B(g11949));
  AND2 AND2_1352(.VSS(VSS),.VDD(VDD),.Y(g16312),.A(g5870),.B(g11950));
  AND2 AND2_1353(.VSS(VSS),.VDD(VDD),.Y(g16321),.A(g1898),.B(g11954));
  AND2 AND2_1354(.VSS(VSS),.VDD(VDD),.Y(g16322),.A(g5877),.B(g11958));
  AND2 AND2_1355(.VSS(VSS),.VDD(VDD),.Y(g16323),.A(g5878),.B(g11959));
  AND2 AND2_1356(.VSS(VSS),.VDD(VDD),.Y(g16324),.A(g5879),.B(g11960));
  AND2 AND2_1357(.VSS(VSS),.VDD(VDD),.Y(g16335),.A(g2591),.B(g11963));
  AND2 AND2_1358(.VSS(VSS),.VDD(VDD),.Y(g16336),.A(g5662),.B(g13300));
  AND2 AND2_1359(.VSS(VSS),.VDD(VDD),.Y(g16342),.A(g5894),.B(g11968));
  AND2 AND2_1360(.VSS(VSS),.VDD(VDD),.Y(g16343),.A(g5895),.B(g11969));
  AND2 AND2_1361(.VSS(VSS),.VDD(VDD),.Y(g16344),.A(g5896),.B(g11970));
  AND2 AND2_1362(.VSS(VSS),.VDD(VDD),.Y(g16345),.A(g5897),.B(g11971));
  AND2 AND2_1363(.VSS(VSS),.VDD(VDD),.Y(g16346),.A(g295),.B(g11972));
  AND2 AND2_1364(.VSS(VSS),.VDD(VDD),.Y(g16347),.A(g5900),.B(g11982));
  AND2 AND2_1365(.VSS(VSS),.VDD(VDD),.Y(g16348),.A(g5901),.B(g11983));
  AND2 AND2_1366(.VSS(VSS),.VDD(VDD),.Y(g16349),.A(g5902),.B(g11984));
  AND2 AND2_1367(.VSS(VSS),.VDD(VDD),.Y(g16350),.A(g981),.B(g11985));
  AND2 AND2_1368(.VSS(VSS),.VDD(VDD),.Y(g16356),.A(g1206),.B(g11989));
  AND2 AND2_1369(.VSS(VSS),.VDD(VDD),.Y(g16357),.A(g5907),.B(g11994));
  AND2 AND2_1370(.VSS(VSS),.VDD(VDD),.Y(g16358),.A(g5908),.B(g11995));
  AND2 AND2_1371(.VSS(VSS),.VDD(VDD),.Y(g16359),.A(g5909),.B(g11996));
  AND2 AND2_1372(.VSS(VSS),.VDD(VDD),.Y(g16367),.A(g1899),.B(g11998));
  AND2 AND2_1373(.VSS(VSS),.VDD(VDD),.Y(g16368),.A(g5915),.B(g12001));
  AND2 AND2_1374(.VSS(VSS),.VDD(VDD),.Y(g16369),.A(g5916),.B(g12002));
  AND2 AND2_1375(.VSS(VSS),.VDD(VDD),.Y(g16370),.A(g5917),.B(g12003));
  AND2 AND2_1376(.VSS(VSS),.VDD(VDD),.Y(g16379),.A(g2592),.B(g12007));
  AND2 AND2_1377(.VSS(VSS),.VDD(VDD),.Y(g16380),.A(g5925),.B(g12020));
  AND2 AND2_1378(.VSS(VSS),.VDD(VDD),.Y(g16381),.A(g5926),.B(g12021));
  AND2 AND2_1379(.VSS(VSS),.VDD(VDD),.Y(g16382),.A(g5927),.B(g12022));
  AND2 AND2_1380(.VSS(VSS),.VDD(VDD),.Y(g16383),.A(g5928),.B(g12023));
  AND2 AND2_1381(.VSS(VSS),.VDD(VDD),.Y(g16384),.A(g296),.B(g12024));
  AND2 AND2_1382(.VSS(VSS),.VDD(VDD),.Y(g16385),.A(g5714),.B(g13336));
  AND2 AND2_1383(.VSS(VSS),.VDD(VDD),.Y(g16386),.A(g5933),.B(g12037));
  AND2 AND2_1384(.VSS(VSS),.VDD(VDD),.Y(g16387),.A(g5934),.B(g12038));
  AND2 AND2_1385(.VSS(VSS),.VDD(VDD),.Y(g16388),.A(g5935),.B(g12039));
  AND2 AND2_1386(.VSS(VSS),.VDD(VDD),.Y(g16389),.A(g5936),.B(g12040));
  AND2 AND2_1387(.VSS(VSS),.VDD(VDD),.Y(g16390),.A(g982),.B(g12041));
  AND2 AND2_1388(.VSS(VSS),.VDD(VDD),.Y(g16391),.A(g5939),.B(g12051));
  AND2 AND2_1389(.VSS(VSS),.VDD(VDD),.Y(g16392),.A(g5940),.B(g12052));
  AND2 AND2_1390(.VSS(VSS),.VDD(VDD),.Y(g16393),.A(g5941),.B(g12053));
  AND2 AND2_1391(.VSS(VSS),.VDD(VDD),.Y(g16394),.A(g1675),.B(g12054));
  AND2 AND2_1392(.VSS(VSS),.VDD(VDD),.Y(g16400),.A(g1900),.B(g12058));
  AND2 AND2_1393(.VSS(VSS),.VDD(VDD),.Y(g16401),.A(g5946),.B(g12063));
  AND2 AND2_1394(.VSS(VSS),.VDD(VDD),.Y(g16402),.A(g5947),.B(g12064));
  AND2 AND2_1395(.VSS(VSS),.VDD(VDD),.Y(g16403),.A(g5948),.B(g12065));
  AND2 AND2_1396(.VSS(VSS),.VDD(VDD),.Y(g16411),.A(g2593),.B(g12067));
  AND2 AND2_1397(.VSS(VSS),.VDD(VDD),.Y(g16413),.A(g5954),.B(g12075));
  AND2 AND2_1398(.VSS(VSS),.VDD(VDD),.Y(g16414),.A(g5955),.B(g12076));
  AND2 AND2_1399(.VSS(VSS),.VDD(VDD),.Y(g16415),.A(g5956),.B(g12077));
  AND2 AND2_1400(.VSS(VSS),.VDD(VDD),.Y(g16416),.A(g5957),.B(g12078));
  AND2 AND2_1401(.VSS(VSS),.VDD(VDD),.Y(g16417),.A(g5759),.B(g13356));
  AND2 AND2_1402(.VSS(VSS),.VDD(VDD),.Y(g16418),.A(g5959),.B(g12084));
  AND2 AND2_1403(.VSS(VSS),.VDD(VDD),.Y(g16419),.A(g5960),.B(g12085));
  AND2 AND2_1404(.VSS(VSS),.VDD(VDD),.Y(g16420),.A(g5961),.B(g12086));
  AND2 AND2_1405(.VSS(VSS),.VDD(VDD),.Y(g16421),.A(g5962),.B(g12087));
  AND2 AND2_1406(.VSS(VSS),.VDD(VDD),.Y(g16422),.A(g983),.B(g12088));
  AND2 AND2_1407(.VSS(VSS),.VDD(VDD),.Y(g16423),.A(g5772),.B(g13361));
  AND2 AND2_1408(.VSS(VSS),.VDD(VDD),.Y(g16424),.A(g5967),.B(g12101));
  AND2 AND2_1409(.VSS(VSS),.VDD(VDD),.Y(g16425),.A(g5968),.B(g12102));
  AND2 AND2_1410(.VSS(VSS),.VDD(VDD),.Y(g16426),.A(g5969),.B(g12103));
  AND2 AND2_1411(.VSS(VSS),.VDD(VDD),.Y(g16427),.A(g5970),.B(g12104));
  AND2 AND2_1412(.VSS(VSS),.VDD(VDD),.Y(g16428),.A(g1676),.B(g12105));
  AND2 AND2_1413(.VSS(VSS),.VDD(VDD),.Y(g16429),.A(g5973),.B(g12115));
  AND2 AND2_1414(.VSS(VSS),.VDD(VDD),.Y(g16430),.A(g5974),.B(g12116));
  AND2 AND2_1415(.VSS(VSS),.VDD(VDD),.Y(g16431),.A(g5975),.B(g12117));
  AND2 AND2_1416(.VSS(VSS),.VDD(VDD),.Y(g16432),.A(g2369),.B(g12118));
  AND2 AND2_1417(.VSS(VSS),.VDD(VDD),.Y(g16438),.A(g2594),.B(g12122));
  AND2 AND2_1418(.VSS(VSS),.VDD(VDD),.Y(g16443),.A(g5980),.B(g12134));
  AND2 AND2_1419(.VSS(VSS),.VDD(VDD),.Y(g16444),.A(g5981),.B(g12135));
  AND2 AND2_1420(.VSS(VSS),.VDD(VDD),.Y(g16445),.A(g5808),.B(g13381));
  AND2 AND2_1421(.VSS(VSS),.VDD(VDD),.Y(g16447),.A(g5983),.B(g12147));
  AND2 AND2_1422(.VSS(VSS),.VDD(VDD),.Y(g16448),.A(g5984),.B(g12148));
  AND2 AND2_1423(.VSS(VSS),.VDD(VDD),.Y(g16449),.A(g5985),.B(g12149));
  AND2 AND2_1424(.VSS(VSS),.VDD(VDD),.Y(g16450),.A(g5986),.B(g12150));
  AND2 AND2_1425(.VSS(VSS),.VDD(VDD),.Y(g16451),.A(g5818),.B(g13386));
  AND2 AND2_1426(.VSS(VSS),.VDD(VDD),.Y(g16452),.A(g5988),.B(g12156));
  AND2 AND2_1427(.VSS(VSS),.VDD(VDD),.Y(g16453),.A(g5989),.B(g12157));
  AND2 AND2_1428(.VSS(VSS),.VDD(VDD),.Y(g16454),.A(g5990),.B(g12158));
  AND2 AND2_1429(.VSS(VSS),.VDD(VDD),.Y(g16455),.A(g5991),.B(g12159));
  AND2 AND2_1430(.VSS(VSS),.VDD(VDD),.Y(g16456),.A(g1677),.B(g12160));
  AND2 AND2_1431(.VSS(VSS),.VDD(VDD),.Y(g16457),.A(g5831),.B(g13391));
  AND2 AND2_1432(.VSS(VSS),.VDD(VDD),.Y(g16458),.A(g5996),.B(g12173));
  AND2 AND2_1433(.VSS(VSS),.VDD(VDD),.Y(g16459),.A(g5997),.B(g12174));
  AND2 AND2_1434(.VSS(VSS),.VDD(VDD),.Y(g16460),.A(g5998),.B(g12175));
  AND2 AND2_1435(.VSS(VSS),.VDD(VDD),.Y(g16461),.A(g5999),.B(g12176));
  AND2 AND2_1436(.VSS(VSS),.VDD(VDD),.Y(g16462),.A(g2370),.B(g12177));
  AND4 AND4_22(.VSS(VSS),.VDD(VDD),.Y(g16505),.A(g14776),.B(g14797),.C(g16142),.D(g16243));
  AND4 AND4_23(.VSS(VSS),.VDD(VDD),.Y(g16513),.A(g15065),.B(g13724),.C(g13764),.D(g13797));
  AND4 AND4_24(.VSS(VSS),.VDD(VDD),.Y(g16527),.A(g14811),.B(g14849),.C(g16201),.D(g16302));
  AND4 AND4_25(.VSS(VSS),.VDD(VDD),.Y(g16535),.A(g15161),.B(g13774),.C(g13805),.D(g13825));
  AND4 AND4_26(.VSS(VSS),.VDD(VDD),.Y(g16558),.A(g14863),.B(g14922),.C(g16266),.D(g16360));
  AND4 AND4_27(.VSS(VSS),.VDD(VDD),.Y(g16590),.A(g14936),.B(g15003),.C(g16325),.D(g16404));
  AND2 AND2_1437(.VSS(VSS),.VDD(VDD),.Y(g16607),.A(g15022),.B(g15096));
  AND2 AND2_1438(.VSS(VSS),.VDD(VDD),.Y(g16625),.A(g15118),.B(g15188));
  AND2 AND2_1439(.VSS(VSS),.VDD(VDD),.Y(g16639),.A(g15210),.B(g15274));
  AND2 AND2_1440(.VSS(VSS),.VDD(VDD),.Y(g16650),.A(g15296),.B(g15366));
  AND2 AND2_1441(.VSS(VSS),.VDD(VDD),.Y(g16850),.A(g6226),.B(g14764));
  AND2 AND2_1442(.VSS(VSS),.VDD(VDD),.Y(g16855),.A(g15722),.B(g8646));
  AND2 AND2_1443(.VSS(VSS),.VDD(VDD),.Y(g16856),.A(g6443),.B(g14794));
  AND2 AND2_1444(.VSS(VSS),.VDD(VDD),.Y(g16859),.A(g15762),.B(g8662));
  AND2 AND2_1445(.VSS(VSS),.VDD(VDD),.Y(g16864),.A(g15790),.B(g8681));
  AND2 AND2_1446(.VSS(VSS),.VDD(VDD),.Y(g16865),.A(g6896),.B(g14881));
  AND2 AND2_1447(.VSS(VSS),.VDD(VDD),.Y(g16879),.A(g15813),.B(g8693));
  AND2 AND2_1448(.VSS(VSS),.VDD(VDD),.Y(g16894),.A(g7156),.B(g14959));
  AND2 AND2_1449(.VSS(VSS),.VDD(VDD),.Y(g16907),.A(g7335),.B(g15017));
  AND2 AND2_1450(.VSS(VSS),.VDD(VDD),.Y(g16908),.A(g7838),.B(g15032));
  AND2 AND2_1451(.VSS(VSS),.VDD(VDD),.Y(g16909),.A(g6908),.B(g15033));
  AND2 AND2_1452(.VSS(VSS),.VDD(VDD),.Y(g16923),.A(g7352),.B(g15048));
  AND2 AND2_1453(.VSS(VSS),.VDD(VDD),.Y(g16938),.A(g7858),.B(g15128));
  AND2 AND2_1454(.VSS(VSS),.VDD(VDD),.Y(g16939),.A(g7158),.B(g15129));
  AND2 AND2_1455(.VSS(VSS),.VDD(VDD),.Y(g16953),.A(g7482),.B(g15144));
  AND2 AND2_1456(.VSS(VSS),.VDD(VDD),.Y(g16964),.A(g7520),.B(g15170));
  AND2 AND2_1457(.VSS(VSS),.VDD(VDD),.Y(g16966),.A(g7529),.B(g15174));
  AND2 AND2_1458(.VSS(VSS),.VDD(VDD),.Y(g16967),.A(g7827),.B(g15175));
  AND2 AND2_1459(.VSS(VSS),.VDD(VDD),.Y(g16968),.A(g6672),.B(g15176));
  AND2 AND2_1460(.VSS(VSS),.VDD(VDD),.Y(g16969),.A(g7888),.B(g15220));
  AND2 AND2_1461(.VSS(VSS),.VDD(VDD),.Y(g16970),.A(g7354),.B(g15221));
  AND2 AND2_1462(.VSS(VSS),.VDD(VDD),.Y(g16984),.A(g7538),.B(g15236));
  AND2 AND2_1463(.VSS(VSS),.VDD(VDD),.Y(g16987),.A(g7555),.B(g15260));
  AND2 AND2_1464(.VSS(VSS),.VDD(VDD),.Y(g16988),.A(g7842),.B(g15261));
  AND2 AND2_1465(.VSS(VSS),.VDD(VDD),.Y(g16989),.A(g6974),.B(g15262));
  AND2 AND2_1466(.VSS(VSS),.VDD(VDD),.Y(g16990),.A(g7912),.B(g15306));
  AND2 AND2_1467(.VSS(VSS),.VDD(VDD),.Y(g16991),.A(g7484),.B(g15307));
  AND2 AND2_1468(.VSS(VSS),.VDD(VDD),.Y(g16993),.A(g7576),.B(g15322));
  AND2 AND2_1469(.VSS(VSS),.VDD(VDD),.Y(g16994),.A(g7819),.B(g15323));
  AND2 AND2_1470(.VSS(VSS),.VDD(VDD),.Y(g16997),.A(g7578),.B(g15352));
  AND2 AND2_1471(.VSS(VSS),.VDD(VDD),.Y(g16998),.A(g7862),.B(g15353));
  AND2 AND2_1472(.VSS(VSS),.VDD(VDD),.Y(g16999),.A(g7224),.B(g15354));
  AND3 AND3_14(.VSS(VSS),.VDD(VDD),.Y(g17001),.A(g3254),.B(g10694),.C(g14144));
  AND2 AND2_1473(.VSS(VSS),.VDD(VDD),.Y(g17015),.A(g7996),.B(g15390));
  AND2 AND2_1474(.VSS(VSS),.VDD(VDD),.Y(g17017),.A(g7590),.B(g15408));
  AND2 AND2_1475(.VSS(VSS),.VDD(VDD),.Y(g17018),.A(g7830),.B(g15409));
  AND2 AND2_1476(.VSS(VSS),.VDD(VDD),.Y(g17021),.A(g7592),.B(g15438));
  AND2 AND2_1477(.VSS(VSS),.VDD(VDD),.Y(g17022),.A(g7892),.B(g15439));
  AND2 AND2_1478(.VSS(VSS),.VDD(VDD),.Y(g17023),.A(g7420),.B(g15440));
  AND2 AND2_1479(.VSS(VSS),.VDD(VDD),.Y(g17028),.A(g7604),.B(g15458));
  AND3 AND3_15(.VSS(VSS),.VDD(VDD),.Y(g17031),.A(g3410),.B(g10714),.C(g14259));
  AND2 AND2_1480(.VSS(VSS),.VDD(VDD),.Y(g17045),.A(g8071),.B(g15474));
  AND2 AND2_1481(.VSS(VSS),.VDD(VDD),.Y(g17047),.A(g7605),.B(g15492));
  AND2 AND2_1482(.VSS(VSS),.VDD(VDD),.Y(g17048),.A(g7845),.B(g15493));
  AND2 AND2_1483(.VSS(VSS),.VDD(VDD),.Y(g17055),.A(g7153),.B(g15524));
  AND2 AND2_1484(.VSS(VSS),.VDD(VDD),.Y(g17056),.A(g7953),.B(g15525));
  AND2 AND2_1485(.VSS(VSS),.VDD(VDD),.Y(g17062),.A(g7613),.B(g15544));
  AND3 AND3_16(.VSS(VSS),.VDD(VDD),.Y(g17065),.A(g3566),.B(g10735),.C(g14381));
  AND2 AND2_1486(.VSS(VSS),.VDD(VDD),.Y(g17079),.A(g8156),.B(g15560));
  AND2 AND2_1487(.VSS(VSS),.VDD(VDD),.Y(g17081),.A(g7614),.B(g15578));
  AND2 AND2_1488(.VSS(VSS),.VDD(VDD),.Y(g17082),.A(g7865),.B(g15579));
  AND2 AND2_1489(.VSS(VSS),.VDD(VDD),.Y(g17084),.A(g7629),.B(g13954));
  AND2 AND2_1490(.VSS(VSS),.VDD(VDD),.Y(g17090),.A(g7349),.B(g15602));
  AND2 AND2_1491(.VSS(VSS),.VDD(VDD),.Y(g17091),.A(g8004),.B(g15603));
  AND2 AND2_1492(.VSS(VSS),.VDD(VDD),.Y(g17097),.A(g7622),.B(g15622));
  AND3 AND3_17(.VSS(VSS),.VDD(VDD),.Y(g17100),.A(g3722),.B(g10754),.C(g14493));
  AND2 AND2_1493(.VSS(VSS),.VDD(VDD),.Y(g17114),.A(g8242),.B(g15638));
  AND2 AND2_1494(.VSS(VSS),.VDD(VDD),.Y(g17116),.A(g7649),.B(g14008));
  AND2 AND2_1495(.VSS(VSS),.VDD(VDD),.Y(g17117),.A(g7906),.B(g15665));
  AND2 AND2_1496(.VSS(VSS),.VDD(VDD),.Y(g17122),.A(g7658),.B(g14024));
  AND2 AND2_1497(.VSS(VSS),.VDD(VDD),.Y(g17128),.A(g7479),.B(g15678));
  AND2 AND2_1498(.VSS(VSS),.VDD(VDD),.Y(g17129),.A(g8079),.B(g15679));
  AND2 AND2_1499(.VSS(VSS),.VDD(VDD),.Y(g17135),.A(g7638),.B(g15698));
  AND2 AND2_1500(.VSS(VSS),.VDD(VDD),.Y(g17138),.A(g7676),.B(g14068));
  AND2 AND2_1501(.VSS(VSS),.VDD(VDD),.Y(g17143),.A(g7685),.B(g14099));
  AND2 AND2_1502(.VSS(VSS),.VDD(VDD),.Y(g17144),.A(g7958),.B(g15724));
  AND2 AND2_1503(.VSS(VSS),.VDD(VDD),.Y(g17149),.A(g7694),.B(g14115));
  AND2 AND2_1504(.VSS(VSS),.VDD(VDD),.Y(g17155),.A(g7535),.B(g15737));
  AND2 AND2_1505(.VSS(VSS),.VDD(VDD),.Y(g17156),.A(g8164),.B(g15738));
  AND2 AND2_1506(.VSS(VSS),.VDD(VDD),.Y(g17161),.A(g7712),.B(g14183));
  AND2 AND2_1507(.VSS(VSS),.VDD(VDD),.Y(g17166),.A(g7721),.B(g14214));
  AND2 AND2_1508(.VSS(VSS),.VDD(VDD),.Y(g17167),.A(g8009),.B(g15764));
  AND2 AND2_1509(.VSS(VSS),.VDD(VDD),.Y(g17172),.A(g7730),.B(g14230));
  AND2 AND2_1510(.VSS(VSS),.VDD(VDD),.Y(g17176),.A(g7742),.B(g14298));
  AND2 AND2_1511(.VSS(VSS),.VDD(VDD),.Y(g17181),.A(g7751),.B(g14329));
  AND2 AND2_1512(.VSS(VSS),.VDD(VDD),.Y(g17182),.A(g8084),.B(g15792));
  AND2 AND2_1513(.VSS(VSS),.VDD(VDD),.Y(g17193),.A(g7766),.B(g14420));
  AND2 AND2_1514(.VSS(VSS),.VDD(VDD),.Y(g17268),.A(g8024),.B(g15991));
  AND2 AND2_1515(.VSS(VSS),.VDD(VDD),.Y(g17301),.A(g8097),.B(g15994));
  AND2 AND2_1516(.VSS(VSS),.VDD(VDD),.Y(g17339),.A(g8176),.B(g15997));
  AND2 AND2_1517(.VSS(VSS),.VDD(VDD),.Y(g17352),.A(g3942),.B(g14960));
  AND2 AND2_1518(.VSS(VSS),.VDD(VDD),.Y(g17353),.A(g3945),.B(g14963));
  AND2 AND2_1519(.VSS(VSS),.VDD(VDD),.Y(g17381),.A(g8250),.B(g16001));
  AND2 AND2_1520(.VSS(VSS),.VDD(VDD),.Y(g17382),.A(g8252),.B(g16002));
  AND2 AND2_1521(.VSS(VSS),.VDD(VDD),.Y(g17393),.A(g3941),.B(g16005));
  AND2 AND2_1522(.VSS(VSS),.VDD(VDD),.Y(g17395),.A(g6177),.B(g15034));
  AND2 AND2_1523(.VSS(VSS),.VDD(VDD),.Y(g17396),.A(g4020),.B(g15037));
  AND2 AND2_1524(.VSS(VSS),.VDD(VDD),.Y(g17397),.A(g4023),.B(g15040));
  AND2 AND2_1525(.VSS(VSS),.VDD(VDD),.Y(g17398),.A(g4026),.B(g15043));
  AND2 AND2_1526(.VSS(VSS),.VDD(VDD),.Y(g17408),.A(g4049),.B(g15049));
  AND2 AND2_1527(.VSS(VSS),.VDD(VDD),.Y(g17409),.A(g4052),.B(g15052));
  AND2 AND2_1528(.VSS(VSS),.VDD(VDD),.Y(g17428),.A(g3994),.B(g16007));
  AND2 AND2_1529(.VSS(VSS),.VDD(VDD),.Y(g17446),.A(g6284),.B(g16011));
  AND2 AND2_1530(.VSS(VSS),.VDD(VDD),.Y(g17447),.A(g4115),.B(g15106));
  AND2 AND2_1531(.VSS(VSS),.VDD(VDD),.Y(g17448),.A(g4118),.B(g15109));
  AND2 AND2_1532(.VSS(VSS),.VDD(VDD),.Y(g17449),.A(g4121),.B(g15112));
  AND2 AND2_1533(.VSS(VSS),.VDD(VDD),.Y(g17450),.A(g4124),.B(g15115));
  AND2 AND2_1534(.VSS(VSS),.VDD(VDD),.Y(g17460),.A(g4048),.B(g16012));
  AND2 AND2_1535(.VSS(VSS),.VDD(VDD),.Y(g17461),.A(g6209),.B(g15130));
  AND2 AND2_1536(.VSS(VSS),.VDD(VDD),.Y(g17462),.A(g4147),.B(g15133));
  AND2 AND2_1537(.VSS(VSS),.VDD(VDD),.Y(g17463),.A(g4150),.B(g15136));
  AND2 AND2_1538(.VSS(VSS),.VDD(VDD),.Y(g17464),.A(g4153),.B(g15139));
  AND2 AND2_1539(.VSS(VSS),.VDD(VDD),.Y(g17474),.A(g4176),.B(g15145));
  AND2 AND2_1540(.VSS(VSS),.VDD(VDD),.Y(g17475),.A(g4179),.B(g15148));
  AND2 AND2_1541(.VSS(VSS),.VDD(VDD),.Y(g17485),.A(g4089),.B(g16013));
  AND2 AND2_1542(.VSS(VSS),.VDD(VDD),.Y(g17486),.A(g4091),.B(g16014));
  AND2 AND2_1543(.VSS(VSS),.VDD(VDD),.Y(g17506),.A(g6675),.B(g16023));
  AND2 AND2_1544(.VSS(VSS),.VDD(VDD),.Y(g17508),.A(g4225),.B(g15179));
  AND2 AND2_1545(.VSS(VSS),.VDD(VDD),.Y(g17509),.A(g4228),.B(g15182));
  AND2 AND2_1546(.VSS(VSS),.VDD(VDD),.Y(g17510),.A(g4231),.B(g15185));
  AND2 AND2_1547(.VSS(VSS),.VDD(VDD),.Y(g17526),.A(g6421),.B(g16025));
  AND2 AND2_1548(.VSS(VSS),.VDD(VDD),.Y(g17527),.A(g4254),.B(g15198));
  AND2 AND2_1549(.VSS(VSS),.VDD(VDD),.Y(g17528),.A(g4257),.B(g15201));
  AND2 AND2_1550(.VSS(VSS),.VDD(VDD),.Y(g17529),.A(g4260),.B(g15204));
  AND2 AND2_1551(.VSS(VSS),.VDD(VDD),.Y(g17530),.A(g4263),.B(g15207));
  AND2 AND2_1552(.VSS(VSS),.VDD(VDD),.Y(g17540),.A(g4175),.B(g16026));
  AND2 AND2_1553(.VSS(VSS),.VDD(VDD),.Y(g17541),.A(g6298),.B(g15222));
  AND2 AND2_1554(.VSS(VSS),.VDD(VDD),.Y(g17542),.A(g4286),.B(g15225));
  AND2 AND2_1555(.VSS(VSS),.VDD(VDD),.Y(g17543),.A(g4289),.B(g15228));
  AND2 AND2_1556(.VSS(VSS),.VDD(VDD),.Y(g17544),.A(g4292),.B(g15231));
  AND2 AND2_1557(.VSS(VSS),.VDD(VDD),.Y(g17554),.A(g4315),.B(g15237));
  AND2 AND2_1558(.VSS(VSS),.VDD(VDD),.Y(g17555),.A(g4318),.B(g15240));
  AND2 AND2_1559(.VSS(VSS),.VDD(VDD),.Y(g17556),.A(g4201),.B(g16027));
  AND2 AND2_1560(.VSS(VSS),.VDD(VDD),.Y(g17576),.A(g4348),.B(g15248));
  AND2 AND2_1561(.VSS(VSS),.VDD(VDD),.Y(g17577),.A(g4351),.B(g15251));
  AND2 AND2_1562(.VSS(VSS),.VDD(VDD),.Y(g17578),.A(g4354),.B(g15254));
  AND2 AND2_1563(.VSS(VSS),.VDD(VDD),.Y(g17597),.A(g6977),.B(g16039));
  AND2 AND2_1564(.VSS(VSS),.VDD(VDD),.Y(g17598),.A(g4380),.B(g15265));
  AND2 AND2_1565(.VSS(VSS),.VDD(VDD),.Y(g17599),.A(g4383),.B(g15268));
  AND2 AND2_1566(.VSS(VSS),.VDD(VDD),.Y(g17600),.A(g4386),.B(g15271));
  AND2 AND2_1567(.VSS(VSS),.VDD(VDD),.Y(g17616),.A(g6626),.B(g16041));
  AND2 AND2_1568(.VSS(VSS),.VDD(VDD),.Y(g17617),.A(g4409),.B(g15284));
  AND2 AND2_1569(.VSS(VSS),.VDD(VDD),.Y(g17618),.A(g4412),.B(g15287));
  AND2 AND2_1570(.VSS(VSS),.VDD(VDD),.Y(g17619),.A(g4415),.B(g15290));
  AND2 AND2_1571(.VSS(VSS),.VDD(VDD),.Y(g17620),.A(g4418),.B(g15293));
  AND2 AND2_1572(.VSS(VSS),.VDD(VDD),.Y(g17630),.A(g4314),.B(g16042));
  AND2 AND2_1573(.VSS(VSS),.VDD(VDD),.Y(g17631),.A(g6435),.B(g15308));
  AND2 AND2_1574(.VSS(VSS),.VDD(VDD),.Y(g17632),.A(g4441),.B(g15311));
  AND2 AND2_1575(.VSS(VSS),.VDD(VDD),.Y(g17633),.A(g4444),.B(g15314));
  AND2 AND2_1576(.VSS(VSS),.VDD(VDD),.Y(g17634),.A(g4447),.B(g15317));
  AND2 AND2_1577(.VSS(VSS),.VDD(VDD),.Y(g17635),.A(g4322),.B(g16043));
  AND2 AND2_1578(.VSS(VSS),.VDD(VDD),.Y(g17636),.A(g4324),.B(g16044));
  AND2 AND2_1579(.VSS(VSS),.VDD(VDD),.Y(g17652),.A(g4480),.B(g15326));
  AND2 AND2_1580(.VSS(VSS),.VDD(VDD),.Y(g17653),.A(g4483),.B(g15329));
  AND2 AND2_1581(.VSS(VSS),.VDD(VDD),.Y(g17654),.A(g4486),.B(g15332));
  AND2 AND2_1582(.VSS(VSS),.VDD(VDD),.Y(g17673),.A(g4517),.B(g15340));
  AND2 AND2_1583(.VSS(VSS),.VDD(VDD),.Y(g17674),.A(g4520),.B(g15343));
  AND2 AND2_1584(.VSS(VSS),.VDD(VDD),.Y(g17675),.A(g4523),.B(g15346));
  AND2 AND2_1585(.VSS(VSS),.VDD(VDD),.Y(g17694),.A(g7227),.B(g16061));
  AND2 AND2_1586(.VSS(VSS),.VDD(VDD),.Y(g17695),.A(g4549),.B(g15357));
  AND2 AND2_1587(.VSS(VSS),.VDD(VDD),.Y(g17696),.A(g4552),.B(g15360));
  AND2 AND2_1588(.VSS(VSS),.VDD(VDD),.Y(g17697),.A(g4555),.B(g15363));
  AND2 AND2_1589(.VSS(VSS),.VDD(VDD),.Y(g17713),.A(g6890),.B(g16063));
  AND2 AND2_1590(.VSS(VSS),.VDD(VDD),.Y(g17714),.A(g4578),.B(g15376));
  AND2 AND2_1591(.VSS(VSS),.VDD(VDD),.Y(g17715),.A(g4581),.B(g15379));
  AND2 AND2_1592(.VSS(VSS),.VDD(VDD),.Y(g17716),.A(g4584),.B(g15382));
  AND2 AND2_1593(.VSS(VSS),.VDD(VDD),.Y(g17717),.A(g4587),.B(g15385));
  AND2 AND2_1594(.VSS(VSS),.VDD(VDD),.Y(g17718),.A(g4451),.B(g16064));
  AND2 AND2_1595(.VSS(VSS),.VDD(VDD),.Y(g17719),.A(g2993),.B(g16065));
  AND2 AND2_1596(.VSS(VSS),.VDD(VDD),.Y(g17734),.A(g4611),.B(g15393));
  AND2 AND2_1597(.VSS(VSS),.VDD(VDD),.Y(g17735),.A(g4614),.B(g15396));
  AND2 AND2_1598(.VSS(VSS),.VDD(VDD),.Y(g17736),.A(g4617),.B(g15399));
  AND2 AND2_1599(.VSS(VSS),.VDD(VDD),.Y(g17737),.A(g4626),.B(g15404));
  AND2 AND2_1600(.VSS(VSS),.VDD(VDD),.Y(g17752),.A(g4656),.B(g15412));
  AND2 AND2_1601(.VSS(VSS),.VDD(VDD),.Y(g17753),.A(g4659),.B(g15415));
  AND2 AND2_1602(.VSS(VSS),.VDD(VDD),.Y(g17754),.A(g4662),.B(g15418));
  AND2 AND2_1603(.VSS(VSS),.VDD(VDD),.Y(g17773),.A(g4693),.B(g15426));
  AND2 AND2_1604(.VSS(VSS),.VDD(VDD),.Y(g17774),.A(g4696),.B(g15429));
  AND2 AND2_1605(.VSS(VSS),.VDD(VDD),.Y(g17775),.A(g4699),.B(g15432));
  AND2 AND2_1606(.VSS(VSS),.VDD(VDD),.Y(g17794),.A(g7423),.B(g16097));
  AND2 AND2_1607(.VSS(VSS),.VDD(VDD),.Y(g17795),.A(g4725),.B(g15443));
  AND2 AND2_1608(.VSS(VSS),.VDD(VDD),.Y(g17796),.A(g4728),.B(g15446));
  AND2 AND2_1609(.VSS(VSS),.VDD(VDD),.Y(g17797),.A(g4731),.B(g15449));
  AND2 AND2_1610(.VSS(VSS),.VDD(VDD),.Y(g17798),.A(g4591),.B(g16099));
  AND2 AND2_1611(.VSS(VSS),.VDD(VDD),.Y(g17812),.A(g4754),.B(g15461));
  AND2 AND2_1612(.VSS(VSS),.VDD(VDD),.Y(g17813),.A(g4757),.B(g15464));
  AND2 AND2_1613(.VSS(VSS),.VDD(VDD),.Y(g17814),.A(g4760),.B(g15467));
  AND2 AND2_1614(.VSS(VSS),.VDD(VDD),.Y(g17824),.A(g4766),.B(g15471));
  AND2 AND2_1615(.VSS(VSS),.VDD(VDD),.Y(g17835),.A(g4788),.B(g15477));
  AND2 AND2_1616(.VSS(VSS),.VDD(VDD),.Y(g17836),.A(g4791),.B(g15480));
  AND2 AND2_1617(.VSS(VSS),.VDD(VDD),.Y(g17837),.A(g4794),.B(g15483));
  AND2 AND2_1618(.VSS(VSS),.VDD(VDD),.Y(g17838),.A(g4803),.B(g15488));
  AND2 AND2_1619(.VSS(VSS),.VDD(VDD),.Y(g17853),.A(g4833),.B(g15496));
  AND2 AND2_1620(.VSS(VSS),.VDD(VDD),.Y(g17854),.A(g4836),.B(g15499));
  AND2 AND2_1621(.VSS(VSS),.VDD(VDD),.Y(g17855),.A(g4839),.B(g15502));
  AND2 AND2_1622(.VSS(VSS),.VDD(VDD),.Y(g17874),.A(g4870),.B(g15510));
  AND2 AND2_1623(.VSS(VSS),.VDD(VDD),.Y(g17875),.A(g4873),.B(g15513));
  AND2 AND2_1624(.VSS(VSS),.VDD(VDD),.Y(g17876),.A(g4876),.B(g15516));
  AND2 AND2_1625(.VSS(VSS),.VDD(VDD),.Y(g17877),.A(g2998),.B(g15521));
  AND2 AND2_1626(.VSS(VSS),.VDD(VDD),.Y(g17900),.A(g4899),.B(g15528));
  AND2 AND2_1627(.VSS(VSS),.VDD(VDD),.Y(g17901),.A(g4902),.B(g15531));
  AND2 AND2_1628(.VSS(VSS),.VDD(VDD),.Y(g17902),.A(g4905),.B(g15534));
  AND2 AND2_1629(.VSS(VSS),.VDD(VDD),.Y(g17912),.A(g4908),.B(g15537));
  AND2 AND2_1630(.VSS(VSS),.VDD(VDD),.Y(g17924),.A(g4930),.B(g15547));
  AND2 AND2_1631(.VSS(VSS),.VDD(VDD),.Y(g17925),.A(g4933),.B(g15550));
  AND2 AND2_1632(.VSS(VSS),.VDD(VDD),.Y(g17926),.A(g4936),.B(g15553));
  AND2 AND2_1633(.VSS(VSS),.VDD(VDD),.Y(g17936),.A(g4942),.B(g15557));
  AND2 AND2_1634(.VSS(VSS),.VDD(VDD),.Y(g17947),.A(g4964),.B(g15563));
  AND2 AND2_1635(.VSS(VSS),.VDD(VDD),.Y(g17948),.A(g4967),.B(g15566));
  AND2 AND2_1636(.VSS(VSS),.VDD(VDD),.Y(g17949),.A(g4970),.B(g15569));
  AND2 AND2_1637(.VSS(VSS),.VDD(VDD),.Y(g17950),.A(g4979),.B(g15574));
  AND2 AND2_1638(.VSS(VSS),.VDD(VDD),.Y(g17965),.A(g5009),.B(g15582));
  AND2 AND2_1639(.VSS(VSS),.VDD(VDD),.Y(g17966),.A(g5012),.B(g15585));
  AND2 AND2_1640(.VSS(VSS),.VDD(VDD),.Y(g17967),.A(g5015),.B(g15588));
  AND2 AND2_1641(.VSS(VSS),.VDD(VDD),.Y(g17989),.A(g5035),.B(g15596));
  AND2 AND2_1642(.VSS(VSS),.VDD(VDD),.Y(g17990),.A(g5038),.B(g15599));
  AND2 AND2_1643(.VSS(VSS),.VDD(VDD),.Y(g18011),.A(g5058),.B(g15606));
  AND2 AND2_1644(.VSS(VSS),.VDD(VDD),.Y(g18012),.A(g5061),.B(g15609));
  AND2 AND2_1645(.VSS(VSS),.VDD(VDD),.Y(g18013),.A(g5064),.B(g15612));
  AND2 AND2_1646(.VSS(VSS),.VDD(VDD),.Y(g18023),.A(g5067),.B(g15615));
  AND2 AND2_1647(.VSS(VSS),.VDD(VDD),.Y(g18035),.A(g5089),.B(g15625));
  AND2 AND2_1648(.VSS(VSS),.VDD(VDD),.Y(g18036),.A(g5092),.B(g15628));
  AND2 AND2_1649(.VSS(VSS),.VDD(VDD),.Y(g18037),.A(g5095),.B(g15631));
  AND2 AND2_1650(.VSS(VSS),.VDD(VDD),.Y(g18047),.A(g5101),.B(g15635));
  AND2 AND2_1651(.VSS(VSS),.VDD(VDD),.Y(g18058),.A(g5123),.B(g15641));
  AND2 AND2_1652(.VSS(VSS),.VDD(VDD),.Y(g18059),.A(g5126),.B(g15644));
  AND2 AND2_1653(.VSS(VSS),.VDD(VDD),.Y(g18060),.A(g5129),.B(g15647));
  AND2 AND2_1654(.VSS(VSS),.VDD(VDD),.Y(g18061),.A(g5138),.B(g15652));
  AND2 AND2_1655(.VSS(VSS),.VDD(VDD),.Y(g18062),.A(g7462),.B(g15655));
  AND2 AND2_1656(.VSS(VSS),.VDD(VDD),.Y(g18088),.A(g5150),.B(g15667));
  AND2 AND2_1657(.VSS(VSS),.VDD(VDD),.Y(g18106),.A(g5164),.B(g15672));
  AND2 AND2_1658(.VSS(VSS),.VDD(VDD),.Y(g18107),.A(g5167),.B(g15675));
  AND2 AND2_1659(.VSS(VSS),.VDD(VDD),.Y(g18128),.A(g5187),.B(g15682));
  AND2 AND2_1660(.VSS(VSS),.VDD(VDD),.Y(g18129),.A(g5190),.B(g15685));
  AND2 AND2_1661(.VSS(VSS),.VDD(VDD),.Y(g18130),.A(g5193),.B(g15688));
  AND2 AND2_1662(.VSS(VSS),.VDD(VDD),.Y(g18140),.A(g5196),.B(g15691));
  AND2 AND2_1663(.VSS(VSS),.VDD(VDD),.Y(g18152),.A(g5218),.B(g15701));
  AND2 AND2_1664(.VSS(VSS),.VDD(VDD),.Y(g18153),.A(g5221),.B(g15704));
  AND2 AND2_1665(.VSS(VSS),.VDD(VDD),.Y(g18154),.A(g5224),.B(g15707));
  AND2 AND2_1666(.VSS(VSS),.VDD(VDD),.Y(g18164),.A(g5230),.B(g15711));
  AND2 AND2_1667(.VSS(VSS),.VDD(VDD),.Y(g18165),.A(g2883),.B(g16287));
  AND2 AND2_1668(.VSS(VSS),.VDD(VDD),.Y(g18169),.A(g7527),.B(g15714));
  AND2 AND2_1669(.VSS(VSS),.VDD(VDD),.Y(g18204),.A(g5243),.B(g15726));
  AND2 AND2_1670(.VSS(VSS),.VDD(VDD),.Y(g18222),.A(g5257),.B(g15731));
  AND2 AND2_1671(.VSS(VSS),.VDD(VDD),.Y(g18223),.A(g5260),.B(g15734));
  AND2 AND2_1672(.VSS(VSS),.VDD(VDD),.Y(g18244),.A(g5280),.B(g15741));
  AND2 AND2_1673(.VSS(VSS),.VDD(VDD),.Y(g18245),.A(g5283),.B(g15744));
  AND2 AND2_1674(.VSS(VSS),.VDD(VDD),.Y(g18246),.A(g5286),.B(g15747));
  AND2 AND2_1675(.VSS(VSS),.VDD(VDD),.Y(g18256),.A(g5289),.B(g15750));
  AND2 AND2_1676(.VSS(VSS),.VDD(VDD),.Y(g18311),.A(g5306),.B(g15766));
  AND2 AND2_1677(.VSS(VSS),.VDD(VDD),.Y(g18329),.A(g5320),.B(g15771));
  AND2 AND2_1678(.VSS(VSS),.VDD(VDD),.Y(g18330),.A(g5323),.B(g15774));
  AND2 AND2_1679(.VSS(VSS),.VDD(VDD),.Y(g18333),.A(g2888),.B(g15777));
  AND2 AND2_1680(.VSS(VSS),.VDD(VDD),.Y(g18404),.A(g5343),.B(g15794));
  AND3 AND3_18(.VSS(VSS),.VDD(VDD),.Y(I24619),.A(g14776),.B(g14837),.C(g16142));
  AND3 AND3_19(.VSS(VSS),.VDD(VDD),.Y(g18547),.A(g13677),.B(g13750),.C(I24619));
  AND3 AND3_20(.VSS(VSS),.VDD(VDD),.Y(I24689),.A(g14811),.B(g14910),.C(g16201));
  AND3 AND3_21(.VSS(VSS),.VDD(VDD),.Y(g18597),.A(g13714),.B(g13791),.C(I24689));
  AND3 AND3_22(.VSS(VSS),.VDD(VDD),.Y(I24738),.A(g14863),.B(g14991),.C(g16266));
  AND3 AND3_23(.VSS(VSS),.VDD(VDD),.Y(g18629),.A(g13764),.B(g13819),.C(I24738));
  AND3 AND3_24(.VSS(VSS),.VDD(VDD),.Y(I24758),.A(g14936),.B(g15080),.C(g16325));
  AND3 AND3_25(.VSS(VSS),.VDD(VDD),.Y(g18638),.A(g13805),.B(g13840),.C(I24758));
  AND4 AND4_28(.VSS(VSS),.VDD(VDD),.Y(g18645),.A(g14776),.B(g14895),.C(g16142),.D(g13750));
  AND3 AND3_26(.VSS(VSS),.VDD(VDD),.Y(g18647),.A(g14895),.B(g16142),.C(g16243));
  AND4 AND4_29(.VSS(VSS),.VDD(VDD),.Y(g18648),.A(g14811),.B(g14976),.C(g16201),.D(g13791));
  AND4 AND4_30(.VSS(VSS),.VDD(VDD),.Y(g18649),.A(g14776),.B(g14837),.C(g13657),.D(g16189));
  AND3 AND3_27(.VSS(VSS),.VDD(VDD),.Y(g18650),.A(g14976),.B(g16201),.C(g16302));
  AND4 AND4_31(.VSS(VSS),.VDD(VDD),.Y(g18651),.A(g14863),.B(g15065),.C(g16266),.D(g13819));
  AND4 AND4_32(.VSS(VSS),.VDD(VDD),.Y(g18652),.A(g14797),.B(g13657),.C(g13677),.D(g16243));
  AND4 AND4_33(.VSS(VSS),.VDD(VDD),.Y(g18653),.A(g14811),.B(g14910),.C(g13687),.D(g16254));
  AND3 AND3_28(.VSS(VSS),.VDD(VDD),.Y(g18654),.A(g15065),.B(g16266),.C(g16360));
  AND4 AND4_34(.VSS(VSS),.VDD(VDD),.Y(g18655),.A(g14936),.B(g15161),.C(g16325),.D(g13840));
  AND4 AND4_35(.VSS(VSS),.VDD(VDD),.Y(g18665),.A(g14776),.B(g14837),.C(g16189),.D(g13706));
  AND4 AND4_36(.VSS(VSS),.VDD(VDD),.Y(g18666),.A(g14849),.B(g13687),.C(g13714),.D(g16302));
  AND4 AND4_37(.VSS(VSS),.VDD(VDD),.Y(g18667),.A(g14863),.B(g14991),.C(g13724),.D(g16313));
  AND3 AND3_29(.VSS(VSS),.VDD(VDD),.Y(g18668),.A(g15161),.B(g16325),.C(g16404));
  AND4 AND4_38(.VSS(VSS),.VDD(VDD),.Y(g18688),.A(g14811),.B(g14910),.C(g16254),.D(g13756));
  AND4 AND4_39(.VSS(VSS),.VDD(VDD),.Y(g18689),.A(g14922),.B(g13724),.C(g13764),.D(g16360));
  AND4 AND4_40(.VSS(VSS),.VDD(VDD),.Y(g18690),.A(g14936),.B(g15080),.C(g13774),.D(g16371));
  AND4 AND4_41(.VSS(VSS),.VDD(VDD),.Y(g18717),.A(g14863),.B(g14991),.C(g16313),.D(g13797));
  AND4 AND4_42(.VSS(VSS),.VDD(VDD),.Y(g18718),.A(g15003),.B(g13774),.C(g13805),.D(g16404));
  AND4 AND4_43(.VSS(VSS),.VDD(VDD),.Y(g18753),.A(g14936),.B(g15080),.C(g16371),.D(g13825));
  AND2 AND2_1681(.VSS(VSS),.VDD(VDD),.Y(g18982),.A(g13519),.B(g16154));
  AND2 AND2_1682(.VSS(VSS),.VDD(VDD),.Y(g18990),.A(g13530),.B(g16213));
  AND4 AND4_44(.VSS(VSS),.VDD(VDD),.Y(g18994),.A(g14895),.B(g13657),.C(g13677),.D(g13706));
  AND2 AND2_1683(.VSS(VSS),.VDD(VDD),.Y(g18997),.A(g13541),.B(g16278));
  AND4 AND4_45(.VSS(VSS),.VDD(VDD),.Y(g19007),.A(g14976),.B(g13687),.C(g13714),.D(g13756));
  AND2 AND2_1684(.VSS(VSS),.VDD(VDD),.Y(g19010),.A(g13552),.B(g16337));
  AND4 AND4_46(.VSS(VSS),.VDD(VDD),.Y(g19063),.A(g18679),.B(g14910),.C(g13687),.D(g16254));
  AND4 AND4_47(.VSS(VSS),.VDD(VDD),.Y(g19079),.A(g14797),.B(g18692),.C(g16142),.D(g16189));
  AND4 AND4_48(.VSS(VSS),.VDD(VDD),.Y(g19080),.A(g18708),.B(g14991),.C(g13724),.D(g16313));
  AND2 AND2_1685(.VSS(VSS),.VDD(VDD),.Y(g19087),.A(g17215),.B(g16540));
  AND4 AND4_49(.VSS(VSS),.VDD(VDD),.Y(g19088),.A(g18656),.B(g14797),.C(g16189),.D(g13706));
  AND4 AND4_50(.VSS(VSS),.VDD(VDD),.Y(g19089),.A(g14849),.B(g18728),.C(g16201),.D(g16254));
  AND4 AND4_51(.VSS(VSS),.VDD(VDD),.Y(g19090),.A(g18744),.B(g15080),.C(g13774),.D(g16371));
  AND4 AND4_52(.VSS(VSS),.VDD(VDD),.Y(g19092),.A(g14776),.B(g18670),.C(g18692),.D(g16293));
  AND2 AND2_1686(.VSS(VSS),.VDD(VDD),.Y(g19093),.A(g17218),.B(g16572));
  AND4 AND4_53(.VSS(VSS),.VDD(VDD),.Y(g19094),.A(g18679),.B(g14849),.C(g16254),.D(g13756));
  AND4 AND4_54(.VSS(VSS),.VDD(VDD),.Y(g19095),.A(g14922),.B(g18765),.C(g16266),.D(g16313));
  AND3 AND3_30(.VSS(VSS),.VDD(VDD),.Y(I25280),.A(g18656),.B(g18670),.C(g18720));
  AND3 AND3_31(.VSS(VSS),.VDD(VDD),.Y(g19097),.A(g13657),.B(g16243),.C(I25280));
  AND4 AND4_55(.VSS(VSS),.VDD(VDD),.Y(g19099),.A(g14811),.B(g18699),.C(g18728),.D(g16351));
  AND2 AND2_1687(.VSS(VSS),.VDD(VDD),.Y(g19100),.A(g17220),.B(g16596));
  AND4 AND4_56(.VSS(VSS),.VDD(VDD),.Y(g19101),.A(g18708),.B(g14922),.C(g16313),.D(g13797));
  AND4 AND4_57(.VSS(VSS),.VDD(VDD),.Y(g19102),.A(g15003),.B(g18796),.C(g16325),.D(g16371));
  AND3 AND3_32(.VSS(VSS),.VDD(VDD),.Y(I25291),.A(g18679),.B(g18699),.C(g18758));
  AND3 AND3_33(.VSS(VSS),.VDD(VDD),.Y(g19104),.A(g13687),.B(g16302),.C(I25291));
  AND4 AND4_58(.VSS(VSS),.VDD(VDD),.Y(g19106),.A(g14863),.B(g18735),.C(g18765),.D(g16395));
  AND2 AND2_1688(.VSS(VSS),.VDD(VDD),.Y(g19107),.A(g17223),.B(g16616));
  AND4 AND4_59(.VSS(VSS),.VDD(VDD),.Y(g19108),.A(g18744),.B(g15003),.C(g16371),.D(g13825));
  AND3 AND3_34(.VSS(VSS),.VDD(VDD),.Y(I25300),.A(g18708),.B(g18735),.C(g18789));
  AND3 AND3_35(.VSS(VSS),.VDD(VDD),.Y(g19109),.A(g13724),.B(g16360),.C(I25300));
  AND4 AND4_60(.VSS(VSS),.VDD(VDD),.Y(g19111),.A(g14936),.B(g18772),.C(g18796),.D(g16433));
  AND2 AND2_1689(.VSS(VSS),.VDD(VDD),.Y(g19112),.A(g14657),.B(g16633));
  AND3 AND3_36(.VSS(VSS),.VDD(VDD),.Y(I25311),.A(g18744),.B(g18772),.C(g18815));
  AND3 AND3_37(.VSS(VSS),.VDD(VDD),.Y(g19116),.A(g13774),.B(g16404),.C(I25311));
  AND2 AND2_1690(.VSS(VSS),.VDD(VDD),.Y(g19117),.A(g14691),.B(g16644));
  AND2 AND2_1691(.VSS(VSS),.VDD(VDD),.Y(g19124),.A(g14725),.B(g16656));
  AND2 AND2_1692(.VSS(VSS),.VDD(VDD),.Y(g19131),.A(g14753),.B(g16673));
  AND2 AND2_1693(.VSS(VSS),.VDD(VDD),.Y(g19142),.A(g17159),.B(g16719));
  AND2 AND2_1694(.VSS(VSS),.VDD(VDD),.Y(g19143),.A(g17174),.B(g16761));
  AND2 AND2_1695(.VSS(VSS),.VDD(VDD),.Y(g19146),.A(g17191),.B(g16788));
  AND2 AND2_1696(.VSS(VSS),.VDD(VDD),.Y(g19148),.A(g17202),.B(g16817));
  AND2 AND2_1697(.VSS(VSS),.VDD(VDD),.Y(g19150),.A(g17189),.B(g8602));
  AND2 AND2_1698(.VSS(VSS),.VDD(VDD),.Y(g19155),.A(g17200),.B(g8614));
  AND2 AND2_1699(.VSS(VSS),.VDD(VDD),.Y(g19161),.A(g17207),.B(g8627));
  AND2 AND2_1700(.VSS(VSS),.VDD(VDD),.Y(g19166),.A(g17212),.B(g8637));
  AND2 AND2_1701(.VSS(VSS),.VDD(VDD),.Y(g19228),.A(g16662),.B(g12125));
  AND2 AND2_1702(.VSS(VSS),.VDD(VDD),.Y(g19236),.A(g16935),.B(g8802));
  AND3 AND3_38(.VSS(VSS),.VDD(VDD),.Y(g19241),.A(g16867),.B(g14158),.C(g14071));
  AND2 AND2_1703(.VSS(VSS),.VDD(VDD),.Y(g19248),.A(g16662),.B(g8817));
  AND2 AND2_1704(.VSS(VSS),.VDD(VDD),.Y(g19252),.A(g18725),.B(g9527));
  AND3 AND3_39(.VSS(VSS),.VDD(VDD),.Y(g19254),.A(g16895),.B(g14273),.C(g14186));
  AND2 AND2_1705(.VSS(VSS),.VDD(VDD),.Y(g19260),.A(g16749),.B(g3124));
  AND3 AND3_40(.VSS(VSS),.VDD(VDD),.Y(g19267),.A(g16924),.B(g14395),.C(g14301));
  AND3 AND3_41(.VSS(VSS),.VDD(VDD),.Y(g19282),.A(g16954),.B(g14507),.C(g14423));
  AND2 AND2_1706(.VSS(VSS),.VDD(VDD),.Y(g19284),.A(g18063),.B(g3111));
  AND2 AND2_1707(.VSS(VSS),.VDD(VDD),.Y(g19285),.A(g16749),.B(g7642));
  AND2 AND2_1708(.VSS(VSS),.VDD(VDD),.Y(g19289),.A(g17029),.B(g8580));
  AND3 AND3_42(.VSS(VSS),.VDD(VDD),.Y(g19303),.A(g16867),.B(g16543),.C(g14071));
  AND2 AND2_1709(.VSS(VSS),.VDD(VDD),.Y(g19307),.A(g17063),.B(g8587));
  AND2 AND2_1710(.VSS(VSS),.VDD(VDD),.Y(g19316),.A(g18063),.B(g3110));
  AND2 AND2_1711(.VSS(VSS),.VDD(VDD),.Y(g19317),.A(g16749),.B(g3126));
  AND3 AND3_43(.VSS(VSS),.VDD(VDD),.Y(g19320),.A(g16867),.B(g16515),.C(g14158));
  AND3 AND3_44(.VSS(VSS),.VDD(VDD),.Y(g19324),.A(g16895),.B(g16575),.C(g14186));
  AND2 AND2_1712(.VSS(VSS),.VDD(VDD),.Y(g19328),.A(g17098),.B(g8594));
  AND3 AND3_45(.VSS(VSS),.VDD(VDD),.Y(g19347),.A(g16895),.B(g16546),.C(g14273));
  AND3 AND3_46(.VSS(VSS),.VDD(VDD),.Y(g19351),.A(g16924),.B(g16599),.C(g14301));
  AND2 AND2_1713(.VSS(VSS),.VDD(VDD),.Y(g19355),.A(g17136),.B(g8605));
  AND2 AND2_1714(.VSS(VSS),.VDD(VDD),.Y(g19356),.A(g18063),.B(g3112));
  AND3 AND3_47(.VSS(VSS),.VDD(VDD),.Y(g19381),.A(g16924),.B(g16578),.C(g14395));
  AND3 AND3_48(.VSS(VSS),.VDD(VDD),.Y(g19385),.A(g16954),.B(g16619),.C(g14423));
  AND3 AND3_49(.VSS(VSS),.VDD(VDD),.Y(g19413),.A(g16954),.B(g16602),.C(g14507));
  AND3 AND3_50(.VSS(VSS),.VDD(VDD),.Y(g19449),.A(g16884),.B(g14797),.C(g14776));
  AND3 AND3_51(.VSS(VSS),.VDD(VDD),.Y(g19476),.A(g16913),.B(g14849),.C(g14811));
  AND3 AND3_52(.VSS(VSS),.VDD(VDD),.Y(g19499),.A(g16943),.B(g14922),.C(g14863));
  AND3 AND3_53(.VSS(VSS),.VDD(VDD),.Y(g19520),.A(g16974),.B(g15003),.C(g14936));
  AND3 AND3_54(.VSS(VSS),.VDD(VDD),.Y(g19531),.A(g16884),.B(g16722),.C(g14776));
  AND3 AND3_55(.VSS(VSS),.VDD(VDD),.Y(g19540),.A(g16884),.B(g16697),.C(g14797));
  AND3 AND3_56(.VSS(VSS),.VDD(VDD),.Y(g19541),.A(g16913),.B(g16764),.C(g14811));
  AND3 AND3_57(.VSS(VSS),.VDD(VDD),.Y(g19544),.A(g16913),.B(g16728),.C(g14849));
  AND3 AND3_58(.VSS(VSS),.VDD(VDD),.Y(g19545),.A(g16943),.B(g16791),.C(g14863));
  AND3 AND3_59(.VSS(VSS),.VDD(VDD),.Y(g19547),.A(g16943),.B(g16770),.C(g14922));
  AND3 AND3_60(.VSS(VSS),.VDD(VDD),.Y(g19548),.A(g16974),.B(g16820),.C(g14936));
  AND2 AND2_1715(.VSS(VSS),.VDD(VDD),.Y(g19549),.A(g7950),.B(g17230));
  AND3 AND3_61(.VSS(VSS),.VDD(VDD),.Y(g19551),.A(g16974),.B(g16797),.C(g15003));
  AND2 AND2_1716(.VSS(VSS),.VDD(VDD),.Y(g19552),.A(g16829),.B(g6048));
  AND2 AND2_1717(.VSS(VSS),.VDD(VDD),.Y(g19553),.A(g7990),.B(g17237));
  AND2 AND2_1718(.VSS(VSS),.VDD(VDD),.Y(g19554),.A(g7993),.B(g17240));
  AND2 AND2_1719(.VSS(VSS),.VDD(VDD),.Y(g19555),.A(g8001),.B(g17243));
  AND2 AND2_1720(.VSS(VSS),.VDD(VDD),.Y(g19557),.A(g8053),.B(g17249));
  AND2 AND2_1721(.VSS(VSS),.VDD(VDD),.Y(g19558),.A(g8056),.B(g17252));
  AND2 AND2_1722(.VSS(VSS),.VDD(VDD),.Y(g19559),.A(g8059),.B(g17255));
  AND2 AND2_1723(.VSS(VSS),.VDD(VDD),.Y(g19560),.A(g8065),.B(g17259));
  AND2 AND2_1724(.VSS(VSS),.VDD(VDD),.Y(g19561),.A(g8068),.B(g17262));
  AND2 AND2_1725(.VSS(VSS),.VDD(VDD),.Y(g19562),.A(g8076),.B(g17265));
  AND2 AND2_1726(.VSS(VSS),.VDD(VDD),.Y(g19564),.A(g8123),.B(g17272));
  AND2 AND2_1727(.VSS(VSS),.VDD(VDD),.Y(g19565),.A(g8126),.B(g17275));
  AND2 AND2_1728(.VSS(VSS),.VDD(VDD),.Y(g19566),.A(g8129),.B(g17278));
  AND2 AND2_1729(.VSS(VSS),.VDD(VDD),.Y(g19567),.A(g8138),.B(g17282));
  AND2 AND2_1730(.VSS(VSS),.VDD(VDD),.Y(g19568),.A(g8141),.B(g17285));
  AND2 AND2_1731(.VSS(VSS),.VDD(VDD),.Y(g19569),.A(g8144),.B(g17288));
  AND2 AND2_1732(.VSS(VSS),.VDD(VDD),.Y(g19570),.A(g8150),.B(g17291));
  AND2 AND2_1733(.VSS(VSS),.VDD(VDD),.Y(g19571),.A(g8153),.B(g17294));
  AND2 AND2_1734(.VSS(VSS),.VDD(VDD),.Y(g19572),.A(g8161),.B(g17297));
  AND2 AND2_1735(.VSS(VSS),.VDD(VDD),.Y(g19574),.A(g8191),.B(g17304));
  AND2 AND2_1736(.VSS(VSS),.VDD(VDD),.Y(g19575),.A(g8194),.B(g17307));
  AND2 AND2_1737(.VSS(VSS),.VDD(VDD),.Y(g19576),.A(g8197),.B(g17310));
  AND2 AND2_1738(.VSS(VSS),.VDD(VDD),.Y(g19584),.A(g640),.B(g18756));
  AND2 AND2_1739(.VSS(VSS),.VDD(VDD),.Y(g19585),.A(g692),.B(g18757));
  AND2 AND2_1740(.VSS(VSS),.VDD(VDD),.Y(g19586),.A(g8209),.B(g17315));
  AND2 AND2_1741(.VSS(VSS),.VDD(VDD),.Y(g19587),.A(g8212),.B(g17318));
  AND2 AND2_1742(.VSS(VSS),.VDD(VDD),.Y(g19588),.A(g8215),.B(g17321));
  AND2 AND2_1743(.VSS(VSS),.VDD(VDD),.Y(g19589),.A(g8224),.B(g17324));
  AND2 AND2_1744(.VSS(VSS),.VDD(VDD),.Y(g19590),.A(g8227),.B(g17327));
  AND2 AND2_1745(.VSS(VSS),.VDD(VDD),.Y(g19591),.A(g8230),.B(g17330));
  AND2 AND2_1746(.VSS(VSS),.VDD(VDD),.Y(g19592),.A(g8236),.B(g17333));
  AND2 AND2_1747(.VSS(VSS),.VDD(VDD),.Y(g19593),.A(g8239),.B(g17336));
  AND2 AND2_1748(.VSS(VSS),.VDD(VDD),.Y(g19594),.A(g16935),.B(g12555));
  AND2 AND2_1749(.VSS(VSS),.VDD(VDD),.Y(g19597),.A(g3922),.B(g17342));
  AND2 AND2_1750(.VSS(VSS),.VDD(VDD),.Y(g19598),.A(g3925),.B(g17345));
  AND2 AND2_1751(.VSS(VSS),.VDD(VDD),.Y(g19599),.A(g3928),.B(g17348));
  AND2 AND2_1752(.VSS(VSS),.VDD(VDD),.Y(g19600),.A(g633),.B(g18783));
  AND2 AND2_1753(.VSS(VSS),.VDD(VDD),.Y(g19601),.A(g640),.B(g18784));
  AND2 AND2_1754(.VSS(VSS),.VDD(VDD),.Y(g19602),.A(g633),.B(g18785));
  AND2 AND2_1755(.VSS(VSS),.VDD(VDD),.Y(g19603),.A(g692),.B(g18786));
  AND2 AND2_1756(.VSS(VSS),.VDD(VDD),.Y(g19604),.A(g3948),.B(g17354));
  AND2 AND2_1757(.VSS(VSS),.VDD(VDD),.Y(g19605),.A(g3951),.B(g17357));
  AND2 AND2_1758(.VSS(VSS),.VDD(VDD),.Y(g19606),.A(g3954),.B(g17360));
  AND2 AND2_1759(.VSS(VSS),.VDD(VDD),.Y(g19614),.A(g1326),.B(g18787));
  AND2 AND2_1760(.VSS(VSS),.VDD(VDD),.Y(g19615),.A(g1378),.B(g18788));
  AND2 AND2_1761(.VSS(VSS),.VDD(VDD),.Y(g19616),.A(g3966),.B(g17363));
  AND2 AND2_1762(.VSS(VSS),.VDD(VDD),.Y(g19617),.A(g3969),.B(g17366));
  AND2 AND2_1763(.VSS(VSS),.VDD(VDD),.Y(g19618),.A(g3972),.B(g17369));
  AND2 AND2_1764(.VSS(VSS),.VDD(VDD),.Y(g19619),.A(g3981),.B(g17372));
  AND2 AND2_1765(.VSS(VSS),.VDD(VDD),.Y(g19620),.A(g3984),.B(g17375));
  AND2 AND2_1766(.VSS(VSS),.VDD(VDD),.Y(g19621),.A(g3987),.B(g17378));
  AND2 AND2_1767(.VSS(VSS),.VDD(VDD),.Y(g19623),.A(g4000),.B(g17384));
  AND2 AND2_1768(.VSS(VSS),.VDD(VDD),.Y(g19624),.A(g4003),.B(g17387));
  AND2 AND2_1769(.VSS(VSS),.VDD(VDD),.Y(g19625),.A(g4006),.B(g17390));
  AND2 AND2_1770(.VSS(VSS),.VDD(VDD),.Y(g19626),.A(g640),.B(g18805));
  AND2 AND2_1771(.VSS(VSS),.VDD(VDD),.Y(g19627),.A(g633),.B(g18806));
  AND2 AND2_1772(.VSS(VSS),.VDD(VDD),.Y(g19628),.A(g653),.B(g18807));
  AND2 AND2_1773(.VSS(VSS),.VDD(VDD),.Y(g19629),.A(g692),.B(g18808));
  AND2 AND2_1774(.VSS(VSS),.VDD(VDD),.Y(g19630),.A(g4029),.B(g17399));
  AND2 AND2_1775(.VSS(VSS),.VDD(VDD),.Y(g19631),.A(g4032),.B(g17402));
  AND2 AND2_1776(.VSS(VSS),.VDD(VDD),.Y(g19632),.A(g4035),.B(g17405));
  AND2 AND2_1777(.VSS(VSS),.VDD(VDD),.Y(g19633),.A(g1319),.B(g18809));
  AND2 AND2_1778(.VSS(VSS),.VDD(VDD),.Y(g19634),.A(g1326),.B(g18810));
  AND2 AND2_1779(.VSS(VSS),.VDD(VDD),.Y(g19635),.A(g1319),.B(g18811));
  AND2 AND2_1780(.VSS(VSS),.VDD(VDD),.Y(g19636),.A(g1378),.B(g18812));
  AND2 AND2_1781(.VSS(VSS),.VDD(VDD),.Y(g19637),.A(g4055),.B(g17410));
  AND2 AND2_1782(.VSS(VSS),.VDD(VDD),.Y(g19638),.A(g4058),.B(g17413));
  AND2 AND2_1783(.VSS(VSS),.VDD(VDD),.Y(g19639),.A(g4061),.B(g17416));
  AND2 AND2_1784(.VSS(VSS),.VDD(VDD),.Y(g19647),.A(g2020),.B(g18813));
  AND2 AND2_1785(.VSS(VSS),.VDD(VDD),.Y(g19648),.A(g2072),.B(g18814));
  AND2 AND2_1786(.VSS(VSS),.VDD(VDD),.Y(g19649),.A(g4073),.B(g17419));
  AND2 AND2_1787(.VSS(VSS),.VDD(VDD),.Y(g19650),.A(g4076),.B(g17422));
  AND2 AND2_1788(.VSS(VSS),.VDD(VDD),.Y(g19651),.A(g4079),.B(g17425));
  AND2 AND2_1789(.VSS(VSS),.VDD(VDD),.Y(g19653),.A(g4095),.B(g17430));
  AND2 AND2_1790(.VSS(VSS),.VDD(VDD),.Y(g19654),.A(g4098),.B(g17433));
  AND2 AND2_1791(.VSS(VSS),.VDD(VDD),.Y(g19655),.A(g4101),.B(g17436));
  AND2 AND2_1792(.VSS(VSS),.VDD(VDD),.Y(g19656),.A(g4104),.B(g17439));
  AND2 AND2_1793(.VSS(VSS),.VDD(VDD),.Y(g19660),.A(g633),.B(g18822));
  AND2 AND2_1794(.VSS(VSS),.VDD(VDD),.Y(g19661),.A(g653),.B(g18823));
  AND2 AND2_1795(.VSS(VSS),.VDD(VDD),.Y(g19662),.A(g646),.B(g18824));
  AND2 AND2_1796(.VSS(VSS),.VDD(VDD),.Y(g19663),.A(g4127),.B(g17451));
  AND2 AND2_1797(.VSS(VSS),.VDD(VDD),.Y(g19664),.A(g4130),.B(g17454));
  AND2 AND2_1798(.VSS(VSS),.VDD(VDD),.Y(g19665),.A(g4133),.B(g17457));
  AND2 AND2_1799(.VSS(VSS),.VDD(VDD),.Y(g19666),.A(g1326),.B(g18825));
  AND2 AND2_1800(.VSS(VSS),.VDD(VDD),.Y(g19667),.A(g1319),.B(g18826));
  AND2 AND2_1801(.VSS(VSS),.VDD(VDD),.Y(g19668),.A(g1339),.B(g18827));
  AND2 AND2_1802(.VSS(VSS),.VDD(VDD),.Y(g19669),.A(g1378),.B(g18828));
  AND2 AND2_1803(.VSS(VSS),.VDD(VDD),.Y(g19670),.A(g4156),.B(g17465));
  AND2 AND2_1804(.VSS(VSS),.VDD(VDD),.Y(g19671),.A(g4159),.B(g17468));
  AND2 AND2_1805(.VSS(VSS),.VDD(VDD),.Y(g19672),.A(g4162),.B(g17471));
  AND2 AND2_1806(.VSS(VSS),.VDD(VDD),.Y(g19673),.A(g2013),.B(g18829));
  AND2 AND2_1807(.VSS(VSS),.VDD(VDD),.Y(g19674),.A(g2020),.B(g18830));
  AND2 AND2_1808(.VSS(VSS),.VDD(VDD),.Y(g19675),.A(g2013),.B(g18831));
  AND2 AND2_1809(.VSS(VSS),.VDD(VDD),.Y(g19676),.A(g2072),.B(g18832));
  AND2 AND2_1810(.VSS(VSS),.VDD(VDD),.Y(g19677),.A(g4182),.B(g17476));
  AND2 AND2_1811(.VSS(VSS),.VDD(VDD),.Y(g19678),.A(g4185),.B(g17479));
  AND2 AND2_1812(.VSS(VSS),.VDD(VDD),.Y(g19679),.A(g4188),.B(g17482));
  AND2 AND2_1813(.VSS(VSS),.VDD(VDD),.Y(g19687),.A(g2714),.B(g18833));
  AND2 AND2_1814(.VSS(VSS),.VDD(VDD),.Y(g19688),.A(g2766),.B(g18834));
  AND2 AND2_1815(.VSS(VSS),.VDD(VDD),.Y(g19691),.A(g16841),.B(g10865));
  AND2 AND2_1816(.VSS(VSS),.VDD(VDD),.Y(g19692),.A(g4205),.B(g17487));
  AND2 AND2_1817(.VSS(VSS),.VDD(VDD),.Y(g19693),.A(g4208),.B(g17490));
  AND2 AND2_1818(.VSS(VSS),.VDD(VDD),.Y(g19694),.A(g4211),.B(g17493));
  AND2 AND2_1819(.VSS(VSS),.VDD(VDD),.Y(g19695),.A(g4214),.B(g17496));
  AND2 AND2_1820(.VSS(VSS),.VDD(VDD),.Y(g19697),.A(g653),.B(g18838));
  AND2 AND2_1821(.VSS(VSS),.VDD(VDD),.Y(g19698),.A(g646),.B(g18839));
  AND2 AND2_1822(.VSS(VSS),.VDD(VDD),.Y(g19699),.A(g660),.B(g18840));
  AND2 AND2_1823(.VSS(VSS),.VDD(VDD),.Y(g19700),.A(g17815),.B(g16024));
  AND2 AND2_1824(.VSS(VSS),.VDD(VDD),.Y(g19701),.A(g4234),.B(g17511));
  AND2 AND2_1825(.VSS(VSS),.VDD(VDD),.Y(g19702),.A(g4237),.B(g17514));
  AND2 AND2_1826(.VSS(VSS),.VDD(VDD),.Y(g19703),.A(g4240),.B(g17517));
  AND2 AND2_1827(.VSS(VSS),.VDD(VDD),.Y(g19704),.A(g4243),.B(g17520));
  AND2 AND2_1828(.VSS(VSS),.VDD(VDD),.Y(g19708),.A(g1319),.B(g18841));
  AND2 AND2_1829(.VSS(VSS),.VDD(VDD),.Y(g19709),.A(g1339),.B(g18842));
  AND2 AND2_1830(.VSS(VSS),.VDD(VDD),.Y(g19710),.A(g1332),.B(g18843));
  AND2 AND2_1831(.VSS(VSS),.VDD(VDD),.Y(g19711),.A(g4266),.B(g17531));
  AND2 AND2_1832(.VSS(VSS),.VDD(VDD),.Y(g19712),.A(g4269),.B(g17534));
  AND2 AND2_1833(.VSS(VSS),.VDD(VDD),.Y(g19713),.A(g4272),.B(g17537));
  AND2 AND2_1834(.VSS(VSS),.VDD(VDD),.Y(g19714),.A(g2020),.B(g18844));
  AND2 AND2_1835(.VSS(VSS),.VDD(VDD),.Y(g19715),.A(g2013),.B(g18845));
  AND2 AND2_1836(.VSS(VSS),.VDD(VDD),.Y(g19716),.A(g2033),.B(g18846));
  AND2 AND2_1837(.VSS(VSS),.VDD(VDD),.Y(g19717),.A(g2072),.B(g18847));
  AND2 AND2_1838(.VSS(VSS),.VDD(VDD),.Y(g19718),.A(g4295),.B(g17545));
  AND2 AND2_1839(.VSS(VSS),.VDD(VDD),.Y(g19719),.A(g4298),.B(g17548));
  AND2 AND2_1840(.VSS(VSS),.VDD(VDD),.Y(g19720),.A(g4301),.B(g17551));
  AND2 AND2_1841(.VSS(VSS),.VDD(VDD),.Y(g19721),.A(g2707),.B(g18848));
  AND2 AND2_1842(.VSS(VSS),.VDD(VDD),.Y(g19722),.A(g2714),.B(g18849));
  AND2 AND2_1843(.VSS(VSS),.VDD(VDD),.Y(g19723),.A(g2707),.B(g18850));
  AND2 AND2_1844(.VSS(VSS),.VDD(VDD),.Y(g19724),.A(g2766),.B(g18851));
  AND2 AND2_1845(.VSS(VSS),.VDD(VDD),.Y(g19726),.A(g16847),.B(g6131));
  AND2 AND2_1846(.VSS(VSS),.VDD(VDD),.Y(g19727),.A(g4329),.B(g17557));
  AND2 AND2_1847(.VSS(VSS),.VDD(VDD),.Y(g19728),.A(g4332),.B(g17560));
  AND2 AND2_1848(.VSS(VSS),.VDD(VDD),.Y(g19729),.A(g4335),.B(g17563));
  AND2 AND2_1849(.VSS(VSS),.VDD(VDD),.Y(g19730),.A(g653),.B(g17573));
  AND2 AND2_1850(.VSS(VSS),.VDD(VDD),.Y(g19731),.A(g646),.B(g18853));
  AND2 AND2_1851(.VSS(VSS),.VDD(VDD),.Y(g19732),.A(g660),.B(g18854));
  AND2 AND2_1852(.VSS(VSS),.VDD(VDD),.Y(g19733),.A(g672),.B(g18855));
  AND2 AND2_1853(.VSS(VSS),.VDD(VDD),.Y(g19734),.A(g17815),.B(g16034));
  AND2 AND2_1854(.VSS(VSS),.VDD(VDD),.Y(g19735),.A(g17903),.B(g16035));
  AND2 AND2_1855(.VSS(VSS),.VDD(VDD),.Y(g19736),.A(g4360),.B(g17579));
  AND2 AND2_1856(.VSS(VSS),.VDD(VDD),.Y(g19737),.A(g4363),.B(g17582));
  AND2 AND2_1857(.VSS(VSS),.VDD(VDD),.Y(g19738),.A(g4366),.B(g17585));
  AND2 AND2_1858(.VSS(VSS),.VDD(VDD),.Y(g19739),.A(g4369),.B(g17588));
  AND2 AND2_1859(.VSS(VSS),.VDD(VDD),.Y(g19741),.A(g1339),.B(g18856));
  AND2 AND2_1860(.VSS(VSS),.VDD(VDD),.Y(g19742),.A(g1332),.B(g18857));
  AND2 AND2_1861(.VSS(VSS),.VDD(VDD),.Y(g19743),.A(g1346),.B(g18858));
  AND2 AND2_1862(.VSS(VSS),.VDD(VDD),.Y(g19744),.A(g17927),.B(g16040));
  AND2 AND2_1863(.VSS(VSS),.VDD(VDD),.Y(g19745),.A(g4389),.B(g17601));
  AND2 AND2_1864(.VSS(VSS),.VDD(VDD),.Y(g19746),.A(g4392),.B(g17604));
  AND2 AND2_1865(.VSS(VSS),.VDD(VDD),.Y(g19747),.A(g4395),.B(g17607));
  AND2 AND2_1866(.VSS(VSS),.VDD(VDD),.Y(g19748),.A(g4398),.B(g17610));
  AND2 AND2_1867(.VSS(VSS),.VDD(VDD),.Y(g19752),.A(g2013),.B(g18859));
  AND2 AND2_1868(.VSS(VSS),.VDD(VDD),.Y(g19753),.A(g2033),.B(g18860));
  AND2 AND2_1869(.VSS(VSS),.VDD(VDD),.Y(g19754),.A(g2026),.B(g18861));
  AND2 AND2_1870(.VSS(VSS),.VDD(VDD),.Y(g19755),.A(g4421),.B(g17621));
  AND2 AND2_1871(.VSS(VSS),.VDD(VDD),.Y(g19756),.A(g4424),.B(g17624));
  AND2 AND2_1872(.VSS(VSS),.VDD(VDD),.Y(g19757),.A(g4427),.B(g17627));
  AND2 AND2_1873(.VSS(VSS),.VDD(VDD),.Y(g19758),.A(g2714),.B(g18862));
  AND2 AND2_1874(.VSS(VSS),.VDD(VDD),.Y(g19759),.A(g2707),.B(g18863));
  AND2 AND2_1875(.VSS(VSS),.VDD(VDD),.Y(g19760),.A(g2727),.B(g18864));
  AND2 AND2_1876(.VSS(VSS),.VDD(VDD),.Y(g19761),.A(g2766),.B(g18865));
  AND2 AND2_1877(.VSS(VSS),.VDD(VDD),.Y(g19764),.A(g4453),.B(g17637));
  AND2 AND2_1878(.VSS(VSS),.VDD(VDD),.Y(g19765),.A(g660),.B(g18870));
  AND2 AND2_1879(.VSS(VSS),.VDD(VDD),.Y(g19766),.A(g672),.B(g18871));
  AND2 AND2_1880(.VSS(VSS),.VDD(VDD),.Y(g19767),.A(g666),.B(g18872));
  AND2 AND2_1881(.VSS(VSS),.VDD(VDD),.Y(g19768),.A(g17815),.B(g16054));
  AND2 AND2_1882(.VSS(VSS),.VDD(VDD),.Y(g19769),.A(g17903),.B(g16055));
  AND2 AND2_1883(.VSS(VSS),.VDD(VDD),.Y(g19770),.A(g4498),.B(g17655));
  AND2 AND2_1884(.VSS(VSS),.VDD(VDD),.Y(g19771),.A(g4501),.B(g17658));
  AND2 AND2_1885(.VSS(VSS),.VDD(VDD),.Y(g19772),.A(g4504),.B(g17661));
  AND2 AND2_1886(.VSS(VSS),.VDD(VDD),.Y(g19773),.A(g1339),.B(g17670));
  AND2 AND2_1887(.VSS(VSS),.VDD(VDD),.Y(g19774),.A(g1332),.B(g18874));
  AND2 AND2_1888(.VSS(VSS),.VDD(VDD),.Y(g19775),.A(g1346),.B(g18875));
  AND2 AND2_1889(.VSS(VSS),.VDD(VDD),.Y(g19776),.A(g1358),.B(g18876));
  AND2 AND2_1890(.VSS(VSS),.VDD(VDD),.Y(g19777),.A(g17927),.B(g16056));
  AND2 AND2_1891(.VSS(VSS),.VDD(VDD),.Y(g19778),.A(g18014),.B(g16057));
  AND2 AND2_1892(.VSS(VSS),.VDD(VDD),.Y(g19779),.A(g4529),.B(g17676));
  AND2 AND2_1893(.VSS(VSS),.VDD(VDD),.Y(g19780),.A(g4532),.B(g17679));
  AND2 AND2_1894(.VSS(VSS),.VDD(VDD),.Y(g19781),.A(g4535),.B(g17682));
  AND2 AND2_1895(.VSS(VSS),.VDD(VDD),.Y(g19782),.A(g4538),.B(g17685));
  AND2 AND2_1896(.VSS(VSS),.VDD(VDD),.Y(g19784),.A(g2033),.B(g18877));
  AND2 AND2_1897(.VSS(VSS),.VDD(VDD),.Y(g19785),.A(g2026),.B(g18878));
  AND2 AND2_1898(.VSS(VSS),.VDD(VDD),.Y(g19786),.A(g2040),.B(g18879));
  AND2 AND2_1899(.VSS(VSS),.VDD(VDD),.Y(g19787),.A(g18038),.B(g16062));
  AND2 AND2_1900(.VSS(VSS),.VDD(VDD),.Y(g19788),.A(g4558),.B(g17698));
  AND2 AND2_1901(.VSS(VSS),.VDD(VDD),.Y(g19789),.A(g4561),.B(g17701));
  AND2 AND2_1902(.VSS(VSS),.VDD(VDD),.Y(g19790),.A(g4564),.B(g17704));
  AND2 AND2_1903(.VSS(VSS),.VDD(VDD),.Y(g19791),.A(g4567),.B(g17707));
  AND2 AND2_1904(.VSS(VSS),.VDD(VDD),.Y(g19795),.A(g2707),.B(g18880));
  AND2 AND2_1905(.VSS(VSS),.VDD(VDD),.Y(g19796),.A(g2727),.B(g18881));
  AND2 AND2_1906(.VSS(VSS),.VDD(VDD),.Y(g19797),.A(g2720),.B(g18882));
  AND3 AND3_62(.VSS(VSS),.VDD(VDD),.Y(I26240),.A(g18174),.B(g18341),.C(g17974));
  AND3 AND3_63(.VSS(VSS),.VDD(VDD),.Y(g19799),.A(g17640),.B(g18074),.C(I26240));
  AND2 AND2_1907(.VSS(VSS),.VDD(VDD),.Y(g19802),.A(g672),.B(g18891));
  AND2 AND2_1908(.VSS(VSS),.VDD(VDD),.Y(g19803),.A(g666),.B(g18892));
  AND2 AND2_1909(.VSS(VSS),.VDD(VDD),.Y(g19804),.A(g679),.B(g18893));
  AND2 AND2_1910(.VSS(VSS),.VDD(VDD),.Y(g19805),.A(g17903),.B(g16088));
  AND2 AND2_1911(.VSS(VSS),.VDD(VDD),.Y(g19806),.A(g4629),.B(g17738));
  AND2 AND2_1912(.VSS(VSS),.VDD(VDD),.Y(g19807),.A(g1346),.B(g18896));
  AND2 AND2_1913(.VSS(VSS),.VDD(VDD),.Y(g19808),.A(g1358),.B(g18897));
  AND2 AND2_1914(.VSS(VSS),.VDD(VDD),.Y(g19809),.A(g1352),.B(g18898));
  AND2 AND2_1915(.VSS(VSS),.VDD(VDD),.Y(g19810),.A(g17927),.B(g16090));
  AND2 AND2_1916(.VSS(VSS),.VDD(VDD),.Y(g19811),.A(g18014),.B(g16091));
  AND2 AND2_1917(.VSS(VSS),.VDD(VDD),.Y(g19812),.A(g4674),.B(g17755));
  AND2 AND2_1918(.VSS(VSS),.VDD(VDD),.Y(g19813),.A(g4677),.B(g17758));
  AND2 AND2_1919(.VSS(VSS),.VDD(VDD),.Y(g19814),.A(g4680),.B(g17761));
  AND2 AND2_1920(.VSS(VSS),.VDD(VDD),.Y(g19815),.A(g2033),.B(g17770));
  AND2 AND2_1921(.VSS(VSS),.VDD(VDD),.Y(g19816),.A(g2026),.B(g18900));
  AND2 AND2_1922(.VSS(VSS),.VDD(VDD),.Y(g19817),.A(g2040),.B(g18901));
  AND2 AND2_1923(.VSS(VSS),.VDD(VDD),.Y(g19818),.A(g2052),.B(g18902));
  AND2 AND2_1924(.VSS(VSS),.VDD(VDD),.Y(g19819),.A(g18038),.B(g16092));
  AND2 AND2_1925(.VSS(VSS),.VDD(VDD),.Y(g19820),.A(g18131),.B(g16093));
  AND2 AND2_1926(.VSS(VSS),.VDD(VDD),.Y(g19821),.A(g4705),.B(g17776));
  AND2 AND2_1927(.VSS(VSS),.VDD(VDD),.Y(g19822),.A(g4708),.B(g17779));
  AND2 AND2_1928(.VSS(VSS),.VDD(VDD),.Y(g19823),.A(g4711),.B(g17782));
  AND2 AND2_1929(.VSS(VSS),.VDD(VDD),.Y(g19824),.A(g4714),.B(g17785));
  AND2 AND2_1930(.VSS(VSS),.VDD(VDD),.Y(g19826),.A(g2727),.B(g18903));
  AND2 AND2_1931(.VSS(VSS),.VDD(VDD),.Y(g19827),.A(g2720),.B(g18904));
  AND2 AND2_1932(.VSS(VSS),.VDD(VDD),.Y(g19828),.A(g2734),.B(g18905));
  AND2 AND2_1933(.VSS(VSS),.VDD(VDD),.Y(g19829),.A(g18155),.B(g16098));
  AND2 AND2_1934(.VSS(VSS),.VDD(VDD),.Y(g19836),.A(g7143),.B(g18908));
  AND2 AND2_1935(.VSS(VSS),.VDD(VDD),.Y(g19837),.A(g6901),.B(g17799));
  AND2 AND2_1936(.VSS(VSS),.VDD(VDD),.Y(g19839),.A(g666),.B(g18909));
  AND2 AND2_1937(.VSS(VSS),.VDD(VDD),.Y(g19840),.A(g679),.B(g18910));
  AND2 AND2_1938(.VSS(VSS),.VDD(VDD),.Y(g19841),.A(g686),.B(g18911));
  AND3 AND3_64(.VSS(VSS),.VDD(VDD),.Y(I26282),.A(g18188),.B(g18089),.C(g17991));
  AND3 AND3_65(.VSS(VSS),.VDD(VDD),.Y(g19842),.A(g14525),.B(g13922),.C(I26282));
  AND3 AND3_66(.VSS(VSS),.VDD(VDD),.Y(I26285),.A(g18281),.B(g18436),.C(g18091));
  AND3 AND3_67(.VSS(VSS),.VDD(VDD),.Y(g19843),.A(g17741),.B(g18190),.C(I26285));
  AND2 AND2_1939(.VSS(VSS),.VDD(VDD),.Y(g19846),.A(g1358),.B(g18914));
  AND2 AND2_1940(.VSS(VSS),.VDD(VDD),.Y(g19847),.A(g1352),.B(g18915));
  AND2 AND2_1941(.VSS(VSS),.VDD(VDD),.Y(g19848),.A(g1365),.B(g18916));
  AND2 AND2_1942(.VSS(VSS),.VDD(VDD),.Y(g19849),.A(g18014),.B(g16126));
  AND2 AND2_1943(.VSS(VSS),.VDD(VDD),.Y(g19850),.A(g4806),.B(g17839));
  AND2 AND2_1944(.VSS(VSS),.VDD(VDD),.Y(g19851),.A(g2040),.B(g18919));
  AND2 AND2_1945(.VSS(VSS),.VDD(VDD),.Y(g19852),.A(g2052),.B(g18920));
  AND2 AND2_1946(.VSS(VSS),.VDD(VDD),.Y(g19853),.A(g2046),.B(g18921));
  AND2 AND2_1947(.VSS(VSS),.VDD(VDD),.Y(g19854),.A(g18038),.B(g16128));
  AND2 AND2_1948(.VSS(VSS),.VDD(VDD),.Y(g19855),.A(g18131),.B(g16129));
  AND2 AND2_1949(.VSS(VSS),.VDD(VDD),.Y(g19856),.A(g4851),.B(g17856));
  AND2 AND2_1950(.VSS(VSS),.VDD(VDD),.Y(g19857),.A(g4854),.B(g17859));
  AND2 AND2_1951(.VSS(VSS),.VDD(VDD),.Y(g19858),.A(g4857),.B(g17862));
  AND2 AND2_1952(.VSS(VSS),.VDD(VDD),.Y(g19859),.A(g2727),.B(g17871));
  AND2 AND2_1953(.VSS(VSS),.VDD(VDD),.Y(g19860),.A(g2720),.B(g18923));
  AND2 AND2_1954(.VSS(VSS),.VDD(VDD),.Y(g19861),.A(g2734),.B(g18924));
  AND2 AND2_1955(.VSS(VSS),.VDD(VDD),.Y(g19862),.A(g2746),.B(g18925));
  AND2 AND2_1956(.VSS(VSS),.VDD(VDD),.Y(g19863),.A(g18155),.B(g16130));
  AND2 AND2_1957(.VSS(VSS),.VDD(VDD),.Y(g19864),.A(g18247),.B(g16131));
  AND3 AND3_68(.VSS(VSS),.VDD(VDD),.Y(g19868),.A(g16498),.B(g16867),.C(g19001));
  AND2 AND2_1958(.VSS(VSS),.VDD(VDD),.Y(g19869),.A(g679),.B(g18926));
  AND2 AND2_1959(.VSS(VSS),.VDD(VDD),.Y(g19870),.A(g686),.B(g18927));
  AND3 AND3_69(.VSS(VSS),.VDD(VDD),.Y(I26311),.A(g18353),.B(g13958),.C(g14011));
  AND3 AND3_70(.VSS(VSS),.VDD(VDD),.Y(g19871),.A(g14086),.B(g18275),.C(I26311));
  AND2 AND2_1960(.VSS(VSS),.VDD(VDD),.Y(g19872),.A(g1352),.B(g18928));
  AND2 AND2_1961(.VSS(VSS),.VDD(VDD),.Y(g19873),.A(g1365),.B(g18929));
  AND2 AND2_1962(.VSS(VSS),.VDD(VDD),.Y(g19874),.A(g1372),.B(g18930));
  AND3 AND3_71(.VSS(VSS),.VDD(VDD),.Y(I26317),.A(g18295),.B(g18205),.C(g18108));
  AND3 AND3_72(.VSS(VSS),.VDD(VDD),.Y(g19875),.A(g14580),.B(g13978),.C(I26317));
  AND3 AND3_73(.VSS(VSS),.VDD(VDD),.Y(I26320),.A(g18374),.B(g18509),.C(g18207));
  AND3 AND3_74(.VSS(VSS),.VDD(VDD),.Y(g19876),.A(g17842),.B(g18297),.C(I26320));
  AND2 AND2_1963(.VSS(VSS),.VDD(VDD),.Y(g19879),.A(g2052),.B(g18933));
  AND2 AND2_1964(.VSS(VSS),.VDD(VDD),.Y(g19880),.A(g2046),.B(g18934));
  AND2 AND2_1965(.VSS(VSS),.VDD(VDD),.Y(g19881),.A(g2059),.B(g18935));
  AND2 AND2_1966(.VSS(VSS),.VDD(VDD),.Y(g19882),.A(g18131),.B(g16177));
  AND2 AND2_1967(.VSS(VSS),.VDD(VDD),.Y(g19883),.A(g4982),.B(g17951));
  AND2 AND2_1968(.VSS(VSS),.VDD(VDD),.Y(g19884),.A(g2734),.B(g18938));
  AND2 AND2_1969(.VSS(VSS),.VDD(VDD),.Y(g19885),.A(g2746),.B(g18939));
  AND2 AND2_1970(.VSS(VSS),.VDD(VDD),.Y(g19886),.A(g2740),.B(g18940));
  AND2 AND2_1971(.VSS(VSS),.VDD(VDD),.Y(g19887),.A(g18155),.B(g16179));
  AND2 AND2_1972(.VSS(VSS),.VDD(VDD),.Y(g19888),.A(g18247),.B(g16180));
  AND2 AND2_1973(.VSS(VSS),.VDD(VDD),.Y(g19889),.A(g2912),.B(g18943));
  AND2 AND2_1974(.VSS(VSS),.VDD(VDD),.Y(g19895),.A(g686),.B(g18945));
  AND3 AND3_75(.VSS(VSS),.VDD(VDD),.Y(g19899),.A(g16520),.B(g16895),.C(g16507));
  AND2 AND2_1975(.VSS(VSS),.VDD(VDD),.Y(g19900),.A(g1365),.B(g18946));
  AND2 AND2_1976(.VSS(VSS),.VDD(VDD),.Y(g19901),.A(g1372),.B(g18947));
  AND3 AND3_76(.VSS(VSS),.VDD(VDD),.Y(I26348),.A(g18448),.B(g14028),.C(g14102));
  AND3 AND3_77(.VSS(VSS),.VDD(VDD),.Y(g19902),.A(g14201),.B(g18368),.C(I26348));
  AND2 AND2_1977(.VSS(VSS),.VDD(VDD),.Y(g19903),.A(g2046),.B(g18948));
  AND2 AND2_1978(.VSS(VSS),.VDD(VDD),.Y(g19904),.A(g2059),.B(g18949));
  AND2 AND2_1979(.VSS(VSS),.VDD(VDD),.Y(g19905),.A(g2066),.B(g18950));
  AND3 AND3_78(.VSS(VSS),.VDD(VDD),.Y(I26354),.A(g18388),.B(g18312),.C(g18224));
  AND3 AND3_79(.VSS(VSS),.VDD(VDD),.Y(g19906),.A(g14614),.B(g14048),.C(I26354));
  AND3 AND3_80(.VSS(VSS),.VDD(VDD),.Y(I26357),.A(g18469),.B(g18573),.C(g18314));
  AND3 AND3_81(.VSS(VSS),.VDD(VDD),.Y(g19907),.A(g17954),.B(g18390),.C(I26357));
  AND2 AND2_1980(.VSS(VSS),.VDD(VDD),.Y(g19910),.A(g2746),.B(g18953));
  AND2 AND2_1981(.VSS(VSS),.VDD(VDD),.Y(g19911),.A(g2740),.B(g18954));
  AND2 AND2_1982(.VSS(VSS),.VDD(VDD),.Y(g19912),.A(g2753),.B(g18955));
  AND2 AND2_1983(.VSS(VSS),.VDD(VDD),.Y(g19913),.A(g18247),.B(g16236));
  AND2 AND2_1984(.VSS(VSS),.VDD(VDD),.Y(g19914),.A(g3018),.B(g18958));
  AND2 AND2_1985(.VSS(VSS),.VDD(VDD),.Y(g19920),.A(g1372),.B(g18961));
  AND3 AND3_82(.VSS(VSS),.VDD(VDD),.Y(g19924),.A(g16551),.B(g16924),.C(g16529));
  AND2 AND2_1986(.VSS(VSS),.VDD(VDD),.Y(g19925),.A(g2059),.B(g18962));
  AND2 AND2_1987(.VSS(VSS),.VDD(VDD),.Y(g19926),.A(g2066),.B(g18963));
  AND3 AND3_83(.VSS(VSS),.VDD(VDD),.Y(I26377),.A(g18521),.B(g14119),.C(g14217));
  AND3 AND3_84(.VSS(VSS),.VDD(VDD),.Y(g19927),.A(g14316),.B(g18463),.C(I26377));
  AND2 AND2_1988(.VSS(VSS),.VDD(VDD),.Y(g19928),.A(g2740),.B(g18964));
  AND2 AND2_1989(.VSS(VSS),.VDD(VDD),.Y(g19929),.A(g2753),.B(g18965));
  AND2 AND2_1990(.VSS(VSS),.VDD(VDD),.Y(g19930),.A(g2760),.B(g18966));
  AND3 AND3_85(.VSS(VSS),.VDD(VDD),.Y(I26383),.A(g18483),.B(g18405),.C(g18331));
  AND3 AND3_86(.VSS(VSS),.VDD(VDD),.Y(g19931),.A(g14637),.B(g14139),.C(I26383));
  AND2 AND2_1991(.VSS(VSS),.VDD(VDD),.Y(g19932),.A(g2917),.B(g18166));
  AND2 AND2_1992(.VSS(VSS),.VDD(VDD),.Y(g19935),.A(g2066),.B(g18972));
  AND3 AND3_87(.VSS(VSS),.VDD(VDD),.Y(g19939),.A(g16583),.B(g16954),.C(g16560));
  AND2 AND2_1993(.VSS(VSS),.VDD(VDD),.Y(g19940),.A(g2753),.B(g18973));
  AND2 AND2_1994(.VSS(VSS),.VDD(VDD),.Y(g19941),.A(g2760),.B(g18974));
  AND3 AND3_88(.VSS(VSS),.VDD(VDD),.Y(I26396),.A(g18585),.B(g14234),.C(g14332));
  AND3 AND3_89(.VSS(VSS),.VDD(VDD),.Y(g19942),.A(g14438),.B(g18536),.C(I26396));
  AND2 AND2_1995(.VSS(VSS),.VDD(VDD),.Y(g19943),.A(g7562),.B(g18976));
  AND2 AND2_1996(.VSS(VSS),.VDD(VDD),.Y(g19944),.A(g3028),.B(g18258));
  AND2 AND2_1997(.VSS(VSS),.VDD(VDD),.Y(g19949),.A(g5293),.B(g18278));
  AND2 AND2_1998(.VSS(VSS),.VDD(VDD),.Y(g19952),.A(g2760),.B(g18987));
  AND2 AND2_1999(.VSS(VSS),.VDD(VDD),.Y(g19953),.A(g7566),.B(g18334));
  AND3 AND3_90(.VSS(VSS),.VDD(VDD),.Y(I26416),.A(g18553),.B(g18491),.C(g18431));
  AND3 AND3_91(.VSS(VSS),.VDD(VDD),.Y(g19970),.A(g18354),.B(g18276),.C(I26416));
  AND2 AND2_2000(.VSS(VSS),.VDD(VDD),.Y(g19971),.A(g5327),.B(g18355));
  AND2 AND2_2001(.VSS(VSS),.VDD(VDD),.Y(g19976),.A(g5330),.B(g18371));
  AND3 AND3_92(.VSS(VSS),.VDD(VDD),.Y(I26432),.A(g18277),.B(g18189),.C(g18090));
  AND3 AND3_93(.VSS(VSS),.VDD(VDD),.Y(g19982),.A(g17992),.B(g17913),.C(I26432));
  AND2 AND2_2002(.VSS(VSS),.VDD(VDD),.Y(g19983),.A(g5352),.B(g18432));
  AND3 AND3_94(.VSS(VSS),.VDD(VDD),.Y(I26440),.A(g18603),.B(g18555),.C(g18504));
  AND3 AND3_95(.VSS(VSS),.VDD(VDD),.Y(g20000),.A(g18449),.B(g18369),.C(I26440));
  AND2 AND2_2003(.VSS(VSS),.VDD(VDD),.Y(g20001),.A(g5355),.B(g18450));
  AND2 AND2_2004(.VSS(VSS),.VDD(VDD),.Y(g20006),.A(g5358),.B(g18466));
  AND2 AND2_2005(.VSS(VSS),.VDD(VDD),.Y(g20011),.A(g18063),.B(g3113));
  AND2 AND2_2006(.VSS(VSS),.VDD(VDD),.Y(g20012),.A(g16804),.B(g3135));
  AND2 AND2_2007(.VSS(VSS),.VDD(VDD),.Y(g20013),.A(g17720),.B(g12848));
  AND2 AND2_2008(.VSS(VSS),.VDD(VDD),.Y(g20014),.A(g7615),.B(g16749));
  AND3 AND3_96(.VSS(VSS),.VDD(VDD),.Y(I26464),.A(g18370),.B(g18296),.C(g18206));
  AND3 AND3_97(.VSS(VSS),.VDD(VDD),.Y(g20020),.A(g18109),.B(g18024),.C(I26464));
  AND2 AND2_2009(.VSS(VSS),.VDD(VDD),.Y(g20021),.A(g5369),.B(g18505));
  AND3 AND3_98(.VSS(VSS),.VDD(VDD),.Y(I26472),.A(g18635),.B(g18605),.C(g18568));
  AND3 AND3_99(.VSS(VSS),.VDD(VDD),.Y(g20038),.A(g18522),.B(g18464),.C(I26472));
  AND2 AND2_2010(.VSS(VSS),.VDD(VDD),.Y(g20039),.A(g5372),.B(g18523));
  AND2 AND2_2011(.VSS(VSS),.VDD(VDD),.Y(g20044),.A(g5375),.B(g18539));
  AND2 AND2_2012(.VSS(VSS),.VDD(VDD),.Y(g20048),.A(g16749),.B(g3127));
  AND2 AND2_2013(.VSS(VSS),.VDD(VDD),.Y(g20049),.A(g17878),.B(g3155));
  AND2 AND2_2014(.VSS(VSS),.VDD(VDD),.Y(g20050),.A(g18070),.B(g3161));
  AND2 AND2_2015(.VSS(VSS),.VDD(VDD),.Y(g20051),.A(g18063),.B(g3114));
  AND2 AND2_2016(.VSS(VSS),.VDD(VDD),.Y(g20052),.A(g16804),.B(g3134));
  AND2 AND2_2017(.VSS(VSS),.VDD(VDD),.Y(g20053),.A(g17720),.B(g12875));
  AND3 AND3_100(.VSS(VSS),.VDD(VDD),.Y(I26500),.A(g18465),.B(g18389),.C(g18313));
  AND3 AND3_101(.VSS(VSS),.VDD(VDD),.Y(g20062),.A(g18225),.B(g18141),.C(I26500));
  AND2 AND2_2018(.VSS(VSS),.VDD(VDD),.Y(g20063),.A(g5382),.B(g18569));
  AND3 AND3_102(.VSS(VSS),.VDD(VDD),.Y(I26508),.A(g18644),.B(g18637),.C(g18618));
  AND3 AND3_103(.VSS(VSS),.VDD(VDD),.Y(g20080),.A(g18586),.B(g18537),.C(I26508));
  AND2 AND2_2019(.VSS(VSS),.VDD(VDD),.Y(g20081),.A(g5385),.B(g18587));
  AND2 AND2_2020(.VSS(VSS),.VDD(VDD),.Y(g20084),.A(g17969),.B(g3158));
  AND2 AND2_2021(.VSS(VSS),.VDD(VDD),.Y(g20085),.A(g18170),.B(g3164));
  AND2 AND2_2022(.VSS(VSS),.VDD(VDD),.Y(g20086),.A(g18337),.B(g3170));
  AND2 AND2_2023(.VSS(VSS),.VDD(VDD),.Y(g20087),.A(g16749),.B(g7574));
  AND2 AND2_2024(.VSS(VSS),.VDD(VDD),.Y(g20088),.A(g16836),.B(g3147));
  AND2 AND2_2025(.VSS(VSS),.VDD(VDD),.Y(g20089),.A(g17969),.B(g9160));
  AND2 AND2_2026(.VSS(VSS),.VDD(VDD),.Y(g20090),.A(g18063),.B(g3120));
  AND2 AND2_2027(.VSS(VSS),.VDD(VDD),.Y(g20091),.A(g16804),.B(g3136));
  AND2 AND2_2028(.VSS(VSS),.VDD(VDD),.Y(g20092),.A(g16749),.B(g7603));
  AND3 AND3_104(.VSS(VSS),.VDD(VDD),.Y(I26525),.A(g18656),.B(g18670),.C(g18692));
  AND4 AND4_61(.VSS(VSS),.VDD(VDD),.Y(g20093),.A(g13657),.B(g13677),.C(g13750),.D(I26525));
  AND3 AND3_105(.VSS(VSS),.VDD(VDD),.Y(I26528),.A(g18656),.B(g14837),.C(g13657));
  AND3 AND3_106(.VSS(VSS),.VDD(VDD),.Y(g20094),.A(g13677),.B(g13706),.C(I26528));
  AND3 AND3_107(.VSS(VSS),.VDD(VDD),.Y(I26541),.A(g18538),.B(g18484),.C(g18406));
  AND3 AND3_108(.VSS(VSS),.VDD(VDD),.Y(g20103),.A(g18332),.B(g18257),.C(I26541));
  AND2 AND2_2029(.VSS(VSS),.VDD(VDD),.Y(g20104),.A(g5391),.B(g18619));
  AND2 AND2_2030(.VSS(VSS),.VDD(VDD),.Y(g20106),.A(g18261),.B(g3167));
  AND2 AND2_2031(.VSS(VSS),.VDD(VDD),.Y(g20107),.A(g18415),.B(g3173));
  AND2 AND2_2032(.VSS(VSS),.VDD(VDD),.Y(g20108),.A(g18543),.B(g3179));
  AND2 AND2_2033(.VSS(VSS),.VDD(VDD),.Y(g20109),.A(g17878),.B(g9504));
  AND2 AND2_2034(.VSS(VSS),.VDD(VDD),.Y(g20110),.A(g18070),.B(g9286));
  AND2 AND2_2035(.VSS(VSS),.VDD(VDD),.Y(g20111),.A(g18261),.B(g9884));
  AND2 AND2_2036(.VSS(VSS),.VDD(VDD),.Y(g20112),.A(g16749),.B(g3132));
  AND2 AND2_2037(.VSS(VSS),.VDD(VDD),.Y(g20113),.A(g16836),.B(g3142));
  AND2 AND2_2038(.VSS(VSS),.VDD(VDD),.Y(g20114),.A(g17969),.B(g9755));
  AND2 AND2_2039(.VSS(VSS),.VDD(VDD),.Y(g20115),.A(g16804),.B(g3139));
  AND3 AND3_109(.VSS(VSS),.VDD(VDD),.Y(I26558),.A(g14776),.B(g18670),.C(g18720));
  AND4 AND4_62(.VSS(VSS),.VDD(VDD),.Y(g20116),.A(g16142),.B(g13677),.C(g13706),.D(I26558));
  AND3 AND3_110(.VSS(VSS),.VDD(VDD),.Y(I26561),.A(g14776),.B(g18720),.C(g13657));
  AND3 AND3_111(.VSS(VSS),.VDD(VDD),.Y(g20117),.A(g16189),.B(g13706),.C(I26561));
  AND3 AND3_112(.VSS(VSS),.VDD(VDD),.Y(I26564),.A(g18679),.B(g18699),.C(g18728));
  AND4 AND4_63(.VSS(VSS),.VDD(VDD),.Y(g20118),.A(g13687),.B(g13714),.C(g13791),.D(I26564));
  AND3 AND3_113(.VSS(VSS),.VDD(VDD),.Y(I26567),.A(g18679),.B(g14910),.C(g13687));
  AND3 AND3_114(.VSS(VSS),.VDD(VDD),.Y(g20119),.A(g13714),.B(g13756),.C(I26567));
  AND2 AND2_2040(.VSS(VSS),.VDD(VDD),.Y(g20131),.A(g18486),.B(g3176));
  AND2 AND2_2041(.VSS(VSS),.VDD(VDD),.Y(g20132),.A(g18593),.B(g3182));
  AND2 AND2_2042(.VSS(VSS),.VDD(VDD),.Y(g20133),.A(g18170),.B(g9505));
  AND2 AND2_2043(.VSS(VSS),.VDD(VDD),.Y(g20134),.A(g18337),.B(g9506));
  AND2 AND2_2044(.VSS(VSS),.VDD(VDD),.Y(g20135),.A(g18486),.B(g9885));
  AND2 AND2_2045(.VSS(VSS),.VDD(VDD),.Y(g20136),.A(g17878),.B(g9423));
  AND2 AND2_2046(.VSS(VSS),.VDD(VDD),.Y(g20137),.A(g18070),.B(g9226));
  AND2 AND2_2047(.VSS(VSS),.VDD(VDD),.Y(g20138),.A(g18261),.B(g9756));
  AND2 AND2_2048(.VSS(VSS),.VDD(VDD),.Y(g20139),.A(g16836),.B(g3151));
  AND3 AND3_115(.VSS(VSS),.VDD(VDD),.Y(g20144),.A(g16679),.B(g16884),.C(g16665));
  AND4 AND4_64(.VSS(VSS),.VDD(VDD),.Y(g20145),.A(g14776),.B(g18670),.C(g16142),.D(g16189));
  AND3 AND3_116(.VSS(VSS),.VDD(VDD),.Y(I26590),.A(g14811),.B(g18699),.C(g18758));
  AND4 AND4_65(.VSS(VSS),.VDD(VDD),.Y(g20146),.A(g16201),.B(g13714),.C(g13756),.D(I26590));
  AND3 AND3_117(.VSS(VSS),.VDD(VDD),.Y(I26593),.A(g14811),.B(g18758),.C(g13687));
  AND3 AND3_118(.VSS(VSS),.VDD(VDD),.Y(g20147),.A(g16254),.B(g13756),.C(I26593));
  AND3 AND3_119(.VSS(VSS),.VDD(VDD),.Y(I26596),.A(g18708),.B(g18735),.C(g18765));
  AND4 AND4_66(.VSS(VSS),.VDD(VDD),.Y(g20148),.A(g13724),.B(g13764),.C(g13819),.D(I26596));
  AND3 AND3_120(.VSS(VSS),.VDD(VDD),.Y(I26599),.A(g18708),.B(g14991),.C(g13724));
  AND3 AND3_121(.VSS(VSS),.VDD(VDD),.Y(g20149),.A(g13764),.B(g13797),.C(I26599));
  AND2 AND2_2049(.VSS(VSS),.VDD(VDD),.Y(g20156),.A(g16809),.B(g3185));
  AND2 AND2_2050(.VSS(VSS),.VDD(VDD),.Y(g20157),.A(g18415),.B(g9287));
  AND2 AND2_2051(.VSS(VSS),.VDD(VDD),.Y(g20158),.A(g18543),.B(g9886));
  AND2 AND2_2052(.VSS(VSS),.VDD(VDD),.Y(g20159),.A(g16809),.B(g9288));
  AND2 AND2_2053(.VSS(VSS),.VDD(VDD),.Y(g20160),.A(g18170),.B(g9424));
  AND2 AND2_2054(.VSS(VSS),.VDD(VDD),.Y(g20161),.A(g18337),.B(g9426));
  AND2 AND2_2055(.VSS(VSS),.VDD(VDD),.Y(g20162),.A(g18486),.B(g9757));
  AND3 AND3_122(.VSS(VSS),.VDD(VDD),.Y(I26615),.A(g14797),.B(g18692),.C(g13657));
  AND3 AND3_123(.VSS(VSS),.VDD(VDD),.Y(g20177),.A(g13677),.B(g13750),.C(I26615));
  AND3 AND3_124(.VSS(VSS),.VDD(VDD),.Y(g20182),.A(g16705),.B(g16913),.C(g16686));
  AND4 AND4_67(.VSS(VSS),.VDD(VDD),.Y(g20183),.A(g14811),.B(g18699),.C(g16201),.D(g16254));
  AND3 AND3_125(.VSS(VSS),.VDD(VDD),.Y(I26621),.A(g14863),.B(g18735),.C(g18789));
  AND4 AND4_68(.VSS(VSS),.VDD(VDD),.Y(g20184),.A(g16266),.B(g13764),.C(g13797),.D(I26621));
  AND3 AND3_126(.VSS(VSS),.VDD(VDD),.Y(I26624),.A(g14863),.B(g18789),.C(g13724));
  AND3 AND3_127(.VSS(VSS),.VDD(VDD),.Y(g20185),.A(g16313),.B(g13797),.C(I26624));
  AND3 AND3_128(.VSS(VSS),.VDD(VDD),.Y(I26627),.A(g18744),.B(g18772),.C(g18796));
  AND4 AND4_69(.VSS(VSS),.VDD(VDD),.Y(g20186),.A(g13774),.B(g13805),.C(g13840),.D(I26627));
  AND3 AND3_129(.VSS(VSS),.VDD(VDD),.Y(I26630),.A(g18744),.B(g15080),.C(g13774));
  AND3 AND3_130(.VSS(VSS),.VDD(VDD),.Y(g20187),.A(g13805),.B(g13825),.C(I26630));
  AND2 AND2_2056(.VSS(VSS),.VDD(VDD),.Y(g20188),.A(g18593),.B(g9425));
  AND2 AND2_2057(.VSS(VSS),.VDD(VDD),.Y(g20189),.A(g16825),.B(g9289));
  AND2 AND2_2058(.VSS(VSS),.VDD(VDD),.Y(g20190),.A(g18415),.B(g9227));
  AND2 AND2_2059(.VSS(VSS),.VDD(VDD),.Y(g20191),.A(g18543),.B(g9758));
  AND2 AND2_2060(.VSS(VSS),.VDD(VDD),.Y(g20192),.A(g16809),.B(g9228));
  AND3 AND3_131(.VSS(VSS),.VDD(VDD),.Y(I26639),.A(g18656),.B(g18670),.C(g16142));
  AND3 AND3_132(.VSS(VSS),.VDD(VDD),.Y(g20197),.A(g13677),.B(g13706),.C(I26639));
  AND3 AND3_133(.VSS(VSS),.VDD(VDD),.Y(I26645),.A(g14849),.B(g18728),.C(g13687));
  AND3 AND3_134(.VSS(VSS),.VDD(VDD),.Y(g20211),.A(g13714),.B(g13791),.C(I26645));
  AND3 AND3_135(.VSS(VSS),.VDD(VDD),.Y(g20216),.A(g16736),.B(g16943),.C(g16712));
  AND4 AND4_70(.VSS(VSS),.VDD(VDD),.Y(g20217),.A(g14863),.B(g18735),.C(g16266),.D(g16313));
  AND3 AND3_136(.VSS(VSS),.VDD(VDD),.Y(I26651),.A(g14936),.B(g18772),.C(g18815));
  AND4 AND4_71(.VSS(VSS),.VDD(VDD),.Y(g20218),.A(g16325),.B(g13805),.C(g13825),.D(I26651));
  AND3 AND3_137(.VSS(VSS),.VDD(VDD),.Y(I26654),.A(g14936),.B(g18815),.C(g13774));
  AND3 AND3_138(.VSS(VSS),.VDD(VDD),.Y(g20219),.A(g16371),.B(g13825),.C(I26654));
  AND2 AND2_2061(.VSS(VSS),.VDD(VDD),.Y(g20220),.A(g18593),.B(g9355));
  AND2 AND2_2062(.VSS(VSS),.VDD(VDD),.Y(g20221),.A(g16825),.B(g10099));
  AND4 AND4_72(.VSS(VSS),.VDD(VDD),.Y(g20222),.A(g18656),.B(g18720),.C(g13657),.D(g16293));
  AND3 AND3_139(.VSS(VSS),.VDD(VDD),.Y(I26661),.A(g18679),.B(g18699),.C(g16201));
  AND3 AND3_140(.VSS(VSS),.VDD(VDD),.Y(g20227),.A(g13714),.B(g13756),.C(I26661));
  AND3 AND3_141(.VSS(VSS),.VDD(VDD),.Y(I26667),.A(g14922),.B(g18765),.C(g13724));
  AND3 AND3_142(.VSS(VSS),.VDD(VDD),.Y(g20241),.A(g13764),.B(g13819),.C(I26667));
  AND3 AND3_143(.VSS(VSS),.VDD(VDD),.Y(g20246),.A(g16778),.B(g16974),.C(g16743));
  AND4 AND4_73(.VSS(VSS),.VDD(VDD),.Y(g20247),.A(g14936),.B(g18772),.C(g16325),.D(g16371));
  AND3 AND3_144(.VSS(VSS),.VDD(VDD),.Y(g20248),.A(g18656),.B(g14837),.C(g16293));
  AND4 AND4_74(.VSS(VSS),.VDD(VDD),.Y(g20249),.A(g18679),.B(g18758),.C(g13687),.D(g16351));
  AND3 AND3_145(.VSS(VSS),.VDD(VDD),.Y(I26676),.A(g18708),.B(g18735),.C(g16266));
  AND3 AND3_146(.VSS(VSS),.VDD(VDD),.Y(g20254),.A(g13764),.B(g13797),.C(I26676));
  AND3 AND3_147(.VSS(VSS),.VDD(VDD),.Y(I26682),.A(g15003),.B(g18796),.C(g13774));
  AND3 AND3_148(.VSS(VSS),.VDD(VDD),.Y(g20268),.A(g13805),.B(g13840),.C(I26682));
  AND4 AND4_75(.VSS(VSS),.VDD(VDD),.Y(g20270),.A(g14797),.B(g18692),.C(g13657),.D(g16243));
  AND3 AND3_149(.VSS(VSS),.VDD(VDD),.Y(g20271),.A(g18679),.B(g14910),.C(g16351));
  AND4 AND4_76(.VSS(VSS),.VDD(VDD),.Y(g20272),.A(g18708),.B(g18789),.C(g13724),.D(g16395));
  AND3 AND3_150(.VSS(VSS),.VDD(VDD),.Y(I26690),.A(g18744),.B(g18772),.C(g16325));
  AND3 AND3_151(.VSS(VSS),.VDD(VDD),.Y(g20277),.A(g13805),.B(g13825),.C(I26690));
  AND3 AND3_152(.VSS(VSS),.VDD(VDD),.Y(I26695),.A(g18670),.B(g18692),.C(g16142));
  AND3 AND3_153(.VSS(VSS),.VDD(VDD),.Y(g20280),.A(g13677),.B(g16243),.C(I26695));
  AND4 AND4_77(.VSS(VSS),.VDD(VDD),.Y(g20282),.A(g14849),.B(g18728),.C(g13687),.D(g16302));
  AND3 AND3_154(.VSS(VSS),.VDD(VDD),.Y(g20283),.A(g18708),.B(g14991),.C(g16395));
  AND4 AND4_78(.VSS(VSS),.VDD(VDD),.Y(g20284),.A(g18744),.B(g18815),.C(g13774),.D(g16433));
  AND2 AND2_2063(.VSS(VSS),.VDD(VDD),.Y(g20285),.A(g16846),.B(g8103));
  AND3 AND3_155(.VSS(VSS),.VDD(VDD),.Y(I26708),.A(g18699),.B(g18728),.C(g16201));
  AND3 AND3_156(.VSS(VSS),.VDD(VDD),.Y(g20291),.A(g13714),.B(g16302),.C(I26708));
  AND4 AND4_79(.VSS(VSS),.VDD(VDD),.Y(g20293),.A(g14922),.B(g18765),.C(g13724),.D(g16360));
  AND3 AND3_157(.VSS(VSS),.VDD(VDD),.Y(g20294),.A(g18744),.B(g15080),.C(g16433));
  AND3 AND3_158(.VSS(VSS),.VDD(VDD),.Y(I26726),.A(g18735),.B(g18765),.C(g16266));
  AND3 AND3_159(.VSS(VSS),.VDD(VDD),.Y(g20307),.A(g13764),.B(g16360),.C(I26726));
  AND4 AND4_80(.VSS(VSS),.VDD(VDD),.Y(g20309),.A(g15003),.B(g18796),.C(g13774),.D(g16404));
  AND3 AND3_160(.VSS(VSS),.VDD(VDD),.Y(I26745),.A(g18772),.B(g18796),.C(g16325));
  AND3 AND3_161(.VSS(VSS),.VDD(VDD),.Y(g20326),.A(g13805),.B(g16404),.C(I26745));
  AND2 AND2_2064(.VSS(VSS),.VDD(VDD),.Y(g20460),.A(g17351),.B(g13644));
  AND2 AND2_2065(.VSS(VSS),.VDD(VDD),.Y(g20472),.A(g17314),.B(g13669));
  AND2 AND2_2066(.VSS(VSS),.VDD(VDD),.Y(g20480),.A(g17313),.B(g11827));
  AND2 AND2_2067(.VSS(VSS),.VDD(VDD),.Y(g20486),.A(g17281),.B(g11859));
  AND2 AND2_2068(.VSS(VSS),.VDD(VDD),.Y(g20492),.A(g17258),.B(g11894));
  AND2 AND2_2069(.VSS(VSS),.VDD(VDD),.Y(g20499),.A(g17648),.B(g11933));
  AND2 AND2_2070(.VSS(VSS),.VDD(VDD),.Y(g20502),.A(g17566),.B(g11973));
  AND2 AND2_2071(.VSS(VSS),.VDD(VDD),.Y(g20503),.A(g17507),.B(g13817));
  AND2 AND2_2072(.VSS(VSS),.VDD(VDD),.Y(g20506),.A(g17499),.B(g12025));
  AND2 AND2_2073(.VSS(VSS),.VDD(VDD),.Y(g20512),.A(g17445),.B(g13836));
  AND2 AND2_2074(.VSS(VSS),.VDD(VDD),.Y(g20525),.A(g17394),.B(g13849));
  AND4 AND4_81(.VSS(VSS),.VDD(VDD),.Y(g20538),.A(g18656),.B(g14837),.C(g13657),.D(g16189));
  AND2 AND2_2075(.VSS(VSS),.VDD(VDD),.Y(g20640),.A(g4809),.B(g19064));
  AND2 AND2_2076(.VSS(VSS),.VDD(VDD),.Y(g20647),.A(g5888),.B(g19075));
  AND2 AND2_2077(.VSS(VSS),.VDD(VDD),.Y(g20665),.A(g4985),.B(g19081));
  AND2 AND2_2078(.VSS(VSS),.VDD(VDD),.Y(g20809),.A(g5712),.B(g19113));
  AND2 AND2_2079(.VSS(VSS),.VDD(VDD),.Y(g20826),.A(g5770),.B(g19118));
  AND2 AND2_2080(.VSS(VSS),.VDD(VDD),.Y(g20836),.A(g5829),.B(g19125));
  AND2 AND2_2081(.VSS(VSS),.VDD(VDD),.Y(g20840),.A(g5885),.B(g19132));
  AND3 AND3_162(.VSS(VSS),.VDD(VDD),.Y(g21049),.A(g20016),.B(g14079),.C(g14165));
  AND2 AND2_2082(.VSS(VSS),.VDD(VDD),.Y(g21067),.A(g20193),.B(g12030));
  AND3 AND3_163(.VSS(VSS),.VDD(VDD),.Y(g21068),.A(g20058),.B(g14194),.C(g14280));
  AND2 AND2_2083(.VSS(VSS),.VDD(VDD),.Y(g21077),.A(g20223),.B(g12094));
  AND3 AND3_164(.VSS(VSS),.VDD(VDD),.Y(g21078),.A(g20099),.B(g14309),.C(g14402));
  AND3 AND3_165(.VSS(VSS),.VDD(VDD),.Y(g21085),.A(g19484),.B(g14158),.C(g19001));
  AND2 AND2_2084(.VSS(VSS),.VDD(VDD),.Y(g21086),.A(g20193),.B(g12142));
  AND2 AND2_2085(.VSS(VSS),.VDD(VDD),.Y(g21091),.A(g20250),.B(g12166));
  AND3 AND3_166(.VSS(VSS),.VDD(VDD),.Y(g21092),.A(g20124),.B(g14431),.C(g14514));
  AND3 AND3_167(.VSS(VSS),.VDD(VDD),.Y(g21097),.A(g19505),.B(g14273),.C(g16507));
  AND2 AND2_2086(.VSS(VSS),.VDD(VDD),.Y(g21098),.A(g20223),.B(g12204));
  AND2 AND2_2087(.VSS(VSS),.VDD(VDD),.Y(g21103),.A(g20273),.B(g12228));
  AND3 AND3_168(.VSS(VSS),.VDD(VDD),.Y(g21107),.A(g19444),.B(g17893),.C(g14079));
  AND3 AND3_169(.VSS(VSS),.VDD(VDD),.Y(g21111),.A(g19524),.B(g14395),.C(g16529));
  AND2 AND2_2088(.VSS(VSS),.VDD(VDD),.Y(g21112),.A(g20250),.B(g12259));
  AND2 AND2_2089(.VSS(VSS),.VDD(VDD),.Y(g21121),.A(g20054),.B(g14244));
  AND2 AND2_2090(.VSS(VSS),.VDD(VDD),.Y(g21122),.A(g20140),.B(g12279));
  AND2 AND2_2091(.VSS(VSS),.VDD(VDD),.Y(g21123),.A(g19970),.B(g19982));
  AND3 AND3_170(.VSS(VSS),.VDD(VDD),.Y(g21124),.A(g19471),.B(g18004),.C(g14194));
  AND3 AND3_171(.VSS(VSS),.VDD(VDD),.Y(g21128),.A(g19534),.B(g14507),.C(g16560));
  AND2 AND2_2092(.VSS(VSS),.VDD(VDD),.Y(g21129),.A(g20273),.B(g12302));
  AND3 AND3_172(.VSS(VSS),.VDD(VDD),.Y(I27695),.A(g19318),.B(g19300),.C(g19286));
  AND3 AND3_173(.VSS(VSS),.VDD(VDD),.Y(g21136),.A(g19271),.B(g19261),.C(I27695));
  AND2 AND2_2093(.VSS(VSS),.VDD(VDD),.Y(g21137),.A(g5750),.B(g19272));
  AND2 AND2_2094(.VSS(VSS),.VDD(VDD),.Y(g21138),.A(g19484),.B(g14347));
  AND2 AND2_2095(.VSS(VSS),.VDD(VDD),.Y(g21140),.A(g20095),.B(g14366));
  AND2 AND2_2096(.VSS(VSS),.VDD(VDD),.Y(g21141),.A(g20178),.B(g12315));
  AND2 AND2_2097(.VSS(VSS),.VDD(VDD),.Y(g21142),.A(g20000),.B(g20020));
  AND3 AND3_174(.VSS(VSS),.VDD(VDD),.Y(g21143),.A(g19494),.B(g18121),.C(g14309));
  AND3 AND3_175(.VSS(VSS),.VDD(VDD),.Y(I27711),.A(g19262),.B(g19414),.C(g19386));
  AND3 AND3_176(.VSS(VSS),.VDD(VDD),.Y(g21152),.A(g19357),.B(g19334),.C(I27711));
  AND3 AND3_177(.VSS(VSS),.VDD(VDD),.Y(g21153),.A(g20054),.B(g16543),.C(g16501));
  AND2 AND2_2098(.VSS(VSS),.VDD(VDD),.Y(g21154),.A(g20193),.B(g12333));
  AND2 AND2_2099(.VSS(VSS),.VDD(VDD),.Y(g21155),.A(g20140),.B(g12336));
  AND3 AND3_178(.VSS(VSS),.VDD(VDD),.Y(I27717),.A(g19345),.B(g19321),.C(g19304));
  AND3 AND3_179(.VSS(VSS),.VDD(VDD),.Y(g21156),.A(g19290),.B(g19276),.C(I27717));
  AND2 AND2_2100(.VSS(VSS),.VDD(VDD),.Y(g21157),.A(g5809),.B(g19291));
  AND2 AND2_2101(.VSS(VSS),.VDD(VDD),.Y(g21158),.A(g19505),.B(g14459));
  AND2 AND2_2102(.VSS(VSS),.VDD(VDD),.Y(g21160),.A(g20120),.B(g14478));
  AND2 AND2_2103(.VSS(VSS),.VDD(VDD),.Y(g21161),.A(g20212),.B(g12343));
  AND2 AND2_2104(.VSS(VSS),.VDD(VDD),.Y(g21162),.A(g20038),.B(g20062));
  AND3 AND3_180(.VSS(VSS),.VDD(VDD),.Y(g21163),.A(g19515),.B(g18237),.C(g14431));
  AND3 AND3_181(.VSS(VSS),.VDD(VDD),.Y(I27733),.A(g19277),.B(g19451),.C(g19416));
  AND3 AND3_182(.VSS(VSS),.VDD(VDD),.Y(g21172),.A(g19389),.B(g19368),.C(I27733));
  AND3 AND3_183(.VSS(VSS),.VDD(VDD),.Y(g21173),.A(g20095),.B(g16575),.C(g16523));
  AND2 AND2_2105(.VSS(VSS),.VDD(VDD),.Y(g21174),.A(g20223),.B(g12363));
  AND2 AND2_2106(.VSS(VSS),.VDD(VDD),.Y(g21175),.A(g20178),.B(g12366));
  AND3 AND3_184(.VSS(VSS),.VDD(VDD),.Y(I27739),.A(g19379),.B(g19348),.C(g19325));
  AND3 AND3_185(.VSS(VSS),.VDD(VDD),.Y(g21176),.A(g19308),.B(g19295),.C(I27739));
  AND2 AND2_2107(.VSS(VSS),.VDD(VDD),.Y(g21177),.A(g5865),.B(g19309));
  AND2 AND2_2108(.VSS(VSS),.VDD(VDD),.Y(g21178),.A(g19524),.B(g14546));
  AND2 AND2_2109(.VSS(VSS),.VDD(VDD),.Y(g21180),.A(g20150),.B(g14565));
  AND2 AND2_2110(.VSS(VSS),.VDD(VDD),.Y(g21181),.A(g20242),.B(g12373));
  AND2 AND2_2111(.VSS(VSS),.VDD(VDD),.Y(g21182),.A(g20080),.B(g20103));
  AND2 AND2_2112(.VSS(VSS),.VDD(VDD),.Y(g21188),.A(g20140),.B(g12379));
  AND3 AND3_186(.VSS(VSS),.VDD(VDD),.Y(I27755),.A(g19296),.B(g19478),.C(g19453));
  AND3 AND3_187(.VSS(VSS),.VDD(VDD),.Y(g21192),.A(g19419),.B(g19400),.C(I27755));
  AND3 AND3_188(.VSS(VSS),.VDD(VDD),.Y(g21193),.A(g20120),.B(g16599),.C(g16554));
  AND2 AND2_2113(.VSS(VSS),.VDD(VDD),.Y(g21194),.A(g20250),.B(g12382));
  AND2 AND2_2114(.VSS(VSS),.VDD(VDD),.Y(g21195),.A(g20212),.B(g12385));
  AND3 AND3_189(.VSS(VSS),.VDD(VDD),.Y(I27761),.A(g19411),.B(g19382),.C(g19352));
  AND3 AND3_190(.VSS(VSS),.VDD(VDD),.Y(g21196),.A(g19329),.B(g19313),.C(I27761));
  AND2 AND2_2115(.VSS(VSS),.VDD(VDD),.Y(g21197),.A(g5912),.B(g19330));
  AND2 AND2_2116(.VSS(VSS),.VDD(VDD),.Y(g21198),.A(g19534),.B(g14601));
  AND2 AND2_2117(.VSS(VSS),.VDD(VDD),.Y(g21203),.A(g20178),.B(g12409));
  AND3 AND3_191(.VSS(VSS),.VDD(VDD),.Y(I27772),.A(g19314),.B(g19501),.C(g19480));
  AND3 AND3_192(.VSS(VSS),.VDD(VDD),.Y(g21207),.A(g19456),.B(g19430),.C(I27772));
  AND3 AND3_193(.VSS(VSS),.VDD(VDD),.Y(g21208),.A(g20150),.B(g16619),.C(g16586));
  AND2 AND2_2118(.VSS(VSS),.VDD(VDD),.Y(g21209),.A(g20273),.B(g12412));
  AND2 AND2_2119(.VSS(VSS),.VDD(VDD),.Y(g21210),.A(g20242),.B(g12415));
  AND2 AND2_2120(.VSS(VSS),.VDD(VDD),.Y(g21218),.A(g20212),.B(g12421));
  AND2 AND2_2121(.VSS(VSS),.VDD(VDD),.Y(g21226),.A(g20242),.B(g12426));
  AND3 AND3_194(.VSS(VSS),.VDD(VDD),.Y(g21229),.A(g19578),.B(g14797),.C(g16665));
  AND3 AND3_195(.VSS(VSS),.VDD(VDD),.Y(g21234),.A(g19608),.B(g14849),.C(g16686));
  AND3 AND3_196(.VSS(VSS),.VDD(VDD),.Y(g21243),.A(g19641),.B(g14922),.C(g16712));
  AND2 AND2_2122(.VSS(VSS),.VDD(VDD),.Y(g21245),.A(g20299),.B(g14837));
  AND3 AND3_197(.VSS(VSS),.VDD(VDD),.Y(g21251),.A(g19681),.B(g15003),.C(g16743));
  AND2 AND2_2123(.VSS(VSS),.VDD(VDD),.Y(g21252),.A(g19578),.B(g14895));
  AND2 AND2_2124(.VSS(VSS),.VDD(VDD),.Y(g21254),.A(g20318),.B(g14910));
  AND3 AND3_198(.VSS(VSS),.VDD(VDD),.Y(g21259),.A(g20299),.B(g16722),.C(g16682));
  AND2 AND2_2125(.VSS(VSS),.VDD(VDD),.Y(g21260),.A(g19608),.B(g14976));
  AND2 AND2_2126(.VSS(VSS),.VDD(VDD),.Y(g21262),.A(g20337),.B(g14991));
  AND3 AND3_199(.VSS(VSS),.VDD(VDD),.Y(g21267),.A(g20318),.B(g16764),.C(g16708));
  AND2 AND2_2127(.VSS(VSS),.VDD(VDD),.Y(g21268),.A(g19641),.B(g15065));
  AND2 AND2_2128(.VSS(VSS),.VDD(VDD),.Y(g21270),.A(g20357),.B(g15080));
  AND3 AND3_200(.VSS(VSS),.VDD(VDD),.Y(g21276),.A(g20337),.B(g16791),.C(g16739));
  AND2 AND2_2129(.VSS(VSS),.VDD(VDD),.Y(g21277),.A(g19681),.B(g15161));
  AND3 AND3_201(.VSS(VSS),.VDD(VDD),.Y(g21283),.A(g20357),.B(g16820),.C(g16781));
  AND2 AND2_2130(.VSS(VSS),.VDD(VDD),.Y(g21284),.A(g9356),.B(g20269));
  AND2 AND2_2131(.VSS(VSS),.VDD(VDD),.Y(g21290),.A(g9356),.B(g20278));
  AND2 AND2_2132(.VSS(VSS),.VDD(VDD),.Y(g21291),.A(g9293),.B(g20279));
  AND2 AND2_2133(.VSS(VSS),.VDD(VDD),.Y(g21292),.A(g9453),.B(g20281));
  AND2 AND2_2134(.VSS(VSS),.VDD(VDD),.Y(g21298),.A(g9356),.B(g20286));
  AND2 AND2_2135(.VSS(VSS),.VDD(VDD),.Y(g21299),.A(g9293),.B(g20287));
  AND2 AND2_2136(.VSS(VSS),.VDD(VDD),.Y(g21300),.A(g9232),.B(g20288));
  AND2 AND2_2137(.VSS(VSS),.VDD(VDD),.Y(g21301),.A(g9453),.B(g20289));
  AND2 AND2_2138(.VSS(VSS),.VDD(VDD),.Y(g21302),.A(g9374),.B(g20290));
  AND2 AND2_2139(.VSS(VSS),.VDD(VDD),.Y(g21303),.A(g9595),.B(g20292));
  AND2 AND2_2140(.VSS(VSS),.VDD(VDD),.Y(g21304),.A(g9293),.B(g20296));
  AND2 AND2_2141(.VSS(VSS),.VDD(VDD),.Y(g21305),.A(g9232),.B(g20297));
  AND2 AND2_2142(.VSS(VSS),.VDD(VDD),.Y(g21306),.A(g9187),.B(g20298));
  AND2 AND2_2143(.VSS(VSS),.VDD(VDD),.Y(g21307),.A(g9453),.B(g20302));
  AND2 AND2_2144(.VSS(VSS),.VDD(VDD),.Y(g21308),.A(g9374),.B(g20303));
  AND2 AND2_2145(.VSS(VSS),.VDD(VDD),.Y(g21309),.A(g9310),.B(g20304));
  AND2 AND2_2146(.VSS(VSS),.VDD(VDD),.Y(g21310),.A(g9595),.B(g20305));
  AND2 AND2_2147(.VSS(VSS),.VDD(VDD),.Y(g21311),.A(g9471),.B(g20306));
  AND2 AND2_2148(.VSS(VSS),.VDD(VDD),.Y(g21312),.A(g9737),.B(g20308));
  AND2 AND2_2149(.VSS(VSS),.VDD(VDD),.Y(g21313),.A(g9232),.B(g20311));
  AND2 AND2_2150(.VSS(VSS),.VDD(VDD),.Y(g21314),.A(g9187),.B(g20312));
  AND2 AND2_2151(.VSS(VSS),.VDD(VDD),.Y(g21315),.A(g9161),.B(g20313));
  AND2 AND2_2152(.VSS(VSS),.VDD(VDD),.Y(g21319),.A(g9374),.B(g20315));
  AND2 AND2_2153(.VSS(VSS),.VDD(VDD),.Y(g21320),.A(g9310),.B(g20316));
  AND2 AND2_2154(.VSS(VSS),.VDD(VDD),.Y(g21321),.A(g9248),.B(g20317));
  AND2 AND2_2155(.VSS(VSS),.VDD(VDD),.Y(g21322),.A(g9595),.B(g20321));
  AND2 AND2_2156(.VSS(VSS),.VDD(VDD),.Y(g21323),.A(g9471),.B(g20322));
  AND2 AND2_2157(.VSS(VSS),.VDD(VDD),.Y(g21324),.A(g9391),.B(g20323));
  AND2 AND2_2158(.VSS(VSS),.VDD(VDD),.Y(g21325),.A(g9737),.B(g20324));
  AND2 AND2_2159(.VSS(VSS),.VDD(VDD),.Y(g21326),.A(g9613),.B(g20325));
  AND2 AND2_2160(.VSS(VSS),.VDD(VDD),.Y(g21328),.A(g9187),.B(g20327));
  AND2 AND2_2161(.VSS(VSS),.VDD(VDD),.Y(g21329),.A(g9161),.B(g20328));
  AND2 AND2_2162(.VSS(VSS),.VDD(VDD),.Y(g21330),.A(g9150),.B(g20329));
  AND2 AND2_2163(.VSS(VSS),.VDD(VDD),.Y(g21334),.A(g9310),.B(g20330));
  AND2 AND2_2164(.VSS(VSS),.VDD(VDD),.Y(g21335),.A(g9248),.B(g20331));
  AND2 AND2_2165(.VSS(VSS),.VDD(VDD),.Y(g21336),.A(g9203),.B(g20332));
  AND2 AND2_2166(.VSS(VSS),.VDD(VDD),.Y(g21337),.A(g9471),.B(g20334));
  AND2 AND2_2167(.VSS(VSS),.VDD(VDD),.Y(g21338),.A(g9391),.B(g20335));
  AND2 AND2_2168(.VSS(VSS),.VDD(VDD),.Y(g21339),.A(g9326),.B(g20336));
  AND2 AND2_2169(.VSS(VSS),.VDD(VDD),.Y(g21340),.A(g9737),.B(g20340));
  AND2 AND2_2170(.VSS(VSS),.VDD(VDD),.Y(g21341),.A(g9613),.B(g20341));
  AND2 AND2_2171(.VSS(VSS),.VDD(VDD),.Y(g21342),.A(g9488),.B(g20342));
  AND2 AND2_2172(.VSS(VSS),.VDD(VDD),.Y(g21343),.A(g9161),.B(g20344));
  AND2 AND2_2173(.VSS(VSS),.VDD(VDD),.Y(g21344),.A(g9150),.B(g20345));
  AND2 AND2_2174(.VSS(VSS),.VDD(VDD),.Y(g21345),.A(g15096),.B(g20346));
  AND2 AND2_2175(.VSS(VSS),.VDD(VDD),.Y(g21349),.A(g9248),.B(g20347));
  AND2 AND2_2176(.VSS(VSS),.VDD(VDD),.Y(g21350),.A(g9203),.B(g20348));
  AND2 AND2_2177(.VSS(VSS),.VDD(VDD),.Y(g21351),.A(g9174),.B(g20349));
  AND2 AND2_2178(.VSS(VSS),.VDD(VDD),.Y(g21352),.A(g9391),.B(g20350));
  AND2 AND2_2179(.VSS(VSS),.VDD(VDD),.Y(g21353),.A(g9326),.B(g20351));
  AND2 AND2_2180(.VSS(VSS),.VDD(VDD),.Y(g21354),.A(g9264),.B(g20352));
  AND2 AND2_2181(.VSS(VSS),.VDD(VDD),.Y(g21355),.A(g9613),.B(g20354));
  AND2 AND2_2182(.VSS(VSS),.VDD(VDD),.Y(g21356),.A(g9488),.B(g20355));
  AND2 AND2_2183(.VSS(VSS),.VDD(VDD),.Y(g21357),.A(g9407),.B(g20356));
  AND2 AND2_2184(.VSS(VSS),.VDD(VDD),.Y(g21360),.A(g9507),.B(g20361));
  AND2 AND2_2185(.VSS(VSS),.VDD(VDD),.Y(g21361),.A(g9150),.B(g20362));
  AND2 AND2_2186(.VSS(VSS),.VDD(VDD),.Y(g21362),.A(g15096),.B(g20363));
  AND2 AND2_2187(.VSS(VSS),.VDD(VDD),.Y(g21363),.A(g15022),.B(g20364));
  AND2 AND2_2188(.VSS(VSS),.VDD(VDD),.Y(g21367),.A(g9203),.B(g20366));
  AND2 AND2_2189(.VSS(VSS),.VDD(VDD),.Y(g21368),.A(g9174),.B(g20367));
  AND2 AND2_2190(.VSS(VSS),.VDD(VDD),.Y(g21369),.A(g15188),.B(g20368));
  AND2 AND2_2191(.VSS(VSS),.VDD(VDD),.Y(g21370),.A(g9326),.B(g20369));
  AND2 AND2_2192(.VSS(VSS),.VDD(VDD),.Y(g21371),.A(g9264),.B(g20370));
  AND2 AND2_2193(.VSS(VSS),.VDD(VDD),.Y(g21372),.A(g9216),.B(g20371));
  AND2 AND2_2194(.VSS(VSS),.VDD(VDD),.Y(g21373),.A(g9488),.B(g20372));
  AND2 AND2_2195(.VSS(VSS),.VDD(VDD),.Y(g21374),.A(g9407),.B(g20373));
  AND2 AND2_2196(.VSS(VSS),.VDD(VDD),.Y(g21375),.A(g9342),.B(g20374));
  AND2 AND2_2197(.VSS(VSS),.VDD(VDD),.Y(g21378),.A(g9507),.B(g20378));
  AND2 AND2_2198(.VSS(VSS),.VDD(VDD),.Y(g21379),.A(g9427),.B(g20379));
  AND2 AND2_2199(.VSS(VSS),.VDD(VDD),.Y(g21380),.A(g15096),.B(g20380));
  AND2 AND2_2200(.VSS(VSS),.VDD(VDD),.Y(g21381),.A(g15022),.B(g20381));
  AND2 AND2_2201(.VSS(VSS),.VDD(VDD),.Y(g21388),.A(g6201),.B(g19657));
  AND2 AND2_2202(.VSS(VSS),.VDD(VDD),.Y(g21389),.A(g9649),.B(g20384));
  AND2 AND2_2203(.VSS(VSS),.VDD(VDD),.Y(g21390),.A(g9174),.B(g20385));
  AND2 AND2_2204(.VSS(VSS),.VDD(VDD),.Y(g21391),.A(g15188),.B(g20386));
  AND2 AND2_2205(.VSS(VSS),.VDD(VDD),.Y(g21392),.A(g15118),.B(g20387));
  AND2 AND2_2206(.VSS(VSS),.VDD(VDD),.Y(g21393),.A(g9264),.B(g20389));
  AND2 AND2_2207(.VSS(VSS),.VDD(VDD),.Y(g21394),.A(g9216),.B(g20390));
  AND2 AND2_2208(.VSS(VSS),.VDD(VDD),.Y(g21395),.A(g15274),.B(g20391));
  AND2 AND2_2209(.VSS(VSS),.VDD(VDD),.Y(g21396),.A(g9407),.B(g20392));
  AND2 AND2_2210(.VSS(VSS),.VDD(VDD),.Y(g21397),.A(g9342),.B(g20393));
  AND2 AND2_2211(.VSS(VSS),.VDD(VDD),.Y(g21398),.A(g9277),.B(g20394));
  AND2 AND2_2212(.VSS(VSS),.VDD(VDD),.Y(g21401),.A(g9507),.B(g20397));
  AND2 AND2_2213(.VSS(VSS),.VDD(VDD),.Y(g21402),.A(g9427),.B(g20398));
  AND2 AND2_2214(.VSS(VSS),.VDD(VDD),.Y(g21403),.A(g15022),.B(g20399));
  AND2 AND2_2215(.VSS(VSS),.VDD(VDD),.Y(g21410),.A(g6363),.B(g20402));
  AND2 AND2_2216(.VSS(VSS),.VDD(VDD),.Y(g21411),.A(g9649),.B(g20403));
  AND2 AND2_2217(.VSS(VSS),.VDD(VDD),.Y(g21412),.A(g9569),.B(g20404));
  AND2 AND2_2218(.VSS(VSS),.VDD(VDD),.Y(g21413),.A(g15188),.B(g20405));
  AND2 AND2_2219(.VSS(VSS),.VDD(VDD),.Y(g21414),.A(g15118),.B(g20406));
  AND2 AND2_2220(.VSS(VSS),.VDD(VDD),.Y(g21418),.A(g6290),.B(g19705));
  AND2 AND2_2221(.VSS(VSS),.VDD(VDD),.Y(g21419),.A(g9795),.B(g20409));
  AND2 AND2_2222(.VSS(VSS),.VDD(VDD),.Y(g21420),.A(g9216),.B(g20410));
  AND2 AND2_2223(.VSS(VSS),.VDD(VDD),.Y(g21421),.A(g15274),.B(g20411));
  AND2 AND2_2224(.VSS(VSS),.VDD(VDD),.Y(g21422),.A(g15210),.B(g20412));
  AND2 AND2_2225(.VSS(VSS),.VDD(VDD),.Y(g21423),.A(g9342),.B(g20414));
  AND2 AND2_2226(.VSS(VSS),.VDD(VDD),.Y(g21424),.A(g9277),.B(g20415));
  AND2 AND2_2227(.VSS(VSS),.VDD(VDD),.Y(g21425),.A(g15366),.B(g20416));
  AND2 AND2_2228(.VSS(VSS),.VDD(VDD),.Y(g21428),.A(g9427),.B(g20420));
  AND2 AND2_2229(.VSS(VSS),.VDD(VDD),.Y(g21438),.A(g9649),.B(g20422));
  AND2 AND2_2230(.VSS(VSS),.VDD(VDD),.Y(g21439),.A(g9569),.B(g20423));
  AND2 AND2_2231(.VSS(VSS),.VDD(VDD),.Y(g21440),.A(g15118),.B(g20424));
  AND2 AND2_2232(.VSS(VSS),.VDD(VDD),.Y(g21444),.A(g6568),.B(g20427));
  AND2 AND2_2233(.VSS(VSS),.VDD(VDD),.Y(g21445),.A(g9795),.B(g20428));
  AND2 AND2_2234(.VSS(VSS),.VDD(VDD),.Y(g21446),.A(g9711),.B(g20429));
  AND2 AND2_2235(.VSS(VSS),.VDD(VDD),.Y(g21447),.A(g15274),.B(g20430));
  AND2 AND2_2236(.VSS(VSS),.VDD(VDD),.Y(g21448),.A(g15210),.B(g20431));
  AND2 AND2_2237(.VSS(VSS),.VDD(VDD),.Y(g21452),.A(g6427),.B(g19749));
  AND2 AND2_2238(.VSS(VSS),.VDD(VDD),.Y(g21453),.A(g9941),.B(g20434));
  AND2 AND2_2239(.VSS(VSS),.VDD(VDD),.Y(g21454),.A(g9277),.B(g20435));
  AND2 AND2_2240(.VSS(VSS),.VDD(VDD),.Y(g21455),.A(g15366),.B(g20436));
  AND2 AND2_2241(.VSS(VSS),.VDD(VDD),.Y(g21456),.A(g15296),.B(g20437));
  AND2 AND2_2242(.VSS(VSS),.VDD(VDD),.Y(g21476),.A(g9569),.B(g20442));
  AND2 AND2_2243(.VSS(VSS),.VDD(VDD),.Y(g21480),.A(g9795),.B(g20444));
  AND2 AND2_2244(.VSS(VSS),.VDD(VDD),.Y(g21481),.A(g9711),.B(g20445));
  AND2 AND2_2245(.VSS(VSS),.VDD(VDD),.Y(g21482),.A(g15210),.B(g20446));
  AND2 AND2_2246(.VSS(VSS),.VDD(VDD),.Y(g21486),.A(g6832),.B(g20449));
  AND2 AND2_2247(.VSS(VSS),.VDD(VDD),.Y(g21487),.A(g9941),.B(g20450));
  AND2 AND2_2248(.VSS(VSS),.VDD(VDD),.Y(g21488),.A(g9857),.B(g20451));
  AND2 AND2_2249(.VSS(VSS),.VDD(VDD),.Y(g21489),.A(g15366),.B(g20452));
  AND2 AND2_2250(.VSS(VSS),.VDD(VDD),.Y(g21490),.A(g15296),.B(g20453));
  AND2 AND2_2251(.VSS(VSS),.VDD(VDD),.Y(g21494),.A(g6632),.B(g19792));
  AND2 AND2_2252(.VSS(VSS),.VDD(VDD),.Y(g21497),.A(g3006),.B(g20456));
  AND2 AND2_2253(.VSS(VSS),.VDD(VDD),.Y(g21517),.A(g9711),.B(g20461));
  AND2 AND2_2254(.VSS(VSS),.VDD(VDD),.Y(g21521),.A(g9941),.B(g20463));
  AND2 AND2_2255(.VSS(VSS),.VDD(VDD),.Y(g21522),.A(g9857),.B(g20464));
  AND2 AND2_2256(.VSS(VSS),.VDD(VDD),.Y(g21523),.A(g15296),.B(g20465));
  AND2 AND2_2257(.VSS(VSS),.VDD(VDD),.Y(g21527),.A(g7134),.B(g20468));
  AND3 AND3_202(.VSS(VSS),.VDD(VDD),.Y(I28068),.A(g17802),.B(g18265),.C(g17882));
  AND4 AND4_82(.VSS(VSS),.VDD(VDD),.Y(g21533),.A(g17724),.B(g18179),.C(g19799),.D(I28068));
  AND2 AND2_2258(.VSS(VSS),.VDD(VDD),.Y(g21553),.A(g9857),.B(g20476));
  AND3 AND3_203(.VSS(VSS),.VDD(VDD),.Y(I28096),.A(g13907),.B(g14238),.C(g13946));
  AND4 AND4_83(.VSS(VSS),.VDD(VDD),.Y(g21564),.A(g13886),.B(g14153),.C(g19799),.D(I28096));
  AND3 AND3_204(.VSS(VSS),.VDD(VDD),.Y(I28103),.A(g17914),.B(g18358),.C(g17993));
  AND4 AND4_84(.VSS(VSS),.VDD(VDD),.Y(g21569),.A(g17825),.B(g18286),.C(g19843),.D(I28103));
  AND2 AND2_2259(.VSS(VSS),.VDD(VDD),.Y(g21589),.A(g3002),.B(g19890));
  AND3 AND3_205(.VSS(VSS),.VDD(VDD),.Y(g21593),.A(g16498),.B(g19484),.C(g14071));
  AND3 AND3_206(.VSS(VSS),.VDD(VDD),.Y(I28126),.A(g13963),.B(g14360),.C(g14016));
  AND4 AND4_85(.VSS(VSS),.VDD(VDD),.Y(g21597),.A(g13927),.B(g14268),.C(g19843),.D(I28126));
  AND3 AND3_207(.VSS(VSS),.VDD(VDD),.Y(I28133),.A(g18025),.B(g18453),.C(g18110));
  AND4 AND4_86(.VSS(VSS),.VDD(VDD),.Y(g21602),.A(g17937),.B(g18379),.C(g19876),.D(I28133));
  AND2 AND2_2260(.VSS(VSS),.VDD(VDD),.Y(g21610),.A(g7522),.B(g20490));
  AND2 AND2_2261(.VSS(VSS),.VDD(VDD),.Y(g21611),.A(g7471),.B(g19915));
  AND3 AND3_208(.VSS(VSS),.VDD(VDD),.Y(g21622),.A(g16520),.B(g19505),.C(g14186));
  AND3 AND3_209(.VSS(VSS),.VDD(VDD),.Y(I28155),.A(g14033),.B(g14472),.C(g14107));
  AND4 AND4_87(.VSS(VSS),.VDD(VDD),.Y(g21626),.A(g13983),.B(g14390),.C(g19876),.D(I28155));
  AND3 AND3_210(.VSS(VSS),.VDD(VDD),.Y(I28162),.A(g18142),.B(g18526),.C(g18226));
  AND4 AND4_88(.VSS(VSS),.VDD(VDD),.Y(g21631),.A(g18048),.B(g18474),.C(g19907),.D(I28162));
  AND2 AND2_2262(.VSS(VSS),.VDD(VDD),.Y(g21635),.A(g7549),.B(g20496));
  AND2 AND2_2263(.VSS(VSS),.VDD(VDD),.Y(g21639),.A(g3398),.B(g20500));
  AND3 AND3_211(.VSS(VSS),.VDD(VDD),.Y(g21650),.A(g16551),.B(g19524),.C(g14301));
  AND3 AND3_212(.VSS(VSS),.VDD(VDD),.Y(I28181),.A(g14124),.B(g14559),.C(g14222));
  AND4 AND4_89(.VSS(VSS),.VDD(VDD),.Y(g21654),.A(g14053),.B(g14502),.C(g19907),.D(I28181));
  AND2 AND2_2264(.VSS(VSS),.VDD(VDD),.Y(g21658),.A(g2896),.B(g20501));
  AND2 AND2_2265(.VSS(VSS),.VDD(VDD),.Y(g21666),.A(g3398),.B(g20504));
  AND2 AND2_2266(.VSS(VSS),.VDD(VDD),.Y(g21670),.A(g3554),.B(g20505));
  AND3 AND3_213(.VSS(VSS),.VDD(VDD),.Y(g21681),.A(g16583),.B(g19534),.C(g14423));
  AND2 AND2_2267(.VSS(VSS),.VDD(VDD),.Y(g21687),.A(g3398),.B(g20516));
  AND2 AND2_2268(.VSS(VSS),.VDD(VDD),.Y(g21695),.A(g3554),.B(g20517));
  AND2 AND2_2269(.VSS(VSS),.VDD(VDD),.Y(g21699),.A(g3710),.B(g20518));
  AND2 AND2_2270(.VSS(VSS),.VDD(VDD),.Y(g21707),.A(g2892),.B(g19978));
  AND2 AND2_2271(.VSS(VSS),.VDD(VDD),.Y(g21723),.A(g3554),.B(g20534));
  AND2 AND2_2272(.VSS(VSS),.VDD(VDD),.Y(g21731),.A(g3710),.B(g20535));
  AND2 AND2_2273(.VSS(VSS),.VDD(VDD),.Y(g21735),.A(g3866),.B(g20536));
  AND2 AND2_2274(.VSS(VSS),.VDD(VDD),.Y(g21749),.A(g3710),.B(g20553));
  AND2 AND2_2275(.VSS(VSS),.VDD(VDD),.Y(g21757),.A(g3866),.B(g20554));
  AND2 AND2_2276(.VSS(VSS),.VDD(VDD),.Y(g21758),.A(g7607),.B(g20045));
  AND2 AND2_2277(.VSS(VSS),.VDD(VDD),.Y(g21773),.A(g3866),.B(g19078));
  AND3 AND3_214(.VSS(VSS),.VDD(VDD),.Y(g21805),.A(g16679),.B(g19578),.C(g14776));
  AND3 AND3_215(.VSS(VSS),.VDD(VDD),.Y(g21812),.A(g16705),.B(g19608),.C(g14811));
  AND3 AND3_216(.VSS(VSS),.VDD(VDD),.Y(g21818),.A(g16736),.B(g19641),.C(g14863));
  AND3 AND3_217(.VSS(VSS),.VDD(VDD),.Y(g21822),.A(g16778),.B(g19681),.C(g14936));
  AND2 AND2_2278(.VSS(VSS),.VDD(VDD),.Y(g21891),.A(g19302),.B(g11749));
  AND2 AND2_2279(.VSS(VSS),.VDD(VDD),.Y(g21892),.A(g19288),.B(g13011));
  AND2 AND2_2280(.VSS(VSS),.VDD(VDD),.Y(g21899),.A(g19323),.B(g11749));
  AND2 AND2_2281(.VSS(VSS),.VDD(VDD),.Y(g21900),.A(g19306),.B(g13011));
  AND2 AND2_2282(.VSS(VSS),.VDD(VDD),.Y(g21906),.A(g5715),.B(g20513));
  AND2 AND2_2283(.VSS(VSS),.VDD(VDD),.Y(g21911),.A(g19350),.B(g11749));
  AND2 AND2_2284(.VSS(VSS),.VDD(VDD),.Y(g21912),.A(g19327),.B(g13011));
  AND2 AND2_2285(.VSS(VSS),.VDD(VDD),.Y(g21913),.A(g4456),.B(g20519));
  AND2 AND2_2286(.VSS(VSS),.VDD(VDD),.Y(g21920),.A(g5773),.B(g20531));
  AND2 AND2_2287(.VSS(VSS),.VDD(VDD),.Y(g21925),.A(g19384),.B(g11749));
  AND2 AND2_2288(.VSS(VSS),.VDD(VDD),.Y(g21926),.A(g19354),.B(g13011));
  AND2 AND2_2289(.VSS(VSS),.VDD(VDD),.Y(g21931),.A(g4632),.B(g20539));
  AND2 AND2_2290(.VSS(VSS),.VDD(VDD),.Y(g21938),.A(g5832),.B(g20550));
  AND2 AND2_2291(.VSS(VSS),.VDD(VDD),.Y(g21990),.A(g291),.B(g21187));
  AND2 AND2_2292(.VSS(VSS),.VDD(VDD),.Y(g22004),.A(g978),.B(g21202));
  AND2 AND2_2293(.VSS(VSS),.VDD(VDD),.Y(g22015),.A(g1672),.B(g21217));
  AND2 AND2_2294(.VSS(VSS),.VDD(VDD),.Y(g22020),.A(g2366),.B(g21225));
  AND3 AND3_218(.VSS(VSS),.VDD(VDD),.Y(I28582),.A(g19141),.B(g21133),.C(g21116));
  AND4 AND4_90(.VSS(VSS),.VDD(VDD),.Y(g22036),.A(g21104),.B(g21095),.C(g21084),.D(I28582));
  AND3 AND3_219(.VSS(VSS),.VDD(VDD),.Y(I28594),.A(g21167),.B(g21147),.C(g21134));
  AND4 AND4_91(.VSS(VSS),.VDD(VDD),.Y(g22046),.A(g21117),.B(g21105),.C(g21096),.D(I28594));
  AND3 AND3_220(.VSS(VSS),.VDD(VDD),.Y(I28609),.A(g21183),.B(g21168),.C(g21148));
  AND4 AND4_92(.VSS(VSS),.VDD(VDD),.Y(g22062),.A(g21135),.B(g21118),.C(g21106),.D(I28609));
  AND2 AND2_2295(.VSS(VSS),.VDD(VDD),.Y(g22187),.A(g21564),.B(g20986));
  AND2 AND2_2296(.VSS(VSS),.VDD(VDD),.Y(g22196),.A(g21597),.B(g21012));
  AND2 AND2_2297(.VSS(VSS),.VDD(VDD),.Y(g22201),.A(g21271),.B(g16881));
  AND2 AND2_2298(.VSS(VSS),.VDD(VDD),.Y(g22202),.A(g21626),.B(g21036));
  AND2 AND2_2299(.VSS(VSS),.VDD(VDD),.Y(g22206),.A(g21895),.B(g11976));
  AND2 AND2_2300(.VSS(VSS),.VDD(VDD),.Y(g22207),.A(g21278),.B(g16910));
  AND2 AND2_2301(.VSS(VSS),.VDD(VDD),.Y(g22208),.A(g21654),.B(g21057));
  AND2 AND2_2302(.VSS(VSS),.VDD(VDD),.Y(g22211),.A(g21661),.B(g12027));
  AND2 AND2_2303(.VSS(VSS),.VDD(VDD),.Y(g22214),.A(g21907),.B(g12045));
  AND2 AND2_2304(.VSS(VSS),.VDD(VDD),.Y(g22215),.A(g21285),.B(g16940));
  AND2 AND2_2305(.VSS(VSS),.VDD(VDD),.Y(g22220),.A(g21690),.B(g12091));
  AND2 AND2_2306(.VSS(VSS),.VDD(VDD),.Y(g22223),.A(g21921),.B(g12109));
  AND2 AND2_2307(.VSS(VSS),.VDD(VDD),.Y(g22224),.A(g21293),.B(g16971));
  AND2 AND2_2308(.VSS(VSS),.VDD(VDD),.Y(g22228),.A(g21716),.B(g12136));
  AND2 AND2_2309(.VSS(VSS),.VDD(VDD),.Y(g22229),.A(g21661),.B(g12139));
  AND2 AND2_2310(.VSS(VSS),.VDD(VDD),.Y(g22235),.A(g21726),.B(g12163));
  AND2 AND2_2311(.VSS(VSS),.VDD(VDD),.Y(g22238),.A(g21939),.B(g12181));
  AND2 AND2_2312(.VSS(VSS),.VDD(VDD),.Y(g22244),.A(g21742),.B(g12198));
  AND2 AND2_2313(.VSS(VSS),.VDD(VDD),.Y(g22245),.A(g21690),.B(g12201));
  AND2 AND2_2314(.VSS(VSS),.VDD(VDD),.Y(g22250),.A(g21752),.B(g12225));
  AND2 AND2_2315(.VSS(VSS),.VDD(VDD),.Y(g22254),.A(g21716),.B(g12239));
  AND2 AND2_2316(.VSS(VSS),.VDD(VDD),.Y(g22255),.A(g21661),.B(g12242));
  AND2 AND2_2317(.VSS(VSS),.VDD(VDD),.Y(g22264),.A(g21766),.B(g12253));
  AND2 AND2_2318(.VSS(VSS),.VDD(VDD),.Y(g22265),.A(g21726),.B(g12256));
  AND2 AND2_2319(.VSS(VSS),.VDD(VDD),.Y(g22270),.A(g92),.B(g21529));
  AND2 AND2_2320(.VSS(VSS),.VDD(VDD),.Y(g22272),.A(g21742),.B(g12282));
  AND2 AND2_2321(.VSS(VSS),.VDD(VDD),.Y(g22273),.A(g21690),.B(g12285));
  AND2 AND2_2322(.VSS(VSS),.VDD(VDD),.Y(g22281),.A(g21782),.B(g12296));
  AND2 AND2_2323(.VSS(VSS),.VDD(VDD),.Y(g22282),.A(g21752),.B(g12299));
  AND2 AND2_2324(.VSS(VSS),.VDD(VDD),.Y(g22285),.A(g21716),.B(g12312));
  AND2 AND2_2325(.VSS(VSS),.VDD(VDD),.Y(g22289),.A(g780),.B(g21565));
  AND2 AND2_2326(.VSS(VSS),.VDD(VDD),.Y(g22291),.A(g21766),.B(g12318));
  AND2 AND2_2327(.VSS(VSS),.VDD(VDD),.Y(g22292),.A(g21726),.B(g12321));
  AND2 AND2_2328(.VSS(VSS),.VDD(VDD),.Y(g22305),.A(g21742),.B(g12340));
  AND2 AND2_2329(.VSS(VSS),.VDD(VDD),.Y(g22309),.A(g1466),.B(g21598));
  AND2 AND2_2330(.VSS(VSS),.VDD(VDD),.Y(g22311),.A(g21782),.B(g12346));
  AND2 AND2_2331(.VSS(VSS),.VDD(VDD),.Y(g22312),.A(g21752),.B(g12349));
  AND2 AND2_2332(.VSS(VSS),.VDD(VDD),.Y(g22333),.A(g21766),.B(g12370));
  AND2 AND2_2333(.VSS(VSS),.VDD(VDD),.Y(g22337),.A(g2160),.B(g21627));
  AND2 AND2_2334(.VSS(VSS),.VDD(VDD),.Y(g22340),.A(g88),.B(g21184));
  AND2 AND2_2335(.VSS(VSS),.VDD(VDD),.Y(g22358),.A(g21782),.B(g12389));
  AND2 AND2_2336(.VSS(VSS),.VDD(VDD),.Y(g22363),.A(g776),.B(g21199));
  AND2 AND2_2337(.VSS(VSS),.VDD(VDD),.Y(g22383),.A(g1462),.B(g21214));
  AND2 AND2_2338(.VSS(VSS),.VDD(VDD),.Y(g22398),.A(g2156),.B(g21222));
  AND2 AND2_2339(.VSS(VSS),.VDD(VDD),.Y(g22483),.A(g646),.B(g21861));
  AND2 AND2_2340(.VSS(VSS),.VDD(VDD),.Y(g22515),.A(g13873),.B(g21382));
  AND2 AND2_2341(.VSS(VSS),.VDD(VDD),.Y(g22516),.A(g20885),.B(g17442));
  AND2 AND2_2342(.VSS(VSS),.VDD(VDD),.Y(g22517),.A(g21895),.B(g12608));
  AND2 AND2_2343(.VSS(VSS),.VDD(VDD),.Y(g22526),.A(g1332),.B(g21867));
  AND2 AND2_2344(.VSS(VSS),.VDD(VDD),.Y(g22546),.A(g13886),.B(g21404));
  AND2 AND2_2345(.VSS(VSS),.VDD(VDD),.Y(g22555),.A(g13895),.B(g21415));
  AND2 AND2_2346(.VSS(VSS),.VDD(VDD),.Y(g22556),.A(g20904),.B(g17523));
  AND2 AND2_2347(.VSS(VSS),.VDD(VDD),.Y(g22557),.A(g21907),.B(g12654));
  AND2 AND2_2348(.VSS(VSS),.VDD(VDD),.Y(g22566),.A(g2026),.B(g21872));
  AND2 AND2_2349(.VSS(VSS),.VDD(VDD),.Y(g22577),.A(g13907),.B(g21429));
  AND2 AND2_2350(.VSS(VSS),.VDD(VDD),.Y(g22581),.A(g21895),.B(g12699));
  AND2 AND2_2351(.VSS(VSS),.VDD(VDD),.Y(g22587),.A(g13927),.B(g21441));
  AND2 AND2_2352(.VSS(VSS),.VDD(VDD),.Y(g22595),.A(g13936),.B(g21449));
  AND2 AND2_2353(.VSS(VSS),.VDD(VDD),.Y(g22596),.A(g20928),.B(g17613));
  AND2 AND2_2354(.VSS(VSS),.VDD(VDD),.Y(g22597),.A(g21921),.B(g12708));
  AND2 AND2_2355(.VSS(VSS),.VDD(VDD),.Y(g22606),.A(g2720),.B(g21876));
  AND2 AND2_2356(.VSS(VSS),.VDD(VDD),.Y(g22607),.A(g13946),.B(g21458));
  AND2 AND2_2357(.VSS(VSS),.VDD(VDD),.Y(g22610),.A(g660),.B(g21473));
  AND2 AND2_2358(.VSS(VSS),.VDD(VDD),.Y(g22614),.A(g13963),.B(g21477));
  AND2 AND2_2359(.VSS(VSS),.VDD(VDD),.Y(g22618),.A(g21907),.B(g12756));
  AND2 AND2_2360(.VSS(VSS),.VDD(VDD),.Y(g22624),.A(g13983),.B(g21483));
  AND2 AND2_2361(.VSS(VSS),.VDD(VDD),.Y(g22632),.A(g13992),.B(g21491));
  AND2 AND2_2362(.VSS(VSS),.VDD(VDD),.Y(g22633),.A(g20956),.B(g17710));
  AND2 AND2_2363(.VSS(VSS),.VDD(VDD),.Y(g22634),.A(g21939),.B(g12765));
  AND2 AND2_2364(.VSS(VSS),.VDD(VDD),.Y(g22637),.A(g20841),.B(g10927));
  AND2 AND2_2365(.VSS(VSS),.VDD(VDD),.Y(g22638),.A(g14001),.B(g21498));
  AND2 AND2_2366(.VSS(VSS),.VDD(VDD),.Y(g22643),.A(g14016),.B(g21505));
  AND2 AND2_2367(.VSS(VSS),.VDD(VDD),.Y(g22646),.A(g1346),.B(g21514));
  AND2 AND2_2368(.VSS(VSS),.VDD(VDD),.Y(g22650),.A(g14033),.B(g21518));
  AND2 AND2_2369(.VSS(VSS),.VDD(VDD),.Y(g22654),.A(g21921),.B(g12798));
  AND2 AND2_2370(.VSS(VSS),.VDD(VDD),.Y(g22660),.A(g14053),.B(g21524));
  AND2 AND2_2371(.VSS(VSS),.VDD(VDD),.Y(g22665),.A(g20920),.B(g6153));
  AND2 AND2_2372(.VSS(VSS),.VDD(VDD),.Y(g22666),.A(g21825),.B(g20014));
  AND2 AND2_2373(.VSS(VSS),.VDD(VDD),.Y(g22667),.A(g14062),.B(g21530));
  AND2 AND2_2374(.VSS(VSS),.VDD(VDD),.Y(g22674),.A(g14092),.B(g21537));
  AND2 AND2_2375(.VSS(VSS),.VDD(VDD),.Y(g22679),.A(g14107),.B(g21541));
  AND2 AND2_2376(.VSS(VSS),.VDD(VDD),.Y(g22682),.A(g2040),.B(g21550));
  AND2 AND2_2377(.VSS(VSS),.VDD(VDD),.Y(g22686),.A(g14124),.B(g21554));
  AND2 AND2_2378(.VSS(VSS),.VDD(VDD),.Y(g22690),.A(g21939),.B(g12837));
  AND2 AND2_2379(.VSS(VSS),.VDD(VDD),.Y(g22699),.A(g7338),.B(g21883));
  AND2 AND2_2380(.VSS(VSS),.VDD(VDD),.Y(g22700),.A(g7146),.B(g21558));
  AND2 AND2_2381(.VSS(VSS),.VDD(VDD),.Y(g22701),.A(g18174),.B(g21561));
  AND2 AND2_2382(.VSS(VSS),.VDD(VDD),.Y(g22707),.A(g14177),.B(g21566));
  AND2 AND2_2383(.VSS(VSS),.VDD(VDD),.Y(g22714),.A(g14207),.B(g21573));
  AND2 AND2_2384(.VSS(VSS),.VDD(VDD),.Y(g22719),.A(g14222),.B(g21577));
  AND2 AND2_2385(.VSS(VSS),.VDD(VDD),.Y(g22722),.A(g2734),.B(g21586));
  AND2 AND2_2386(.VSS(VSS),.VDD(VDD),.Y(g22726),.A(g3036),.B(g21886));
  AND2 AND2_2387(.VSS(VSS),.VDD(VDD),.Y(g22727),.A(g14238),.B(g21590));
  AND2 AND2_2388(.VSS(VSS),.VDD(VDD),.Y(g22732),.A(g18281),.B(g21594));
  AND2 AND2_2389(.VSS(VSS),.VDD(VDD),.Y(g22738),.A(g14292),.B(g21599));
  AND2 AND2_2390(.VSS(VSS),.VDD(VDD),.Y(g22745),.A(g14322),.B(g21606));
  AND2 AND2_2391(.VSS(VSS),.VDD(VDD),.Y(g22754),.A(g14342),.B(g21612));
  AND2 AND2_2392(.VSS(VSS),.VDD(VDD),.Y(g22759),.A(g14360),.B(g21619));
  AND2 AND2_2393(.VSS(VSS),.VDD(VDD),.Y(g22764),.A(g18374),.B(g21623));
  AND2 AND2_2394(.VSS(VSS),.VDD(VDD),.Y(g22770),.A(g14414),.B(g21628));
  AND2 AND2_2395(.VSS(VSS),.VDD(VDD),.Y(g22788),.A(g14454),.B(g21640));
  AND2 AND2_2396(.VSS(VSS),.VDD(VDD),.Y(g22793),.A(g14472),.B(g21647));
  AND2 AND2_2397(.VSS(VSS),.VDD(VDD),.Y(g22798),.A(g18469),.B(g21651));
  AND2 AND2_2398(.VSS(VSS),.VDD(VDD),.Y(g22804),.A(g2920),.B(g21655));
  AND2 AND2_2399(.VSS(VSS),.VDD(VDD),.Y(g22830),.A(g14541),.B(g21671));
  AND2 AND2_2400(.VSS(VSS),.VDD(VDD),.Y(g22835),.A(g14559),.B(g21678));
  AND2 AND2_2401(.VSS(VSS),.VDD(VDD),.Y(g22841),.A(g7583),.B(g21902));
  AND2 AND2_2402(.VSS(VSS),.VDD(VDD),.Y(g22842),.A(g3032),.B(g21682));
  AND2 AND2_2403(.VSS(VSS),.VDD(VDD),.Y(g22869),.A(g14596),.B(g21700));
  AND2 AND2_2404(.VSS(VSS),.VDD(VDD),.Y(g22874),.A(g7587),.B(g21708));
  AND2 AND2_2405(.VSS(VSS),.VDD(VDD),.Y(g22906),.A(g2924),.B(g21927));
  AND2 AND2_2406(.VSS(VSS),.VDD(VDD),.Y(g22984),.A(g16840),.B(g21400));
  AND2 AND2_2407(.VSS(VSS),.VDD(VDD),.Y(g23104),.A(g20842),.B(g15859));
  AND2 AND2_2408(.VSS(VSS),.VDD(VDD),.Y(g23106),.A(g5857),.B(g21050));
  AND2 AND2_2409(.VSS(VSS),.VDD(VDD),.Y(g23118),.A(g20850),.B(g15890));
  AND2 AND2_2410(.VSS(VSS),.VDD(VDD),.Y(g23119),.A(g5904),.B(g21069));
  AND2 AND2_2411(.VSS(VSS),.VDD(VDD),.Y(g23127),.A(g20858),.B(g15923));
  AND2 AND2_2412(.VSS(VSS),.VDD(VDD),.Y(g23128),.A(g5943),.B(g21079));
  AND2 AND2_2413(.VSS(VSS),.VDD(VDD),.Y(g23138),.A(g20866),.B(g15952));
  AND2 AND2_2414(.VSS(VSS),.VDD(VDD),.Y(g23139),.A(g5977),.B(g21093));
  AND2 AND2_2415(.VSS(VSS),.VDD(VDD),.Y(g23409),.A(g21533),.B(g22408));
  AND2 AND2_2416(.VSS(VSS),.VDD(VDD),.Y(g23414),.A(g21569),.B(g22421));
  AND2 AND2_2417(.VSS(VSS),.VDD(VDD),.Y(g23419),.A(g22755),.B(g19577));
  AND2 AND2_2418(.VSS(VSS),.VDD(VDD),.Y(g23423),.A(g21602),.B(g22443));
  AND2 AND2_2419(.VSS(VSS),.VDD(VDD),.Y(g23428),.A(g22789),.B(g19607));
  AND2 AND2_2420(.VSS(VSS),.VDD(VDD),.Y(g23432),.A(g21631),.B(g22476));
  AND2 AND2_2421(.VSS(VSS),.VDD(VDD),.Y(g23434),.A(g22831),.B(g19640));
  AND2 AND2_2422(.VSS(VSS),.VDD(VDD),.Y(g23440),.A(g22870),.B(g19680));
  AND2 AND2_2423(.VSS(VSS),.VDD(VDD),.Y(g23451),.A(g18552),.B(g22547));
  AND2 AND2_2424(.VSS(VSS),.VDD(VDD),.Y(g23458),.A(g18602),.B(g22588));
  AND2 AND2_2425(.VSS(VSS),.VDD(VDD),.Y(g23462),.A(g17988),.B(g22609));
  AND2 AND2_2426(.VSS(VSS),.VDD(VDD),.Y(g23467),.A(g18634),.B(g22625));
  AND2 AND2_2427(.VSS(VSS),.VDD(VDD),.Y(g23471),.A(g18105),.B(g22645));
  AND2 AND2_2428(.VSS(VSS),.VDD(VDD),.Y(g23476),.A(g18643),.B(g22661));
  AND2 AND2_2429(.VSS(VSS),.VDD(VDD),.Y(g23483),.A(g22945),.B(g8847));
  AND2 AND2_2430(.VSS(VSS),.VDD(VDD),.Y(g23484),.A(g18221),.B(g22681));
  AND2 AND2_2431(.VSS(VSS),.VDD(VDD),.Y(g23494),.A(g18328),.B(g22721));
  AND2 AND2_2432(.VSS(VSS),.VDD(VDD),.Y(g23496),.A(g5802),.B(g22300));
  AND2 AND2_2433(.VSS(VSS),.VDD(VDD),.Y(g23510),.A(g5890),.B(g22753));
  AND2 AND2_2434(.VSS(VSS),.VDD(VDD),.Y(g23512),.A(g5858),.B(g22328));
  AND2 AND2_2435(.VSS(VSS),.VDD(VDD),.Y(g23525),.A(g5929),.B(g22787));
  AND2 AND2_2436(.VSS(VSS),.VDD(VDD),.Y(g23527),.A(g5905),.B(g22353));
  AND2 AND2_2437(.VSS(VSS),.VDD(VDD),.Y(g23536),.A(g5963),.B(g22829));
  AND2 AND2_2438(.VSS(VSS),.VDD(VDD),.Y(g23538),.A(g5944),.B(g22376));
  AND2 AND2_2439(.VSS(VSS),.VDD(VDD),.Y(g23544),.A(g5992),.B(g22868));
  AND2 AND2_2440(.VSS(VSS),.VDD(VDD),.Y(g23547),.A(g8062),.B(g22405));
  AND2 AND2_2441(.VSS(VSS),.VDD(VDD),.Y(g23550),.A(g8132),.B(g22409));
  AND2 AND2_2442(.VSS(VSS),.VDD(VDD),.Y(g23551),.A(g8135),.B(g22412));
  AND2 AND2_2443(.VSS(VSS),.VDD(VDD),.Y(g23552),.A(g6136),.B(g22415));
  AND2 AND2_2444(.VSS(VSS),.VDD(VDD),.Y(g23554),.A(g8147),.B(g22418));
  AND2 AND2_2445(.VSS(VSS),.VDD(VDD),.Y(g23558),.A(g8200),.B(g22422));
  AND2 AND2_2446(.VSS(VSS),.VDD(VDD),.Y(g23559),.A(g8203),.B(g22425));
  AND2 AND2_2447(.VSS(VSS),.VDD(VDD),.Y(g23560),.A(g8206),.B(g22428));
  AND2 AND2_2448(.VSS(VSS),.VDD(VDD),.Y(g23563),.A(g8218),.B(g22431));
  AND2 AND2_2449(.VSS(VSS),.VDD(VDD),.Y(g23564),.A(g8221),.B(g22434));
  AND2 AND2_2450(.VSS(VSS),.VDD(VDD),.Y(g23565),.A(g6146),.B(g22437));
  AND2 AND2_2451(.VSS(VSS),.VDD(VDD),.Y(g23567),.A(g8233),.B(g22440));
  AND2 AND2_2452(.VSS(VSS),.VDD(VDD),.Y(g23571),.A(g3931),.B(g22445));
  AND2 AND2_2453(.VSS(VSS),.VDD(VDD),.Y(g23572),.A(g3934),.B(g22448));
  AND2 AND2_2454(.VSS(VSS),.VDD(VDD),.Y(g23573),.A(g3937),.B(g22451));
  AND2 AND2_2455(.VSS(VSS),.VDD(VDD),.Y(g23577),.A(g3957),.B(g22455));
  AND2 AND2_2456(.VSS(VSS),.VDD(VDD),.Y(g23578),.A(g3960),.B(g22458));
  AND2 AND2_2457(.VSS(VSS),.VDD(VDD),.Y(g23579),.A(g3963),.B(g22461));
  AND2 AND2_2458(.VSS(VSS),.VDD(VDD),.Y(g23582),.A(g3975),.B(g22464));
  AND2 AND2_2459(.VSS(VSS),.VDD(VDD),.Y(g23583),.A(g3978),.B(g22467));
  AND2 AND2_2460(.VSS(VSS),.VDD(VDD),.Y(g23584),.A(g6167),.B(g22470));
  AND2 AND2_2461(.VSS(VSS),.VDD(VDD),.Y(g23586),.A(g3990),.B(g22473));
  AND2 AND2_2462(.VSS(VSS),.VDD(VDD),.Y(g23590),.A(g4009),.B(g22477));
  AND2 AND2_2463(.VSS(VSS),.VDD(VDD),.Y(g23591),.A(g4012),.B(g22480));
  AND2 AND2_2464(.VSS(VSS),.VDD(VDD),.Y(g23592),.A(g17640),.B(g22986));
  AND2 AND2_2465(.VSS(VSS),.VDD(VDD),.Y(g23593),.A(g22845),.B(g20365));
  AND2 AND2_2466(.VSS(VSS),.VDD(VDD),.Y(g23598),.A(g4038),.B(g22484));
  AND2 AND2_2467(.VSS(VSS),.VDD(VDD),.Y(g23599),.A(g4041),.B(g22487));
  AND2 AND2_2468(.VSS(VSS),.VDD(VDD),.Y(g23600),.A(g4044),.B(g22490));
  AND2 AND2_2469(.VSS(VSS),.VDD(VDD),.Y(g23604),.A(g4064),.B(g22494));
  AND2 AND2_2470(.VSS(VSS),.VDD(VDD),.Y(g23605),.A(g4067),.B(g22497));
  AND2 AND2_2471(.VSS(VSS),.VDD(VDD),.Y(g23606),.A(g4070),.B(g22500));
  AND2 AND2_2472(.VSS(VSS),.VDD(VDD),.Y(g23609),.A(g4082),.B(g22503));
  AND2 AND2_2473(.VSS(VSS),.VDD(VDD),.Y(g23610),.A(g4085),.B(g22506));
  AND2 AND2_2474(.VSS(VSS),.VDD(VDD),.Y(g23611),.A(g6194),.B(g22509));
  AND2 AND2_2475(.VSS(VSS),.VDD(VDD),.Y(g23615),.A(g4107),.B(g22512));
  AND2 AND2_2476(.VSS(VSS),.VDD(VDD),.Y(g23616),.A(g17724),.B(g22988));
  AND2 AND2_2477(.VSS(VSS),.VDD(VDD),.Y(g23617),.A(g22810),.B(g20382));
  AND2 AND2_2478(.VSS(VSS),.VDD(VDD),.Y(g23618),.A(g22608),.B(g20383));
  AND2 AND2_2479(.VSS(VSS),.VDD(VDD),.Y(g23622),.A(g4136),.B(g22520));
  AND2 AND2_2480(.VSS(VSS),.VDD(VDD),.Y(g23623),.A(g4139),.B(g22523));
  AND2 AND2_2481(.VSS(VSS),.VDD(VDD),.Y(g23624),.A(g17741),.B(g22989));
  AND2 AND2_2482(.VSS(VSS),.VDD(VDD),.Y(g23625),.A(g22880),.B(g20388));
  AND2 AND2_2483(.VSS(VSS),.VDD(VDD),.Y(g23630),.A(g4165),.B(g22527));
  AND2 AND2_2484(.VSS(VSS),.VDD(VDD),.Y(g23631),.A(g4168),.B(g22530));
  AND2 AND2_2485(.VSS(VSS),.VDD(VDD),.Y(g23632),.A(g4171),.B(g22533));
  AND2 AND2_2486(.VSS(VSS),.VDD(VDD),.Y(g23636),.A(g4191),.B(g22537));
  AND2 AND2_2487(.VSS(VSS),.VDD(VDD),.Y(g23637),.A(g4194),.B(g22540));
  AND2 AND2_2488(.VSS(VSS),.VDD(VDD),.Y(g23638),.A(g4197),.B(g22543));
  AND2 AND2_2489(.VSS(VSS),.VDD(VDD),.Y(g23639),.A(g21825),.B(g22805));
  AND2 AND2_2490(.VSS(VSS),.VDD(VDD),.Y(g23643),.A(g17802),.B(g22991));
  AND2 AND2_2491(.VSS(VSS),.VDD(VDD),.Y(g23659),.A(g22784),.B(g17500));
  AND2 AND2_2492(.VSS(VSS),.VDD(VDD),.Y(g23664),.A(g4246),.B(g22552));
  AND2 AND2_2493(.VSS(VSS),.VDD(VDD),.Y(g23665),.A(g17825),.B(g22995));
  AND2 AND2_2494(.VSS(VSS),.VDD(VDD),.Y(g23666),.A(g22851),.B(g20407));
  AND2 AND2_2495(.VSS(VSS),.VDD(VDD),.Y(g23667),.A(g22644),.B(g20408));
  AND2 AND2_2496(.VSS(VSS),.VDD(VDD),.Y(g23671),.A(g4275),.B(g22560));
  AND2 AND2_2497(.VSS(VSS),.VDD(VDD),.Y(g23672),.A(g4278),.B(g22563));
  AND2 AND2_2498(.VSS(VSS),.VDD(VDD),.Y(g23673),.A(g17842),.B(g22996));
  AND2 AND2_2499(.VSS(VSS),.VDD(VDD),.Y(g23674),.A(g22915),.B(g20413));
  AND2 AND2_2500(.VSS(VSS),.VDD(VDD),.Y(g23679),.A(g4304),.B(g22567));
  AND2 AND2_2501(.VSS(VSS),.VDD(VDD),.Y(g23680),.A(g4307),.B(g22570));
  AND2 AND2_2502(.VSS(VSS),.VDD(VDD),.Y(g23681),.A(g4310),.B(g22573));
  AND2 AND2_2503(.VSS(VSS),.VDD(VDD),.Y(g23686),.A(g17882),.B(g22998));
  AND2 AND2_2504(.VSS(VSS),.VDD(VDD),.Y(g23687),.A(g22668),.B(g17570));
  AND2 AND2_2505(.VSS(VSS),.VDD(VDD),.Y(g23689),.A(g6513),.B(g23001));
  AND2 AND2_2506(.VSS(VSS),.VDD(VDD),.Y(g23693),.A(g17914),.B(g23002));
  AND2 AND2_2507(.VSS(VSS),.VDD(VDD),.Y(g23709),.A(g22826),.B(g17591));
  AND2 AND2_2508(.VSS(VSS),.VDD(VDD),.Y(g23714),.A(g4401),.B(g22592));
  AND2 AND2_2509(.VSS(VSS),.VDD(VDD),.Y(g23715),.A(g17937),.B(g23006));
  AND2 AND2_2510(.VSS(VSS),.VDD(VDD),.Y(g23716),.A(g22886),.B(g20432));
  AND2 AND2_2511(.VSS(VSS),.VDD(VDD),.Y(g23717),.A(g22680),.B(g20433));
  AND2 AND2_2512(.VSS(VSS),.VDD(VDD),.Y(g23721),.A(g4430),.B(g22600));
  AND2 AND2_2513(.VSS(VSS),.VDD(VDD),.Y(g23722),.A(g4433),.B(g22603));
  AND2 AND2_2514(.VSS(VSS),.VDD(VDD),.Y(g23723),.A(g17954),.B(g23007));
  AND2 AND2_2515(.VSS(VSS),.VDD(VDD),.Y(g23724),.A(g22940),.B(g20438));
  AND2 AND2_2516(.VSS(VSS),.VDD(VDD),.Y(g23726),.A(g21825),.B(g22843));
  AND2 AND2_2517(.VSS(VSS),.VDD(VDD),.Y(g23734),.A(g17974),.B(g23008));
  AND2 AND2_2518(.VSS(VSS),.VDD(VDD),.Y(g23735),.A(g22949),.B(g9450));
  AND2 AND2_2519(.VSS(VSS),.VDD(VDD),.Y(g23740),.A(g17993),.B(g23012));
  AND2 AND2_2520(.VSS(VSS),.VDD(VDD),.Y(g23741),.A(g22708),.B(g17667));
  AND2 AND2_2521(.VSS(VSS),.VDD(VDD),.Y(g23743),.A(g6777),.B(g23015));
  AND2 AND2_2522(.VSS(VSS),.VDD(VDD),.Y(g23747),.A(g18025),.B(g23016));
  AND2 AND2_2523(.VSS(VSS),.VDD(VDD),.Y(g23763),.A(g22865),.B(g17688));
  AND2 AND2_2524(.VSS(VSS),.VDD(VDD),.Y(g23768),.A(g4570),.B(g22629));
  AND2 AND2_2525(.VSS(VSS),.VDD(VDD),.Y(g23769),.A(g18048),.B(g23020));
  AND2 AND2_2526(.VSS(VSS),.VDD(VDD),.Y(g23770),.A(g22921),.B(g20454));
  AND2 AND2_2527(.VSS(VSS),.VDD(VDD),.Y(g23771),.A(g22720),.B(g20455));
  AND2 AND2_2528(.VSS(VSS),.VDD(VDD),.Y(g23772),.A(g21825),.B(g22875));
  AND2 AND2_2529(.VSS(VSS),.VDD(VDD),.Y(g23776),.A(g18074),.B(g23021));
  AND2 AND2_2530(.VSS(VSS),.VDD(VDD),.Y(g23777),.A(g22949),.B(g9528));
  AND2 AND2_2531(.VSS(VSS),.VDD(VDD),.Y(g23778),.A(g22954),.B(g9531));
  AND2 AND2_2532(.VSS(VSS),.VDD(VDD),.Y(g23789),.A(g18091),.B(g23024));
  AND2 AND2_2533(.VSS(VSS),.VDD(VDD),.Y(g23790),.A(g22958),.B(g9592));
  AND2 AND2_2534(.VSS(VSS),.VDD(VDD),.Y(g23795),.A(g18110),.B(g23028));
  AND2 AND2_2535(.VSS(VSS),.VDD(VDD),.Y(g23796),.A(g22739),.B(g17767));
  AND2 AND2_2536(.VSS(VSS),.VDD(VDD),.Y(g23798),.A(g7079),.B(g23031));
  AND2 AND2_2537(.VSS(VSS),.VDD(VDD),.Y(g23802),.A(g18142),.B(g23032));
  AND2 AND2_2538(.VSS(VSS),.VDD(VDD),.Y(g23818),.A(g22900),.B(g17788));
  AND2 AND2_2539(.VSS(VSS),.VDD(VDD),.Y(g23820),.A(g3013),.B(g23036));
  AND2 AND2_2540(.VSS(VSS),.VDD(VDD),.Y(g23822),.A(g14148),.B(g23037));
  AND2 AND2_2541(.VSS(VSS),.VDD(VDD),.Y(g23824),.A(g22949),.B(g9641));
  AND2 AND2_2542(.VSS(VSS),.VDD(VDD),.Y(g23825),.A(g22954),.B(g9644));
  AND2 AND2_2543(.VSS(VSS),.VDD(VDD),.Y(g23829),.A(g18190),.B(g23038));
  AND2 AND2_2544(.VSS(VSS),.VDD(VDD),.Y(g23830),.A(g22958),.B(g9670));
  AND2 AND2_2545(.VSS(VSS),.VDD(VDD),.Y(g23831),.A(g22962),.B(g9673));
  AND2 AND2_2546(.VSS(VSS),.VDD(VDD),.Y(g23842),.A(g18207),.B(g23041));
  AND2 AND2_2547(.VSS(VSS),.VDD(VDD),.Y(g23843),.A(g22966),.B(g9734));
  AND2 AND2_2548(.VSS(VSS),.VDD(VDD),.Y(g23848),.A(g18226),.B(g23045));
  AND2 AND2_2549(.VSS(VSS),.VDD(VDD),.Y(g23849),.A(g22771),.B(g17868));
  AND2 AND2_2550(.VSS(VSS),.VDD(VDD),.Y(g23851),.A(g7329),.B(g23048));
  AND2 AND2_2551(.VSS(VSS),.VDD(VDD),.Y(g23852),.A(g19179),.B(g22696));
  AND2 AND2_2552(.VSS(VSS),.VDD(VDD),.Y(g23854),.A(g18265),.B(g23049));
  AND2 AND2_2553(.VSS(VSS),.VDD(VDD),.Y(g23855),.A(g22954),.B(g9767));
  AND2 AND2_2554(.VSS(VSS),.VDD(VDD),.Y(g23857),.A(g14263),.B(g23056));
  AND2 AND2_2555(.VSS(VSS),.VDD(VDD),.Y(g23859),.A(g22958),.B(g9787));
  AND2 AND2_2556(.VSS(VSS),.VDD(VDD),.Y(g23860),.A(g22962),.B(g9790));
  AND2 AND2_2557(.VSS(VSS),.VDD(VDD),.Y(g23864),.A(g18297),.B(g23057));
  AND2 AND2_2558(.VSS(VSS),.VDD(VDD),.Y(g23865),.A(g22966),.B(g9816));
  AND2 AND2_2559(.VSS(VSS),.VDD(VDD),.Y(g23866),.A(g22971),.B(g9819));
  AND2 AND2_2560(.VSS(VSS),.VDD(VDD),.Y(g23877),.A(g18314),.B(g23060));
  AND2 AND2_2561(.VSS(VSS),.VDD(VDD),.Y(g23878),.A(g22975),.B(g9880));
  AND2 AND2_2562(.VSS(VSS),.VDD(VDD),.Y(g23886),.A(g18341),.B(g23064));
  AND2 AND2_2563(.VSS(VSS),.VDD(VDD),.Y(g23888),.A(g18358),.B(g23069));
  AND2 AND2_2564(.VSS(VSS),.VDD(VDD),.Y(g23889),.A(g22962),.B(g9913));
  AND2 AND2_2565(.VSS(VSS),.VDD(VDD),.Y(g23891),.A(g14385),.B(g23074));
  AND2 AND2_2566(.VSS(VSS),.VDD(VDD),.Y(g23893),.A(g22966),.B(g9933));
  AND2 AND2_2567(.VSS(VSS),.VDD(VDD),.Y(g23894),.A(g22971),.B(g9936));
  AND2 AND2_2568(.VSS(VSS),.VDD(VDD),.Y(g23898),.A(g18390),.B(g23075));
  AND2 AND2_2569(.VSS(VSS),.VDD(VDD),.Y(g23899),.A(g22975),.B(g9962));
  AND2 AND2_2570(.VSS(VSS),.VDD(VDD),.Y(g23900),.A(g22980),.B(g9965));
  AND2 AND2_2571(.VSS(VSS),.VDD(VDD),.Y(g23904),.A(g3010),.B(g22750));
  AND2 AND2_2572(.VSS(VSS),.VDD(VDD),.Y(g23907),.A(g18436),.B(g23079));
  AND2 AND2_2573(.VSS(VSS),.VDD(VDD),.Y(g23909),.A(g18453),.B(g23082));
  AND2 AND2_2574(.VSS(VSS),.VDD(VDD),.Y(g23910),.A(g22971),.B(g10067));
  AND2 AND2_2575(.VSS(VSS),.VDD(VDD),.Y(g23912),.A(g14497),.B(g23087));
  AND2 AND2_2576(.VSS(VSS),.VDD(VDD),.Y(g23914),.A(g22975),.B(g10087));
  AND2 AND2_2577(.VSS(VSS),.VDD(VDD),.Y(g23915),.A(g22980),.B(g10090));
  AND2 AND2_2578(.VSS(VSS),.VDD(VDD),.Y(g23917),.A(g7545),.B(g23088));
  AND2 AND2_2579(.VSS(VSS),.VDD(VDD),.Y(g23939),.A(g18509),.B(g23095));
  AND2 AND2_2580(.VSS(VSS),.VDD(VDD),.Y(g23941),.A(g18526),.B(g23098));
  AND2 AND2_2581(.VSS(VSS),.VDD(VDD),.Y(g23942),.A(g22980),.B(g10176));
  AND2 AND2_2582(.VSS(VSS),.VDD(VDD),.Y(g23944),.A(g7570),.B(g23103));
  AND2 AND2_2583(.VSS(VSS),.VDD(VDD),.Y(g23971),.A(g18573),.B(g23112));
  AND2 AND2_2584(.VSS(VSS),.VDD(VDD),.Y(g23972),.A(g2903),.B(g23115));
  AND2 AND2_2585(.VSS(VSS),.VDD(VDD),.Y(g24029),.A(g2900),.B(g22903));
  AND2 AND2_2586(.VSS(VSS),.VDD(VDD),.Y(g24211),.A(g22014),.B(g10969));
  AND2 AND2_2587(.VSS(VSS),.VDD(VDD),.Y(g24217),.A(g22825),.B(g10999));
  AND2 AND2_2588(.VSS(VSS),.VDD(VDD),.Y(g24221),.A(g22979),.B(g11042));
  AND2 AND2_2589(.VSS(VSS),.VDD(VDD),.Y(g24224),.A(g22219),.B(g11045));
  AND2 AND2_2590(.VSS(VSS),.VDD(VDD),.Y(g24229),.A(g22232),.B(g11105));
  AND2 AND2_2591(.VSS(VSS),.VDD(VDD),.Y(g24236),.A(g22243),.B(g11157));
  AND2 AND2_2592(.VSS(VSS),.VDD(VDD),.Y(g24241),.A(g22259),.B(g11228));
  AND2 AND2_2593(.VSS(VSS),.VDD(VDD),.Y(g24246),.A(g21982),.B(g11291));
  AND2 AND2_2594(.VSS(VSS),.VDD(VDD),.Y(g24247),.A(g22551),.B(g11297));
  AND2 AND2_2595(.VSS(VSS),.VDD(VDD),.Y(g24253),.A(g21995),.B(g11370));
  AND2 AND2_2596(.VSS(VSS),.VDD(VDD),.Y(g24256),.A(g22003),.B(g11438));
  AND3 AND3_221(.VSS(VSS),.VDD(VDD),.Y(g24427),.A(g17086),.B(g24134),.C(g13626));
  AND2 AND2_2597(.VSS(VSS),.VDD(VDD),.Y(g24429),.A(g24115),.B(g13614));
  AND3 AND3_222(.VSS(VSS),.VDD(VDD),.Y(g24431),.A(g17124),.B(g24153),.C(g13637));
  AND3 AND3_223(.VSS(VSS),.VDD(VDD),.Y(g24432),.A(g14642),.B(g15904),.C(g24115));
  AND2 AND2_2598(.VSS(VSS),.VDD(VDD),.Y(g24433),.A(g24134),.B(g13626));
  AND3 AND3_224(.VSS(VSS),.VDD(VDD),.Y(g24435),.A(g17151),.B(g24168),.C(g13649));
  AND3 AND3_225(.VSS(VSS),.VDD(VDD),.Y(g24436),.A(g14669),.B(g15933),.C(g24134));
  AND2 AND2_2599(.VSS(VSS),.VDD(VDD),.Y(g24437),.A(g24153),.B(g13637));
  AND3 AND3_226(.VSS(VSS),.VDD(VDD),.Y(g24439),.A(g14703),.B(g15962),.C(g24153));
  AND2 AND2_2600(.VSS(VSS),.VDD(VDD),.Y(g24440),.A(g24168),.B(g13649));
  AND3 AND3_227(.VSS(VSS),.VDD(VDD),.Y(g24441),.A(g14737),.B(g15981),.C(g24168));
  AND3 AND3_228(.VSS(VSS),.VDD(VDD),.Y(g24478),.A(g23545),.B(g21119),.C(g21227));
  AND3 AND3_229(.VSS(VSS),.VDD(VDD),.Y(g24529),.A(g19933),.B(g17896),.C(g23403));
  AND3 AND3_230(.VSS(VSS),.VDD(VDD),.Y(g24540),.A(g18548),.B(g23089),.C(g23403));
  AND3 AND3_231(.VSS(VSS),.VDD(VDD),.Y(g24541),.A(g23420),.B(g17896),.C(g23052));
  AND3 AND3_232(.VSS(VSS),.VDD(VDD),.Y(g24542),.A(g19950),.B(g18007),.C(g23410));
  AND3 AND3_233(.VSS(VSS),.VDD(VDD),.Y(g24550),.A(g18548),.B(g23420),.C(g19948));
  AND3 AND3_234(.VSS(VSS),.VDD(VDD),.Y(g24552),.A(g18598),.B(g23107),.C(g23410));
  AND3 AND3_235(.VSS(VSS),.VDD(VDD),.Y(g24553),.A(g23429),.B(g18007),.C(g23071));
  AND3 AND3_236(.VSS(VSS),.VDD(VDD),.Y(g24554),.A(g19977),.B(g18124),.C(g23415));
  AND2 AND2_2601(.VSS(VSS),.VDD(VDD),.Y(g24559),.A(g79),.B(g23448));
  AND3 AND3_237(.VSS(VSS),.VDD(VDD),.Y(g24561),.A(g18598),.B(g23429),.C(g19975));
  AND3 AND3_238(.VSS(VSS),.VDD(VDD),.Y(g24563),.A(g18630),.B(g23120),.C(g23415));
  AND3 AND3_239(.VSS(VSS),.VDD(VDD),.Y(g24564),.A(g23435),.B(g18124),.C(g23084));
  AND3 AND3_240(.VSS(VSS),.VDD(VDD),.Y(g24565),.A(g20007),.B(g18240),.C(g23424));
  AND2 AND2_2602(.VSS(VSS),.VDD(VDD),.Y(g24569),.A(g767),.B(g23455));
  AND3 AND3_241(.VSS(VSS),.VDD(VDD),.Y(g24571),.A(g18630),.B(g23435),.C(g20005));
  AND3 AND3_242(.VSS(VSS),.VDD(VDD),.Y(g24573),.A(g18639),.B(g23129),.C(g23424));
  AND3 AND3_243(.VSS(VSS),.VDD(VDD),.Y(g24574),.A(g23441),.B(g18240),.C(g23100));
  AND2 AND2_2603(.VSS(VSS),.VDD(VDD),.Y(g24578),.A(g1453),.B(g23464));
  AND3 AND3_244(.VSS(VSS),.VDD(VDD),.Y(g24580),.A(g18639),.B(g23441),.C(g20043));
  AND2 AND2_2604(.VSS(VSS),.VDD(VDD),.Y(g24585),.A(g2147),.B(g23473));
  AND2 AND2_2605(.VSS(VSS),.VDD(VDD),.Y(g24590),.A(g23486),.B(g23478));
  AND2 AND2_2606(.VSS(VSS),.VDD(VDD),.Y(g24591),.A(g83),.B(g23853));
  AND2 AND2_2607(.VSS(VSS),.VDD(VDD),.Y(g24595),.A(g23502),.B(g23489));
  AND2 AND2_2608(.VSS(VSS),.VDD(VDD),.Y(g24596),.A(g771),.B(g23887));
  AND2 AND2_2609(.VSS(VSS),.VDD(VDD),.Y(g24603),.A(g23518),.B(g23505));
  AND2 AND2_2610(.VSS(VSS),.VDD(VDD),.Y(g24604),.A(g1457),.B(g23908));
  AND2 AND2_2611(.VSS(VSS),.VDD(VDD),.Y(g24610),.A(g23533),.B(g23521));
  AND2 AND2_2612(.VSS(VSS),.VDD(VDD),.Y(g24611),.A(g2151),.B(g23940));
  AND2 AND2_2613(.VSS(VSS),.VDD(VDD),.Y(g24644),.A(g17203),.B(g24115));
  AND2 AND2_2614(.VSS(VSS),.VDD(VDD),.Y(g24664),.A(g17208),.B(g24134));
  AND2 AND2_2615(.VSS(VSS),.VDD(VDD),.Y(g24676),.A(g13568),.B(g24115));
  AND2 AND2_2616(.VSS(VSS),.VDD(VDD),.Y(g24683),.A(g17214),.B(g24153));
  AND2 AND2_2617(.VSS(VSS),.VDD(VDD),.Y(g24695),.A(g13576),.B(g24134));
  AND2 AND2_2618(.VSS(VSS),.VDD(VDD),.Y(g24700),.A(g17217),.B(g24168));
  AND2 AND2_2619(.VSS(VSS),.VDD(VDD),.Y(g24712),.A(g13585),.B(g24153));
  AND2 AND2_2620(.VSS(VSS),.VDD(VDD),.Y(g24723),.A(g13605),.B(g24168));
  AND2 AND2_2621(.VSS(VSS),.VDD(VDD),.Y(g24745),.A(g15454),.B(g24096));
  AND2 AND2_2622(.VSS(VSS),.VDD(VDD),.Y(g24746),.A(g15454),.B(g24098));
  AND2 AND2_2623(.VSS(VSS),.VDD(VDD),.Y(g24747),.A(g9427),.B(g24099));
  AND2 AND2_2624(.VSS(VSS),.VDD(VDD),.Y(g24748),.A(g672),.B(g24101));
  AND2 AND2_2625(.VSS(VSS),.VDD(VDD),.Y(g24749),.A(g15540),.B(g24102));
  AND2 AND2_2626(.VSS(VSS),.VDD(VDD),.Y(g24750),.A(g15454),.B(g24104));
  AND2 AND2_2627(.VSS(VSS),.VDD(VDD),.Y(g24751),.A(g9427),.B(g24105));
  AND2 AND2_2628(.VSS(VSS),.VDD(VDD),.Y(g24752),.A(g9507),.B(g24106));
  AND2 AND2_2629(.VSS(VSS),.VDD(VDD),.Y(g24754),.A(g15540),.B(g24107));
  AND2 AND2_2630(.VSS(VSS),.VDD(VDD),.Y(g24755),.A(g9569),.B(g24108));
  AND2 AND2_2631(.VSS(VSS),.VDD(VDD),.Y(g24757),.A(g1358),.B(g24110));
  AND2 AND2_2632(.VSS(VSS),.VDD(VDD),.Y(g24758),.A(g15618),.B(g24111));
  AND2 AND2_2633(.VSS(VSS),.VDD(VDD),.Y(g24759),.A(g21825),.B(g23885));
  AND2 AND2_2634(.VSS(VSS),.VDD(VDD),.Y(g24760),.A(g9427),.B(g24112));
  AND2 AND2_2635(.VSS(VSS),.VDD(VDD),.Y(g24761),.A(g9507),.B(g24113));
  AND2 AND2_2636(.VSS(VSS),.VDD(VDD),.Y(g24762),.A(g12876),.B(g24114));
  AND2 AND2_2637(.VSS(VSS),.VDD(VDD),.Y(g24767),.A(g15540),.B(g24121));
  AND2 AND2_2638(.VSS(VSS),.VDD(VDD),.Y(g24768),.A(g9569),.B(g24122));
  AND2 AND2_2639(.VSS(VSS),.VDD(VDD),.Y(g24769),.A(g9649),.B(g24123));
  AND2 AND2_2640(.VSS(VSS),.VDD(VDD),.Y(g24772),.A(g15618),.B(g24124));
  AND2 AND2_2641(.VSS(VSS),.VDD(VDD),.Y(g24773),.A(g9711),.B(g24125));
  AND2 AND2_2642(.VSS(VSS),.VDD(VDD),.Y(g24774),.A(g2052),.B(g24127));
  AND2 AND2_2643(.VSS(VSS),.VDD(VDD),.Y(g24775),.A(g15694),.B(g24128));
  AND2 AND2_2644(.VSS(VSS),.VDD(VDD),.Y(g24776),.A(g9507),.B(g24129));
  AND2 AND2_2645(.VSS(VSS),.VDD(VDD),.Y(g24777),.A(g12876),.B(g24130));
  AND2 AND2_2646(.VSS(VSS),.VDD(VDD),.Y(g24779),.A(g9569),.B(g24131));
  AND2 AND2_2647(.VSS(VSS),.VDD(VDD),.Y(g24780),.A(g9649),.B(g24132));
  AND2 AND2_2648(.VSS(VSS),.VDD(VDD),.Y(g24781),.A(g12916),.B(g24133));
  AND2 AND2_2649(.VSS(VSS),.VDD(VDD),.Y(g24788),.A(g15618),.B(g24140));
  AND2 AND2_2650(.VSS(VSS),.VDD(VDD),.Y(g24789),.A(g9711),.B(g24141));
  AND2 AND2_2651(.VSS(VSS),.VDD(VDD),.Y(g24790),.A(g9795),.B(g24142));
  AND2 AND2_2652(.VSS(VSS),.VDD(VDD),.Y(g24792),.A(g15694),.B(g24143));
  AND2 AND2_2653(.VSS(VSS),.VDD(VDD),.Y(g24793),.A(g9857),.B(g24144));
  AND2 AND2_2654(.VSS(VSS),.VDD(VDD),.Y(g24794),.A(g2746),.B(g24146));
  AND2 AND2_2655(.VSS(VSS),.VDD(VDD),.Y(g24795),.A(g12017),.B(g24232));
  AND2 AND2_2656(.VSS(VSS),.VDD(VDD),.Y(g24796),.A(g12876),.B(g24147));
  AND2 AND2_2657(.VSS(VSS),.VDD(VDD),.Y(g24798),.A(g9649),.B(g24148));
  AND2 AND2_2658(.VSS(VSS),.VDD(VDD),.Y(g24799),.A(g12916),.B(g24149));
  AND2 AND2_2659(.VSS(VSS),.VDD(VDD),.Y(g24802),.A(g9711),.B(g24150));
  AND2 AND2_2660(.VSS(VSS),.VDD(VDD),.Y(g24803),.A(g9795),.B(g24151));
  AND2 AND2_2661(.VSS(VSS),.VDD(VDD),.Y(g24804),.A(g12945),.B(g24152));
  AND2 AND2_2662(.VSS(VSS),.VDD(VDD),.Y(g24809),.A(g15694),.B(g24159));
  AND2 AND2_2663(.VSS(VSS),.VDD(VDD),.Y(g24810),.A(g9857),.B(g24160));
  AND2 AND2_2664(.VSS(VSS),.VDD(VDD),.Y(g24811),.A(g9941),.B(g24161));
  AND2 AND2_2665(.VSS(VSS),.VDD(VDD),.Y(g24813),.A(g21825),.B(g23905));
  AND2 AND2_2666(.VSS(VSS),.VDD(VDD),.Y(g24818),.A(g12916),.B(g24162));
  AND2 AND2_2667(.VSS(VSS),.VDD(VDD),.Y(g24821),.A(g9795),.B(g24163));
  AND2 AND2_2668(.VSS(VSS),.VDD(VDD),.Y(g24822),.A(g12945),.B(g24164));
  AND2 AND2_2669(.VSS(VSS),.VDD(VDD),.Y(g24824),.A(g9857),.B(g24165));
  AND2 AND2_2670(.VSS(VSS),.VDD(VDD),.Y(g24825),.A(g9941),.B(g24166));
  AND2 AND2_2671(.VSS(VSS),.VDD(VDD),.Y(g24826),.A(g12974),.B(g24167));
  AND2 AND2_2672(.VSS(VSS),.VDD(VDD),.Y(g24831),.A(g24100),.B(g20401));
  AND2 AND2_2673(.VSS(VSS),.VDD(VDD),.Y(g24838),.A(g12945),.B(g24175));
  AND2 AND2_2674(.VSS(VSS),.VDD(VDD),.Y(g24840),.A(g9941),.B(g24176));
  AND2 AND2_2675(.VSS(VSS),.VDD(VDD),.Y(g24841),.A(g12974),.B(g24177));
  AND2 AND2_2676(.VSS(VSS),.VDD(VDD),.Y(g24843),.A(g21825),.B(g23918));
  AND2 AND2_2677(.VSS(VSS),.VDD(VDD),.Y(g24846),.A(g24109),.B(g20426));
  AND2 AND2_2678(.VSS(VSS),.VDD(VDD),.Y(g24853),.A(g12974),.B(g24180));
  AND2 AND2_2679(.VSS(VSS),.VDD(VDD),.Y(g24855),.A(g18174),.B(g23731));
  AND2 AND2_2680(.VSS(VSS),.VDD(VDD),.Y(g24858),.A(g24047),.B(g18873));
  AND2 AND2_2681(.VSS(VSS),.VDD(VDD),.Y(g24861),.A(g24126),.B(g20448));
  AND2 AND2_2682(.VSS(VSS),.VDD(VDD),.Y(g24867),.A(g666),.B(g23779));
  AND2 AND2_2683(.VSS(VSS),.VDD(VDD),.Y(g24869),.A(g24047),.B(g18894));
  AND2 AND2_2684(.VSS(VSS),.VDD(VDD),.Y(g24870),.A(g18281),.B(g23786));
  AND2 AND2_2685(.VSS(VSS),.VDD(VDD),.Y(g24874),.A(g24060),.B(g18899));
  AND2 AND2_2686(.VSS(VSS),.VDD(VDD),.Y(g24876),.A(g24145),.B(g20467));
  AND2 AND2_2687(.VSS(VSS),.VDD(VDD),.Y(g24878),.A(g19830),.B(g24210));
  AND2 AND2_2688(.VSS(VSS),.VDD(VDD),.Y(g24881),.A(g24047),.B(g18912));
  AND2 AND2_2689(.VSS(VSS),.VDD(VDD),.Y(g24882),.A(g1352),.B(g23832));
  AND2 AND2_2690(.VSS(VSS),.VDD(VDD),.Y(g24884),.A(g24060),.B(g18917));
  AND2 AND2_2691(.VSS(VSS),.VDD(VDD),.Y(g24885),.A(g18374),.B(g23839));
  AND2 AND2_2692(.VSS(VSS),.VDD(VDD),.Y(g24888),.A(g24073),.B(g18922));
  AND2 AND2_2693(.VSS(VSS),.VDD(VDD),.Y(g24898),.A(g24060),.B(g18931));
  AND2 AND2_2694(.VSS(VSS),.VDD(VDD),.Y(g24899),.A(g2046),.B(g23867));
  AND2 AND2_2695(.VSS(VSS),.VDD(VDD),.Y(g24901),.A(g24073),.B(g18936));
  AND2 AND2_2696(.VSS(VSS),.VDD(VDD),.Y(g24902),.A(g18469),.B(g23874));
  AND2 AND2_2697(.VSS(VSS),.VDD(VDD),.Y(g24905),.A(g24084),.B(g18941));
  AND2 AND2_2698(.VSS(VSS),.VDD(VDD),.Y(g24906),.A(g18886),.B(g23879));
  AND2 AND2_2699(.VSS(VSS),.VDD(VDD),.Y(g24907),.A(g7466),.B(g24220));
  AND2 AND2_2700(.VSS(VSS),.VDD(VDD),.Y(g24908),.A(g7342),.B(g23882));
  AND2 AND2_2701(.VSS(VSS),.VDD(VDD),.Y(g24921),.A(g24073),.B(g18951));
  AND2 AND2_2702(.VSS(VSS),.VDD(VDD),.Y(g24922),.A(g2740),.B(g23901));
  AND2 AND2_2703(.VSS(VSS),.VDD(VDD),.Y(g24924),.A(g24084),.B(g18956));
  AND2 AND2_2704(.VSS(VSS),.VDD(VDD),.Y(g24938),.A(g24084),.B(g18967));
  AND2 AND2_2705(.VSS(VSS),.VDD(VDD),.Y(g24964),.A(g7595),.B(g24251));
  AND2 AND2_2706(.VSS(VSS),.VDD(VDD),.Y(g24974),.A(g7600),.B(g24030));
  AND2 AND2_2707(.VSS(VSS),.VDD(VDD),.Y(g25086),.A(g23444),.B(g10880));
  AND2 AND2_2708(.VSS(VSS),.VDD(VDD),.Y(g25102),.A(g23444),.B(g10915));
  AND2 AND2_2709(.VSS(VSS),.VDD(VDD),.Y(g25117),.A(g23444),.B(g10974));
  AND3 AND3_245(.VSS(VSS),.VDD(VDD),.Y(g25128),.A(g17051),.B(g24115),.C(g13614));
  AND2 AND2_2710(.VSS(VSS),.VDD(VDD),.Y(g25178),.A(g24623),.B(g20634));
  AND2 AND2_2711(.VSS(VSS),.VDD(VDD),.Y(g25181),.A(g24636),.B(g20673));
  AND2 AND2_2712(.VSS(VSS),.VDD(VDD),.Y(g25182),.A(g24681),.B(g20676));
  AND2 AND2_2713(.VSS(VSS),.VDD(VDD),.Y(g25184),.A(g24694),.B(g20735));
  AND2 AND2_2714(.VSS(VSS),.VDD(VDD),.Y(g25187),.A(g24633),.B(g16608));
  AND2 AND2_2715(.VSS(VSS),.VDD(VDD),.Y(g25188),.A(g24652),.B(g20763));
  AND2 AND2_2716(.VSS(VSS),.VDD(VDD),.Y(g25192),.A(g24711),.B(g20790));
  AND2 AND2_2717(.VSS(VSS),.VDD(VDD),.Y(g25193),.A(g24653),.B(g16626));
  AND2 AND2_2718(.VSS(VSS),.VDD(VDD),.Y(g25196),.A(g24672),.B(g16640));
  AND2 AND2_2719(.VSS(VSS),.VDD(VDD),.Y(g25198),.A(g24691),.B(g16651));
  AND2 AND2_2720(.VSS(VSS),.VDD(VDD),.Y(g25269),.A(g24648),.B(g8700));
  AND2 AND2_2721(.VSS(VSS),.VDD(VDD),.Y(g25277),.A(g24648),.B(g8714));
  AND2 AND2_2722(.VSS(VSS),.VDD(VDD),.Y(g25278),.A(g24668),.B(g8719));
  AND2 AND2_2723(.VSS(VSS),.VDD(VDD),.Y(g25281),.A(g5606),.B(g24815));
  AND2 AND2_2724(.VSS(VSS),.VDD(VDD),.Y(g25282),.A(g24648),.B(g8748));
  AND2 AND2_2725(.VSS(VSS),.VDD(VDD),.Y(g25286),.A(g24668),.B(g8752));
  AND2 AND2_2726(.VSS(VSS),.VDD(VDD),.Y(g25287),.A(g24687),.B(g8757));
  AND2 AND2_2727(.VSS(VSS),.VDD(VDD),.Y(g25289),.A(g5631),.B(g24834));
  AND2 AND2_2728(.VSS(VSS),.VDD(VDD),.Y(g25290),.A(g24668),.B(g8771));
  AND2 AND2_2729(.VSS(VSS),.VDD(VDD),.Y(g25294),.A(g24687),.B(g8775));
  AND2 AND2_2730(.VSS(VSS),.VDD(VDD),.Y(g25295),.A(g24704),.B(g8780));
  AND2 AND2_2731(.VSS(VSS),.VDD(VDD),.Y(g25299),.A(g5659),.B(g24850));
  AND2 AND2_2732(.VSS(VSS),.VDD(VDD),.Y(g25300),.A(g24687),.B(g8794));
  AND2 AND2_2733(.VSS(VSS),.VDD(VDD),.Y(g25304),.A(g24704),.B(g8798));
  AND2 AND2_2734(.VSS(VSS),.VDD(VDD),.Y(g25309),.A(g5697),.B(g24864));
  AND2 AND2_2735(.VSS(VSS),.VDD(VDD),.Y(g25310),.A(g24704),.B(g8813));
  AND3 AND3_246(.VSS(VSS),.VDD(VDD),.Y(g25318),.A(g24682),.B(g19358),.C(g19335));
  AND2 AND2_2736(.VSS(VSS),.VDD(VDD),.Y(g25321),.A(g25075),.B(g9669));
  AND2 AND2_2737(.VSS(VSS),.VDD(VDD),.Y(g25328),.A(g24644),.B(g17892));
  AND2 AND2_2738(.VSS(VSS),.VDD(VDD),.Y(g25334),.A(g24644),.B(g17984));
  AND2 AND2_2739(.VSS(VSS),.VDD(VDD),.Y(g25337),.A(g24664),.B(g18003));
  AND2 AND2_2740(.VSS(VSS),.VDD(VDD),.Y(g25342),.A(g5851),.B(g24600));
  AND2 AND2_2741(.VSS(VSS),.VDD(VDD),.Y(g25346),.A(g24644),.B(g18084));
  AND2 AND2_2742(.VSS(VSS),.VDD(VDD),.Y(g25348),.A(g24664),.B(g18101));
  AND2 AND2_2743(.VSS(VSS),.VDD(VDD),.Y(g25351),.A(g24683),.B(g18120));
  AND2 AND2_2744(.VSS(VSS),.VDD(VDD),.Y(g25356),.A(g5898),.B(g24607));
  AND2 AND2_2745(.VSS(VSS),.VDD(VDD),.Y(g25360),.A(g24664),.B(g18200));
  AND2 AND2_2746(.VSS(VSS),.VDD(VDD),.Y(g25362),.A(g24683),.B(g18217));
  AND2 AND2_2747(.VSS(VSS),.VDD(VDD),.Y(g25365),.A(g24700),.B(g18236));
  AND2 AND2_2748(.VSS(VSS),.VDD(VDD),.Y(g25371),.A(g5937),.B(g24619));
  AND2 AND2_2749(.VSS(VSS),.VDD(VDD),.Y(g25375),.A(g24683),.B(g18307));
  AND2 AND2_2750(.VSS(VSS),.VDD(VDD),.Y(g25377),.A(g24700),.B(g18324));
  AND2 AND2_2751(.VSS(VSS),.VDD(VDD),.Y(g25388),.A(g5971),.B(g24630));
  AND2 AND2_2752(.VSS(VSS),.VDD(VDD),.Y(g25392),.A(g24700),.B(g18400));
  AND2 AND2_2753(.VSS(VSS),.VDD(VDD),.Y(g25453),.A(g6142),.B(g24763));
  AND2 AND2_2754(.VSS(VSS),.VDD(VDD),.Y(g25457),.A(g6163),.B(g24784));
  AND2 AND2_2755(.VSS(VSS),.VDD(VDD),.Y(g25461),.A(g6190),.B(g24805));
  AND2 AND2_2756(.VSS(VSS),.VDD(VDD),.Y(g25466),.A(g6222),.B(g24827));
  AND2 AND2_2757(.VSS(VSS),.VDD(VDD),.Y(g25470),.A(g24479),.B(g20400));
  AND2 AND2_2758(.VSS(VSS),.VDD(VDD),.Y(g25475),.A(g14148),.B(g25087));
  AND2 AND2_2759(.VSS(VSS),.VDD(VDD),.Y(g25482),.A(g24480),.B(g17567));
  AND2 AND2_2760(.VSS(VSS),.VDD(VDD),.Y(g25483),.A(g24481),.B(g20421));
  AND2 AND2_2761(.VSS(VSS),.VDD(VDD),.Y(g25487),.A(g24485),.B(g20425));
  AND2 AND2_2762(.VSS(VSS),.VDD(VDD),.Y(g25505),.A(g6707),.B(g25094));
  AND2 AND2_2763(.VSS(VSS),.VDD(VDD),.Y(g25506),.A(g14263),.B(g25095));
  AND2 AND2_2764(.VSS(VSS),.VDD(VDD),.Y(g25513),.A(g24487),.B(g17664));
  AND2 AND2_2765(.VSS(VSS),.VDD(VDD),.Y(g25514),.A(g24488),.B(g20443));
  AND2 AND2_2766(.VSS(VSS),.VDD(VDD),.Y(g25518),.A(g24489),.B(g20447));
  AND2 AND2_2767(.VSS(VSS),.VDD(VDD),.Y(g25552),.A(g7009),.B(g25104));
  AND2 AND2_2768(.VSS(VSS),.VDD(VDD),.Y(g25553),.A(g14385),.B(g25105));
  AND2 AND2_2769(.VSS(VSS),.VDD(VDD),.Y(g25560),.A(g24494),.B(g17764));
  AND2 AND2_2770(.VSS(VSS),.VDD(VDD),.Y(g25561),.A(g24495),.B(g20462));
  AND2 AND2_2771(.VSS(VSS),.VDD(VDD),.Y(g25565),.A(g24496),.B(g20466));
  AND2 AND2_2772(.VSS(VSS),.VDD(VDD),.Y(g25618),.A(g7259),.B(g25110));
  AND2 AND2_2773(.VSS(VSS),.VDD(VDD),.Y(g25619),.A(g14497),.B(g25111));
  AND2 AND2_2774(.VSS(VSS),.VDD(VDD),.Y(g25626),.A(g24504),.B(g17865));
  AND2 AND2_2775(.VSS(VSS),.VDD(VDD),.Y(g25627),.A(g24505),.B(g20477));
  AND2 AND2_2776(.VSS(VSS),.VDD(VDD),.Y(g25628),.A(g21008),.B(g25115));
  AND2 AND2_2777(.VSS(VSS),.VDD(VDD),.Y(g25629),.A(g3024),.B(g25116));
  AND2 AND2_2778(.VSS(VSS),.VDD(VDD),.Y(g25697),.A(g7455),.B(g25120));
  AND2 AND2_2779(.VSS(VSS),.VDD(VDD),.Y(g25881),.A(g2908),.B(g25126));
  AND2 AND2_2780(.VSS(VSS),.VDD(VDD),.Y(g25951),.A(g24800),.B(g13670));
  AND2 AND2_2781(.VSS(VSS),.VDD(VDD),.Y(g25953),.A(g24783),.B(g13699));
  AND2 AND2_2782(.VSS(VSS),.VDD(VDD),.Y(g25957),.A(g24782),.B(g11869));
  AND2 AND2_2783(.VSS(VSS),.VDD(VDD),.Y(g25961),.A(g24770),.B(g11901));
  AND2 AND2_2784(.VSS(VSS),.VDD(VDD),.Y(g25963),.A(g24756),.B(g11944));
  AND2 AND2_2785(.VSS(VSS),.VDD(VDD),.Y(g25968),.A(g24871),.B(g11986));
  AND2 AND2_2786(.VSS(VSS),.VDD(VDD),.Y(g25972),.A(g24859),.B(g12042));
  AND2 AND2_2787(.VSS(VSS),.VDD(VDD),.Y(g25973),.A(g24847),.B(g13838));
  AND2 AND2_2788(.VSS(VSS),.VDD(VDD),.Y(g25975),.A(g24606),.B(g21917));
  AND2 AND2_2789(.VSS(VSS),.VDD(VDD),.Y(g25977),.A(g24845),.B(g12089));
  AND2 AND2_2790(.VSS(VSS),.VDD(VDD),.Y(g25978),.A(g24836),.B(g13850));
  AND2 AND2_2791(.VSS(VSS),.VDD(VDD),.Y(g25980),.A(g24663),.B(g21928));
  AND2 AND2_2792(.VSS(VSS),.VDD(VDD),.Y(g25981),.A(g24819),.B(g13858));
  AND2 AND2_2793(.VSS(VSS),.VDD(VDD),.Y(g26023),.A(g25422),.B(g24912));
  AND2 AND2_2794(.VSS(VSS),.VDD(VDD),.Y(g26024),.A(g25301),.B(g21102));
  AND2 AND2_2795(.VSS(VSS),.VDD(VDD),.Y(g26026),.A(g25431),.B(g24929));
  AND2 AND2_2796(.VSS(VSS),.VDD(VDD),.Y(g26027),.A(g25418),.B(g22271));
  AND2 AND2_2797(.VSS(VSS),.VDD(VDD),.Y(g26028),.A(g25438),.B(g24941));
  AND2 AND2_2798(.VSS(VSS),.VDD(VDD),.Y(g26029),.A(g25445),.B(g24952));
  AND2 AND2_2799(.VSS(VSS),.VDD(VDD),.Y(g26030),.A(g25429),.B(g22304));
  AND2 AND2_2800(.VSS(VSS),.VDD(VDD),.Y(g26032),.A(g25379),.B(g19415));
  AND2 AND2_2801(.VSS(VSS),.VDD(VDD),.Y(g26033),.A(g25395),.B(g19452));
  AND2 AND2_2802(.VSS(VSS),.VDD(VDD),.Y(g26034),.A(g25405),.B(g19479));
  AND2 AND2_2803(.VSS(VSS),.VDD(VDD),.Y(g26035),.A(g25523),.B(g19483));
  AND2 AND2_2804(.VSS(VSS),.VDD(VDD),.Y(g26036),.A(g25413),.B(g19502));
  AND2 AND2_2805(.VSS(VSS),.VDD(VDD),.Y(g26038),.A(g25589),.B(g19504));
  AND2 AND2_2806(.VSS(VSS),.VDD(VDD),.Y(g26039),.A(g25668),.B(g19523));
  AND2 AND2_2807(.VSS(VSS),.VDD(VDD),.Y(g26040),.A(g25745),.B(g19533));
  AND2 AND2_2808(.VSS(VSS),.VDD(VDD),.Y(g26051),.A(g70),.B(g25296));
  AND2 AND2_2809(.VSS(VSS),.VDD(VDD),.Y(g26052),.A(g25941),.B(g21087));
  AND2 AND2_2810(.VSS(VSS),.VDD(VDD),.Y(g26053),.A(g758),.B(g25306));
  AND2 AND2_2811(.VSS(VSS),.VDD(VDD),.Y(g26054),.A(g25944),.B(g21099));
  AND2 AND2_2812(.VSS(VSS),.VDD(VDD),.Y(g26060),.A(g25943),.B(g21108));
  AND2 AND2_2813(.VSS(VSS),.VDD(VDD),.Y(g26061),.A(g1444),.B(g25315));
  AND2 AND2_2814(.VSS(VSS),.VDD(VDD),.Y(g26062),.A(g25947),.B(g21113));
  AND2 AND2_2815(.VSS(VSS),.VDD(VDD),.Y(g26067),.A(g25946),.B(g21125));
  AND2 AND2_2816(.VSS(VSS),.VDD(VDD),.Y(g26068),.A(g2138),.B(g25324));
  AND2 AND2_2817(.VSS(VSS),.VDD(VDD),.Y(g26069),.A(g25949),.B(g21130));
  AND2 AND2_2818(.VSS(VSS),.VDD(VDD),.Y(g26074),.A(g25948),.B(g21144));
  AND2 AND2_2819(.VSS(VSS),.VDD(VDD),.Y(g26075),.A(g74),.B(g25698));
  AND2 AND2_2820(.VSS(VSS),.VDD(VDD),.Y(g26080),.A(g25950),.B(g21164));
  AND2 AND2_2821(.VSS(VSS),.VDD(VDD),.Y(g26082),.A(g762),.B(g25771));
  AND2 AND2_2822(.VSS(VSS),.VDD(VDD),.Y(g26085),.A(g1448),.B(g25825));
  AND2 AND2_2823(.VSS(VSS),.VDD(VDD),.Y(g26091),.A(g2142),.B(g25860));
  AND2 AND2_2824(.VSS(VSS),.VDD(VDD),.Y(g26157),.A(g21825),.B(g25630));
  AND2 AND2_2825(.VSS(VSS),.VDD(VDD),.Y(g26158),.A(g679),.B(g25937));
  AND2 AND2_2826(.VSS(VSS),.VDD(VDD),.Y(g26163),.A(g1365),.B(g25939));
  AND2 AND2_2827(.VSS(VSS),.VDD(VDD),.Y(g26166),.A(g686),.B(g25454));
  AND2 AND2_2828(.VSS(VSS),.VDD(VDD),.Y(g26171),.A(g2059),.B(g25942));
  AND2 AND2_2829(.VSS(VSS),.VDD(VDD),.Y(g26186),.A(g1372),.B(g25458));
  AND2 AND2_2830(.VSS(VSS),.VDD(VDD),.Y(g26188),.A(g2753),.B(g25945));
  AND2 AND2_2831(.VSS(VSS),.VDD(VDD),.Y(g26207),.A(g2066),.B(g25463));
  AND2 AND2_2832(.VSS(VSS),.VDD(VDD),.Y(g26212),.A(g4217),.B(g25467));
  AND2 AND2_2833(.VSS(VSS),.VDD(VDD),.Y(g26213),.A(g25895),.B(g9306));
  AND2 AND2_2834(.VSS(VSS),.VDD(VDD),.Y(g26231),.A(g2760),.B(g25472));
  AND2 AND2_2835(.VSS(VSS),.VDD(VDD),.Y(g26233),.A(g4340),.B(g25476));
  AND2 AND2_2836(.VSS(VSS),.VDD(VDD),.Y(g26234),.A(g4343),.B(g25479));
  AND2 AND2_2837(.VSS(VSS),.VDD(VDD),.Y(g26235),.A(g25895),.B(g9368));
  AND2 AND2_2838(.VSS(VSS),.VDD(VDD),.Y(g26236),.A(g25899),.B(g9371));
  AND2 AND2_2839(.VSS(VSS),.VDD(VDD),.Y(g26243),.A(g4372),.B(g25484));
  AND2 AND2_2840(.VSS(VSS),.VDD(VDD),.Y(g26244),.A(g25903),.B(g9387));
  AND2 AND2_2841(.VSS(VSS),.VDD(VDD),.Y(g26257),.A(g4465),.B(g25493));
  AND2 AND2_2842(.VSS(VSS),.VDD(VDD),.Y(g26258),.A(g4468),.B(g25496));
  AND2 AND2_2843(.VSS(VSS),.VDD(VDD),.Y(g26259),.A(g4471),.B(g25499));
  AND2 AND2_2844(.VSS(VSS),.VDD(VDD),.Y(g26260),.A(g25254),.B(g17649));
  AND2 AND2_2845(.VSS(VSS),.VDD(VDD),.Y(g26261),.A(g25895),.B(g9443));
  AND2 AND2_2846(.VSS(VSS),.VDD(VDD),.Y(g26262),.A(g25899),.B(g9446));
  AND2 AND2_2847(.VSS(VSS),.VDD(VDD),.Y(g26263),.A(g4476),.B(g25502));
  AND2 AND2_2848(.VSS(VSS),.VDD(VDD),.Y(g26268),.A(g4509),.B(g25507));
  AND2 AND2_2849(.VSS(VSS),.VDD(VDD),.Y(g26269),.A(g4512),.B(g25510));
  AND2 AND2_2850(.VSS(VSS),.VDD(VDD),.Y(g26270),.A(g25903),.B(g9465));
  AND2 AND2_2851(.VSS(VSS),.VDD(VDD),.Y(g26271),.A(g25907),.B(g9468));
  AND2 AND2_2852(.VSS(VSS),.VDD(VDD),.Y(g26278),.A(g4541),.B(g25515));
  AND2 AND2_2853(.VSS(VSS),.VDD(VDD),.Y(g26279),.A(g25911),.B(g9484));
  AND2 AND2_2854(.VSS(VSS),.VDD(VDD),.Y(g26288),.A(g4592),.B(g25524));
  AND2 AND2_2855(.VSS(VSS),.VDD(VDD),.Y(g26289),.A(g4595),.B(g25527));
  AND2 AND2_2856(.VSS(VSS),.VDD(VDD),.Y(g26290),.A(g4598),.B(g25530));
  AND2 AND2_2857(.VSS(VSS),.VDD(VDD),.Y(g26291),.A(g25899),.B(g9524));
  AND2 AND2_2858(.VSS(VSS),.VDD(VDD),.Y(g26292),.A(g4603),.B(g25533));
  AND2 AND2_2859(.VSS(VSS),.VDD(VDD),.Y(g26293),.A(g4606),.B(g25536));
  AND2 AND2_2860(.VSS(VSS),.VDD(VDD),.Y(g26298),.A(g4641),.B(g25540));
  AND2 AND2_2861(.VSS(VSS),.VDD(VDD),.Y(g26299),.A(g4644),.B(g25543));
  AND2 AND2_2862(.VSS(VSS),.VDD(VDD),.Y(g26300),.A(g4647),.B(g25546));
  AND2 AND2_2863(.VSS(VSS),.VDD(VDD),.Y(g26301),.A(g25258),.B(g17749));
  AND2 AND2_2864(.VSS(VSS),.VDD(VDD),.Y(g26302),.A(g25903),.B(g9585));
  AND2 AND2_2865(.VSS(VSS),.VDD(VDD),.Y(g26303),.A(g25907),.B(g9588));
  AND2 AND2_2866(.VSS(VSS),.VDD(VDD),.Y(g26307),.A(g4652),.B(g25549));
  AND2 AND2_2867(.VSS(VSS),.VDD(VDD),.Y(g26309),.A(g4685),.B(g25554));
  AND2 AND2_2868(.VSS(VSS),.VDD(VDD),.Y(g26310),.A(g4688),.B(g25557));
  AND2 AND2_2869(.VSS(VSS),.VDD(VDD),.Y(g26311),.A(g25911),.B(g9607));
  AND2 AND2_2870(.VSS(VSS),.VDD(VDD),.Y(g26312),.A(g25915),.B(g9610));
  AND2 AND2_2871(.VSS(VSS),.VDD(VDD),.Y(g26316),.A(g4717),.B(g25562));
  AND2 AND2_2872(.VSS(VSS),.VDD(VDD),.Y(g26317),.A(g25919),.B(g9626));
  AND2 AND2_2873(.VSS(VSS),.VDD(VDD),.Y(g26318),.A(g4737),.B(g25573));
  AND2 AND2_2874(.VSS(VSS),.VDD(VDD),.Y(g26319),.A(g4740),.B(g25576));
  AND2 AND2_2875(.VSS(VSS),.VDD(VDD),.Y(g26324),.A(g4743),.B(g25579));
  AND2 AND2_2876(.VSS(VSS),.VDD(VDD),.Y(g26325),.A(g4746),.B(g25582));
  AND2 AND2_2877(.VSS(VSS),.VDD(VDD),.Y(g26326),.A(g4749),.B(g25585));
  AND2 AND2_2878(.VSS(VSS),.VDD(VDD),.Y(g26332),.A(g4769),.B(g25590));
  AND2 AND2_2879(.VSS(VSS),.VDD(VDD),.Y(g26333),.A(g4772),.B(g25593));
  AND2 AND2_2880(.VSS(VSS),.VDD(VDD),.Y(g26334),.A(g4775),.B(g25596));
  AND2 AND2_2881(.VSS(VSS),.VDD(VDD),.Y(g26335),.A(g25907),.B(g9666));
  AND2 AND2_2882(.VSS(VSS),.VDD(VDD),.Y(g26339),.A(g4780),.B(g25599));
  AND2 AND2_2883(.VSS(VSS),.VDD(VDD),.Y(g26340),.A(g4783),.B(g25602));
  AND2 AND2_2884(.VSS(VSS),.VDD(VDD),.Y(g26342),.A(g4818),.B(g25606));
  AND2 AND2_2885(.VSS(VSS),.VDD(VDD),.Y(g26343),.A(g4821),.B(g25609));
  AND2 AND2_2886(.VSS(VSS),.VDD(VDD),.Y(g26344),.A(g4824),.B(g25612));
  AND2 AND2_2887(.VSS(VSS),.VDD(VDD),.Y(g26345),.A(g25261),.B(g17850));
  AND2 AND2_2888(.VSS(VSS),.VDD(VDD),.Y(g26346),.A(g25911),.B(g9727));
  AND2 AND2_2889(.VSS(VSS),.VDD(VDD),.Y(g26347),.A(g25915),.B(g9730));
  AND2 AND2_2890(.VSS(VSS),.VDD(VDD),.Y(g26348),.A(g4829),.B(g25615));
  AND2 AND2_2891(.VSS(VSS),.VDD(VDD),.Y(g26350),.A(g4862),.B(g25620));
  AND2 AND2_2892(.VSS(VSS),.VDD(VDD),.Y(g26351),.A(g4865),.B(g25623));
  AND2 AND2_2893(.VSS(VSS),.VDD(VDD),.Y(g26352),.A(g25919),.B(g9749));
  AND2 AND2_2894(.VSS(VSS),.VDD(VDD),.Y(g26353),.A(g25923),.B(g9752));
  AND2 AND2_2895(.VSS(VSS),.VDD(VDD),.Y(g26357),.A(g4882),.B(g25634));
  AND2 AND2_2896(.VSS(VSS),.VDD(VDD),.Y(g26361),.A(g4888),.B(g25637));
  AND2 AND2_2897(.VSS(VSS),.VDD(VDD),.Y(g26362),.A(g4891),.B(g25640));
  AND2 AND2_2898(.VSS(VSS),.VDD(VDD),.Y(g26363),.A(g4894),.B(g25643));
  AND2 AND2_2899(.VSS(VSS),.VDD(VDD),.Y(g26365),.A(g4913),.B(g25652));
  AND2 AND2_2900(.VSS(VSS),.VDD(VDD),.Y(g26366),.A(g4916),.B(g25655));
  AND2 AND2_2901(.VSS(VSS),.VDD(VDD),.Y(g26371),.A(g4919),.B(g25658));
  AND2 AND2_2902(.VSS(VSS),.VDD(VDD),.Y(g26372),.A(g4922),.B(g25661));
  AND2 AND2_2903(.VSS(VSS),.VDD(VDD),.Y(g26373),.A(g4925),.B(g25664));
  AND2 AND2_2904(.VSS(VSS),.VDD(VDD),.Y(g26379),.A(g4945),.B(g25669));
  AND2 AND2_2905(.VSS(VSS),.VDD(VDD),.Y(g26380),.A(g4948),.B(g25672));
  AND2 AND2_2906(.VSS(VSS),.VDD(VDD),.Y(g26381),.A(g4951),.B(g25675));
  AND2 AND2_2907(.VSS(VSS),.VDD(VDD),.Y(g26382),.A(g25915),.B(g9812));
  AND2 AND2_2908(.VSS(VSS),.VDD(VDD),.Y(g26383),.A(g4956),.B(g25678));
  AND2 AND2_2909(.VSS(VSS),.VDD(VDD),.Y(g26384),.A(g4959),.B(g25681));
  AND2 AND2_2910(.VSS(VSS),.VDD(VDD),.Y(g26386),.A(g4994),.B(g25685));
  AND2 AND2_2911(.VSS(VSS),.VDD(VDD),.Y(g26387),.A(g4997),.B(g25688));
  AND2 AND2_2912(.VSS(VSS),.VDD(VDD),.Y(g26388),.A(g5000),.B(g25691));
  AND2 AND2_2913(.VSS(VSS),.VDD(VDD),.Y(g26389),.A(g25264),.B(g17962));
  AND2 AND2_2914(.VSS(VSS),.VDD(VDD),.Y(g26390),.A(g25919),.B(g9873));
  AND2 AND2_2915(.VSS(VSS),.VDD(VDD),.Y(g26391),.A(g25923),.B(g9876));
  AND2 AND2_2916(.VSS(VSS),.VDD(VDD),.Y(g26392),.A(g5005),.B(g25694));
  AND2 AND2_2917(.VSS(VSS),.VDD(VDD),.Y(g26396),.A(g5027),.B(g25700));
  AND2 AND2_2918(.VSS(VSS),.VDD(VDD),.Y(g26397),.A(g5030),.B(g25703));
  AND2 AND2_2919(.VSS(VSS),.VDD(VDD),.Y(g26400),.A(g5041),.B(g25711));
  AND2 AND2_2920(.VSS(VSS),.VDD(VDD),.Y(g26404),.A(g5047),.B(g25714));
  AND2 AND2_2921(.VSS(VSS),.VDD(VDD),.Y(g26405),.A(g5050),.B(g25717));
  AND2 AND2_2922(.VSS(VSS),.VDD(VDD),.Y(g26406),.A(g5053),.B(g25720));
  AND2 AND2_2923(.VSS(VSS),.VDD(VDD),.Y(g26408),.A(g5072),.B(g25729));
  AND2 AND2_2924(.VSS(VSS),.VDD(VDD),.Y(g26409),.A(g5075),.B(g25732));
  AND2 AND2_2925(.VSS(VSS),.VDD(VDD),.Y(g26414),.A(g5078),.B(g25735));
  AND2 AND2_2926(.VSS(VSS),.VDD(VDD),.Y(g26415),.A(g5081),.B(g25738));
  AND2 AND2_2927(.VSS(VSS),.VDD(VDD),.Y(g26416),.A(g5084),.B(g25741));
  AND2 AND2_2928(.VSS(VSS),.VDD(VDD),.Y(g26422),.A(g5104),.B(g25746));
  AND2 AND2_2929(.VSS(VSS),.VDD(VDD),.Y(g26423),.A(g5107),.B(g25749));
  AND2 AND2_2930(.VSS(VSS),.VDD(VDD),.Y(g26424),.A(g5110),.B(g25752));
  AND2 AND2_2931(.VSS(VSS),.VDD(VDD),.Y(g26425),.A(g25923),.B(g9958));
  AND2 AND2_2932(.VSS(VSS),.VDD(VDD),.Y(g26426),.A(g5115),.B(g25755));
  AND2 AND2_2933(.VSS(VSS),.VDD(VDD),.Y(g26427),.A(g5118),.B(g25758));
  AND2 AND2_2934(.VSS(VSS),.VDD(VDD),.Y(g26432),.A(g5145),.B(g25767));
  AND2 AND2_2935(.VSS(VSS),.VDD(VDD),.Y(g26437),.A(g5156),.B(g25773));
  AND2 AND2_2936(.VSS(VSS),.VDD(VDD),.Y(g26438),.A(g5159),.B(g25776));
  AND2 AND2_2937(.VSS(VSS),.VDD(VDD),.Y(g26441),.A(g5170),.B(g25784));
  AND2 AND2_2938(.VSS(VSS),.VDD(VDD),.Y(g26445),.A(g5176),.B(g25787));
  AND2 AND2_2939(.VSS(VSS),.VDD(VDD),.Y(g26446),.A(g5179),.B(g25790));
  AND2 AND2_2940(.VSS(VSS),.VDD(VDD),.Y(g26447),.A(g5182),.B(g25793));
  AND2 AND2_2941(.VSS(VSS),.VDD(VDD),.Y(g26449),.A(g5201),.B(g25802));
  AND2 AND2_2942(.VSS(VSS),.VDD(VDD),.Y(g26450),.A(g5204),.B(g25805));
  AND2 AND2_2943(.VSS(VSS),.VDD(VDD),.Y(g26455),.A(g5207),.B(g25808));
  AND2 AND2_2944(.VSS(VSS),.VDD(VDD),.Y(g26456),.A(g5210),.B(g25811));
  AND2 AND2_2945(.VSS(VSS),.VDD(VDD),.Y(g26457),.A(g5213),.B(g25814));
  AND2 AND2_2946(.VSS(VSS),.VDD(VDD),.Y(g26464),.A(g5238),.B(g25821));
  AND2 AND2_2947(.VSS(VSS),.VDD(VDD),.Y(g26469),.A(g5249),.B(g25827));
  AND2 AND2_2948(.VSS(VSS),.VDD(VDD),.Y(g26470),.A(g5252),.B(g25830));
  AND2 AND2_2949(.VSS(VSS),.VDD(VDD),.Y(g26473),.A(g5263),.B(g25838));
  AND2 AND2_2950(.VSS(VSS),.VDD(VDD),.Y(g26477),.A(g5269),.B(g25841));
  AND2 AND2_2951(.VSS(VSS),.VDD(VDD),.Y(g26478),.A(g5272),.B(g25844));
  AND2 AND2_2952(.VSS(VSS),.VDD(VDD),.Y(g26479),.A(g5275),.B(g25847));
  AND2 AND2_2953(.VSS(VSS),.VDD(VDD),.Y(g26488),.A(g5301),.B(g25856));
  AND2 AND2_2954(.VSS(VSS),.VDD(VDD),.Y(g26493),.A(g5312),.B(g25862));
  AND2 AND2_2955(.VSS(VSS),.VDD(VDD),.Y(g26494),.A(g5315),.B(g25865));
  AND2 AND2_2956(.VSS(VSS),.VDD(VDD),.Y(g26504),.A(g5338),.B(g25877));
  AND2 AND2_2957(.VSS(VSS),.VDD(VDD),.Y(g26663),.A(g25274),.B(g21066));
  AND2 AND2_2958(.VSS(VSS),.VDD(VDD),.Y(g26668),.A(g25283),.B(g21076));
  AND2 AND2_2959(.VSS(VSS),.VDD(VDD),.Y(g26673),.A(g12431),.B(g25318));
  AND2 AND2_2960(.VSS(VSS),.VDD(VDD),.Y(g26674),.A(g25291),.B(g21090));
  AND2 AND2_2961(.VSS(VSS),.VDD(VDD),.Y(g26754),.A(g14657),.B(g26508));
  AND2 AND2_2962(.VSS(VSS),.VDD(VDD),.Y(g26755),.A(g26083),.B(g22239));
  AND2 AND2_2963(.VSS(VSS),.VDD(VDD),.Y(g26756),.A(g26113),.B(g22240));
  AND3 AND3_247(.VSS(VSS),.VDD(VDD),.Y(g26758),.A(g16614),.B(g26521),.C(g13637));
  AND2 AND2_2964(.VSS(VSS),.VDD(VDD),.Y(g26759),.A(g26356),.B(g19251));
  AND2 AND2_2965(.VSS(VSS),.VDD(VDD),.Y(g26760),.A(g26137),.B(g22256));
  AND2 AND2_2966(.VSS(VSS),.VDD(VDD),.Y(g26761),.A(g26154),.B(g22257));
  AND2 AND2_2967(.VSS(VSS),.VDD(VDD),.Y(g26763),.A(g14691),.B(g26516));
  AND3 AND3_248(.VSS(VSS),.VDD(VDD),.Y(g26764),.A(g16632),.B(g26525),.C(g13649));
  AND2 AND2_2968(.VSS(VSS),.VDD(VDD),.Y(g26765),.A(g26399),.B(g19265));
  AND2 AND2_2969(.VSS(VSS),.VDD(VDD),.Y(g26766),.A(g14725),.B(g26521));
  AND2 AND2_2970(.VSS(VSS),.VDD(VDD),.Y(g26767),.A(g26087),.B(g22287));
  AND2 AND2_2971(.VSS(VSS),.VDD(VDD),.Y(g26768),.A(g26440),.B(g19280));
  AND2 AND2_2972(.VSS(VSS),.VDD(VDD),.Y(g26769),.A(g14753),.B(g26525));
  AND2 AND2_2973(.VSS(VSS),.VDD(VDD),.Y(g26770),.A(g26059),.B(g19287));
  AND3 AND3_249(.VSS(VSS),.VDD(VDD),.Y(g26771),.A(g24912),.B(g26508),.C(g13614));
  AND2 AND2_2974(.VSS(VSS),.VDD(VDD),.Y(g26773),.A(g26145),.B(g22303));
  AND2 AND2_2975(.VSS(VSS),.VDD(VDD),.Y(g26774),.A(g26472),.B(g19299));
  AND2 AND2_2976(.VSS(VSS),.VDD(VDD),.Y(g26775),.A(g26099),.B(g22318));
  AND2 AND2_2977(.VSS(VSS),.VDD(VDD),.Y(g26777),.A(g26066),.B(g19305));
  AND3 AND3_250(.VSS(VSS),.VDD(VDD),.Y(g26778),.A(g24929),.B(g26516),.C(g13626));
  AND2 AND2_2978(.VSS(VSS),.VDD(VDD),.Y(g26780),.A(g26119),.B(g16622));
  AND2 AND2_2979(.VSS(VSS),.VDD(VDD),.Y(g26783),.A(g26073),.B(g19326));
  AND3 AND3_251(.VSS(VSS),.VDD(VDD),.Y(g26784),.A(g24941),.B(g26521),.C(g13637));
  AND2 AND2_2980(.VSS(VSS),.VDD(VDD),.Y(g26787),.A(g26129),.B(g16636));
  AND2 AND2_2981(.VSS(VSS),.VDD(VDD),.Y(g26790),.A(g26079),.B(g19353));
  AND3 AND3_252(.VSS(VSS),.VDD(VDD),.Y(g26791),.A(g24952),.B(g26525),.C(g13649));
  AND2 AND2_2982(.VSS(VSS),.VDD(VDD),.Y(g26794),.A(g26143),.B(g16647));
  AND2 AND2_2983(.VSS(VSS),.VDD(VDD),.Y(g26797),.A(g26148),.B(g16659));
  AND2 AND2_2984(.VSS(VSS),.VDD(VDD),.Y(g26829),.A(g5623),.B(g26209));
  AND2 AND2_2985(.VSS(VSS),.VDD(VDD),.Y(g26833),.A(g5651),.B(g26237));
  AND2 AND2_2986(.VSS(VSS),.VDD(VDD),.Y(g26842),.A(g5689),.B(g26275));
  AND2 AND2_2987(.VSS(VSS),.VDD(VDD),.Y(g26845),.A(g5664),.B(g26056));
  AND2 AND2_2988(.VSS(VSS),.VDD(VDD),.Y(g26851),.A(g5741),.B(g26313));
  AND2 AND2_2989(.VSS(VSS),.VDD(VDD),.Y(g26853),.A(g5716),.B(g26063));
  AND2 AND2_2990(.VSS(VSS),.VDD(VDD),.Y(g26860),.A(g5774),.B(g26070));
  AND2 AND2_2991(.VSS(VSS),.VDD(VDD),.Y(g26866),.A(g5833),.B(g26076));
  AND2 AND2_2992(.VSS(VSS),.VDD(VDD),.Y(g26955),.A(g6157),.B(g26533));
  AND2 AND2_2993(.VSS(VSS),.VDD(VDD),.Y(g26958),.A(g6184),.B(g26538));
  AND2 AND2_2994(.VSS(VSS),.VDD(VDD),.Y(g26961),.A(g13907),.B(g26175));
  AND2 AND2_2995(.VSS(VSS),.VDD(VDD),.Y(g26962),.A(g6180),.B(g26178));
  AND2 AND2_2996(.VSS(VSS),.VDD(VDD),.Y(g26963),.A(g6216),.B(g26539));
  AND2 AND2_2997(.VSS(VSS),.VDD(VDD),.Y(g26965),.A(g23320),.B(g26540));
  AND2 AND2_2998(.VSS(VSS),.VDD(VDD),.Y(g26966),.A(g13963),.B(g26196));
  AND2 AND2_2999(.VSS(VSS),.VDD(VDD),.Y(g26967),.A(g6212),.B(g26202));
  AND2 AND2_3000(.VSS(VSS),.VDD(VDD),.Y(g26968),.A(g6305),.B(g26542));
  AND2 AND2_3001(.VSS(VSS),.VDD(VDD),.Y(g26969),.A(g23320),.B(g26543));
  AND2 AND2_3002(.VSS(VSS),.VDD(VDD),.Y(g26970),.A(g21976),.B(g26544));
  AND2 AND2_3003(.VSS(VSS),.VDD(VDD),.Y(g26971),.A(g23325),.B(g26546));
  AND2 AND2_3004(.VSS(VSS),.VDD(VDD),.Y(g26972),.A(g14033),.B(g26223));
  AND2 AND2_3005(.VSS(VSS),.VDD(VDD),.Y(g26973),.A(g6301),.B(g26226));
  AND2 AND2_3006(.VSS(VSS),.VDD(VDD),.Y(g26977),.A(g23320),.B(g26550));
  AND2 AND2_3007(.VSS(VSS),.VDD(VDD),.Y(g26978),.A(g21976),.B(g26551));
  AND2 AND2_3008(.VSS(VSS),.VDD(VDD),.Y(g26979),.A(g23331),.B(g26552));
  AND2 AND2_3009(.VSS(VSS),.VDD(VDD),.Y(g26980),.A(g23360),.B(g26554));
  AND2 AND2_3010(.VSS(VSS),.VDD(VDD),.Y(g26981),.A(g23325),.B(g26555));
  AND2 AND2_3011(.VSS(VSS),.VDD(VDD),.Y(g26982),.A(g21983),.B(g26556));
  AND2 AND2_3012(.VSS(VSS),.VDD(VDD),.Y(g26984),.A(g23335),.B(g26558));
  AND2 AND2_3013(.VSS(VSS),.VDD(VDD),.Y(g26985),.A(g14124),.B(g26251));
  AND2 AND2_3014(.VSS(VSS),.VDD(VDD),.Y(g26986),.A(g6438),.B(g26254));
  AND2 AND2_3015(.VSS(VSS),.VDD(VDD),.Y(g26993),.A(g21976),.B(g26561));
  AND2 AND2_3016(.VSS(VSS),.VDD(VDD),.Y(g26994),.A(g23331),.B(g26562));
  AND2 AND2_3017(.VSS(VSS),.VDD(VDD),.Y(g26995),.A(g21991),.B(g26563));
  AND2 AND2_3018(.VSS(VSS),.VDD(VDD),.Y(g26996),.A(g23360),.B(g26564));
  AND2 AND2_3019(.VSS(VSS),.VDD(VDD),.Y(g26997),.A(g22050),.B(g26565));
  AND2 AND2_3020(.VSS(VSS),.VDD(VDD),.Y(g26998),.A(g23325),.B(g26566));
  AND2 AND2_3021(.VSS(VSS),.VDD(VDD),.Y(g26999),.A(g21983),.B(g26567));
  AND2 AND2_3022(.VSS(VSS),.VDD(VDD),.Y(g27000),.A(g23340),.B(g26568));
  AND2 AND2_3023(.VSS(VSS),.VDD(VDD),.Y(g27001),.A(g23364),.B(g26570));
  AND2 AND2_3024(.VSS(VSS),.VDD(VDD),.Y(g27002),.A(g23335),.B(g26571));
  AND2 AND2_3025(.VSS(VSS),.VDD(VDD),.Y(g27003),.A(g21996),.B(g26572));
  AND2 AND2_3026(.VSS(VSS),.VDD(VDD),.Y(g27004),.A(g23344),.B(g26574));
  AND2 AND2_3027(.VSS(VSS),.VDD(VDD),.Y(g27005),.A(g23331),.B(g26578));
  AND2 AND2_3028(.VSS(VSS),.VDD(VDD),.Y(g27006),.A(g21991),.B(g26579));
  AND2 AND2_3029(.VSS(VSS),.VDD(VDD),.Y(g27007),.A(g23360),.B(g26580));
  AND2 AND2_3030(.VSS(VSS),.VDD(VDD),.Y(g27008),.A(g22050),.B(g26581));
  AND2 AND2_3031(.VSS(VSS),.VDD(VDD),.Y(g27009),.A(g23368),.B(g26582));
  AND2 AND2_3032(.VSS(VSS),.VDD(VDD),.Y(g27016),.A(g21983),.B(g26584));
  AND2 AND2_3033(.VSS(VSS),.VDD(VDD),.Y(g27017),.A(g23340),.B(g26585));
  AND2 AND2_3034(.VSS(VSS),.VDD(VDD),.Y(g27018),.A(g22005),.B(g26586));
  AND2 AND2_3035(.VSS(VSS),.VDD(VDD),.Y(g27019),.A(g23364),.B(g26587));
  AND2 AND2_3036(.VSS(VSS),.VDD(VDD),.Y(g27020),.A(g22069),.B(g26588));
  AND2 AND2_3037(.VSS(VSS),.VDD(VDD),.Y(g27021),.A(g23335),.B(g26589));
  AND2 AND2_3038(.VSS(VSS),.VDD(VDD),.Y(g27022),.A(g21996),.B(g26590));
  AND2 AND2_3039(.VSS(VSS),.VDD(VDD),.Y(g27023),.A(g23349),.B(g26591));
  AND2 AND2_3040(.VSS(VSS),.VDD(VDD),.Y(g27024),.A(g23372),.B(g26593));
  AND2 AND2_3041(.VSS(VSS),.VDD(VDD),.Y(g27025),.A(g23344),.B(g26594));
  AND2 AND2_3042(.VSS(VSS),.VDD(VDD),.Y(g27026),.A(g22009),.B(g26595));
  AND2 AND2_3043(.VSS(VSS),.VDD(VDD),.Y(g27027),.A(g21991),.B(g26598));
  AND2 AND2_3044(.VSS(VSS),.VDD(VDD),.Y(g27028),.A(g22050),.B(g26599));
  AND2 AND2_3045(.VSS(VSS),.VDD(VDD),.Y(g27029),.A(g23368),.B(g26600));
  AND2 AND2_3046(.VSS(VSS),.VDD(VDD),.Y(g27030),.A(g22083),.B(g26601));
  AND2 AND2_3047(.VSS(VSS),.VDD(VDD),.Y(g27031),.A(g23340),.B(g26602));
  AND2 AND2_3048(.VSS(VSS),.VDD(VDD),.Y(g27032),.A(g22005),.B(g26603));
  AND2 AND2_3049(.VSS(VSS),.VDD(VDD),.Y(g27033),.A(g23364),.B(g26604));
  AND2 AND2_3050(.VSS(VSS),.VDD(VDD),.Y(g27034),.A(g22069),.B(g26605));
  AND2 AND2_3051(.VSS(VSS),.VDD(VDD),.Y(g27035),.A(g23377),.B(g26606));
  AND2 AND2_3052(.VSS(VSS),.VDD(VDD),.Y(g27042),.A(g21996),.B(g26608));
  AND2 AND2_3053(.VSS(VSS),.VDD(VDD),.Y(g27043),.A(g23349),.B(g26609));
  AND2 AND2_3054(.VSS(VSS),.VDD(VDD),.Y(g27044),.A(g22016),.B(g26610));
  AND2 AND2_3055(.VSS(VSS),.VDD(VDD),.Y(g27045),.A(g23372),.B(g26611));
  AND2 AND2_3056(.VSS(VSS),.VDD(VDD),.Y(g27046),.A(g22093),.B(g26612));
  AND2 AND2_3057(.VSS(VSS),.VDD(VDD),.Y(g27047),.A(g23344),.B(g26613));
  AND2 AND2_3058(.VSS(VSS),.VDD(VDD),.Y(g27048),.A(g22009),.B(g26614));
  AND2 AND2_3059(.VSS(VSS),.VDD(VDD),.Y(g27049),.A(g23353),.B(g26615));
  AND2 AND2_3060(.VSS(VSS),.VDD(VDD),.Y(g27050),.A(g23381),.B(g26617));
  AND2 AND2_3061(.VSS(VSS),.VDD(VDD),.Y(g27052),.A(g4885),.B(g26358));
  AND2 AND2_3062(.VSS(VSS),.VDD(VDD),.Y(g27053),.A(g23368),.B(g26619));
  AND2 AND2_3063(.VSS(VSS),.VDD(VDD),.Y(g27054),.A(g22083),.B(g26620));
  AND2 AND2_3064(.VSS(VSS),.VDD(VDD),.Y(g27055),.A(g22005),.B(g26621));
  AND2 AND2_3065(.VSS(VSS),.VDD(VDD),.Y(g27056),.A(g22069),.B(g26622));
  AND2 AND2_3066(.VSS(VSS),.VDD(VDD),.Y(g27057),.A(g23377),.B(g26623));
  AND2 AND2_3067(.VSS(VSS),.VDD(VDD),.Y(g27058),.A(g22108),.B(g26624));
  AND2 AND2_3068(.VSS(VSS),.VDD(VDD),.Y(g27059),.A(g23349),.B(g26625));
  AND2 AND2_3069(.VSS(VSS),.VDD(VDD),.Y(g27060),.A(g22016),.B(g26626));
  AND2 AND2_3070(.VSS(VSS),.VDD(VDD),.Y(g27061),.A(g23372),.B(g26627));
  AND2 AND2_3071(.VSS(VSS),.VDD(VDD),.Y(g27062),.A(g22093),.B(g26628));
  AND2 AND2_3072(.VSS(VSS),.VDD(VDD),.Y(g27063),.A(g23388),.B(g26629));
  AND2 AND2_3073(.VSS(VSS),.VDD(VDD),.Y(g27070),.A(g22009),.B(g26631));
  AND2 AND2_3074(.VSS(VSS),.VDD(VDD),.Y(g27071),.A(g23353),.B(g26632));
  AND2 AND2_3075(.VSS(VSS),.VDD(VDD),.Y(g27072),.A(g22021),.B(g26633));
  AND2 AND2_3076(.VSS(VSS),.VDD(VDD),.Y(g27073),.A(g23381),.B(g26634));
  AND2 AND2_3077(.VSS(VSS),.VDD(VDD),.Y(g27074),.A(g22118),.B(g26635));
  AND2 AND2_3078(.VSS(VSS),.VDD(VDD),.Y(g27076),.A(g5024),.B(g26393));
  AND2 AND2_3079(.VSS(VSS),.VDD(VDD),.Y(g27077),.A(g22083),.B(g26636));
  AND2 AND2_3080(.VSS(VSS),.VDD(VDD),.Y(g27079),.A(g5044),.B(g26401));
  AND2 AND2_3081(.VSS(VSS),.VDD(VDD),.Y(g27080),.A(g23377),.B(g26637));
  AND2 AND2_3082(.VSS(VSS),.VDD(VDD),.Y(g27081),.A(g22108),.B(g26638));
  AND2 AND2_3083(.VSS(VSS),.VDD(VDD),.Y(g27082),.A(g22016),.B(g26639));
  AND2 AND2_3084(.VSS(VSS),.VDD(VDD),.Y(g27083),.A(g22093),.B(g26640));
  AND2 AND2_3085(.VSS(VSS),.VDD(VDD),.Y(g27084),.A(g23388),.B(g26641));
  AND2 AND2_3086(.VSS(VSS),.VDD(VDD),.Y(g27085),.A(g22134),.B(g26642));
  AND2 AND2_3087(.VSS(VSS),.VDD(VDD),.Y(g27086),.A(g23353),.B(g26643));
  AND2 AND2_3088(.VSS(VSS),.VDD(VDD),.Y(g27087),.A(g22021),.B(g26644));
  AND2 AND2_3089(.VSS(VSS),.VDD(VDD),.Y(g27088),.A(g23381),.B(g26645));
  AND2 AND2_3090(.VSS(VSS),.VDD(VDD),.Y(g27089),.A(g22118),.B(g26646));
  AND2 AND2_3091(.VSS(VSS),.VDD(VDD),.Y(g27090),.A(g23395),.B(g26647));
  AND2 AND2_3092(.VSS(VSS),.VDD(VDD),.Y(g27091),.A(g5142),.B(g26429));
  AND2 AND2_3093(.VSS(VSS),.VDD(VDD),.Y(g27092),.A(g5153),.B(g26434));
  AND2 AND2_3094(.VSS(VSS),.VDD(VDD),.Y(g27093),.A(g22108),.B(g26648));
  AND2 AND2_3095(.VSS(VSS),.VDD(VDD),.Y(g27095),.A(g5173),.B(g26442));
  AND2 AND2_3096(.VSS(VSS),.VDD(VDD),.Y(g27096),.A(g23388),.B(g26649));
  AND2 AND2_3097(.VSS(VSS),.VDD(VDD),.Y(g27097),.A(g22134),.B(g26650));
  AND2 AND2_3098(.VSS(VSS),.VDD(VDD),.Y(g27098),.A(g22021),.B(g26651));
  AND2 AND2_3099(.VSS(VSS),.VDD(VDD),.Y(g27099),.A(g22118),.B(g26652));
  AND2 AND2_3100(.VSS(VSS),.VDD(VDD),.Y(g27100),.A(g23395),.B(g26653));
  AND2 AND2_3101(.VSS(VSS),.VDD(VDD),.Y(g27101),.A(g22157),.B(g26654));
  AND2 AND2_3102(.VSS(VSS),.VDD(VDD),.Y(g27103),.A(g5235),.B(g26461));
  AND2 AND2_3103(.VSS(VSS),.VDD(VDD),.Y(g27104),.A(g5246),.B(g26466));
  AND2 AND2_3104(.VSS(VSS),.VDD(VDD),.Y(g27105),.A(g22134),.B(g26656));
  AND2 AND2_3105(.VSS(VSS),.VDD(VDD),.Y(g27107),.A(g5266),.B(g26474));
  AND2 AND2_3106(.VSS(VSS),.VDD(VDD),.Y(g27108),.A(g23395),.B(g26657));
  AND2 AND2_3107(.VSS(VSS),.VDD(VDD),.Y(g27109),.A(g22157),.B(g26658));
  AND2 AND2_3108(.VSS(VSS),.VDD(VDD),.Y(g27110),.A(g5298),.B(g26485));
  AND2 AND2_3109(.VSS(VSS),.VDD(VDD),.Y(g27111),.A(g5309),.B(g26490));
  AND2 AND2_3110(.VSS(VSS),.VDD(VDD),.Y(g27112),.A(g22157),.B(g26662));
  AND2 AND2_3111(.VSS(VSS),.VDD(VDD),.Y(g27115),.A(g5335),.B(g26501));
  AND2 AND2_3112(.VSS(VSS),.VDD(VDD),.Y(g27178),.A(g26110),.B(g22213));
  AND3 AND3_253(.VSS(VSS),.VDD(VDD),.Y(g27181),.A(g16570),.B(g26508),.C(g13614));
  AND2 AND2_3113(.VSS(VSS),.VDD(VDD),.Y(g27182),.A(g26151),.B(g22217));
  AND2 AND2_3114(.VSS(VSS),.VDD(VDD),.Y(g27185),.A(g26126),.B(g22230));
  AND3 AND3_254(.VSS(VSS),.VDD(VDD),.Y(g27187),.A(g16594),.B(g26516),.C(g13626));
  AND2 AND2_3115(.VSS(VSS),.VDD(VDD),.Y(g27240),.A(g26905),.B(g22241));
  AND2 AND2_3116(.VSS(VSS),.VDD(VDD),.Y(g27241),.A(g10730),.B(g26934));
  AND2 AND2_3117(.VSS(VSS),.VDD(VDD),.Y(g27242),.A(g26793),.B(g8357));
  AND2 AND2_3118(.VSS(VSS),.VDD(VDD),.Y(g27244),.A(g26914),.B(g22258));
  AND2 AND2_3119(.VSS(VSS),.VDD(VDD),.Y(g27245),.A(g26877),.B(g22286));
  AND2 AND2_3120(.VSS(VSS),.VDD(VDD),.Y(g27246),.A(g26988),.B(g16676));
  AND2 AND2_3121(.VSS(VSS),.VDD(VDD),.Y(g27247),.A(g27011),.B(g16702));
  AND2 AND2_3122(.VSS(VSS),.VDD(VDD),.Y(g27248),.A(g27037),.B(g16733));
  AND2 AND2_3123(.VSS(VSS),.VDD(VDD),.Y(g27249),.A(g27065),.B(g16775));
  AND2 AND2_3124(.VSS(VSS),.VDD(VDD),.Y(g27355),.A(g61),.B(g26837));
  AND2 AND2_3125(.VSS(VSS),.VDD(VDD),.Y(g27356),.A(g65),.B(g26987));
  AND2 AND2_3126(.VSS(VSS),.VDD(VDD),.Y(g27358),.A(g749),.B(g26846));
  AND2 AND2_3127(.VSS(VSS),.VDD(VDD),.Y(g27359),.A(g753),.B(g27010));
  AND2 AND2_3128(.VSS(VSS),.VDD(VDD),.Y(g27364),.A(g1435),.B(g26855));
  AND2 AND2_3129(.VSS(VSS),.VDD(VDD),.Y(g27365),.A(g1439),.B(g27036));
  AND2 AND2_3130(.VSS(VSS),.VDD(VDD),.Y(g27370),.A(g27126),.B(g8874));
  AND2 AND2_3131(.VSS(VSS),.VDD(VDD),.Y(g27371),.A(g2129),.B(g26861));
  AND2 AND2_3132(.VSS(VSS),.VDD(VDD),.Y(g27372),.A(g2133),.B(g27064));
  AND2 AND2_3133(.VSS(VSS),.VDD(VDD),.Y(g27394),.A(g17802),.B(g27134));
  AND2 AND2_3134(.VSS(VSS),.VDD(VDD),.Y(g27396),.A(g692),.B(g27135));
  AND2 AND2_3135(.VSS(VSS),.VDD(VDD),.Y(g27407),.A(g17914),.B(g27136));
  AND2 AND2_3136(.VSS(VSS),.VDD(VDD),.Y(g27409),.A(g1378),.B(g27137));
  AND2 AND2_3137(.VSS(VSS),.VDD(VDD),.Y(g27425),.A(g18025),.B(g27138));
  AND2 AND2_3138(.VSS(VSS),.VDD(VDD),.Y(g27427),.A(g2072),.B(g27139));
  AND2 AND2_3139(.VSS(VSS),.VDD(VDD),.Y(g27446),.A(g18142),.B(g27141));
  AND2 AND2_3140(.VSS(VSS),.VDD(VDD),.Y(g27448),.A(g2766),.B(g27142));
  AND2 AND2_3141(.VSS(VSS),.VDD(VDD),.Y(g27495),.A(g23945),.B(g27146));
  AND2 AND2_3142(.VSS(VSS),.VDD(VDD),.Y(g27509),.A(g23945),.B(g27148));
  AND2 AND2_3143(.VSS(VSS),.VDD(VDD),.Y(g27516),.A(g23974),.B(g27151));
  AND2 AND2_3144(.VSS(VSS),.VDD(VDD),.Y(g27530),.A(g23945),.B(g27153));
  AND2 AND2_3145(.VSS(VSS),.VDD(VDD),.Y(g27534),.A(g23974),.B(g27155));
  AND2 AND2_3146(.VSS(VSS),.VDD(VDD),.Y(g27541),.A(g24004),.B(g27159));
  AND2 AND2_3147(.VSS(VSS),.VDD(VDD),.Y(g27552),.A(g23974),.B(g27162));
  AND2 AND2_3148(.VSS(VSS),.VDD(VDD),.Y(g27554),.A(g24004),.B(g27164));
  AND2 AND2_3149(.VSS(VSS),.VDD(VDD),.Y(g27561),.A(g24038),.B(g27167));
  AND2 AND2_3150(.VSS(VSS),.VDD(VDD),.Y(g27568),.A(g24004),.B(g27172));
  AND2 AND2_3151(.VSS(VSS),.VDD(VDD),.Y(g27570),.A(g24038),.B(g27173));
  AND2 AND2_3152(.VSS(VSS),.VDD(VDD),.Y(g27578),.A(g24038),.B(g27177));
  AND2 AND2_3153(.VSS(VSS),.VDD(VDD),.Y(g27656),.A(g26796),.B(g11004));
  AND2 AND2_3154(.VSS(VSS),.VDD(VDD),.Y(g27657),.A(g27114),.B(g11051));
  AND2 AND2_3155(.VSS(VSS),.VDD(VDD),.Y(g27659),.A(g27132),.B(g11114));
  AND2 AND2_3156(.VSS(VSS),.VDD(VDD),.Y(g27660),.A(g26835),.B(g11117));
  AND2 AND2_3157(.VSS(VSS),.VDD(VDD),.Y(g27661),.A(g26841),.B(g11173));
  AND2 AND2_3158(.VSS(VSS),.VDD(VDD),.Y(g27666),.A(g26849),.B(g11243));
  AND2 AND2_3159(.VSS(VSS),.VDD(VDD),.Y(g27671),.A(g26885),.B(g22212));
  AND2 AND2_3160(.VSS(VSS),.VDD(VDD),.Y(g27673),.A(g26854),.B(g11312));
  AND2 AND2_3161(.VSS(VSS),.VDD(VDD),.Y(g27679),.A(g26782),.B(g11386));
  AND2 AND2_3162(.VSS(VSS),.VDD(VDD),.Y(g27680),.A(g26983),.B(g11392));
  AND2 AND2_3163(.VSS(VSS),.VDD(VDD),.Y(g27681),.A(g26788),.B(g11456));
  AND2 AND2_3164(.VSS(VSS),.VDD(VDD),.Y(g27719),.A(g27496),.B(g20649));
  AND2 AND2_3165(.VSS(VSS),.VDD(VDD),.Y(g27720),.A(g27481),.B(g20652));
  AND2 AND2_3166(.VSS(VSS),.VDD(VDD),.Y(g27721),.A(g27579),.B(g20655));
  AND2 AND2_3167(.VSS(VSS),.VDD(VDD),.Y(g27723),.A(g27464),.B(g20679));
  AND2 AND2_3168(.VSS(VSS),.VDD(VDD),.Y(g27725),.A(g27532),.B(g20704));
  AND2 AND2_3169(.VSS(VSS),.VDD(VDD),.Y(g27726),.A(g27531),.B(g20732));
  AND2 AND2_3170(.VSS(VSS),.VDD(VDD),.Y(g27727),.A(g27414),.B(g19301));
  AND2 AND2_3171(.VSS(VSS),.VDD(VDD),.Y(g27728),.A(g27564),.B(g20766));
  AND2 AND2_3172(.VSS(VSS),.VDD(VDD),.Y(g27729),.A(g27435),.B(g19322));
  AND2 AND2_3173(.VSS(VSS),.VDD(VDD),.Y(g27730),.A(g27454),.B(g19349));
  AND2 AND2_3174(.VSS(VSS),.VDD(VDD),.Y(g27731),.A(g27470),.B(g19383));
  AND2 AND2_3175(.VSS(VSS),.VDD(VDD),.Y(g27732),.A(g27492),.B(g16758));
  AND2 AND2_3176(.VSS(VSS),.VDD(VDD),.Y(g27733),.A(g27513),.B(g16785));
  AND2 AND2_3177(.VSS(VSS),.VDD(VDD),.Y(g27734),.A(g27538),.B(g16814));
  AND2 AND2_3178(.VSS(VSS),.VDD(VDD),.Y(g27737),.A(g27558),.B(g16832));
  AND2 AND2_3179(.VSS(VSS),.VDD(VDD),.Y(g27770),.A(g5642),.B(g27449));
  AND2 AND2_3180(.VSS(VSS),.VDD(VDD),.Y(g27772),.A(g5680),.B(g27465));
  AND2 AND2_3181(.VSS(VSS),.VDD(VDD),.Y(g27773),.A(g5732),.B(g27484));
  AND2 AND2_3182(.VSS(VSS),.VDD(VDD),.Y(g27774),.A(g5702),.B(g27361));
  AND2 AND2_3183(.VSS(VSS),.VDD(VDD),.Y(g27775),.A(g5790),.B(g27506));
  AND2 AND2_3184(.VSS(VSS),.VDD(VDD),.Y(g27779),.A(g5760),.B(g27367));
  AND2 AND2_3185(.VSS(VSS),.VDD(VDD),.Y(g27783),.A(g5819),.B(g27373));
  AND2 AND2_3186(.VSS(VSS),.VDD(VDD),.Y(g27790),.A(g5875),.B(g27376));
  AND2 AND2_3187(.VSS(VSS),.VDD(VDD),.Y(g27904),.A(g13873),.B(g27387));
  AND2 AND2_3188(.VSS(VSS),.VDD(VDD),.Y(g27908),.A(g13886),.B(g27391));
  AND2 AND2_3189(.VSS(VSS),.VDD(VDD),.Y(g27909),.A(g13895),.B(g27397));
  AND2 AND2_3190(.VSS(VSS),.VDD(VDD),.Y(g27913),.A(g4017),.B(g27401));
  AND2 AND2_3191(.VSS(VSS),.VDD(VDD),.Y(g27914),.A(g13927),.B(g27404));
  AND2 AND2_3192(.VSS(VSS),.VDD(VDD),.Y(g27915),.A(g13936),.B(g27410));
  AND2 AND2_3193(.VSS(VSS),.VDD(VDD),.Y(g27922),.A(g4112),.B(g27416));
  AND2 AND2_3194(.VSS(VSS),.VDD(VDD),.Y(g27923),.A(g4144),.B(g27419));
  AND2 AND2_3195(.VSS(VSS),.VDD(VDD),.Y(g27924),.A(g13983),.B(g27422));
  AND2 AND2_3196(.VSS(VSS),.VDD(VDD),.Y(g27926),.A(g13992),.B(g27428));
  AND2 AND2_3197(.VSS(VSS),.VDD(VDD),.Y(g27931),.A(g4221),.B(g27432));
  AND2 AND2_3198(.VSS(VSS),.VDD(VDD),.Y(g27935),.A(g4251),.B(g27437));
  AND2 AND2_3199(.VSS(VSS),.VDD(VDD),.Y(g27936),.A(g4283),.B(g27440));
  AND2 AND2_3200(.VSS(VSS),.VDD(VDD),.Y(g27938),.A(g14053),.B(g27443));
  AND2 AND2_3201(.VSS(VSS),.VDD(VDD),.Y(g27945),.A(g4376),.B(g27451));
  AND2 AND2_3202(.VSS(VSS),.VDD(VDD),.Y(g27949),.A(g4406),.B(g27456));
  AND2 AND2_3203(.VSS(VSS),.VDD(VDD),.Y(g27951),.A(g4438),.B(g27459));
  AND2 AND2_3204(.VSS(VSS),.VDD(VDD),.Y(g27963),.A(g4545),.B(g27467));
  AND2 AND2_3205(.VSS(VSS),.VDD(VDD),.Y(g27968),.A(g4575),.B(g27472));
  AND2 AND2_3206(.VSS(VSS),.VDD(VDD),.Y(g27970),.A(g14238),.B(g27475));
  AND2 AND2_3207(.VSS(VSS),.VDD(VDD),.Y(g27984),.A(g4721),.B(g27486));
  AND2 AND2_3208(.VSS(VSS),.VDD(VDD),.Y(g27985),.A(g14342),.B(g27489));
  AND2 AND2_3209(.VSS(VSS),.VDD(VDD),.Y(g27991),.A(g14360),.B(g27498));
  AND2 AND2_3210(.VSS(VSS),.VDD(VDD),.Y(g28008),.A(g27590),.B(g9770));
  AND2 AND2_3211(.VSS(VSS),.VDD(VDD),.Y(g28009),.A(g14454),.B(g27510));
  AND2 AND2_3212(.VSS(VSS),.VDD(VDD),.Y(g28015),.A(g14472),.B(g27518));
  AND2 AND2_3213(.VSS(VSS),.VDD(VDD),.Y(g28027),.A(g27590),.B(g9895));
  AND2 AND2_3214(.VSS(VSS),.VDD(VDD),.Y(g28028),.A(g27595),.B(g9898));
  AND2 AND2_3215(.VSS(VSS),.VDD(VDD),.Y(g28035),.A(g27599),.B(g9916));
  AND2 AND2_3216(.VSS(VSS),.VDD(VDD),.Y(g28036),.A(g14541),.B(g27535));
  AND2 AND2_3217(.VSS(VSS),.VDD(VDD),.Y(g28042),.A(g14559),.B(g27543));
  AND2 AND2_3218(.VSS(VSS),.VDD(VDD),.Y(g28050),.A(g27590),.B(g10018));
  AND2 AND2_3219(.VSS(VSS),.VDD(VDD),.Y(g28051),.A(g27595),.B(g10021));
  AND2 AND2_3220(.VSS(VSS),.VDD(VDD),.Y(g28057),.A(g27599),.B(g10049));
  AND2 AND2_3221(.VSS(VSS),.VDD(VDD),.Y(g28058),.A(g27604),.B(g10052));
  AND2 AND2_3222(.VSS(VSS),.VDD(VDD),.Y(g28065),.A(g27608),.B(g10070));
  AND2 AND2_3223(.VSS(VSS),.VDD(VDD),.Y(g28066),.A(g14596),.B(g27555));
  AND2 AND2_3224(.VSS(VSS),.VDD(VDD),.Y(g28073),.A(g27595),.B(g10109));
  AND2 AND2_3225(.VSS(VSS),.VDD(VDD),.Y(g28079),.A(g27599),.B(g10127));
  AND2 AND2_3226(.VSS(VSS),.VDD(VDD),.Y(g28080),.A(g27604),.B(g10130));
  AND2 AND2_3227(.VSS(VSS),.VDD(VDD),.Y(g28086),.A(g27608),.B(g10158));
  AND2 AND2_3228(.VSS(VSS),.VDD(VDD),.Y(g28087),.A(g27613),.B(g10161));
  AND2 AND2_3229(.VSS(VSS),.VDD(VDD),.Y(g28094),.A(g27617),.B(g10179));
  AND2 AND2_3230(.VSS(VSS),.VDD(VDD),.Y(g28098),.A(g27604),.B(g10214));
  AND2 AND2_3231(.VSS(VSS),.VDD(VDD),.Y(g28104),.A(g27608),.B(g10232));
  AND2 AND2_3232(.VSS(VSS),.VDD(VDD),.Y(g28105),.A(g27613),.B(g10235));
  AND2 AND2_3233(.VSS(VSS),.VDD(VDD),.Y(g28111),.A(g27617),.B(g10263));
  AND2 AND2_3234(.VSS(VSS),.VDD(VDD),.Y(g28112),.A(g27622),.B(g10266));
  AND2 AND2_3235(.VSS(VSS),.VDD(VDD),.Y(g28116),.A(g27613),.B(g10316));
  AND2 AND2_3236(.VSS(VSS),.VDD(VDD),.Y(g28122),.A(g27617),.B(g10334));
  AND2 AND2_3237(.VSS(VSS),.VDD(VDD),.Y(g28123),.A(g27622),.B(g10337));
  AND2 AND2_3238(.VSS(VSS),.VDD(VDD),.Y(g28127),.A(g27622),.B(g10409));
  AND2 AND2_3239(.VSS(VSS),.VDD(VDD),.Y(g28171),.A(g27349),.B(g10898));
  AND2 AND2_3240(.VSS(VSS),.VDD(VDD),.Y(g28176),.A(g27349),.B(g10940));
  AND2 AND2_3241(.VSS(VSS),.VDD(VDD),.Y(g28188),.A(g27349),.B(g11008));
  AND2 AND2_3242(.VSS(VSS),.VDD(VDD),.Y(g28193),.A(g27573),.B(g21914));
  AND2 AND2_3243(.VSS(VSS),.VDD(VDD),.Y(g28319),.A(g27855),.B(g22246));
  AND2 AND2_3244(.VSS(VSS),.VDD(VDD),.Y(g28320),.A(g27854),.B(g20637));
  AND2 AND2_3245(.VSS(VSS),.VDD(VDD),.Y(g28322),.A(g27937),.B(g13868));
  AND2 AND2_3246(.VSS(VSS),.VDD(VDD),.Y(g28323),.A(g8580),.B(g27838));
  AND2 AND2_3247(.VSS(VSS),.VDD(VDD),.Y(g28324),.A(g27810),.B(g20659));
  AND2 AND2_3248(.VSS(VSS),.VDD(VDD),.Y(g28326),.A(g27865),.B(g22274));
  AND2 AND2_3249(.VSS(VSS),.VDD(VDD),.Y(g28327),.A(g27900),.B(g22275));
  AND2 AND2_3250(.VSS(VSS),.VDD(VDD),.Y(g28329),.A(g27823),.B(g20708));
  AND2 AND2_3251(.VSS(VSS),.VDD(VDD),.Y(g28330),.A(g27864),.B(g20711));
  AND2 AND2_3252(.VSS(VSS),.VDD(VDD),.Y(g28331),.A(g27802),.B(g22307));
  AND2 AND2_3253(.VSS(VSS),.VDD(VDD),.Y(g28332),.A(g27883),.B(g22331));
  AND2 AND2_3254(.VSS(VSS),.VDD(VDD),.Y(g28333),.A(g27882),.B(g20772));
  AND2 AND2_3255(.VSS(VSS),.VDD(VDD),.Y(g28334),.A(g27842),.B(g20793));
  AND2 AND2_3256(.VSS(VSS),.VDD(VDD),.Y(g28335),.A(g27814),.B(g22343));
  AND2 AND2_3257(.VSS(VSS),.VDD(VDD),.Y(g28336),.A(g27896),.B(g20810));
  AND2 AND2_3258(.VSS(VSS),.VDD(VDD),.Y(g28337),.A(g28002),.B(g19448));
  AND2 AND2_3259(.VSS(VSS),.VDD(VDD),.Y(g28338),.A(g28029),.B(g19475));
  AND2 AND2_3260(.VSS(VSS),.VDD(VDD),.Y(g28339),.A(g28059),.B(g19498));
  AND2 AND2_3261(.VSS(VSS),.VDD(VDD),.Y(g28340),.A(g28088),.B(g19519));
  AND2 AND2_3262(.VSS(VSS),.VDD(VDD),.Y(g28373),.A(g56),.B(g27969));
  AND2 AND2_3263(.VSS(VSS),.VDD(VDD),.Y(g28376),.A(g744),.B(g27990));
  AND2 AND2_3264(.VSS(VSS),.VDD(VDD),.Y(g28378),.A(g52),.B(g27776));
  AND3 AND3_255(.VSS(VSS),.VDD(VDD),.Y(g28379),.A(g27868),.B(g19390),.C(g19369));
  AND2 AND2_3265(.VSS(VSS),.VDD(VDD),.Y(g28380),.A(g1430),.B(g28014));
  AND2 AND2_3266(.VSS(VSS),.VDD(VDD),.Y(g28381),.A(g28157),.B(g9815));
  AND2 AND2_3267(.VSS(VSS),.VDD(VDD),.Y(g28383),.A(g740),.B(g27780));
  AND2 AND2_3268(.VSS(VSS),.VDD(VDD),.Y(g28385),.A(g2124),.B(g28041));
  AND2 AND2_3269(.VSS(VSS),.VDD(VDD),.Y(g28387),.A(g1426),.B(g27787));
  AND2 AND2_3270(.VSS(VSS),.VDD(VDD),.Y(g28389),.A(g2120),.B(g27794));
  AND2 AND2_3271(.VSS(VSS),.VDD(VDD),.Y(g28396),.A(g7754),.B(g27806));
  AND2 AND2_3272(.VSS(VSS),.VDD(VDD),.Y(g28398),.A(g7769),.B(g27817));
  AND2 AND2_3273(.VSS(VSS),.VDD(VDD),.Y(g28399),.A(g7776),.B(g27820));
  AND2 AND2_3274(.VSS(VSS),.VDD(VDD),.Y(g28401),.A(g7782),.B(g27831));
  AND2 AND2_3275(.VSS(VSS),.VDD(VDD),.Y(g28402),.A(g7785),.B(g27839));
  AND2 AND2_3276(.VSS(VSS),.VDD(VDD),.Y(g28404),.A(g7792),.B(g27843));
  AND2 AND2_3277(.VSS(VSS),.VDD(VDD),.Y(g28405),.A(g7796),.B(g27847));
  AND2 AND2_3278(.VSS(VSS),.VDD(VDD),.Y(g28407),.A(g7799),.B(g27858));
  AND2 AND2_3279(.VSS(VSS),.VDD(VDD),.Y(g28408),.A(g7806),.B(g27861));
  AND2 AND2_3280(.VSS(VSS),.VDD(VDD),.Y(g28411),.A(g7809),.B(g27872));
  AND2 AND2_3281(.VSS(VSS),.VDD(VDD),.Y(g28412),.A(g7812),.B(g27879));
  AND2 AND2_3282(.VSS(VSS),.VDD(VDD),.Y(g28416),.A(g7823),.B(g27889));
  AND2 AND2_3283(.VSS(VSS),.VDD(VDD),.Y(g28422),.A(g17640),.B(g28150));
  AND2 AND2_3284(.VSS(VSS),.VDD(VDD),.Y(g28423),.A(g17724),.B(g28152));
  AND2 AND2_3285(.VSS(VSS),.VDD(VDD),.Y(g28424),.A(g17741),.B(g28153));
  AND2 AND2_3286(.VSS(VSS),.VDD(VDD),.Y(g28426),.A(g28128),.B(g9170));
  AND2 AND2_3287(.VSS(VSS),.VDD(VDD),.Y(g28427),.A(g26092),.B(g28154));
  AND2 AND2_3288(.VSS(VSS),.VDD(VDD),.Y(g28428),.A(g17825),.B(g28155));
  AND2 AND2_3289(.VSS(VSS),.VDD(VDD),.Y(g28429),.A(g17842),.B(g28156));
  AND2 AND2_3290(.VSS(VSS),.VDD(VDD),.Y(g28430),.A(g28128),.B(g9196));
  AND2 AND2_3291(.VSS(VSS),.VDD(VDD),.Y(g28431),.A(g26092),.B(g28158));
  AND2 AND2_3292(.VSS(VSS),.VDD(VDD),.Y(g28433),.A(g28133),.B(g9212));
  AND2 AND2_3293(.VSS(VSS),.VDD(VDD),.Y(g28434),.A(g26114),.B(g28159));
  AND2 AND2_3294(.VSS(VSS),.VDD(VDD),.Y(g28435),.A(g17937),.B(g28160));
  AND2 AND2_3295(.VSS(VSS),.VDD(VDD),.Y(g28436),.A(g17954),.B(g28161));
  AND2 AND2_3296(.VSS(VSS),.VDD(VDD),.Y(g28438),.A(g17882),.B(g27919));
  AND2 AND2_3297(.VSS(VSS),.VDD(VDD),.Y(g28439),.A(g28128),.B(g9242));
  AND2 AND2_3298(.VSS(VSS),.VDD(VDD),.Y(g28440),.A(g26092),.B(g28162));
  AND2 AND2_3299(.VSS(VSS),.VDD(VDD),.Y(g28441),.A(g28133),.B(g9257));
  AND2 AND2_3300(.VSS(VSS),.VDD(VDD),.Y(g28442),.A(g26114),.B(g28163));
  AND2 AND2_3301(.VSS(VSS),.VDD(VDD),.Y(g28444),.A(g28137),.B(g9273));
  AND2 AND2_3302(.VSS(VSS),.VDD(VDD),.Y(g28445),.A(g26121),.B(g28164));
  AND2 AND2_3303(.VSS(VSS),.VDD(VDD),.Y(g28446),.A(g18048),.B(g28165));
  AND2 AND2_3304(.VSS(VSS),.VDD(VDD),.Y(g28448),.A(g17974),.B(g27928));
  AND2 AND2_3305(.VSS(VSS),.VDD(VDD),.Y(g28450),.A(g17993),.B(g27932));
  AND2 AND2_3306(.VSS(VSS),.VDD(VDD),.Y(g28451),.A(g28133),.B(g9320));
  AND2 AND2_3307(.VSS(VSS),.VDD(VDD),.Y(g28452),.A(g26114),.B(g28166));
  AND2 AND2_3308(.VSS(VSS),.VDD(VDD),.Y(g28453),.A(g28137),.B(g9335));
  AND2 AND2_3309(.VSS(VSS),.VDD(VDD),.Y(g28454),.A(g26121),.B(g28167));
  AND2 AND2_3310(.VSS(VSS),.VDD(VDD),.Y(g28456),.A(g28141),.B(g9351));
  AND2 AND2_3311(.VSS(VSS),.VDD(VDD),.Y(g28457),.A(g26131),.B(g28168));
  AND2 AND2_3312(.VSS(VSS),.VDD(VDD),.Y(g28459),.A(g18074),.B(g27939));
  AND2 AND2_3313(.VSS(VSS),.VDD(VDD),.Y(g28460),.A(g18091),.B(g27942));
  AND2 AND2_3314(.VSS(VSS),.VDD(VDD),.Y(g28462),.A(g18110),.B(g27946));
  AND2 AND2_3315(.VSS(VSS),.VDD(VDD),.Y(g28463),.A(g28137),.B(g9401));
  AND2 AND2_3316(.VSS(VSS),.VDD(VDD),.Y(g28464),.A(g26121),.B(g28169));
  AND2 AND2_3317(.VSS(VSS),.VDD(VDD),.Y(g28465),.A(g28141),.B(g9416));
  AND2 AND2_3318(.VSS(VSS),.VDD(VDD),.Y(g28466),.A(g26131),.B(g28170));
  AND2 AND2_3319(.VSS(VSS),.VDD(VDD),.Y(g28468),.A(g18265),.B(g28172));
  AND2 AND2_3320(.VSS(VSS),.VDD(VDD),.Y(g28469),.A(g18179),.B(g27952));
  AND2 AND2_3321(.VSS(VSS),.VDD(VDD),.Y(g28471),.A(g18190),.B(g27956));
  AND2 AND2_3322(.VSS(VSS),.VDD(VDD),.Y(g28472),.A(g18207),.B(g27959));
  AND2 AND2_3323(.VSS(VSS),.VDD(VDD),.Y(g28474),.A(g18226),.B(g27965));
  AND2 AND2_3324(.VSS(VSS),.VDD(VDD),.Y(g28475),.A(g28141),.B(g9498));
  AND2 AND2_3325(.VSS(VSS),.VDD(VDD),.Y(g28476),.A(g26131),.B(g28173));
  AND2 AND2_3326(.VSS(VSS),.VDD(VDD),.Y(g28477),.A(g18341),.B(g28174));
  AND2 AND2_3327(.VSS(VSS),.VDD(VDD),.Y(g28478),.A(g18358),.B(g28175));
  AND2 AND2_3328(.VSS(VSS),.VDD(VDD),.Y(g28479),.A(g18286),.B(g27973));
  AND2 AND2_3329(.VSS(VSS),.VDD(VDD),.Y(g28480),.A(g18297),.B(g27977));
  AND2 AND2_3330(.VSS(VSS),.VDD(VDD),.Y(g28481),.A(g18314),.B(g27981));
  AND2 AND2_3331(.VSS(VSS),.VDD(VDD),.Y(g28484),.A(g18436),.B(g28177));
  AND2 AND2_3332(.VSS(VSS),.VDD(VDD),.Y(g28485),.A(g18453),.B(g28178));
  AND2 AND2_3333(.VSS(VSS),.VDD(VDD),.Y(g28486),.A(g18379),.B(g27994));
  AND2 AND2_3334(.VSS(VSS),.VDD(VDD),.Y(g28487),.A(g18390),.B(g27999));
  AND2 AND2_3335(.VSS(VSS),.VDD(VDD),.Y(g28492),.A(g18509),.B(g28186));
  AND2 AND2_3336(.VSS(VSS),.VDD(VDD),.Y(g28493),.A(g18526),.B(g28187));
  AND2 AND2_3337(.VSS(VSS),.VDD(VDD),.Y(g28494),.A(g18474),.B(g28018));
  AND2 AND2_3338(.VSS(VSS),.VDD(VDD),.Y(g28497),.A(g18573),.B(g28190));
  AND2 AND2_3339(.VSS(VSS),.VDD(VDD),.Y(g28657),.A(g27925),.B(g13700));
  AND2 AND2_3340(.VSS(VSS),.VDD(VDD),.Y(g28659),.A(g27917),.B(g13736));
  AND2 AND2_3341(.VSS(VSS),.VDD(VDD),.Y(g28660),.A(g27916),.B(g11911));
  AND2 AND2_3342(.VSS(VSS),.VDD(VDD),.Y(g28662),.A(g27911),.B(g11951));
  AND2 AND2_3343(.VSS(VSS),.VDD(VDD),.Y(g28663),.A(g27906),.B(g11997));
  AND2 AND2_3344(.VSS(VSS),.VDD(VDD),.Y(g28664),.A(g27997),.B(g12055));
  AND2 AND2_3345(.VSS(VSS),.VDD(VDD),.Y(g28665),.A(g27827),.B(g22222));
  AND2 AND2_3346(.VSS(VSS),.VDD(VDD),.Y(g28666),.A(g27980),.B(g12106));
  AND2 AND2_3347(.VSS(VSS),.VDD(VDD),.Y(g28667),.A(g27964),.B(g13852));
  AND2 AND2_3348(.VSS(VSS),.VDD(VDD),.Y(g28669),.A(g27897),.B(g22233));
  AND2 AND2_3349(.VSS(VSS),.VDD(VDD),.Y(g28670),.A(g27798),.B(g21935));
  AND2 AND2_3350(.VSS(VSS),.VDD(VDD),.Y(g28671),.A(g27962),.B(g12161));
  AND2 AND2_3351(.VSS(VSS),.VDD(VDD),.Y(g28672),.A(g27950),.B(g13859));
  AND2 AND2_3352(.VSS(VSS),.VDD(VDD),.Y(g28707),.A(g12436),.B(g28379));
  AND2 AND2_3353(.VSS(VSS),.VDD(VDD),.Y(g28708),.A(g28392),.B(g22260));
  AND2 AND2_3354(.VSS(VSS),.VDD(VDD),.Y(g28709),.A(g28400),.B(g22261));
  AND2 AND2_3355(.VSS(VSS),.VDD(VDD),.Y(g28710),.A(g28403),.B(g22262));
  AND2 AND2_3356(.VSS(VSS),.VDD(VDD),.Y(g28711),.A(g10749),.B(g28415));
  AND2 AND2_3357(.VSS(VSS),.VDD(VDD),.Y(g28712),.A(g28406),.B(g22276));
  AND2 AND2_3358(.VSS(VSS),.VDD(VDD),.Y(g28713),.A(g28410),.B(g22290));
  AND2 AND2_3359(.VSS(VSS),.VDD(VDD),.Y(g28714),.A(g28394),.B(g22306));
  AND2 AND2_3360(.VSS(VSS),.VDD(VDD),.Y(g28715),.A(g28414),.B(g22332));
  AND2 AND2_3361(.VSS(VSS),.VDD(VDD),.Y(g28716),.A(g28449),.B(g19319));
  AND2 AND2_3362(.VSS(VSS),.VDD(VDD),.Y(g28717),.A(g28461),.B(g19346));
  AND2 AND2_3363(.VSS(VSS),.VDD(VDD),.Y(g28718),.A(g28473),.B(g19380));
  AND2 AND2_3364(.VSS(VSS),.VDD(VDD),.Y(g28719),.A(g28482),.B(g19412));
  AND2 AND2_3365(.VSS(VSS),.VDD(VDD),.Y(g28722),.A(g28523),.B(g16694));
  AND2 AND2_3366(.VSS(VSS),.VDD(VDD),.Y(g28724),.A(g28551),.B(g16725));
  AND2 AND2_3367(.VSS(VSS),.VDD(VDD),.Y(g28726),.A(g28578),.B(g16767));
  AND2 AND2_3368(.VSS(VSS),.VDD(VDD),.Y(g28729),.A(g28606),.B(g16794));
  AND2 AND2_3369(.VSS(VSS),.VDD(VDD),.Y(g28834),.A(g5751),.B(g28483));
  AND2 AND2_3370(.VSS(VSS),.VDD(VDD),.Y(g28836),.A(g5810),.B(g28491));
  AND2 AND2_3371(.VSS(VSS),.VDD(VDD),.Y(g28838),.A(g5866),.B(g28496));
  AND2 AND2_3372(.VSS(VSS),.VDD(VDD),.Y(g28840),.A(g5913),.B(g28500));
  AND2 AND2_3373(.VSS(VSS),.VDD(VDD),.Y(g28841),.A(g27834),.B(g28554));
  AND2 AND2_3374(.VSS(VSS),.VDD(VDD),.Y(g28843),.A(g27834),.B(g28581));
  AND2 AND2_3375(.VSS(VSS),.VDD(VDD),.Y(g28844),.A(g27850),.B(g28582));
  AND2 AND2_3376(.VSS(VSS),.VDD(VDD),.Y(g28846),.A(g27834),.B(g28608));
  AND2 AND2_3377(.VSS(VSS),.VDD(VDD),.Y(g28847),.A(g27850),.B(g28609));
  AND2 AND2_3378(.VSS(VSS),.VDD(VDD),.Y(g28848),.A(g27875),.B(g28610));
  AND2 AND2_3379(.VSS(VSS),.VDD(VDD),.Y(g28849),.A(g27850),.B(g28616));
  AND2 AND2_3380(.VSS(VSS),.VDD(VDD),.Y(g28850),.A(g27875),.B(g28617));
  AND2 AND2_3381(.VSS(VSS),.VDD(VDD),.Y(g28851),.A(g27892),.B(g28618));
  AND2 AND2_3382(.VSS(VSS),.VDD(VDD),.Y(g28852),.A(g27875),.B(g28623));
  AND2 AND2_3383(.VSS(VSS),.VDD(VDD),.Y(g28853),.A(g27892),.B(g28624));
  AND2 AND2_3384(.VSS(VSS),.VDD(VDD),.Y(g28854),.A(g27892),.B(g28629));
  AND2 AND2_3385(.VSS(VSS),.VDD(VDD),.Y(g28880),.A(g13946),.B(g28639));
  AND2 AND2_3386(.VSS(VSS),.VDD(VDD),.Y(g28881),.A(g28612),.B(g9199));
  AND2 AND2_3387(.VSS(VSS),.VDD(VDD),.Y(g28892),.A(g14001),.B(g28640));
  AND2 AND2_3388(.VSS(VSS),.VDD(VDD),.Y(g28893),.A(g28612),.B(g9245));
  AND2 AND2_3389(.VSS(VSS),.VDD(VDD),.Y(g28897),.A(g14016),.B(g28641));
  AND2 AND2_3390(.VSS(VSS),.VDD(VDD),.Y(g28898),.A(g28619),.B(g9260));
  AND2 AND2_3391(.VSS(VSS),.VDD(VDD),.Y(g28909),.A(g14062),.B(g28642));
  AND2 AND2_3392(.VSS(VSS),.VDD(VDD),.Y(g28910),.A(g28612),.B(g9303));
  AND2 AND2_3393(.VSS(VSS),.VDD(VDD),.Y(g28914),.A(g14092),.B(g28643));
  AND2 AND2_3394(.VSS(VSS),.VDD(VDD),.Y(g28915),.A(g28619),.B(g9323));
  AND2 AND2_3395(.VSS(VSS),.VDD(VDD),.Y(g28919),.A(g14107),.B(g28644));
  AND2 AND2_3396(.VSS(VSS),.VDD(VDD),.Y(g28923),.A(g28625),.B(g9338));
  AND2 AND2_3397(.VSS(VSS),.VDD(VDD),.Y(g28931),.A(g14153),.B(g28645));
  AND2 AND2_3398(.VSS(VSS),.VDD(VDD),.Y(g28935),.A(g14177),.B(g28646));
  AND2 AND2_3399(.VSS(VSS),.VDD(VDD),.Y(g28936),.A(g28619),.B(g9384));
  AND2 AND2_3400(.VSS(VSS),.VDD(VDD),.Y(g28940),.A(g14207),.B(g28647));
  AND2 AND2_3401(.VSS(VSS),.VDD(VDD),.Y(g28944),.A(g28625),.B(g9404));
  AND2 AND2_3402(.VSS(VSS),.VDD(VDD),.Y(g28948),.A(g14222),.B(g28648));
  AND2 AND2_3403(.VSS(VSS),.VDD(VDD),.Y(g28949),.A(g28630),.B(g9419));
  AND2 AND2_3404(.VSS(VSS),.VDD(VDD),.Y(g28958),.A(g14268),.B(g28649));
  AND2 AND2_3405(.VSS(VSS),.VDD(VDD),.Y(g28962),.A(g14292),.B(g28650));
  AND2 AND2_3406(.VSS(VSS),.VDD(VDD),.Y(g28966),.A(g28625),.B(g9481));
  AND2 AND2_3407(.VSS(VSS),.VDD(VDD),.Y(g28970),.A(g14322),.B(g28651));
  AND2 AND2_3408(.VSS(VSS),.VDD(VDD),.Y(g28971),.A(g28630),.B(g9501));
  AND2 AND2_3409(.VSS(VSS),.VDD(VDD),.Y(g28986),.A(g14390),.B(g28652));
  AND2 AND2_3410(.VSS(VSS),.VDD(VDD),.Y(g28996),.A(g14414),.B(g28653));
  AND2 AND2_3411(.VSS(VSS),.VDD(VDD),.Y(g28997),.A(g28630),.B(g9623));
  AND2 AND2_3412(.VSS(VSS),.VDD(VDD),.Y(g29022),.A(g14502),.B(g28655));
  AND2 AND2_3413(.VSS(VSS),.VDD(VDD),.Y(g29130),.A(g28397),.B(g22221));
  AND2 AND2_3414(.VSS(VSS),.VDD(VDD),.Y(g29174),.A(g29031),.B(g20684));
  AND2 AND2_3415(.VSS(VSS),.VDD(VDD),.Y(g29175),.A(g29009),.B(g20687));
  AND2 AND2_3416(.VSS(VSS),.VDD(VDD),.Y(g29176),.A(g29097),.B(g20690));
  AND2 AND2_3417(.VSS(VSS),.VDD(VDD),.Y(g29180),.A(g28982),.B(g20714));
  AND2 AND2_3418(.VSS(VSS),.VDD(VDD),.Y(g29183),.A(g29064),.B(g20739));
  AND2 AND2_3419(.VSS(VSS),.VDD(VDD),.Y(g29186),.A(g29063),.B(g20769));
  AND2 AND2_3420(.VSS(VSS),.VDD(VDD),.Y(g29188),.A(g29083),.B(g20796));
  AND2 AND2_3421(.VSS(VSS),.VDD(VDD),.Y(g29196),.A(g15022),.B(g28741));
  AND2 AND2_3422(.VSS(VSS),.VDD(VDD),.Y(g29200),.A(g15096),.B(g28751));
  AND2 AND2_3423(.VSS(VSS),.VDD(VDD),.Y(g29203),.A(g15118),.B(g28755));
  AND2 AND2_3424(.VSS(VSS),.VDD(VDD),.Y(g29208),.A(g15188),.B(g28764));
  AND2 AND2_3425(.VSS(VSS),.VDD(VDD),.Y(g29211),.A(g15210),.B(g28768));
  AND2 AND2_3426(.VSS(VSS),.VDD(VDD),.Y(g29217),.A(g15274),.B(g28775));
  AND2 AND2_3427(.VSS(VSS),.VDD(VDD),.Y(g29220),.A(g15296),.B(g28779));
  AND2 AND2_3428(.VSS(VSS),.VDD(VDD),.Y(g29225),.A(g15366),.B(g28785));
  AND2 AND2_3429(.VSS(VSS),.VDD(VDD),.Y(g29229),.A(g9293),.B(g28791));
  AND2 AND2_3430(.VSS(VSS),.VDD(VDD),.Y(g29232),.A(g9356),.B(g28796));
  AND2 AND2_3431(.VSS(VSS),.VDD(VDD),.Y(g29233),.A(g9374),.B(g28799));
  AND2 AND2_3432(.VSS(VSS),.VDD(VDD),.Y(g29234),.A(g9427),.B(g28804));
  AND2 AND2_3433(.VSS(VSS),.VDD(VDD),.Y(g29235),.A(g9453),.B(g28807));
  AND2 AND2_3434(.VSS(VSS),.VDD(VDD),.Y(g29236),.A(g9471),.B(g28810));
  AND2 AND2_3435(.VSS(VSS),.VDD(VDD),.Y(g29238),.A(g9569),.B(g28814));
  AND2 AND2_3436(.VSS(VSS),.VDD(VDD),.Y(g29239),.A(g9595),.B(g28817));
  AND2 AND2_3437(.VSS(VSS),.VDD(VDD),.Y(g29240),.A(g9613),.B(g28820));
  AND2 AND2_3438(.VSS(VSS),.VDD(VDD),.Y(g29241),.A(g9711),.B(g28823));
  AND2 AND2_3439(.VSS(VSS),.VDD(VDD),.Y(g29242),.A(g9737),.B(g28826));
  AND2 AND2_3440(.VSS(VSS),.VDD(VDD),.Y(g29243),.A(g9857),.B(g28829));
  AND2 AND2_3441(.VSS(VSS),.VDD(VDD),.Y(g29248),.A(g28855),.B(g8836));
  AND2 AND2_3442(.VSS(VSS),.VDD(VDD),.Y(g29251),.A(g28855),.B(g8856));
  AND2 AND2_3443(.VSS(VSS),.VDD(VDD),.Y(g29252),.A(g28859),.B(g8863));
  AND2 AND2_3444(.VSS(VSS),.VDD(VDD),.Y(g29255),.A(g28855),.B(g8885));
  AND2 AND2_3445(.VSS(VSS),.VDD(VDD),.Y(g29256),.A(g28859),.B(g8894));
  AND2 AND2_3446(.VSS(VSS),.VDD(VDD),.Y(g29257),.A(g28863),.B(g8901));
  AND2 AND2_3447(.VSS(VSS),.VDD(VDD),.Y(g29259),.A(g28859),.B(g8925));
  AND2 AND2_3448(.VSS(VSS),.VDD(VDD),.Y(g29260),.A(g28863),.B(g8934));
  AND2 AND2_3449(.VSS(VSS),.VDD(VDD),.Y(g29261),.A(g28867),.B(g8941));
  AND2 AND2_3450(.VSS(VSS),.VDD(VDD),.Y(g29262),.A(g28863),.B(g8965));
  AND2 AND2_3451(.VSS(VSS),.VDD(VDD),.Y(g29263),.A(g28867),.B(g8974));
  AND2 AND2_3452(.VSS(VSS),.VDD(VDD),.Y(g29264),.A(g28867),.B(g8997));
  AND2 AND2_3453(.VSS(VSS),.VDD(VDD),.Y(g29284),.A(g29001),.B(g28871));
  AND2 AND2_3454(.VSS(VSS),.VDD(VDD),.Y(g29289),.A(g29030),.B(g28883));
  AND2 AND2_3455(.VSS(VSS),.VDD(VDD),.Y(g29294),.A(g29053),.B(g28900));
  AND2 AND2_3456(.VSS(VSS),.VDD(VDD),.Y(g29300),.A(g29072),.B(g28925));
  AND2 AND2_3457(.VSS(VSS),.VDD(VDD),.Y(g29302),.A(g29026),.B(g28928));
  AND2 AND2_3458(.VSS(VSS),.VDD(VDD),.Y(g29310),.A(g28978),.B(g28951));
  AND2 AND2_3459(.VSS(VSS),.VDD(VDD),.Y(g29312),.A(g29049),.B(g28955));
  AND2 AND2_3460(.VSS(VSS),.VDD(VDD),.Y(g29320),.A(g29088),.B(g28972));
  AND2 AND2_3461(.VSS(VSS),.VDD(VDD),.Y(g29321),.A(g29008),.B(g28979));
  AND2 AND2_3462(.VSS(VSS),.VDD(VDD),.Y(g29323),.A(g29068),.B(g28983));
  AND2 AND2_3463(.VSS(VSS),.VDD(VDD),.Y(g29329),.A(g29096),.B(g29002));
  AND2 AND2_3464(.VSS(VSS),.VDD(VDD),.Y(g29330),.A(g29038),.B(g29010));
  AND2 AND2_3465(.VSS(VSS),.VDD(VDD),.Y(g29332),.A(g29080),.B(g29019));
  AND2 AND2_3466(.VSS(VSS),.VDD(VDD),.Y(g29336),.A(g29045),.B(g29023));
  AND2 AND2_3467(.VSS(VSS),.VDD(VDD),.Y(g29337),.A(g29103),.B(g29032));
  AND2 AND2_3468(.VSS(VSS),.VDD(VDD),.Y(g29338),.A(g29060),.B(g29042));
  AND2 AND2_3469(.VSS(VSS),.VDD(VDD),.Y(g29341),.A(g29062),.B(g29046));
  AND2 AND2_3470(.VSS(VSS),.VDD(VDD),.Y(g29342),.A(g29107),.B(g29054));
  AND2 AND2_3471(.VSS(VSS),.VDD(VDD),.Y(g29344),.A(g29076),.B(g29065));
  AND2 AND2_3472(.VSS(VSS),.VDD(VDD),.Y(g29346),.A(g29087),.B(g29077));
  AND2 AND2_3473(.VSS(VSS),.VDD(VDD),.Y(g29411),.A(g29090),.B(g21932));
  AND2 AND2_3474(.VSS(VSS),.VDD(VDD),.Y(g29464),.A(g29190),.B(g8375));
  AND2 AND2_3475(.VSS(VSS),.VDD(VDD),.Y(g29465),.A(g29191),.B(g8424));
  AND2 AND2_3476(.VSS(VSS),.VDD(VDD),.Y(g29466),.A(g8587),.B(g29265));
  AND2 AND2_3477(.VSS(VSS),.VDD(VDD),.Y(g29467),.A(g29340),.B(g19467));
  AND2 AND2_3478(.VSS(VSS),.VDD(VDD),.Y(g29468),.A(g29343),.B(g19490));
  AND2 AND2_3479(.VSS(VSS),.VDD(VDD),.Y(g29469),.A(g29345),.B(g19511));
  AND2 AND2_3480(.VSS(VSS),.VDD(VDD),.Y(g29470),.A(g29347),.B(g19530));
  AND2 AND2_3481(.VSS(VSS),.VDD(VDD),.Y(g29471),.A(g21461),.B(g29266));
  AND2 AND2_3482(.VSS(VSS),.VDD(VDD),.Y(g29472),.A(g21461),.B(g29268));
  AND2 AND2_3483(.VSS(VSS),.VDD(VDD),.Y(g29473),.A(g21508),.B(g29269));
  AND2 AND2_3484(.VSS(VSS),.VDD(VDD),.Y(g29474),.A(g21508),.B(g29271));
  AND2 AND2_3485(.VSS(VSS),.VDD(VDD),.Y(g29475),.A(g21544),.B(g29272));
  AND2 AND2_3486(.VSS(VSS),.VDD(VDD),.Y(g29476),.A(g21544),.B(g29274));
  AND2 AND2_3487(.VSS(VSS),.VDD(VDD),.Y(g29477),.A(g21580),.B(g29275));
  AND2 AND2_3488(.VSS(VSS),.VDD(VDD),.Y(g29478),.A(g21580),.B(g29277));
  AND2 AND2_3489(.VSS(VSS),.VDD(VDD),.Y(g29479),.A(g21461),.B(g29280));
  AND2 AND2_3490(.VSS(VSS),.VDD(VDD),.Y(g29480),.A(g21461),.B(g29282));
  AND2 AND2_3491(.VSS(VSS),.VDD(VDD),.Y(g29481),.A(g21508),.B(g29283));
  AND2 AND2_3492(.VSS(VSS),.VDD(VDD),.Y(g29482),.A(g21461),.B(g29285));
  AND2 AND2_3493(.VSS(VSS),.VDD(VDD),.Y(g29483),.A(g21508),.B(g29286));
  AND2 AND2_3494(.VSS(VSS),.VDD(VDD),.Y(g29484),.A(g21544),.B(g29287));
  AND2 AND2_3495(.VSS(VSS),.VDD(VDD),.Y(g29485),.A(g21508),.B(g29290));
  AND2 AND2_3496(.VSS(VSS),.VDD(VDD),.Y(g29486),.A(g21544),.B(g29291));
  AND2 AND2_3497(.VSS(VSS),.VDD(VDD),.Y(g29487),.A(g21580),.B(g29292));
  AND2 AND2_3498(.VSS(VSS),.VDD(VDD),.Y(g29488),.A(g21544),.B(g29295));
  AND2 AND2_3499(.VSS(VSS),.VDD(VDD),.Y(g29489),.A(g21580),.B(g29296));
  AND2 AND2_3500(.VSS(VSS),.VDD(VDD),.Y(g29490),.A(g21580),.B(g29301));
  AND2 AND2_3501(.VSS(VSS),.VDD(VDD),.Y(g29502),.A(g29350),.B(g8912));
  AND2 AND2_3502(.VSS(VSS),.VDD(VDD),.Y(g29518),.A(g28728),.B(g29360));
  AND2 AND2_3503(.VSS(VSS),.VDD(VDD),.Y(g29520),.A(g28731),.B(g29361));
  AND2 AND2_3504(.VSS(VSS),.VDD(VDD),.Y(g29521),.A(g28733),.B(g29362));
  AND2 AND2_3505(.VSS(VSS),.VDD(VDD),.Y(g29522),.A(g27735),.B(g29363));
  AND2 AND2_3506(.VSS(VSS),.VDD(VDD),.Y(g29523),.A(g28737),.B(g29364));
  AND2 AND2_3507(.VSS(VSS),.VDD(VDD),.Y(g29524),.A(g28739),.B(g29365));
  AND2 AND2_3508(.VSS(VSS),.VDD(VDD),.Y(g29525),.A(g29195),.B(g29366));
  AND2 AND2_3509(.VSS(VSS),.VDD(VDD),.Y(g29526),.A(g27741),.B(g29367));
  AND2 AND2_3510(.VSS(VSS),.VDD(VDD),.Y(g29527),.A(g28748),.B(g29368));
  AND2 AND2_3511(.VSS(VSS),.VDD(VDD),.Y(g29528),.A(g28750),.B(g29369));
  AND2 AND2_3512(.VSS(VSS),.VDD(VDD),.Y(g29529),.A(g29199),.B(g29370));
  AND2 AND2_3513(.VSS(VSS),.VDD(VDD),.Y(g29531),.A(g29202),.B(g29371));
  AND2 AND2_3514(.VSS(VSS),.VDD(VDD),.Y(g29532),.A(g27746),.B(g29372));
  AND2 AND2_3515(.VSS(VSS),.VDD(VDD),.Y(g29533),.A(g28762),.B(g29373));
  AND2 AND2_3516(.VSS(VSS),.VDD(VDD),.Y(g29534),.A(g29206),.B(g29374));
  AND2 AND2_3517(.VSS(VSS),.VDD(VDD),.Y(g29536),.A(g29207),.B(g29375));
  AND2 AND2_3518(.VSS(VSS),.VDD(VDD),.Y(g29538),.A(g29210),.B(g29376));
  AND2 AND2_3519(.VSS(VSS),.VDD(VDD),.Y(g29539),.A(g27754),.B(g29377));
  AND2 AND2_3520(.VSS(VSS),.VDD(VDD),.Y(g29540),.A(g26041),.B(g29378));
  AND2 AND2_3521(.VSS(VSS),.VDD(VDD),.Y(g29541),.A(g29214),.B(g29379));
  AND2 AND2_3522(.VSS(VSS),.VDD(VDD),.Y(g29543),.A(g29215),.B(g29380));
  AND2 AND2_3523(.VSS(VSS),.VDD(VDD),.Y(g29545),.A(g29216),.B(g29381));
  AND2 AND2_3524(.VSS(VSS),.VDD(VDD),.Y(g29547),.A(g29219),.B(g29382));
  AND2 AND2_3525(.VSS(VSS),.VDD(VDD),.Y(g29548),.A(g28784),.B(g29383));
  AND2 AND2_3526(.VSS(VSS),.VDD(VDD),.Y(g29549),.A(g26043),.B(g29384));
  AND2 AND2_3527(.VSS(VSS),.VDD(VDD),.Y(g29550),.A(g29222),.B(g29385));
  AND2 AND2_3528(.VSS(VSS),.VDD(VDD),.Y(g29553),.A(g29223),.B(g29386));
  AND2 AND2_3529(.VSS(VSS),.VDD(VDD),.Y(g29555),.A(g29224),.B(g29387));
  AND2 AND2_3530(.VSS(VSS),.VDD(VDD),.Y(g29557),.A(g28789),.B(g29388));
  AND2 AND2_3531(.VSS(VSS),.VDD(VDD),.Y(g29558),.A(g28790),.B(g29389));
  AND2 AND2_3532(.VSS(VSS),.VDD(VDD),.Y(g29559),.A(g26045),.B(g29390));
  AND2 AND2_3533(.VSS(VSS),.VDD(VDD),.Y(g29560),.A(g29227),.B(g29391));
  AND2 AND2_3534(.VSS(VSS),.VDD(VDD),.Y(g29562),.A(g29228),.B(g29392));
  AND2 AND2_3535(.VSS(VSS),.VDD(VDD),.Y(g29564),.A(g28794),.B(g29393));
  AND2 AND2_3536(.VSS(VSS),.VDD(VDD),.Y(g29565),.A(g28795),.B(g29394));
  AND2 AND2_3537(.VSS(VSS),.VDD(VDD),.Y(g29566),.A(g26047),.B(g29395));
  AND2 AND2_3538(.VSS(VSS),.VDD(VDD),.Y(g29567),.A(g29231),.B(g29396));
  AND2 AND2_3539(.VSS(VSS),.VDD(VDD),.Y(g29572),.A(g28802),.B(g29397));
  AND2 AND2_3540(.VSS(VSS),.VDD(VDD),.Y(g29573),.A(g28803),.B(g29398));
  AND2 AND2_3541(.VSS(VSS),.VDD(VDD),.Y(g29575),.A(g28813),.B(g29402));
  AND2 AND2_3542(.VSS(VSS),.VDD(VDD),.Y(g29607),.A(g29193),.B(g11056));
  AND2 AND2_3543(.VSS(VSS),.VDD(VDD),.Y(g29610),.A(g29349),.B(g11123));
  AND2 AND2_3544(.VSS(VSS),.VDD(VDD),.Y(g29614),.A(g29359),.B(g11182));
  AND2 AND2_3545(.VSS(VSS),.VDD(VDD),.Y(g29615),.A(g29245),.B(g11185));
  AND2 AND2_3546(.VSS(VSS),.VDD(VDD),.Y(g29619),.A(g29247),.B(g11259));
  AND2 AND2_3547(.VSS(VSS),.VDD(VDD),.Y(g29622),.A(g29250),.B(g11327));
  AND2 AND2_3548(.VSS(VSS),.VDD(VDD),.Y(g29624),.A(g29254),.B(g11407));
  AND2 AND2_3549(.VSS(VSS),.VDD(VDD),.Y(g29625),.A(g29189),.B(g11472));
  AND2 AND2_3550(.VSS(VSS),.VDD(VDD),.Y(g29626),.A(g29318),.B(g11478));
  AND2 AND2_3551(.VSS(VSS),.VDD(VDD),.Y(g29790),.A(g29491),.B(g10918));
  AND2 AND2_3552(.VSS(VSS),.VDD(VDD),.Y(g29792),.A(g29491),.B(g10977));
  AND2 AND2_3553(.VSS(VSS),.VDD(VDD),.Y(g29793),.A(g29491),.B(g11063));
  AND2 AND2_3554(.VSS(VSS),.VDD(VDD),.Y(g29810),.A(g29748),.B(g22248));
  AND2 AND2_3555(.VSS(VSS),.VDD(VDD),.Y(g29811),.A(g29703),.B(g20644));
  AND2 AND2_3556(.VSS(VSS),.VDD(VDD),.Y(g29812),.A(g29762),.B(g12223));
  AND2 AND2_3557(.VSS(VSS),.VDD(VDD),.Y(g29813),.A(g29760),.B(g13869));
  AND2 AND2_3558(.VSS(VSS),.VDD(VDD),.Y(g29814),.A(g29728),.B(g22266));
  AND2 AND2_3559(.VSS(VSS),.VDD(VDD),.Y(g29815),.A(g29727),.B(g20662));
  AND2 AND2_3560(.VSS(VSS),.VDD(VDD),.Y(g29816),.A(g29759),.B(g13883));
  AND2 AND2_3561(.VSS(VSS),.VDD(VDD),.Y(g29817),.A(g29709),.B(g20694));
  AND2 AND2_3562(.VSS(VSS),.VDD(VDD),.Y(g29818),.A(g29732),.B(g22293));
  AND2 AND2_3563(.VSS(VSS),.VDD(VDD),.Y(g29819),.A(g29751),.B(g22294));
  AND2 AND2_3564(.VSS(VSS),.VDD(VDD),.Y(g29820),.A(g29717),.B(g20743));
  AND2 AND2_3565(.VSS(VSS),.VDD(VDD),.Y(g29821),.A(g29731),.B(g20746));
  AND2 AND2_3566(.VSS(VSS),.VDD(VDD),.Y(g29822),.A(g29705),.B(g22335));
  AND2 AND2_3567(.VSS(VSS),.VDD(VDD),.Y(g29827),.A(g29741),.B(g22356));
  AND2 AND2_3568(.VSS(VSS),.VDD(VDD),.Y(g29828),.A(g29740),.B(g20802));
  AND2 AND2_3569(.VSS(VSS),.VDD(VDD),.Y(g29833),.A(g29725),.B(g20813));
  AND2 AND2_3570(.VSS(VSS),.VDD(VDD),.Y(g29834),.A(g29713),.B(g22366));
  AND2 AND2_3571(.VSS(VSS),.VDD(VDD),.Y(g29839),.A(g29747),.B(g20827));
  AND3 AND3_256(.VSS(VSS),.VDD(VDD),.Y(g29909),.A(g29735),.B(g19420),.C(g19401));
  AND2 AND2_3572(.VSS(VSS),.VDD(VDD),.Y(g29910),.A(g29779),.B(g9961));
  AND2 AND2_3573(.VSS(VSS),.VDD(VDD),.Y(g29942),.A(g29771),.B(g28877));
  AND2 AND2_3574(.VSS(VSS),.VDD(VDD),.Y(g29944),.A(g29782),.B(g28889));
  AND2 AND2_3575(.VSS(VSS),.VDD(VDD),.Y(g29945),.A(g29773),.B(g28894));
  AND2 AND2_3576(.VSS(VSS),.VDD(VDD),.Y(g29946),.A(g29778),.B(g28906));
  AND2 AND2_3577(.VSS(VSS),.VDD(VDD),.Y(g29947),.A(g29785),.B(g28911));
  AND2 AND2_3578(.VSS(VSS),.VDD(VDD),.Y(g29948),.A(g29775),.B(g28916));
  AND2 AND2_3579(.VSS(VSS),.VDD(VDD),.Y(g29949),.A(g29781),.B(g28932));
  AND2 AND2_3580(.VSS(VSS),.VDD(VDD),.Y(g29950),.A(g29788),.B(g28937));
  AND2 AND2_3581(.VSS(VSS),.VDD(VDD),.Y(g29951),.A(g29777),.B(g28945));
  AND2 AND2_3582(.VSS(VSS),.VDD(VDD),.Y(g29952),.A(g29784),.B(g28959));
  AND2 AND2_3583(.VSS(VSS),.VDD(VDD),.Y(g29953),.A(g29791),.B(g28967));
  AND2 AND2_3584(.VSS(VSS),.VDD(VDD),.Y(g29954),.A(g29770),.B(g28975));
  AND2 AND2_3585(.VSS(VSS),.VDD(VDD),.Y(g29955),.A(g29787),.B(g28993));
  AND2 AND2_3586(.VSS(VSS),.VDD(VDD),.Y(g29956),.A(g29780),.B(g28998));
  AND2 AND2_3587(.VSS(VSS),.VDD(VDD),.Y(g29957),.A(g29772),.B(g29005));
  AND2 AND2_3588(.VSS(VSS),.VDD(VDD),.Y(g29958),.A(g29783),.B(g29027));
  AND2 AND2_3589(.VSS(VSS),.VDD(VDD),.Y(g29959),.A(g29774),.B(g29035));
  AND2 AND2_3590(.VSS(VSS),.VDD(VDD),.Y(g29960),.A(g29786),.B(g29050));
  AND2 AND2_3591(.VSS(VSS),.VDD(VDD),.Y(g29961),.A(g29776),.B(g29057));
  AND2 AND2_3592(.VSS(VSS),.VDD(VDD),.Y(g29962),.A(g29789),.B(g29069));
  AND2 AND2_3593(.VSS(VSS),.VDD(VDD),.Y(g29963),.A(g29758),.B(g13737));
  AND2 AND2_3594(.VSS(VSS),.VDD(VDD),.Y(g29964),.A(g29757),.B(g13786));
  AND2 AND2_3595(.VSS(VSS),.VDD(VDD),.Y(g29965),.A(g29756),.B(g11961));
  AND2 AND2_3596(.VSS(VSS),.VDD(VDD),.Y(g29966),.A(g29755),.B(g12004));
  AND2 AND2_3597(.VSS(VSS),.VDD(VDD),.Y(g29967),.A(g29754),.B(g12066));
  AND2 AND2_3598(.VSS(VSS),.VDD(VDD),.Y(g29968),.A(g29765),.B(g12119));
  AND2 AND2_3599(.VSS(VSS),.VDD(VDD),.Y(g29969),.A(g29721),.B(g22237));
  AND2 AND2_3600(.VSS(VSS),.VDD(VDD),.Y(g29970),.A(g29764),.B(g12178));
  AND2 AND2_3601(.VSS(VSS),.VDD(VDD),.Y(g29971),.A(g29763),.B(g13861));
  AND2 AND2_3602(.VSS(VSS),.VDD(VDD),.Y(g29980),.A(g29881),.B(g8324));
  AND2 AND2_3603(.VSS(VSS),.VDD(VDD),.Y(g29981),.A(g29869),.B(g8330));
  AND2 AND2_3604(.VSS(VSS),.VDD(VDD),.Y(g29982),.A(g29893),.B(g8336));
  AND2 AND2_3605(.VSS(VSS),.VDD(VDD),.Y(g29983),.A(g29885),.B(g8344));
  AND2 AND2_3606(.VSS(VSS),.VDD(VDD),.Y(g29984),.A(g29873),.B(g8351));
  AND2 AND2_3607(.VSS(VSS),.VDD(VDD),.Y(g29985),.A(g29897),.B(g8363));
  AND2 AND2_3608(.VSS(VSS),.VDD(VDD),.Y(g29986),.A(g29877),.B(g8366));
  AND2 AND2_3609(.VSS(VSS),.VDD(VDD),.Y(g29987),.A(g29889),.B(g8369));
  AND2 AND2_3610(.VSS(VSS),.VDD(VDD),.Y(g29988),.A(g29881),.B(g8382));
  AND2 AND2_3611(.VSS(VSS),.VDD(VDD),.Y(g29989),.A(g29893),.B(g8391));
  AND2 AND2_3612(.VSS(VSS),.VDD(VDD),.Y(g29990),.A(g29885),.B(g8397));
  AND2 AND2_3613(.VSS(VSS),.VDD(VDD),.Y(g29991),.A(g29901),.B(g8403));
  AND2 AND2_3614(.VSS(VSS),.VDD(VDD),.Y(g29992),.A(g12441),.B(g29909));
  AND2 AND2_3615(.VSS(VSS),.VDD(VDD),.Y(g29993),.A(g29897),.B(g8411));
  AND2 AND2_3616(.VSS(VSS),.VDD(VDD),.Y(g29994),.A(g29889),.B(g8418));
  AND2 AND2_3617(.VSS(VSS),.VDD(VDD),.Y(g29995),.A(g29893),.B(g8434));
  AND2 AND2_3618(.VSS(VSS),.VDD(VDD),.Y(g29996),.A(g29901),.B(g8443));
  AND2 AND2_3619(.VSS(VSS),.VDD(VDD),.Y(g29997),.A(g29918),.B(g22277));
  AND2 AND2_3620(.VSS(VSS),.VDD(VDD),.Y(g29998),.A(g29922),.B(g22278));
  AND2 AND2_3621(.VSS(VSS),.VDD(VDD),.Y(g29999),.A(g29924),.B(g22279));
  AND2 AND2_3622(.VSS(VSS),.VDD(VDD),.Y(g30000),.A(g10767),.B(g29930));
  AND2 AND2_3623(.VSS(VSS),.VDD(VDD),.Y(g30001),.A(g29897),.B(g8449));
  AND2 AND2_3624(.VSS(VSS),.VDD(VDD),.Y(g30002),.A(g29905),.B(g8455));
  AND2 AND2_3625(.VSS(VSS),.VDD(VDD),.Y(g30003),.A(g29901),.B(g8469));
  AND2 AND2_3626(.VSS(VSS),.VDD(VDD),.Y(g30004),.A(g29926),.B(g22295));
  AND2 AND2_3627(.VSS(VSS),.VDD(VDD),.Y(g30005),.A(g29905),.B(g8478));
  AND2 AND2_3628(.VSS(VSS),.VDD(VDD),.Y(g30006),.A(g29928),.B(g22310));
  AND2 AND2_3629(.VSS(VSS),.VDD(VDD),.Y(g30007),.A(g29905),.B(g8494));
  AND2 AND2_3630(.VSS(VSS),.VDD(VDD),.Y(g30008),.A(g29919),.B(g22334));
  AND2 AND2_3631(.VSS(VSS),.VDD(VDD),.Y(g30009),.A(g29929),.B(g22357));
  AND2 AND2_3632(.VSS(VSS),.VDD(VDD),.Y(g30077),.A(g29823),.B(g10963));
  AND2 AND2_3633(.VSS(VSS),.VDD(VDD),.Y(g30079),.A(g29823),.B(g10988));
  AND2 AND2_3634(.VSS(VSS),.VDD(VDD),.Y(g30080),.A(g29829),.B(g10996));
  AND2 AND2_3635(.VSS(VSS),.VDD(VDD),.Y(g30081),.A(g29823),.B(g11022));
  AND2 AND2_3636(.VSS(VSS),.VDD(VDD),.Y(g30082),.A(g29829),.B(g11036));
  AND2 AND2_3637(.VSS(VSS),.VDD(VDD),.Y(g30083),.A(g29835),.B(g11048));
  AND2 AND2_3638(.VSS(VSS),.VDD(VDD),.Y(g30085),.A(g29829),.B(g11092));
  AND2 AND2_3639(.VSS(VSS),.VDD(VDD),.Y(g30086),.A(g29835),.B(g11108));
  AND2 AND2_3640(.VSS(VSS),.VDD(VDD),.Y(g30087),.A(g29840),.B(g11120));
  AND2 AND2_3641(.VSS(VSS),.VDD(VDD),.Y(g30088),.A(g29844),.B(g11138));
  AND2 AND2_3642(.VSS(VSS),.VDD(VDD),.Y(g30089),.A(g29835),.B(g11160));
  AND2 AND2_3643(.VSS(VSS),.VDD(VDD),.Y(g30090),.A(g29840),.B(g11176));
  AND2 AND2_3644(.VSS(VSS),.VDD(VDD),.Y(g30091),.A(g29844),.B(g11202));
  AND2 AND2_3645(.VSS(VSS),.VDD(VDD),.Y(g30092),.A(g29849),.B(g11205));
  AND2 AND2_3646(.VSS(VSS),.VDD(VDD),.Y(g30093),.A(g29853),.B(g11222));
  AND2 AND2_3647(.VSS(VSS),.VDD(VDD),.Y(g30094),.A(g29840),.B(g11246));
  AND2 AND2_3648(.VSS(VSS),.VDD(VDD),.Y(g30095),.A(g29857),.B(g11265));
  AND2 AND2_3649(.VSS(VSS),.VDD(VDD),.Y(g30096),.A(g29844),.B(g11268));
  AND2 AND2_3650(.VSS(VSS),.VDD(VDD),.Y(g30097),.A(g29849),.B(g11271));
  AND2 AND2_3651(.VSS(VSS),.VDD(VDD),.Y(g30098),.A(g29853),.B(g11284));
  AND2 AND2_3652(.VSS(VSS),.VDD(VDD),.Y(g30099),.A(g29861),.B(g11287));
  AND2 AND2_3653(.VSS(VSS),.VDD(VDD),.Y(g30100),.A(g29865),.B(g11306));
  AND2 AND2_3654(.VSS(VSS),.VDD(VDD),.Y(g30101),.A(g29857),.B(g11341));
  AND2 AND2_3655(.VSS(VSS),.VDD(VDD),.Y(g30102),.A(g29849),.B(g11348));
  AND2 AND2_3656(.VSS(VSS),.VDD(VDD),.Y(g30103),.A(g29869),.B(g11358));
  AND2 AND2_3657(.VSS(VSS),.VDD(VDD),.Y(g30104),.A(g29853),.B(g11361));
  AND2 AND2_3658(.VSS(VSS),.VDD(VDD),.Y(g30105),.A(g29861),.B(g11364));
  AND2 AND2_3659(.VSS(VSS),.VDD(VDD),.Y(g30106),.A(g29865),.B(g11379));
  AND2 AND2_3660(.VSS(VSS),.VDD(VDD),.Y(g30107),.A(g29873),.B(g11382));
  AND2 AND2_3661(.VSS(VSS),.VDD(VDD),.Y(g30108),.A(g29877),.B(g11401));
  AND2 AND2_3662(.VSS(VSS),.VDD(VDD),.Y(g30109),.A(g29857),.B(g11411));
  AND2 AND2_3663(.VSS(VSS),.VDD(VDD),.Y(g30110),.A(g29881),.B(g11417));
  AND2 AND2_3664(.VSS(VSS),.VDD(VDD),.Y(g30111),.A(g29869),.B(g11425));
  AND2 AND2_3665(.VSS(VSS),.VDD(VDD),.Y(g30112),.A(g29861),.B(g11432));
  AND2 AND2_3666(.VSS(VSS),.VDD(VDD),.Y(g30113),.A(g29885),.B(g11444));
  AND2 AND2_3667(.VSS(VSS),.VDD(VDD),.Y(g30114),.A(g29865),.B(g11447));
  AND2 AND2_3668(.VSS(VSS),.VDD(VDD),.Y(g30115),.A(g29873),.B(g11450));
  AND2 AND2_3669(.VSS(VSS),.VDD(VDD),.Y(g30116),.A(g29921),.B(g22236));
  AND2 AND2_3670(.VSS(VSS),.VDD(VDD),.Y(g30117),.A(g29877),.B(g11465));
  AND2 AND2_3671(.VSS(VSS),.VDD(VDD),.Y(g30118),.A(g29889),.B(g11468));
  AND2 AND2_3672(.VSS(VSS),.VDD(VDD),.Y(g30123),.A(g30070),.B(g20641));
  AND2 AND2_3673(.VSS(VSS),.VDD(VDD),.Y(g30127),.A(g30065),.B(g20719));
  AND2 AND2_3674(.VSS(VSS),.VDD(VDD),.Y(g30128),.A(g30062),.B(g20722));
  AND2 AND2_3675(.VSS(VSS),.VDD(VDD),.Y(g30129),.A(g30071),.B(g20725));
  AND2 AND2_3676(.VSS(VSS),.VDD(VDD),.Y(g30131),.A(g30059),.B(g20749));
  AND2 AND2_3677(.VSS(VSS),.VDD(VDD),.Y(g30132),.A(g30068),.B(g20776));
  AND2 AND2_3678(.VSS(VSS),.VDD(VDD),.Y(g30133),.A(g30067),.B(g20799));
  AND2 AND2_3679(.VSS(VSS),.VDD(VDD),.Y(g30138),.A(g30069),.B(g20816));
  AND2 AND2_3680(.VSS(VSS),.VDD(VDD),.Y(g30216),.A(g30036),.B(g8921));
  AND2 AND2_3681(.VSS(VSS),.VDD(VDD),.Y(g30217),.A(g30036),.B(g8955));
  AND2 AND2_3682(.VSS(VSS),.VDD(VDD),.Y(g30218),.A(g30040),.B(g8961));
  AND2 AND2_3683(.VSS(VSS),.VDD(VDD),.Y(g30219),.A(g30036),.B(g8980));
  AND2 AND2_3684(.VSS(VSS),.VDD(VDD),.Y(g30220),.A(g30040),.B(g8987));
  AND2 AND2_3685(.VSS(VSS),.VDD(VDD),.Y(g30221),.A(g30044),.B(g8993));
  AND2 AND2_3686(.VSS(VSS),.VDD(VDD),.Y(g30222),.A(g30040),.B(g9010));
  AND2 AND2_3687(.VSS(VSS),.VDD(VDD),.Y(g30223),.A(g30044),.B(g9016));
  AND2 AND2_3688(.VSS(VSS),.VDD(VDD),.Y(g30224),.A(g30048),.B(g9022));
  AND2 AND2_3689(.VSS(VSS),.VDD(VDD),.Y(g30225),.A(g30044),.B(g9035));
  AND2 AND2_3690(.VSS(VSS),.VDD(VDD),.Y(g30226),.A(g30048),.B(g9041));
  AND2 AND2_3691(.VSS(VSS),.VDD(VDD),.Y(g30227),.A(g30048),.B(g9058));
  AND2 AND2_3692(.VSS(VSS),.VDD(VDD),.Y(g30327),.A(g30187),.B(g8321));
  AND2 AND2_3693(.VSS(VSS),.VDD(VDD),.Y(g30330),.A(g30195),.B(g8333));
  AND2 AND2_3694(.VSS(VSS),.VDD(VDD),.Y(g30333),.A(g30191),.B(g8341));
  AND2 AND2_3695(.VSS(VSS),.VDD(VDD),.Y(g30334),.A(g30203),.B(g8347));
  AND2 AND2_3696(.VSS(VSS),.VDD(VDD),.Y(g30337),.A(g30199),.B(g8354));
  AND2 AND2_3697(.VSS(VSS),.VDD(VDD),.Y(g30340),.A(g30207),.B(g8372));
  AND2 AND2_3698(.VSS(VSS),.VDD(VDD),.Y(g30345),.A(g30195),.B(g8388));
  AND2 AND2_3699(.VSS(VSS),.VDD(VDD),.Y(g30348),.A(g30203),.B(g8400));
  AND2 AND2_3700(.VSS(VSS),.VDD(VDD),.Y(g30351),.A(g30199),.B(g8408));
  AND2 AND2_3701(.VSS(VSS),.VDD(VDD),.Y(g30352),.A(g30211),.B(g8414));
  AND2 AND2_3702(.VSS(VSS),.VDD(VDD),.Y(g30355),.A(g30207),.B(g8421));
  AND2 AND2_3703(.VSS(VSS),.VDD(VDD),.Y(g30361),.A(g30203),.B(g8440));
  AND2 AND2_3704(.VSS(VSS),.VDD(VDD),.Y(g30364),.A(g30211),.B(g8452));
  AND2 AND2_3705(.VSS(VSS),.VDD(VDD),.Y(g30367),.A(g30207),.B(g8460));
  AND2 AND2_3706(.VSS(VSS),.VDD(VDD),.Y(g30372),.A(g8594),.B(g30228));
  AND2 AND2_3707(.VSS(VSS),.VDD(VDD),.Y(g30374),.A(g30211),.B(g8475));
  AND2 AND2_3708(.VSS(VSS),.VDD(VDD),.Y(g30387),.A(g30229),.B(g8888));
  AND2 AND2_3709(.VSS(VSS),.VDD(VDD),.Y(g30388),.A(g30229),.B(g8918));
  AND2 AND2_3710(.VSS(VSS),.VDD(VDD),.Y(g30389),.A(g30233),.B(g8928));
  AND2 AND2_3711(.VSS(VSS),.VDD(VDD),.Y(g30390),.A(g30229),.B(g8952));
  AND2 AND2_3712(.VSS(VSS),.VDD(VDD),.Y(g30391),.A(g30233),.B(g8958));
  AND2 AND2_3713(.VSS(VSS),.VDD(VDD),.Y(g30392),.A(g30237),.B(g8968));
  AND2 AND2_3714(.VSS(VSS),.VDD(VDD),.Y(g30393),.A(g30233),.B(g8984));
  AND2 AND2_3715(.VSS(VSS),.VDD(VDD),.Y(g30394),.A(g30237),.B(g8990));
  AND2 AND2_3716(.VSS(VSS),.VDD(VDD),.Y(g30395),.A(g30241),.B(g9000));
  AND2 AND2_3717(.VSS(VSS),.VDD(VDD),.Y(g30396),.A(g30237),.B(g9013));
  AND2 AND2_3718(.VSS(VSS),.VDD(VDD),.Y(g30397),.A(g30241),.B(g9019));
  AND2 AND2_3719(.VSS(VSS),.VDD(VDD),.Y(g30398),.A(g30241),.B(g9038));
  AND2 AND2_3720(.VSS(VSS),.VDD(VDD),.Y(g30407),.A(g30134),.B(g10991));
  AND2 AND2_3721(.VSS(VSS),.VDD(VDD),.Y(g30409),.A(g30134),.B(g11025));
  AND2 AND2_3722(.VSS(VSS),.VDD(VDD),.Y(g30410),.A(g30139),.B(g11028));
  AND2 AND2_3723(.VSS(VSS),.VDD(VDD),.Y(g30411),.A(g30143),.B(g11039));
  AND2 AND2_3724(.VSS(VSS),.VDD(VDD),.Y(g30436),.A(g30134),.B(g11079));
  AND2 AND2_3725(.VSS(VSS),.VDD(VDD),.Y(g30437),.A(g30139),.B(g11082));
  AND2 AND2_3726(.VSS(VSS),.VDD(VDD),.Y(g30438),.A(g30147),.B(g11085));
  AND2 AND2_3727(.VSS(VSS),.VDD(VDD),.Y(g30440),.A(g30143),.B(g11095));
  AND2 AND2_3728(.VSS(VSS),.VDD(VDD),.Y(g30441),.A(g30151),.B(g11098));
  AND2 AND2_3729(.VSS(VSS),.VDD(VDD),.Y(g30442),.A(g30155),.B(g11111));
  AND2 AND2_3730(.VSS(VSS),.VDD(VDD),.Y(g30444),.A(g30139),.B(g11132));
  AND2 AND2_3731(.VSS(VSS),.VDD(VDD),.Y(g30445),.A(g30147),.B(g11135));
  AND2 AND2_3732(.VSS(VSS),.VDD(VDD),.Y(g30447),.A(g30143),.B(g11145));
  AND2 AND2_3733(.VSS(VSS),.VDD(VDD),.Y(g30448),.A(g30151),.B(g11148));
  AND2 AND2_3734(.VSS(VSS),.VDD(VDD),.Y(g30449),.A(g30159),.B(g11151));
  AND2 AND2_3735(.VSS(VSS),.VDD(VDD),.Y(g30451),.A(g30155),.B(g11163));
  AND2 AND2_3736(.VSS(VSS),.VDD(VDD),.Y(g30452),.A(g30163),.B(g11166));
  AND2 AND2_3737(.VSS(VSS),.VDD(VDD),.Y(g30453),.A(g30167),.B(g11179));
  AND2 AND2_3738(.VSS(VSS),.VDD(VDD),.Y(g30454),.A(g30147),.B(g11199));
  AND2 AND2_3739(.VSS(VSS),.VDD(VDD),.Y(g30457),.A(g30151),.B(g11216));
  AND2 AND2_3740(.VSS(VSS),.VDD(VDD),.Y(g30458),.A(g30159),.B(g11219));
  AND2 AND2_3741(.VSS(VSS),.VDD(VDD),.Y(g30460),.A(g30155),.B(g11231));
  AND2 AND2_3742(.VSS(VSS),.VDD(VDD),.Y(g30461),.A(g30163),.B(g11234));
  AND2 AND2_3743(.VSS(VSS),.VDD(VDD),.Y(g30462),.A(g30171),.B(g11237));
  AND2 AND2_3744(.VSS(VSS),.VDD(VDD),.Y(g30464),.A(g30167),.B(g11249));
  AND2 AND2_3745(.VSS(VSS),.VDD(VDD),.Y(g30465),.A(g30175),.B(g11252));
  AND2 AND2_3746(.VSS(VSS),.VDD(VDD),.Y(g30467),.A(g30179),.B(g11274));
  AND2 AND2_3747(.VSS(VSS),.VDD(VDD),.Y(g30469),.A(g30159),.B(g11281));
  AND2 AND2_3748(.VSS(VSS),.VDD(VDD),.Y(g30472),.A(g30163),.B(g11300));
  AND2 AND2_3749(.VSS(VSS),.VDD(VDD),.Y(g30473),.A(g30171),.B(g11303));
  AND2 AND2_3750(.VSS(VSS),.VDD(VDD),.Y(g30475),.A(g30167),.B(g11315));
  AND2 AND2_3751(.VSS(VSS),.VDD(VDD),.Y(g30476),.A(g30175),.B(g11318));
  AND2 AND2_3752(.VSS(VSS),.VDD(VDD),.Y(g30477),.A(g30183),.B(g11321));
  AND2 AND2_3753(.VSS(VSS),.VDD(VDD),.Y(g30478),.A(g30187),.B(g11344));
  AND2 AND2_3754(.VSS(VSS),.VDD(VDD),.Y(g30481),.A(g30179),.B(g11351));
  AND2 AND2_3755(.VSS(VSS),.VDD(VDD),.Y(g30484),.A(g30191),.B(g11367));
  AND2 AND2_3756(.VSS(VSS),.VDD(VDD),.Y(g30486),.A(g30171),.B(g11376));
  AND2 AND2_3757(.VSS(VSS),.VDD(VDD),.Y(g30489),.A(g30175),.B(g11395));
  AND2 AND2_3758(.VSS(VSS),.VDD(VDD),.Y(g30490),.A(g30183),.B(g11398));
  AND2 AND2_3759(.VSS(VSS),.VDD(VDD),.Y(g30492),.A(g30187),.B(g11414));
  AND2 AND2_3760(.VSS(VSS),.VDD(VDD),.Y(g30495),.A(g30179),.B(g11422));
  AND2 AND2_3761(.VSS(VSS),.VDD(VDD),.Y(g30496),.A(g30195),.B(g11428));
  AND2 AND2_3762(.VSS(VSS),.VDD(VDD),.Y(g30499),.A(g30191),.B(g11435));
  AND2 AND2_3763(.VSS(VSS),.VDD(VDD),.Y(g30502),.A(g30199),.B(g11453));
  AND2 AND2_3764(.VSS(VSS),.VDD(VDD),.Y(g30504),.A(g30183),.B(g11462));
  AND2 AND2_3765(.VSS(VSS),.VDD(VDD),.Y(g30696),.A(g30383),.B(g10943));
  AND2 AND2_3766(.VSS(VSS),.VDD(VDD),.Y(g30697),.A(g30383),.B(g11011));
  AND2 AND2_3767(.VSS(VSS),.VDD(VDD),.Y(g30698),.A(g30383),.B(g11126));
  AND2 AND2_3768(.VSS(VSS),.VDD(VDD),.Y(g30728),.A(g30605),.B(g22252));
  AND2 AND2_3769(.VSS(VSS),.VDD(VDD),.Y(g30735),.A(g30629),.B(g22268));
  AND2 AND2_3770(.VSS(VSS),.VDD(VDD),.Y(g30736),.A(g30584),.B(g20669));
  AND2 AND2_3771(.VSS(VSS),.VDD(VDD),.Y(g30743),.A(g30610),.B(g22283));
  AND2 AND2_3772(.VSS(VSS),.VDD(VDD),.Y(g30744),.A(g30609),.B(g20697));
  AND2 AND2_3773(.VSS(VSS),.VDD(VDD),.Y(g30750),.A(g30593),.B(g20729));
  AND2 AND2_3774(.VSS(VSS),.VDD(VDD),.Y(g30754),.A(g30614),.B(g22313));
  AND2 AND2_3775(.VSS(VSS),.VDD(VDD),.Y(g30755),.A(g30632),.B(g22314));
  AND2 AND2_3776(.VSS(VSS),.VDD(VDD),.Y(g30757),.A(g30601),.B(g20780));
  AND2 AND2_3777(.VSS(VSS),.VDD(VDD),.Y(g30758),.A(g30613),.B(g20783));
  AND2 AND2_3778(.VSS(VSS),.VDD(VDD),.Y(g30759),.A(g30588),.B(g22360));
  AND2 AND2_3779(.VSS(VSS),.VDD(VDD),.Y(g30760),.A(g30622),.B(g22379));
  AND2 AND2_3780(.VSS(VSS),.VDD(VDD),.Y(g30761),.A(g30621),.B(g20822));
  AND2 AND2_3781(.VSS(VSS),.VDD(VDD),.Y(g30762),.A(g30608),.B(g20830));
  AND2 AND2_3782(.VSS(VSS),.VDD(VDD),.Y(g30763),.A(g30597),.B(g22386));
  AND2 AND2_3783(.VSS(VSS),.VDD(VDD),.Y(g30764),.A(g30628),.B(g20837));
  AND3 AND3_257(.VSS(VSS),.VDD(VDD),.Y(g30766),.A(g30617),.B(g19457),.C(g19431));
  AND2 AND2_3784(.VSS(VSS),.VDD(VDD),.Y(g30916),.A(g30785),.B(g22251));
  AND2 AND2_3785(.VSS(VSS),.VDD(VDD),.Y(g30917),.A(g12446),.B(g30766));
  AND2 AND2_3786(.VSS(VSS),.VDD(VDD),.Y(g30918),.A(g30780),.B(g22296));
  AND2 AND2_3787(.VSS(VSS),.VDD(VDD),.Y(g30919),.A(g30786),.B(g22297));
  AND2 AND2_3788(.VSS(VSS),.VDD(VDD),.Y(g30920),.A(g30787),.B(g22298));
  AND2 AND2_3789(.VSS(VSS),.VDD(VDD),.Y(g30921),.A(g10773),.B(g30791));
  AND2 AND2_3790(.VSS(VSS),.VDD(VDD),.Y(g30922),.A(g30788),.B(g22315));
  AND2 AND2_3791(.VSS(VSS),.VDD(VDD),.Y(g30923),.A(g30789),.B(g22338));
  AND2 AND2_3792(.VSS(VSS),.VDD(VDD),.Y(g30924),.A(g30783),.B(g22359));
  AND2 AND2_3793(.VSS(VSS),.VDD(VDD),.Y(g30925),.A(g30790),.B(g22380));
  AND2 AND2_3794(.VSS(VSS),.VDD(VDD),.Y(g30944),.A(g30935),.B(g20666));
  AND2 AND2_3795(.VSS(VSS),.VDD(VDD),.Y(g30945),.A(g30931),.B(g20754));
  AND2 AND2_3796(.VSS(VSS),.VDD(VDD),.Y(g30946),.A(g30930),.B(g20757));
  AND2 AND2_3797(.VSS(VSS),.VDD(VDD),.Y(g30947),.A(g30936),.B(g20760));
  AND2 AND2_3798(.VSS(VSS),.VDD(VDD),.Y(g30948),.A(g30929),.B(g20786));
  AND2 AND2_3799(.VSS(VSS),.VDD(VDD),.Y(g30949),.A(g30933),.B(g20806));
  AND2 AND2_3800(.VSS(VSS),.VDD(VDD),.Y(g30950),.A(g30932),.B(g20819));
  AND2 AND2_3801(.VSS(VSS),.VDD(VDD),.Y(g30951),.A(g30934),.B(g20833));
  AND2 AND2_3802(.VSS(VSS),.VDD(VDD),.Y(g30953),.A(g8605),.B(g30952));
//
  OR2 OR2_0(.VSS(VSS),.VDD(VDD),.Y(g9144),.A(g2986),.B(g5389));
  OR2 OR2_1(.VSS(VSS),.VDD(VDD),.Y(g10778),.A(g2929),.B(g8022));
  OR2 OR2_2(.VSS(VSS),.VDD(VDD),.Y(g12377),.A(g7553),.B(g11059));
  OR2 OR2_3(.VSS(VSS),.VDD(VDD),.Y(g12407),.A(g7573),.B(g10779));
  OR2 OR2_4(.VSS(VSS),.VDD(VDD),.Y(g12886),.A(g9534),.B(g3398));
  OR2 OR2_5(.VSS(VSS),.VDD(VDD),.Y(g12926),.A(g9676),.B(g3554));
  OR2 OR2_6(.VSS(VSS),.VDD(VDD),.Y(g12955),.A(g9822),.B(g3710));
  OR2 OR2_7(.VSS(VSS),.VDD(VDD),.Y(g12984),.A(g9968),.B(g3866));
  OR2 OR2_8(.VSS(VSS),.VDD(VDD),.Y(g16539),.A(g15880),.B(g14657));
  OR2 OR2_9(.VSS(VSS),.VDD(VDD),.Y(g16571),.A(g15913),.B(g14691));
  OR2 OR2_10(.VSS(VSS),.VDD(VDD),.Y(g16595),.A(g15942),.B(g14725));
  OR2 OR2_11(.VSS(VSS),.VDD(VDD),.Y(g16615),.A(g15971),.B(g14753));
  OR2 OR2_12(.VSS(VSS),.VDD(VDD),.Y(g17973),.A(g11623),.B(g15659));
  OR2 OR2_13(.VSS(VSS),.VDD(VDD),.Y(g19181),.A(g17729),.B(g17979));
  OR2 OR2_14(.VSS(VSS),.VDD(VDD),.Y(g19186),.A(g18419),.B(g17887));
  OR2 OR2_15(.VSS(VSS),.VDD(VDD),.Y(g19187),.A(g18419),.B(g17729));
  OR2 OR2_16(.VSS(VSS),.VDD(VDD),.Y(g19188),.A(g17830),.B(g18096));
  OR2 OR2_17(.VSS(VSS),.VDD(VDD),.Y(g19191),.A(g17807),.B(g17887));
  OR2 OR2_18(.VSS(VSS),.VDD(VDD),.Y(g19192),.A(g18183),.B(g18270));
  OR2 OR2_19(.VSS(VSS),.VDD(VDD),.Y(g19193),.A(g18492),.B(g17998));
  OR2 OR2_20(.VSS(VSS),.VDD(VDD),.Y(g19194),.A(g18492),.B(g17830));
  OR2 OR2_21(.VSS(VSS),.VDD(VDD),.Y(g19195),.A(g17942),.B(g18212));
  OR2 OR2_22(.VSS(VSS),.VDD(VDD),.Y(g19200),.A(g18346),.B(g18424));
  OR2 OR2_23(.VSS(VSS),.VDD(VDD),.Y(g19201),.A(g18183),.B(g18424));
  OR2 OR2_24(.VSS(VSS),.VDD(VDD),.Y(g19202),.A(g17919),.B(g17998));
  OR2 OR2_25(.VSS(VSS),.VDD(VDD),.Y(g19203),.A(g18290),.B(g18363));
  OR2 OR2_26(.VSS(VSS),.VDD(VDD),.Y(g19204),.A(g18556),.B(g18115));
  OR2 OR2_27(.VSS(VSS),.VDD(VDD),.Y(g19205),.A(g18556),.B(g17942));
  OR2 OR2_28(.VSS(VSS),.VDD(VDD),.Y(g19206),.A(g18053),.B(g18319));
  OR2 OR2_29(.VSS(VSS),.VDD(VDD),.Y(g19209),.A(g18079),.B(g18346));
  OR2 OR2_30(.VSS(VSS),.VDD(VDD),.Y(g19210),.A(g18079),.B(g18183));
  OR2 OR2_31(.VSS(VSS),.VDD(VDD),.Y(g19211),.A(g18441),.B(g18497));
  OR2 OR2_32(.VSS(VSS),.VDD(VDD),.Y(g19212),.A(g18290),.B(g18497));
  OR2 OR2_33(.VSS(VSS),.VDD(VDD),.Y(g19213),.A(g18030),.B(g18115));
  OR2 OR2_34(.VSS(VSS),.VDD(VDD),.Y(g19214),.A(g18383),.B(g18458));
  OR2 OR2_35(.VSS(VSS),.VDD(VDD),.Y(g19215),.A(g18606),.B(g18231));
  OR2 OR2_36(.VSS(VSS),.VDD(VDD),.Y(g19216),.A(g18606),.B(g18053));
  OR2 OR2_37(.VSS(VSS),.VDD(VDD),.Y(g19221),.A(g18270),.B(g18346));
  OR2 OR2_38(.VSS(VSS),.VDD(VDD),.Y(g19222),.A(g18195),.B(g18441));
  OR2 OR2_39(.VSS(VSS),.VDD(VDD),.Y(g19223),.A(g18195),.B(g18290));
  OR2 OR2_40(.VSS(VSS),.VDD(VDD),.Y(g19224),.A(g18514),.B(g18561));
  OR2 OR2_41(.VSS(VSS),.VDD(VDD),.Y(g19225),.A(g18383),.B(g18561));
  OR2 OR2_42(.VSS(VSS),.VDD(VDD),.Y(g19226),.A(g18147),.B(g18231));
  OR2 OR2_43(.VSS(VSS),.VDD(VDD),.Y(g19227),.A(g18478),.B(g18531));
  OR3 OR3_0(.VSS(VSS),.VDD(VDD),.Y(I25477),.A(g17024),.B(g17000),.C(g16992));
  OR3 OR3_1(.VSS(VSS),.VDD(VDD),.Y(g19230),.A(g16985),.B(g16965),.C(I25477));
  OR2 OR2_44(.VSS(VSS),.VDD(VDD),.Y(g19231),.A(g18363),.B(g18441));
  OR2 OR2_45(.VSS(VSS),.VDD(VDD),.Y(g19232),.A(g18302),.B(g18514));
  OR2 OR2_46(.VSS(VSS),.VDD(VDD),.Y(g19233),.A(g18302),.B(g18383));
  OR2 OR2_47(.VSS(VSS),.VDD(VDD),.Y(g19234),.A(g18578),.B(g18611));
  OR2 OR2_48(.VSS(VSS),.VDD(VDD),.Y(g19235),.A(g18478),.B(g18611));
  OR3 OR3_2(.VSS(VSS),.VDD(VDD),.Y(I25495),.A(g17158),.B(g17137),.C(g17115));
  OR3 OR3_3(.VSS(VSS),.VDD(VDD),.Y(g19240),.A(g17083),.B(g17050),.C(I25495));
  OR2 OR2_49(.VSS(VSS),.VDD(VDD),.Y(g19242),.A(g14244),.B(g16501));
  OR3 OR3_4(.VSS(VSS),.VDD(VDD),.Y(I25500),.A(g17058),.B(g17030),.C(g17016));
  OR3 OR3_5(.VSS(VSS),.VDD(VDD),.Y(g19243),.A(g16995),.B(g16986),.C(I25500));
  OR2 OR2_50(.VSS(VSS),.VDD(VDD),.Y(g19244),.A(g18458),.B(g18514));
  OR2 OR2_51(.VSS(VSS),.VDD(VDD),.Y(g19245),.A(g18395),.B(g18578));
  OR2 OR2_52(.VSS(VSS),.VDD(VDD),.Y(g19246),.A(g18395),.B(g18478));
  OR2 OR2_53(.VSS(VSS),.VDD(VDD),.Y(g19250),.A(g17729),.B(g17807));
  OR3 OR3_6(.VSS(VSS),.VDD(VDD),.Y(I25516),.A(g17173),.B(g17160),.C(g17142));
  OR3 OR3_7(.VSS(VSS),.VDD(VDD),.Y(g19253),.A(g17121),.B(g17085),.C(I25516));
  OR2 OR2_54(.VSS(VSS),.VDD(VDD),.Y(g19255),.A(g14366),.B(g16523));
  OR3 OR3_8(.VSS(VSS),.VDD(VDD),.Y(I25521),.A(g17093),.B(g17064),.C(g17046));
  OR3 OR3_9(.VSS(VSS),.VDD(VDD),.Y(g19256),.A(g17019),.B(g16996),.C(I25521));
  OR2 OR2_55(.VSS(VSS),.VDD(VDD),.Y(g19257),.A(g18531),.B(g18578));
  OR2 OR2_56(.VSS(VSS),.VDD(VDD),.Y(g19263),.A(g17887),.B(g17979));
  OR2 OR2_57(.VSS(VSS),.VDD(VDD),.Y(g19264),.A(g17830),.B(g17919));
  OR3 OR3_10(.VSS(VSS),.VDD(VDD),.Y(I25549),.A(g17190),.B(g17175),.C(g17165));
  OR3 OR3_11(.VSS(VSS),.VDD(VDD),.Y(g19266),.A(g17148),.B(g17123),.C(I25549));
  OR2 OR2_58(.VSS(VSS),.VDD(VDD),.Y(g19268),.A(g14478),.B(g16554));
  OR3 OR3_12(.VSS(VSS),.VDD(VDD),.Y(I25554),.A(g17131),.B(g17099),.C(g17080));
  OR3 OR3_13(.VSS(VSS),.VDD(VDD),.Y(g19269),.A(g17049),.B(g17020),.C(I25554));
  OR3 OR3_14(.VSS(VSS),.VDD(VDD),.Y(g19275),.A(g16867),.B(g16515),.C(g19001));
  OR2 OR2_59(.VSS(VSS),.VDD(VDD),.Y(g19278),.A(g17998),.B(g18096));
  OR2 OR2_60(.VSS(VSS),.VDD(VDD),.Y(g19279),.A(g17942),.B(g18030));
  OR3 OR3_15(.VSS(VSS),.VDD(VDD),.Y(I25588),.A(g17201),.B(g17192),.C(g17180));
  OR3 OR3_16(.VSS(VSS),.VDD(VDD),.Y(g19281),.A(g17171),.B(g17150),.C(I25588));
  OR2 OR2_61(.VSS(VSS),.VDD(VDD),.Y(g19283),.A(g14565),.B(g16586));
  OR3 OR3_17(.VSS(VSS),.VDD(VDD),.Y(g19294),.A(g16895),.B(g16546),.C(g16507));
  OR2 OR2_62(.VSS(VSS),.VDD(VDD),.Y(g19297),.A(g18115),.B(g18212));
  OR2 OR2_63(.VSS(VSS),.VDD(VDD),.Y(g19298),.A(g18053),.B(g18147));
  OR3 OR3_18(.VSS(VSS),.VDD(VDD),.Y(g19312),.A(g16924),.B(g16578),.C(g16529));
  OR2 OR2_64(.VSS(VSS),.VDD(VDD),.Y(g19315),.A(g18231),.B(g18319));
  OR3 OR3_19(.VSS(VSS),.VDD(VDD),.Y(g19333),.A(g16954),.B(g16602),.C(g16560));
  OR2 OR2_65(.VSS(VSS),.VDD(VDD),.Y(g19450),.A(g14837),.B(g16682));
  OR2 OR2_66(.VSS(VSS),.VDD(VDD),.Y(g19477),.A(g14910),.B(g16708));
  OR2 OR2_67(.VSS(VSS),.VDD(VDD),.Y(g19500),.A(g14991),.B(g16739));
  OR3 OR3_20(.VSS(VSS),.VDD(VDD),.Y(g19503),.A(g16884),.B(g16697),.C(g16665));
  OR2 OR2_68(.VSS(VSS),.VDD(VDD),.Y(g19521),.A(g15080),.B(g16781));
  OR3 OR3_21(.VSS(VSS),.VDD(VDD),.Y(g19522),.A(g16913),.B(g16728),.C(g16686));
  OR3 OR3_22(.VSS(VSS),.VDD(VDD),.Y(g19532),.A(g16943),.B(g16770),.C(g16712));
  OR3 OR3_23(.VSS(VSS),.VDD(VDD),.Y(g19542),.A(g16974),.B(g16797),.C(g16743));
  OR3 OR3_24(.VSS(VSS),.VDD(VDD),.Y(I26429),.A(g17979),.B(g17887),.C(g17807));
  OR3 OR3_25(.VSS(VSS),.VDD(VDD),.Y(g19981),.A(g17729),.B(g18419),.C(I26429));
  OR3 OR3_26(.VSS(VSS),.VDD(VDD),.Y(I26455),.A(g18424),.B(g18346),.C(g18270));
  OR3 OR3_27(.VSS(VSS),.VDD(VDD),.Y(g20015),.A(g18183),.B(g18079),.C(I26455));
  OR3 OR3_28(.VSS(VSS),.VDD(VDD),.Y(I26461),.A(g18096),.B(g17998),.C(g17919));
  OR3 OR3_29(.VSS(VSS),.VDD(VDD),.Y(g20019),.A(g17830),.B(g18492),.C(I26461));
  OR3 OR3_30(.VSS(VSS),.VDD(VDD),.Y(I26491),.A(g18497),.B(g18441),.C(g18363));
  OR3 OR3_31(.VSS(VSS),.VDD(VDD),.Y(g20057),.A(g18290),.B(g18195),.C(I26491));
  OR3 OR3_32(.VSS(VSS),.VDD(VDD),.Y(I26497),.A(g18212),.B(g18115),.C(g18030));
  OR3 OR3_33(.VSS(VSS),.VDD(VDD),.Y(g20061),.A(g17942),.B(g18556),.C(I26497));
  OR3 OR3_34(.VSS(VSS),.VDD(VDD),.Y(I26532),.A(g18561),.B(g18514),.C(g18458));
  OR3 OR3_35(.VSS(VSS),.VDD(VDD),.Y(g20098),.A(g18383),.B(g18302),.C(I26532));
  OR3 OR3_36(.VSS(VSS),.VDD(VDD),.Y(I26538),.A(g18319),.B(g18231),.C(g18147));
  OR3 OR3_37(.VSS(VSS),.VDD(VDD),.Y(g20102),.A(g18053),.B(g18606),.C(I26538));
  OR3 OR3_38(.VSS(VSS),.VDD(VDD),.Y(I26571),.A(g18611),.B(g18578),.C(g18531));
  OR3 OR3_39(.VSS(VSS),.VDD(VDD),.Y(g20123),.A(g18478),.B(g18395),.C(I26571));
  OR3 OR3_40(.VSS(VSS),.VDD(VDD),.Y(g21120),.A(g19484),.B(g16515),.C(g14071));
  OR3 OR3_41(.VSS(VSS),.VDD(VDD),.Y(g21139),.A(g19505),.B(g16546),.C(g14186));
  OR3 OR3_42(.VSS(VSS),.VDD(VDD),.Y(g21159),.A(g19524),.B(g16578),.C(g14301));
  OR3 OR3_43(.VSS(VSS),.VDD(VDD),.Y(g21179),.A(g19534),.B(g16602),.C(g14423));
  OR3 OR3_44(.VSS(VSS),.VDD(VDD),.Y(g21244),.A(g19578),.B(g16697),.C(g14776));
  OR3 OR3_45(.VSS(VSS),.VDD(VDD),.Y(g21253),.A(g19608),.B(g16728),.C(g14811));
  OR3 OR3_46(.VSS(VSS),.VDD(VDD),.Y(g21261),.A(g19641),.B(g16770),.C(g14863));
  OR3 OR3_47(.VSS(VSS),.VDD(VDD),.Y(g21269),.A(g19681),.B(g16797),.C(g14936));
  OR3 OR3_48(.VSS(VSS),.VDD(VDD),.Y(g21501),.A(g20522),.B(g16867),.C(g14071));
  OR3 OR3_49(.VSS(VSS),.VDD(VDD),.Y(g21536),.A(g20522),.B(g19484),.C(g19001));
  OR3 OR3_50(.VSS(VSS),.VDD(VDD),.Y(g21540),.A(g20542),.B(g16895),.C(g14186));
  OR3 OR3_51(.VSS(VSS),.VDD(VDD),.Y(g21572),.A(g20542),.B(g19505),.C(g16507));
  OR3 OR3_52(.VSS(VSS),.VDD(VDD),.Y(g21576),.A(g19067),.B(g16924),.C(g14301));
  OR3 OR3_53(.VSS(VSS),.VDD(VDD),.Y(g21605),.A(g19067),.B(g19524),.C(g16529));
  OR3 OR3_54(.VSS(VSS),.VDD(VDD),.Y(g21609),.A(g19084),.B(g16954),.C(g14423));
  OR3 OR3_55(.VSS(VSS),.VDD(VDD),.Y(g21634),.A(g19084),.B(g19534),.C(g16560));
  OR3 OR3_56(.VSS(VSS),.VDD(VDD),.Y(g21774),.A(g19121),.B(g16884),.C(g14776));
  OR3 OR3_57(.VSS(VSS),.VDD(VDD),.Y(g21787),.A(g19121),.B(g19578),.C(g16665));
  OR3 OR3_58(.VSS(VSS),.VDD(VDD),.Y(I28305),.A(g20197),.B(g20177),.C(g20145));
  OR3 OR3_59(.VSS(VSS),.VDD(VDD),.Y(g21788),.A(g20117),.B(g20094),.C(I28305));
  OR3 OR3_60(.VSS(VSS),.VDD(VDD),.Y(g21789),.A(g19128),.B(g16913),.C(g14811));
  OR3 OR3_61(.VSS(VSS),.VDD(VDD),.Y(I28318),.A(g19092),.B(g19088),.C(g19079));
  OR4 OR4_0(.VSS(VSS),.VDD(VDD),.Y(g21799),.A(g16505),.B(g20538),.C(g18994),.D(I28318));
  OR4 OR4_1(.VSS(VSS),.VDD(VDD),.Y(g21800),.A(g18665),.B(g20270),.C(g20248),.D(g18647));
  OR3 OR3_62(.VSS(VSS),.VDD(VDD),.Y(g21801),.A(g19128),.B(g19608),.C(g16686));
  OR3 OR3_63(.VSS(VSS),.VDD(VDD),.Y(I28323),.A(g20227),.B(g20211),.C(g20183));
  OR3 OR3_64(.VSS(VSS),.VDD(VDD),.Y(g21802),.A(g20147),.B(g20119),.C(I28323));
  OR3 OR3_65(.VSS(VSS),.VDD(VDD),.Y(g21803),.A(g19135),.B(g16943),.C(g14863));
  OR4 OR4_2(.VSS(VSS),.VDD(VDD),.Y(g21806),.A(g20116),.B(g20093),.C(g18547),.D(g19097));
  OR3 OR3_66(.VSS(VSS),.VDD(VDD),.Y(I28330),.A(g19099),.B(g19094),.C(g19089));
  OR4 OR4_3(.VSS(VSS),.VDD(VDD),.Y(g21807),.A(g16527),.B(g19063),.C(g19007),.D(I28330));
  OR4 OR4_4(.VSS(VSS),.VDD(VDD),.Y(g21808),.A(g18688),.B(g20282),.C(g20271),.D(g18650));
  OR3 OR3_67(.VSS(VSS),.VDD(VDD),.Y(g21809),.A(g19135),.B(g19641),.C(g16712));
  OR3 OR3_68(.VSS(VSS),.VDD(VDD),.Y(I28335),.A(g20254),.B(g20241),.C(g20217));
  OR3 OR3_69(.VSS(VSS),.VDD(VDD),.Y(g21810),.A(g20185),.B(g20149),.C(I28335));
  OR3 OR3_70(.VSS(VSS),.VDD(VDD),.Y(g21811),.A(g19138),.B(g16974),.C(g14936));
  OR4 OR4_5(.VSS(VSS),.VDD(VDD),.Y(g21813),.A(g20146),.B(g20118),.C(g18597),.D(g19104));
  OR3 OR3_71(.VSS(VSS),.VDD(VDD),.Y(I28341),.A(g19106),.B(g19101),.C(g19095));
  OR4 OR4_6(.VSS(VSS),.VDD(VDD),.Y(g21814),.A(g16558),.B(g19080),.C(g16513),.D(I28341));
  OR4 OR4_7(.VSS(VSS),.VDD(VDD),.Y(g21815),.A(g18717),.B(g20293),.C(g20283),.D(g18654));
  OR3 OR3_72(.VSS(VSS),.VDD(VDD),.Y(g21816),.A(g19138),.B(g19681),.C(g16743));
  OR3 OR3_73(.VSS(VSS),.VDD(VDD),.Y(I28346),.A(g20277),.B(g20268),.C(g20247));
  OR3 OR3_74(.VSS(VSS),.VDD(VDD),.Y(g21817),.A(g20219),.B(g20187),.C(I28346));
  OR4 OR4_8(.VSS(VSS),.VDD(VDD),.Y(g21819),.A(g20184),.B(g20148),.C(g18629),.D(g19109));
  OR3 OR3_75(.VSS(VSS),.VDD(VDD),.Y(I28351),.A(g19111),.B(g19108),.C(g19102));
  OR4 OR4_9(.VSS(VSS),.VDD(VDD),.Y(g21820),.A(g16590),.B(g19090),.C(g16535),.D(I28351));
  OR4 OR4_10(.VSS(VSS),.VDD(VDD),.Y(g21821),.A(g18753),.B(g20309),.C(g20294),.D(g18668));
  OR4 OR4_11(.VSS(VSS),.VDD(VDD),.Y(g21823),.A(g20218),.B(g20186),.C(g18638),.D(g19116));
  OR3 OR3_76(.VSS(VSS),.VDD(VDD),.Y(I28365),.A(g20280),.B(g18652),.C(g18649));
  OR3 OR3_77(.VSS(VSS),.VDD(VDD),.Y(g21844),.A(g20222),.B(g18645),.C(I28365));
  OR3 OR3_78(.VSS(VSS),.VDD(VDD),.Y(I28369),.A(g20291),.B(g18666),.C(g18653));
  OR3 OR3_79(.VSS(VSS),.VDD(VDD),.Y(g21846),.A(g20249),.B(g18648),.C(I28369));
  OR3 OR3_80(.VSS(VSS),.VDD(VDD),.Y(I28374),.A(g20307),.B(g18689),.C(g18667));
  OR3 OR3_81(.VSS(VSS),.VDD(VDD),.Y(g21849),.A(g20272),.B(g18651),.C(I28374));
  OR3 OR3_82(.VSS(VSS),.VDD(VDD),.Y(I28380),.A(g20326),.B(g18718),.C(g18690));
  OR3 OR3_83(.VSS(VSS),.VDD(VDD),.Y(g21856),.A(g20284),.B(g18655),.C(I28380));
  OR2 OR2_69(.VSS(VSS),.VDD(VDD),.Y(g22175),.A(g16075),.B(g20842));
  OR2 OR2_70(.VSS(VSS),.VDD(VDD),.Y(g22190),.A(g16113),.B(g20850));
  OR2 OR2_71(.VSS(VSS),.VDD(VDD),.Y(g22199),.A(g16164),.B(g20858));
  OR2 OR2_72(.VSS(VSS),.VDD(VDD),.Y(g22205),.A(g16223),.B(g20866));
  OR4 OR4_12(.VSS(VSS),.VDD(VDD),.Y(g22811),.A(g562),.B(g559),.C(g12451),.D(g21851));
  OR3 OR3_84(.VSS(VSS),.VDD(VDD),.Y(g23052),.A(g21800),.B(g21788),.C(g21844));
  OR3 OR3_85(.VSS(VSS),.VDD(VDD),.Y(g23071),.A(g21808),.B(g21802),.C(g21846));
  OR3 OR3_86(.VSS(VSS),.VDD(VDD),.Y(g23084),.A(g21815),.B(g21810),.C(g21849));
  OR2 OR2_73(.VSS(VSS),.VDD(VDD),.Y(g23089),.A(g21806),.B(g21799));
  OR3 OR3_87(.VSS(VSS),.VDD(VDD),.Y(g23100),.A(g21821),.B(g21817),.C(g21856));
  OR2 OR2_74(.VSS(VSS),.VDD(VDD),.Y(g23107),.A(g21813),.B(g21807));
  OR2 OR2_75(.VSS(VSS),.VDD(VDD),.Y(g23120),.A(g21819),.B(g21814));
  OR2 OR2_76(.VSS(VSS),.VDD(VDD),.Y(g23129),.A(g21823),.B(g21820));
  OR2 OR2_77(.VSS(VSS),.VDD(VDD),.Y(g23319),.A(g14493),.B(g22385));
  OR2 OR2_78(.VSS(VSS),.VDD(VDD),.Y(g23688),.A(g23106),.B(g21906));
  OR2 OR2_79(.VSS(VSS),.VDD(VDD),.Y(g23742),.A(g23119),.B(g21920));
  OR2 OR2_80(.VSS(VSS),.VDD(VDD),.Y(g23797),.A(g23128),.B(g21938));
  OR2 OR2_81(.VSS(VSS),.VDD(VDD),.Y(g23850),.A(g23139),.B(g20647));
  OR2 OR2_82(.VSS(VSS),.VDD(VDD),.Y(g23919),.A(g22666),.B(g23140));
  OR2 OR2_83(.VSS(VSS),.VDD(VDD),.Y(g24239),.A(g19387),.B(g22401));
  OR2 OR2_84(.VSS(VSS),.VDD(VDD),.Y(g24244),.A(g14144),.B(g22317));
  OR2 OR2_85(.VSS(VSS),.VDD(VDD),.Y(g24245),.A(g19417),.B(g22402));
  OR2 OR2_86(.VSS(VSS),.VDD(VDD),.Y(g24252),.A(g14259),.B(g22342));
  OR2 OR2_87(.VSS(VSS),.VDD(VDD),.Y(g24254),.A(g19454),.B(g22403));
  OR2 OR2_88(.VSS(VSS),.VDD(VDD),.Y(g24257),.A(g14381),.B(g22365));
  OR2 OR2_89(.VSS(VSS),.VDD(VDD),.Y(g24258),.A(g19481),.B(g22404));
  OR2 OR2_90(.VSS(VSS),.VDD(VDD),.Y(g24633),.A(g24094),.B(g20842));
  OR2 OR2_91(.VSS(VSS),.VDD(VDD),.Y(g24653),.A(g24095),.B(g20850));
  OR2 OR2_92(.VSS(VSS),.VDD(VDD),.Y(g24672),.A(g24097),.B(g20858));
  OR2 OR2_93(.VSS(VSS),.VDD(VDD),.Y(g24691),.A(g24103),.B(g20866));
  OR2 OR2_94(.VSS(VSS),.VDD(VDD),.Y(g24890),.A(g23639),.B(g23144));
  OR2 OR2_95(.VSS(VSS),.VDD(VDD),.Y(g24909),.A(g23726),.B(g23142));
  OR2 OR2_96(.VSS(VSS),.VDD(VDD),.Y(g24925),.A(g23772),.B(g23141));
  OR2 OR2_97(.VSS(VSS),.VDD(VDD),.Y(g24965),.A(g23922),.B(g23945));
  OR2 OR2_98(.VSS(VSS),.VDD(VDD),.Y(g24978),.A(g23954),.B(g23974));
  OR2 OR2_99(.VSS(VSS),.VDD(VDD),.Y(g24989),.A(g23983),.B(g24004));
  OR2 OR2_100(.VSS(VSS),.VDD(VDD),.Y(g25000),.A(g24013),.B(g24038));
  OR2 OR2_101(.VSS(VSS),.VDD(VDD),.Y(g25183),.A(g24958),.B(g24893));
  OR2 OR2_102(.VSS(VSS),.VDD(VDD),.Y(g25186),.A(g24969),.B(g24916));
  OR2 OR2_103(.VSS(VSS),.VDD(VDD),.Y(g25190),.A(g24982),.B(g24933));
  OR2 OR2_104(.VSS(VSS),.VDD(VDD),.Y(g25195),.A(g24993),.B(g24945));
  OR2 OR2_105(.VSS(VSS),.VDD(VDD),.Y(g25489),.A(g24795),.B(g16466));
  OR2 OR2_106(.VSS(VSS),.VDD(VDD),.Y(g25490),.A(g24759),.B(g23146));
  OR2 OR2_107(.VSS(VSS),.VDD(VDD),.Y(g25520),.A(g24813),.B(g23145));
  OR2 OR2_108(.VSS(VSS),.VDD(VDD),.Y(g25566),.A(g24843),.B(g23143));
  OR2 OR2_109(.VSS(VSS),.VDD(VDD),.Y(g26320),.A(g25852),.B(g25870));
  OR2 OR2_110(.VSS(VSS),.VDD(VDD),.Y(g26367),.A(g25873),.B(g25882));
  OR2 OR2_111(.VSS(VSS),.VDD(VDD),.Y(g26410),.A(g25885),.B(g25887));
  OR2 OR2_112(.VSS(VSS),.VDD(VDD),.Y(g26451),.A(g25890),.B(g25892));
  OR2 OR2_113(.VSS(VSS),.VDD(VDD),.Y(g26974),.A(g26157),.B(g23147));
  OR3 OR3_88(.VSS(VSS),.VDD(VDD),.Y(g27113),.A(g1248),.B(g1245),.C(g26534));
  OR2 OR2_114(.VSS(VSS),.VDD(VDD),.Y(g28501),.A(g27738),.B(g25764));
  OR2 OR2_115(.VSS(VSS),.VDD(VDD),.Y(g28512),.A(g26481),.B(g27738));
  OR2 OR2_116(.VSS(VSS),.VDD(VDD),.Y(g28529),.A(g27743),.B(g25818));
  OR2 OR2_117(.VSS(VSS),.VDD(VDD),.Y(g28540),.A(g26497),.B(g27743));
  OR2 OR2_118(.VSS(VSS),.VDD(VDD),.Y(g28556),.A(g27751),.B(g25853));
  OR2 OR2_119(.VSS(VSS),.VDD(VDD),.Y(g28567),.A(g26512),.B(g27751));
  OR2 OR2_120(.VSS(VSS),.VDD(VDD),.Y(g28584),.A(g27756),.B(g25874));
  OR2 OR2_121(.VSS(VSS),.VDD(VDD),.Y(g28595),.A(g26520),.B(g27756));
  OR3 OR3_89(.VSS(VSS),.VDD(VDD),.Y(g29348),.A(g1942),.B(g1939),.C(g29113));
  OR3 OR3_90(.VSS(VSS),.VDD(VDD),.Y(g30305),.A(g2636),.B(g2633),.C(g30072));
//
  NAND2 NAND2_0(.VSS(VSS),.VDD(VDD),.Y(I15167),.A(g2981),.B(g2874));
  NAND2 NAND2_1(.VSS(VSS),.VDD(VDD),.Y(I15168),.A(g2981),.B(I15167));
  NAND2 NAND2_2(.VSS(VSS),.VDD(VDD),.Y(I15169),.A(g2874),.B(I15167));
  NAND2 NAND2_3(.VSS(VSS),.VDD(VDD),.Y(g7855),.A(I15168),.B(I15169));
  NAND2 NAND2_4(.VSS(VSS),.VDD(VDD),.Y(I15183),.A(g2975),.B(g2978));
  NAND2 NAND2_5(.VSS(VSS),.VDD(VDD),.Y(I15184),.A(g2975),.B(I15183));
  NAND2 NAND2_6(.VSS(VSS),.VDD(VDD),.Y(I15185),.A(g2978),.B(I15183));
  NAND2 NAND2_7(.VSS(VSS),.VDD(VDD),.Y(g7875),.A(I15184),.B(I15185));
  NAND2 NAND2_8(.VSS(VSS),.VDD(VDD),.Y(I15190),.A(g2956),.B(g2959));
  NAND2 NAND2_9(.VSS(VSS),.VDD(VDD),.Y(I15191),.A(g2956),.B(I15190));
  NAND2 NAND2_10(.VSS(VSS),.VDD(VDD),.Y(I15192),.A(g2959),.B(I15190));
  NAND2 NAND2_11(.VSS(VSS),.VDD(VDD),.Y(g7876),.A(I15191),.B(I15192));
  NAND2 NAND2_12(.VSS(VSS),.VDD(VDD),.Y(I15204),.A(g2969),.B(g2972));
  NAND2 NAND2_13(.VSS(VSS),.VDD(VDD),.Y(I15205),.A(g2969),.B(I15204));
  NAND2 NAND2_14(.VSS(VSS),.VDD(VDD),.Y(I15206),.A(g2972),.B(I15204));
  NAND2 NAND2_15(.VSS(VSS),.VDD(VDD),.Y(g7895),.A(I15205),.B(I15206));
  NAND2 NAND2_16(.VSS(VSS),.VDD(VDD),.Y(I15211),.A(g2947),.B(g2953));
  NAND2 NAND2_17(.VSS(VSS),.VDD(VDD),.Y(I15212),.A(g2947),.B(I15211));
  NAND2 NAND2_18(.VSS(VSS),.VDD(VDD),.Y(I15213),.A(g2953),.B(I15211));
  NAND2 NAND2_19(.VSS(VSS),.VDD(VDD),.Y(g7896),.A(I15212),.B(I15213));
  NAND2 NAND2_20(.VSS(VSS),.VDD(VDD),.Y(I15237),.A(g2963),.B(g2966));
  NAND2 NAND2_21(.VSS(VSS),.VDD(VDD),.Y(I15238),.A(g2963),.B(I15237));
  NAND2 NAND2_22(.VSS(VSS),.VDD(VDD),.Y(I15239),.A(g2966),.B(I15237));
  NAND2 NAND2_23(.VSS(VSS),.VDD(VDD),.Y(g7922),.A(I15238),.B(I15239));
  NAND2 NAND2_24(.VSS(VSS),.VDD(VDD),.Y(I15244),.A(g2941),.B(g2944));
  NAND2 NAND2_25(.VSS(VSS),.VDD(VDD),.Y(I15245),.A(g2941),.B(I15244));
  NAND2 NAND2_26(.VSS(VSS),.VDD(VDD),.Y(I15246),.A(g2944),.B(I15244));
  NAND2 NAND2_27(.VSS(VSS),.VDD(VDD),.Y(g7923),.A(I15245),.B(I15246));
  NAND2 NAND2_28(.VSS(VSS),.VDD(VDD),.Y(I15276),.A(g2935),.B(g2938));
  NAND2 NAND2_29(.VSS(VSS),.VDD(VDD),.Y(I15277),.A(g2935),.B(I15276));
  NAND2 NAND2_30(.VSS(VSS),.VDD(VDD),.Y(I15278),.A(g2938),.B(I15276));
  NAND2 NAND2_31(.VSS(VSS),.VDD(VDD),.Y(g7970),.A(I15277),.B(I15278));
  NAND4 NAND4_0(.VSS(VSS),.VDD(VDD),.Y(g8381),.A(g8182),.B(g8120),.C(g8044),.D(g7989));
  NAND2 NAND2_32(.VSS(VSS),.VDD(VDD),.Y(g8533),.A(g3398),.B(g3366));
  NAND2 NAND2_33(.VSS(VSS),.VDD(VDD),.Y(g8547),.A(g3398),.B(g3366));
  NAND2 NAND2_34(.VSS(VSS),.VDD(VDD),.Y(g8550),.A(g3554),.B(g3522));
  NAND2 NAND2_35(.VSS(VSS),.VDD(VDD),.Y(g8560),.A(g3554),.B(g3522));
  NAND2 NAND2_36(.VSS(VSS),.VDD(VDD),.Y(g8563),.A(g3710),.B(g3678));
  NAND2 NAND2_37(.VSS(VSS),.VDD(VDD),.Y(g8571),.A(g3710),.B(g3678));
  NAND2 NAND2_38(.VSS(VSS),.VDD(VDD),.Y(g8574),.A(g3866),.B(g3834));
  NAND2 NAND2_39(.VSS(VSS),.VDD(VDD),.Y(g8577),.A(g3866),.B(g3834));
  NAND2 NAND2_40(.VSS(VSS),.VDD(VDD),.Y(I16879),.A(g4203),.B(g3998));
  NAND2 NAND2_41(.VSS(VSS),.VDD(VDD),.Y(I16880),.A(g4203),.B(I16879));
  NAND2 NAND2_42(.VSS(VSS),.VDD(VDD),.Y(I16881),.A(g3998),.B(I16879));
  NAND2 NAND2_43(.VSS(VSS),.VDD(VDD),.Y(g9883),.A(I16880),.B(I16881));
  NAND2 NAND2_44(.VSS(VSS),.VDD(VDD),.Y(I16965),.A(g4734),.B(g4452));
  NAND2 NAND2_45(.VSS(VSS),.VDD(VDD),.Y(I16966),.A(g4734),.B(I16965));
  NAND2 NAND2_46(.VSS(VSS),.VDD(VDD),.Y(I16967),.A(g4452),.B(I16965));
  NAND2 NAND2_47(.VSS(VSS),.VDD(VDD),.Y(g10003),.A(I16966),.B(I16967));
  NAND2 NAND2_48(.VSS(VSS),.VDD(VDD),.Y(g10038),.A(g7772),.B(g3366));
  NAND2 NAND2_49(.VSS(VSS),.VDD(VDD),.Y(I17059),.A(g6637),.B(g6309));
  NAND2 NAND2_50(.VSS(VSS),.VDD(VDD),.Y(I17060),.A(g6637),.B(I17059));
  NAND2 NAND2_51(.VSS(VSS),.VDD(VDD),.Y(I17061),.A(g6309),.B(I17059));
  NAND2 NAND2_52(.VSS(VSS),.VDD(VDD),.Y(g10095),.A(I17060),.B(I17061));
  NAND2 NAND2_53(.VSS(VSS),.VDD(VDD),.Y(g10147),.A(g7788),.B(g3522));
  NAND2 NAND2_54(.VSS(VSS),.VDD(VDD),.Y(I17149),.A(g7465),.B(g7142));
  NAND2 NAND2_55(.VSS(VSS),.VDD(VDD),.Y(I17150),.A(g7465),.B(I17149));
  NAND2 NAND2_56(.VSS(VSS),.VDD(VDD),.Y(I17151),.A(g7142),.B(I17149));
  NAND2 NAND2_57(.VSS(VSS),.VDD(VDD),.Y(g10185),.A(I17150),.B(I17151));
  NAND2 NAND2_58(.VSS(VSS),.VDD(VDD),.Y(g10252),.A(g7802),.B(g3678));
  NAND2 NAND2_59(.VSS(VSS),.VDD(VDD),.Y(g10354),.A(g7815),.B(g3834));
  NAND2 NAND2_60(.VSS(VSS),.VDD(VDD),.Y(g10649),.A(g3398),.B(g6912));
  NAND2 NAND2_61(.VSS(VSS),.VDD(VDD),.Y(g10676),.A(g3398),.B(g6678));
  NAND2 NAND2_62(.VSS(VSS),.VDD(VDD),.Y(g10677),.A(g3398),.B(g6912));
  NAND2 NAND2_63(.VSS(VSS),.VDD(VDD),.Y(g10679),.A(g3554),.B(g7162));
  NAND2 NAND2_64(.VSS(VSS),.VDD(VDD),.Y(g10703),.A(g3398),.B(g6678));
  NAND2 NAND2_65(.VSS(VSS),.VDD(VDD),.Y(g10705),.A(g3554),.B(g6980));
  NAND2 NAND2_66(.VSS(VSS),.VDD(VDD),.Y(g10706),.A(g3554),.B(g7162));
  NAND2 NAND2_67(.VSS(VSS),.VDD(VDD),.Y(g10708),.A(g3710),.B(g7358));
  NAND2 NAND2_68(.VSS(VSS),.VDD(VDD),.Y(g10723),.A(g3554),.B(g6980));
  NAND2 NAND2_69(.VSS(VSS),.VDD(VDD),.Y(g10725),.A(g3710),.B(g7230));
  NAND2 NAND2_70(.VSS(VSS),.VDD(VDD),.Y(g10726),.A(g3710),.B(g7358));
  NAND2 NAND2_71(.VSS(VSS),.VDD(VDD),.Y(g10728),.A(g3866),.B(g7488));
  NAND2 NAND2_72(.VSS(VSS),.VDD(VDD),.Y(g10744),.A(g3710),.B(g7230));
  NAND2 NAND2_73(.VSS(VSS),.VDD(VDD),.Y(g10746),.A(g3866),.B(g7426));
  NAND2 NAND2_74(.VSS(VSS),.VDD(VDD),.Y(g10747),.A(g3866),.B(g7488));
  NAND2 NAND2_75(.VSS(VSS),.VDD(VDD),.Y(g10763),.A(g3866),.B(g7426));
  NAND2 NAND2_76(.VSS(VSS),.VDD(VDD),.Y(I18106),.A(g7875),.B(g7855));
  NAND2 NAND2_77(.VSS(VSS),.VDD(VDD),.Y(I18107),.A(g7875),.B(I18106));
  NAND2 NAND2_78(.VSS(VSS),.VDD(VDD),.Y(I18108),.A(g7855),.B(I18106));
  NAND2 NAND2_79(.VSS(VSS),.VDD(VDD),.Y(g11188),.A(I18107),.B(I18108));
  NAND2 NAND2_80(.VSS(VSS),.VDD(VDD),.Y(I18113),.A(g3997),.B(g8181));
  NAND2 NAND2_81(.VSS(VSS),.VDD(VDD),.Y(I18114),.A(g3997),.B(I18113));
  NAND2 NAND2_82(.VSS(VSS),.VDD(VDD),.Y(I18115),.A(g8181),.B(I18113));
  NAND2 NAND2_83(.VSS(VSS),.VDD(VDD),.Y(g11189),.A(I18114),.B(I18115));
  NAND2 NAND2_84(.VSS(VSS),.VDD(VDD),.Y(I18190),.A(g7922),.B(g7895));
  NAND2 NAND2_85(.VSS(VSS),.VDD(VDD),.Y(I18191),.A(g7922),.B(I18190));
  NAND2 NAND2_86(.VSS(VSS),.VDD(VDD),.Y(I18192),.A(g7895),.B(I18190));
  NAND2 NAND2_87(.VSS(VSS),.VDD(VDD),.Y(g11262),.A(I18191),.B(I18192));
  NAND2 NAND2_88(.VSS(VSS),.VDD(VDD),.Y(I18197),.A(g7896),.B(g7876));
  NAND2 NAND2_89(.VSS(VSS),.VDD(VDD),.Y(I18198),.A(g7896),.B(I18197));
  NAND2 NAND2_90(.VSS(VSS),.VDD(VDD),.Y(I18199),.A(g7876),.B(I18197));
  NAND2 NAND2_91(.VSS(VSS),.VDD(VDD),.Y(g11263),.A(I18198),.B(I18199));
  NAND2 NAND2_92(.VSS(VSS),.VDD(VDD),.Y(I18204),.A(g7975),.B(g4202));
  NAND2 NAND2_93(.VSS(VSS),.VDD(VDD),.Y(I18205),.A(g7975),.B(I18204));
  NAND2 NAND2_94(.VSS(VSS),.VDD(VDD),.Y(I18206),.A(g4202),.B(I18204));
  NAND2 NAND2_95(.VSS(VSS),.VDD(VDD),.Y(g11264),.A(I18205),.B(I18206));
  NAND2 NAND2_96(.VSS(VSS),.VDD(VDD),.Y(I18280),.A(g7970),.B(g7923));
  NAND2 NAND2_97(.VSS(VSS),.VDD(VDD),.Y(I18281),.A(g7970),.B(I18280));
  NAND2 NAND2_98(.VSS(VSS),.VDD(VDD),.Y(I18282),.A(g7923),.B(I18280));
  NAND2 NAND2_99(.VSS(VSS),.VDD(VDD),.Y(g11330),.A(I18281),.B(I18282));
  NAND2 NAND2_100(.VSS(VSS),.VDD(VDD),.Y(I18287),.A(g8256),.B(g8102));
  NAND2 NAND2_101(.VSS(VSS),.VDD(VDD),.Y(I18288),.A(g8256),.B(I18287));
  NAND2 NAND2_102(.VSS(VSS),.VDD(VDD),.Y(I18289),.A(g8102),.B(I18287));
  NAND2 NAND2_103(.VSS(VSS),.VDD(VDD),.Y(g11331),.A(I18288),.B(I18289));
  NAND2 NAND2_104(.VSS(VSS),.VDD(VDD),.Y(I18368),.A(g4325),.B(g4093));
  NAND2 NAND2_105(.VSS(VSS),.VDD(VDD),.Y(I18369),.A(g4325),.B(I18368));
  NAND2 NAND2_106(.VSS(VSS),.VDD(VDD),.Y(I18370),.A(g4093),.B(I18368));
  NAND2 NAND2_107(.VSS(VSS),.VDD(VDD),.Y(g11410),.A(I18369),.B(I18370));
  NAND2 NAND2_108(.VSS(VSS),.VDD(VDD),.Y(g11617),.A(g8313),.B(g2883));
  NAND2 NAND2_109(.VSS(VSS),.VDD(VDD),.Y(I18799),.A(g11410),.B(g11331));
  NAND2 NAND2_110(.VSS(VSS),.VDD(VDD),.Y(I18800),.A(g11410),.B(I18799));
  NAND2 NAND2_111(.VSS(VSS),.VDD(VDD),.Y(I18801),.A(g11331),.B(I18799));
  NAND2 NAND2_112(.VSS(VSS),.VDD(VDD),.Y(g11621),.A(I18800),.B(I18801));
  NAND2 NAND2_113(.VSS(VSS),.VDD(VDD),.Y(g11661),.A(g9534),.B(g3366));
  NAND2 NAND2_114(.VSS(VSS),.VDD(VDD),.Y(g11662),.A(g9534),.B(g3366));
  NAND2 NAND2_115(.VSS(VSS),.VDD(VDD),.Y(g11672),.A(g9534),.B(g3366));
  NAND2 NAND2_116(.VSS(VSS),.VDD(VDD),.Y(g11673),.A(g9676),.B(g3522));
  NAND2 NAND2_117(.VSS(VSS),.VDD(VDD),.Y(g11674),.A(g9676),.B(g3522));
  NAND2 NAND2_118(.VSS(VSS),.VDD(VDD),.Y(g11683),.A(g9534),.B(g3366));
  NAND2 NAND2_119(.VSS(VSS),.VDD(VDD),.Y(g11684),.A(g9676),.B(g3522));
  NAND2 NAND2_120(.VSS(VSS),.VDD(VDD),.Y(g11685),.A(g9822),.B(g3678));
  NAND2 NAND2_121(.VSS(VSS),.VDD(VDD),.Y(g11686),.A(g9822),.B(g3678));
  NAND2 NAND2_122(.VSS(VSS),.VDD(VDD),.Y(g11691),.A(g9534),.B(g3366));
  NAND2 NAND2_123(.VSS(VSS),.VDD(VDD),.Y(g11692),.A(g9676),.B(g3522));
  NAND2 NAND2_124(.VSS(VSS),.VDD(VDD),.Y(g11693),.A(g9822),.B(g3678));
  NAND2 NAND2_125(.VSS(VSS),.VDD(VDD),.Y(g11694),.A(g9968),.B(g3834));
  NAND2 NAND2_126(.VSS(VSS),.VDD(VDD),.Y(g11695),.A(g9968),.B(g3834));
  NAND2 NAND2_127(.VSS(VSS),.VDD(VDD),.Y(g11696),.A(g9534),.B(g3366));
  NAND2 NAND2_128(.VSS(VSS),.VDD(VDD),.Y(g11698),.A(g9676),.B(g3522));
  NAND2 NAND2_129(.VSS(VSS),.VDD(VDD),.Y(g11699),.A(g9822),.B(g3678));
  NAND2 NAND2_130(.VSS(VSS),.VDD(VDD),.Y(g11700),.A(g9968),.B(g3834));
  NAND2 NAND2_131(.VSS(VSS),.VDD(VDD),.Y(g11701),.A(g9534),.B(g3366));
  NAND2 NAND2_132(.VSS(VSS),.VDD(VDD),.Y(g11702),.A(g9676),.B(g3522));
  NAND2 NAND2_133(.VSS(VSS),.VDD(VDD),.Y(g11704),.A(g9822),.B(g3678));
  NAND2 NAND2_134(.VSS(VSS),.VDD(VDD),.Y(g11705),.A(g9968),.B(g3834));
  NAND2 NAND2_135(.VSS(VSS),.VDD(VDD),.Y(g11707),.A(g9534),.B(g3366));
  NAND2 NAND2_136(.VSS(VSS),.VDD(VDD),.Y(g11708),.A(g9534),.B(g3366));
  NAND2 NAND2_137(.VSS(VSS),.VDD(VDD),.Y(g11709),.A(g9676),.B(g3522));
  NAND2 NAND2_138(.VSS(VSS),.VDD(VDD),.Y(g11710),.A(g9822),.B(g3678));
  NAND2 NAND2_139(.VSS(VSS),.VDD(VDD),.Y(g11712),.A(g9968),.B(g3834));
  NAND2 NAND2_140(.VSS(VSS),.VDD(VDD),.Y(g11713),.A(g10481),.B(g9144));
  NAND2 NAND2_141(.VSS(VSS),.VDD(VDD),.Y(g11716),.A(g9534),.B(g3366));
  NAND2 NAND2_142(.VSS(VSS),.VDD(VDD),.Y(g11717),.A(g9676),.B(g3522));
  NAND2 NAND2_143(.VSS(VSS),.VDD(VDD),.Y(g11718),.A(g9676),.B(g3522));
  NAND2 NAND2_144(.VSS(VSS),.VDD(VDD),.Y(g11719),.A(g9822),.B(g3678));
  NAND2 NAND2_145(.VSS(VSS),.VDD(VDD),.Y(g11720),.A(g9968),.B(g3834));
  NAND2 NAND2_146(.VSS(VSS),.VDD(VDD),.Y(g11721),.A(g9534),.B(g3366));
  NAND2 NAND2_147(.VSS(VSS),.VDD(VDD),.Y(g11722),.A(g9676),.B(g3522));
  NAND2 NAND2_148(.VSS(VSS),.VDD(VDD),.Y(g11723),.A(g9822),.B(g3678));
  NAND2 NAND2_149(.VSS(VSS),.VDD(VDD),.Y(g11724),.A(g9822),.B(g3678));
  NAND2 NAND2_150(.VSS(VSS),.VDD(VDD),.Y(g11725),.A(g9968),.B(g3834));
  NAND2 NAND2_151(.VSS(VSS),.VDD(VDD),.Y(g11726),.A(g9676),.B(g3522));
  NAND2 NAND2_152(.VSS(VSS),.VDD(VDD),.Y(g11727),.A(g9822),.B(g3678));
  NAND2 NAND2_153(.VSS(VSS),.VDD(VDD),.Y(g11728),.A(g9968),.B(g3834));
  NAND2 NAND2_154(.VSS(VSS),.VDD(VDD),.Y(g11729),.A(g9968),.B(g3834));
  NAND2 NAND2_155(.VSS(VSS),.VDD(VDD),.Y(g11730),.A(g9822),.B(g3678));
  NAND2 NAND2_156(.VSS(VSS),.VDD(VDD),.Y(g11731),.A(g9968),.B(g3834));
  NAND2 NAND2_157(.VSS(VSS),.VDD(VDD),.Y(g11733),.A(g9968),.B(g3834));
  NAND2 NAND2_158(.VSS(VSS),.VDD(VDD),.Y(g12433),.A(g2879),.B(g10778));
  NAND2 NAND2_159(.VSS(VSS),.VDD(VDD),.Y(g12486),.A(g8278),.B(g6448));
  NAND2 NAND2_160(.VSS(VSS),.VDD(VDD),.Y(g12503),.A(g8278),.B(g5438));
  NAND2 NAND2_161(.VSS(VSS),.VDD(VDD),.Y(g12506),.A(g8287),.B(g6713));
  NAND2 NAND2_162(.VSS(VSS),.VDD(VDD),.Y(g12520),.A(g8287),.B(g5473));
  NAND2 NAND2_163(.VSS(VSS),.VDD(VDD),.Y(g12523),.A(g8296),.B(g7015));
  NAND2 NAND2_164(.VSS(VSS),.VDD(VDD),.Y(g12535),.A(g8296),.B(g5512));
  NAND2 NAND2_165(.VSS(VSS),.VDD(VDD),.Y(g12538),.A(g8305),.B(g7265));
  NAND2 NAND2_166(.VSS(VSS),.VDD(VDD),.Y(g12544),.A(g8305),.B(g5556));
  NAND2 NAND2_167(.VSS(VSS),.VDD(VDD),.Y(I20031),.A(g10003),.B(g9883));
  NAND2 NAND2_168(.VSS(VSS),.VDD(VDD),.Y(I20032),.A(g10003),.B(I20031));
  NAND2 NAND2_169(.VSS(VSS),.VDD(VDD),.Y(I20033),.A(g9883),.B(I20031));
  NAND2 NAND2_170(.VSS(VSS),.VDD(VDD),.Y(g12988),.A(I20032),.B(I20033));
  NAND2 NAND2_171(.VSS(VSS),.VDD(VDD),.Y(I20048),.A(g10185),.B(g10095));
  NAND2 NAND2_172(.VSS(VSS),.VDD(VDD),.Y(I20049),.A(g10185),.B(I20048));
  NAND2 NAND2_173(.VSS(VSS),.VDD(VDD),.Y(I20050),.A(g10095),.B(I20048));
  NAND2 NAND2_174(.VSS(VSS),.VDD(VDD),.Y(g12999),.A(I20049),.B(I20050));
  NAND2 NAND2_175(.VSS(VSS),.VDD(VDD),.Y(g13020),.A(g9534),.B(g6912));
  NAND2 NAND2_176(.VSS(VSS),.VDD(VDD),.Y(g13021),.A(g9534),.B(g6912));
  NAND2 NAND2_177(.VSS(VSS),.VDD(VDD),.Y(g13026),.A(g9534),.B(g6678));
  NAND2 NAND2_178(.VSS(VSS),.VDD(VDD),.Y(g13027),.A(g9534),.B(g6912));
  NAND2 NAND2_179(.VSS(VSS),.VDD(VDD),.Y(g13028),.A(g9534),.B(g6678));
  NAND2 NAND2_180(.VSS(VSS),.VDD(VDD),.Y(g13029),.A(g9676),.B(g7162));
  NAND2 NAND2_181(.VSS(VSS),.VDD(VDD),.Y(g13030),.A(g9676),.B(g7162));
  NAND2 NAND2_182(.VSS(VSS),.VDD(VDD),.Y(g13034),.A(g9534),.B(g6678));
  NAND2 NAND2_183(.VSS(VSS),.VDD(VDD),.Y(g13035),.A(g9534),.B(g6912));
  NAND2 NAND2_184(.VSS(VSS),.VDD(VDD),.Y(g13037),.A(g9676),.B(g6980));
  NAND2 NAND2_185(.VSS(VSS),.VDD(VDD),.Y(g13038),.A(g9676),.B(g7162));
  NAND2 NAND2_186(.VSS(VSS),.VDD(VDD),.Y(g13039),.A(g9676),.B(g6980));
  NAND2 NAND2_187(.VSS(VSS),.VDD(VDD),.Y(g13040),.A(g9822),.B(g7358));
  NAND2 NAND2_188(.VSS(VSS),.VDD(VDD),.Y(g13041),.A(g9822),.B(g7358));
  NAND2 NAND2_189(.VSS(VSS),.VDD(VDD),.Y(g13044),.A(g9534),.B(g6678));
  NAND2 NAND2_190(.VSS(VSS),.VDD(VDD),.Y(g13045),.A(g9534),.B(g6912));
  NAND2 NAND2_191(.VSS(VSS),.VDD(VDD),.Y(g13047),.A(g9676),.B(g6980));
  NAND2 NAND2_192(.VSS(VSS),.VDD(VDD),.Y(g13048),.A(g9676),.B(g7162));
  NAND2 NAND2_193(.VSS(VSS),.VDD(VDD),.Y(g13050),.A(g9822),.B(g7230));
  NAND2 NAND2_194(.VSS(VSS),.VDD(VDD),.Y(g13051),.A(g9822),.B(g7358));
  NAND2 NAND2_195(.VSS(VSS),.VDD(VDD),.Y(g13052),.A(g9822),.B(g7230));
  NAND2 NAND2_196(.VSS(VSS),.VDD(VDD),.Y(g13053),.A(g9968),.B(g7488));
  NAND2 NAND2_197(.VSS(VSS),.VDD(VDD),.Y(g13054),.A(g9968),.B(g7488));
  NAND2 NAND2_198(.VSS(VSS),.VDD(VDD),.Y(g13058),.A(g9534),.B(g6678));
  NAND2 NAND2_199(.VSS(VSS),.VDD(VDD),.Y(g13059),.A(g9534),.B(g6912));
  NAND2 NAND2_200(.VSS(VSS),.VDD(VDD),.Y(g13061),.A(g9676),.B(g6980));
  NAND2 NAND2_201(.VSS(VSS),.VDD(VDD),.Y(g13062),.A(g9676),.B(g7162));
  NAND2 NAND2_202(.VSS(VSS),.VDD(VDD),.Y(g13064),.A(g9822),.B(g7230));
  NAND2 NAND2_203(.VSS(VSS),.VDD(VDD),.Y(g13065),.A(g9822),.B(g7358));
  NAND2 NAND2_204(.VSS(VSS),.VDD(VDD),.Y(g13067),.A(g9968),.B(g7426));
  NAND2 NAND2_205(.VSS(VSS),.VDD(VDD),.Y(g13068),.A(g9968),.B(g7488));
  NAND2 NAND2_206(.VSS(VSS),.VDD(VDD),.Y(g13069),.A(g9968),.B(g7426));
  NAND2 NAND2_207(.VSS(VSS),.VDD(VDD),.Y(g13071),.A(g9534),.B(g6678));
  NAND2 NAND2_208(.VSS(VSS),.VDD(VDD),.Y(g13072),.A(g9534),.B(g6912));
  NAND2 NAND2_209(.VSS(VSS),.VDD(VDD),.Y(g13074),.A(g9676),.B(g6980));
  NAND2 NAND2_210(.VSS(VSS),.VDD(VDD),.Y(g13075),.A(g9676),.B(g7162));
  NAND2 NAND2_211(.VSS(VSS),.VDD(VDD),.Y(g13077),.A(g9822),.B(g7230));
  NAND2 NAND2_212(.VSS(VSS),.VDD(VDD),.Y(g13078),.A(g9822),.B(g7358));
  NAND2 NAND2_213(.VSS(VSS),.VDD(VDD),.Y(g13080),.A(g9968),.B(g7426));
  NAND2 NAND2_214(.VSS(VSS),.VDD(VDD),.Y(g13081),.A(g9968),.B(g7488));
  NAND2 NAND2_215(.VSS(VSS),.VDD(VDD),.Y(g13087),.A(g9534),.B(g6678));
  NAND2 NAND2_216(.VSS(VSS),.VDD(VDD),.Y(g13088),.A(g9534),.B(g6912));
  NAND2 NAND2_217(.VSS(VSS),.VDD(VDD),.Y(g13089),.A(g9534),.B(g6912));
  NAND2 NAND2_218(.VSS(VSS),.VDD(VDD),.Y(g13090),.A(g9676),.B(g6980));
  NAND2 NAND2_219(.VSS(VSS),.VDD(VDD),.Y(g13091),.A(g9676),.B(g7162));
  NAND2 NAND2_220(.VSS(VSS),.VDD(VDD),.Y(g13093),.A(g9822),.B(g7230));
  NAND2 NAND2_221(.VSS(VSS),.VDD(VDD),.Y(g13094),.A(g9822),.B(g7358));
  NAND2 NAND2_222(.VSS(VSS),.VDD(VDD),.Y(g13096),.A(g9968),.B(g7426));
  NAND2 NAND2_223(.VSS(VSS),.VDD(VDD),.Y(g13097),.A(g9968),.B(g7488));
  NAND2 NAND2_224(.VSS(VSS),.VDD(VDD),.Y(g13098),.A(g9534),.B(g6678));
  NAND2 NAND2_225(.VSS(VSS),.VDD(VDD),.Y(g13099),.A(g9534),.B(g6912));
  NAND2 NAND2_226(.VSS(VSS),.VDD(VDD),.Y(g13100),.A(g9534),.B(g6678));
  NAND2 NAND2_227(.VSS(VSS),.VDD(VDD),.Y(g13102),.A(g9676),.B(g6980));
  NAND2 NAND2_228(.VSS(VSS),.VDD(VDD),.Y(g13103),.A(g9676),.B(g7162));
  NAND2 NAND2_229(.VSS(VSS),.VDD(VDD),.Y(g13104),.A(g9676),.B(g7162));
  NAND2 NAND2_230(.VSS(VSS),.VDD(VDD),.Y(g13105),.A(g9822),.B(g7230));
  NAND2 NAND2_231(.VSS(VSS),.VDD(VDD),.Y(g13106),.A(g9822),.B(g7358));
  NAND2 NAND2_232(.VSS(VSS),.VDD(VDD),.Y(g13108),.A(g9968),.B(g7426));
  NAND2 NAND2_233(.VSS(VSS),.VDD(VDD),.Y(g13109),.A(g9968),.B(g7488));
  NAND2 NAND2_234(.VSS(VSS),.VDD(VDD),.Y(g13112),.A(g9534),.B(g6678));
  NAND2 NAND2_235(.VSS(VSS),.VDD(VDD),.Y(g13113),.A(g9534),.B(g6912));
  NAND2 NAND2_236(.VSS(VSS),.VDD(VDD),.Y(g13114),.A(g9676),.B(g6980));
  NAND2 NAND2_237(.VSS(VSS),.VDD(VDD),.Y(g13115),.A(g9676),.B(g7162));
  NAND2 NAND2_238(.VSS(VSS),.VDD(VDD),.Y(g13116),.A(g9676),.B(g6980));
  NAND2 NAND2_239(.VSS(VSS),.VDD(VDD),.Y(g13118),.A(g9822),.B(g7230));
  NAND2 NAND2_240(.VSS(VSS),.VDD(VDD),.Y(g13119),.A(g9822),.B(g7358));
  NAND2 NAND2_241(.VSS(VSS),.VDD(VDD),.Y(g13120),.A(g9822),.B(g7358));
  NAND2 NAND2_242(.VSS(VSS),.VDD(VDD),.Y(g13121),.A(g9968),.B(g7426));
  NAND2 NAND2_243(.VSS(VSS),.VDD(VDD),.Y(g13122),.A(g9968),.B(g7488));
  NAND2 NAND2_244(.VSS(VSS),.VDD(VDD),.Y(g13123),.A(g9534),.B(g6678));
  NAND2 NAND2_245(.VSS(VSS),.VDD(VDD),.Y(g13125),.A(g9676),.B(g6980));
  NAND2 NAND2_246(.VSS(VSS),.VDD(VDD),.Y(g13126),.A(g9676),.B(g7162));
  NAND2 NAND2_247(.VSS(VSS),.VDD(VDD),.Y(g13127),.A(g9822),.B(g7230));
  NAND2 NAND2_248(.VSS(VSS),.VDD(VDD),.Y(g13128),.A(g9822),.B(g7358));
  NAND2 NAND2_249(.VSS(VSS),.VDD(VDD),.Y(g13129),.A(g9822),.B(g7230));
  NAND2 NAND2_250(.VSS(VSS),.VDD(VDD),.Y(g13131),.A(g9968),.B(g7426));
  NAND2 NAND2_251(.VSS(VSS),.VDD(VDD),.Y(g13132),.A(g9968),.B(g7488));
  NAND2 NAND2_252(.VSS(VSS),.VDD(VDD),.Y(g13133),.A(g9968),.B(g7488));
  NAND2 NAND2_253(.VSS(VSS),.VDD(VDD),.Y(g13134),.A(g9676),.B(g6980));
  NAND2 NAND2_254(.VSS(VSS),.VDD(VDD),.Y(g13136),.A(g9822),.B(g7230));
  NAND2 NAND2_255(.VSS(VSS),.VDD(VDD),.Y(g13137),.A(g9822),.B(g7358));
  NAND2 NAND2_256(.VSS(VSS),.VDD(VDD),.Y(g13138),.A(g9968),.B(g7426));
  NAND2 NAND2_257(.VSS(VSS),.VDD(VDD),.Y(g13139),.A(g9968),.B(g7488));
  NAND2 NAND2_258(.VSS(VSS),.VDD(VDD),.Y(g13140),.A(g9968),.B(g7426));
  NAND2 NAND2_259(.VSS(VSS),.VDD(VDD),.Y(g13142),.A(g9822),.B(g7230));
  NAND2 NAND2_260(.VSS(VSS),.VDD(VDD),.Y(g13144),.A(g9968),.B(g7426));
  NAND2 NAND2_261(.VSS(VSS),.VDD(VDD),.Y(g13145),.A(g9968),.B(g7488));
  NAND2 NAND2_262(.VSS(VSS),.VDD(VDD),.Y(g13146),.A(g9968),.B(g7426));
  NAND2 NAND2_263(.VSS(VSS),.VDD(VDD),.Y(g13147),.A(g8278),.B(g3306));
  NAND2 NAND2_264(.VSS(VSS),.VDD(VDD),.Y(g13150),.A(g8287),.B(g3462));
  NAND2 NAND2_265(.VSS(VSS),.VDD(VDD),.Y(g13156),.A(g8296),.B(g3618));
  NAND2 NAND2_266(.VSS(VSS),.VDD(VDD),.Y(g13165),.A(g8305),.B(g3774));
  NAND2 NAND2_267(.VSS(VSS),.VDD(VDD),.Y(g13245),.A(g10779),.B(g7901));
  NAND2 NAND2_268(.VSS(VSS),.VDD(VDD),.Y(g13305),.A(g8317),.B(g2993));
  NAND2 NAND2_269(.VSS(VSS),.VDD(VDD),.Y(I20429),.A(g11262),.B(g11188));
  NAND2 NAND2_270(.VSS(VSS),.VDD(VDD),.Y(I20430),.A(g11262),.B(I20429));
  NAND2 NAND2_271(.VSS(VSS),.VDD(VDD),.Y(I20431),.A(g11188),.B(I20429));
  NAND2 NAND2_272(.VSS(VSS),.VDD(VDD),.Y(g13348),.A(I20430),.B(I20431));
  NAND2 NAND2_273(.VSS(VSS),.VDD(VDD),.Y(I20465),.A(g11330),.B(g11263));
  NAND2 NAND2_274(.VSS(VSS),.VDD(VDD),.Y(I20466),.A(g11330),.B(I20465));
  NAND2 NAND2_275(.VSS(VSS),.VDD(VDD),.Y(I20467),.A(g11263),.B(I20465));
  NAND2 NAND2_276(.VSS(VSS),.VDD(VDD),.Y(g13370),.A(I20466),.B(I20467));
  NAND2 NAND2_277(.VSS(VSS),.VDD(VDD),.Y(I20504),.A(g11264),.B(g11189));
  NAND2 NAND2_278(.VSS(VSS),.VDD(VDD),.Y(I20505),.A(g11264),.B(I20504));
  NAND2 NAND2_279(.VSS(VSS),.VDD(VDD),.Y(I20506),.A(g11189),.B(I20504));
  NAND2 NAND2_280(.VSS(VSS),.VDD(VDD),.Y(g13399),.A(I20505),.B(I20506));
  NAND2 NAND2_281(.VSS(VSS),.VDD(VDD),.Y(g13476),.A(g12565),.B(g3254));
  NAND2 NAND2_282(.VSS(VSS),.VDD(VDD),.Y(g13478),.A(g12611),.B(g3410));
  NAND2 NAND2_283(.VSS(VSS),.VDD(VDD),.Y(g13482),.A(g12657),.B(g3566));
  NAND2 NAND2_284(.VSS(VSS),.VDD(VDD),.Y(g13494),.A(g12565),.B(g3254));
  NAND2 NAND2_285(.VSS(VSS),.VDD(VDD),.Y(g13495),.A(g12611),.B(g3410));
  NAND2 NAND2_286(.VSS(VSS),.VDD(VDD),.Y(g13497),.A(g12657),.B(g3566));
  NAND2 NAND2_287(.VSS(VSS),.VDD(VDD),.Y(g13501),.A(g12711),.B(g3722));
  NAND2 NAND2_288(.VSS(VSS),.VDD(VDD),.Y(I20743),.A(g11621),.B(g13399));
  NAND2 NAND2_289(.VSS(VSS),.VDD(VDD),.Y(I20744),.A(g11621),.B(I20743));
  NAND2 NAND2_290(.VSS(VSS),.VDD(VDD),.Y(I20745),.A(g13399),.B(I20743));
  NAND2 NAND2_291(.VSS(VSS),.VDD(VDD),.Y(g13507),.A(I20744),.B(I20745));
  NAND2 NAND2_292(.VSS(VSS),.VDD(VDD),.Y(g13510),.A(g12565),.B(g3254));
  NAND2 NAND2_293(.VSS(VSS),.VDD(VDD),.Y(g13511),.A(g12611),.B(g3410));
  NAND2 NAND2_294(.VSS(VSS),.VDD(VDD),.Y(g13512),.A(g12657),.B(g3566));
  NAND2 NAND2_295(.VSS(VSS),.VDD(VDD),.Y(g13514),.A(g12711),.B(g3722));
  NAND2 NAND2_296(.VSS(VSS),.VDD(VDD),.Y(g13518),.A(g12565),.B(g3254));
  NAND2 NAND2_297(.VSS(VSS),.VDD(VDD),.Y(g13524),.A(g12611),.B(g3410));
  NAND2 NAND2_298(.VSS(VSS),.VDD(VDD),.Y(g13525),.A(g12657),.B(g3566));
  NAND2 NAND2_299(.VSS(VSS),.VDD(VDD),.Y(g13526),.A(g12711),.B(g3722));
  NAND2 NAND2_300(.VSS(VSS),.VDD(VDD),.Y(g13528),.A(g12565),.B(g3254));
  NAND2 NAND2_301(.VSS(VSS),.VDD(VDD),.Y(g13529),.A(g12611),.B(g3410));
  NAND2 NAND2_302(.VSS(VSS),.VDD(VDD),.Y(g13535),.A(g12657),.B(g3566));
  NAND2 NAND2_303(.VSS(VSS),.VDD(VDD),.Y(g13536),.A(g12711),.B(g3722));
  NAND2 NAND2_304(.VSS(VSS),.VDD(VDD),.Y(g13537),.A(g12565),.B(g3254));
  NAND2 NAND2_305(.VSS(VSS),.VDD(VDD),.Y(g13538),.A(g12565),.B(g3254));
  NAND2 NAND2_306(.VSS(VSS),.VDD(VDD),.Y(g13539),.A(g12611),.B(g3410));
  NAND2 NAND2_307(.VSS(VSS),.VDD(VDD),.Y(g13540),.A(g12657),.B(g3566));
  NAND2 NAND2_308(.VSS(VSS),.VDD(VDD),.Y(g13546),.A(g12711),.B(g3722));
  NAND2 NAND2_309(.VSS(VSS),.VDD(VDD),.Y(g13547),.A(g12565),.B(g3254));
  NAND2 NAND2_310(.VSS(VSS),.VDD(VDD),.Y(g13548),.A(g12611),.B(g3410));
  NAND2 NAND2_311(.VSS(VSS),.VDD(VDD),.Y(g13549),.A(g12611),.B(g3410));
  NAND2 NAND2_312(.VSS(VSS),.VDD(VDD),.Y(g13550),.A(g12657),.B(g3566));
  NAND2 NAND2_313(.VSS(VSS),.VDD(VDD),.Y(g13551),.A(g12711),.B(g3722));
  NAND2 NAND2_314(.VSS(VSS),.VDD(VDD),.Y(g13557),.A(g12611),.B(g3410));
  NAND2 NAND2_315(.VSS(VSS),.VDD(VDD),.Y(g13558),.A(g12657),.B(g3566));
  NAND2 NAND2_316(.VSS(VSS),.VDD(VDD),.Y(g13559),.A(g12657),.B(g3566));
  NAND2 NAND2_317(.VSS(VSS),.VDD(VDD),.Y(g13560),.A(g12711),.B(g3722));
  NAND2 NAND2_318(.VSS(VSS),.VDD(VDD),.Y(g13561),.A(g12657),.B(g3566));
  NAND2 NAND2_319(.VSS(VSS),.VDD(VDD),.Y(g13562),.A(g12711),.B(g3722));
  NAND2 NAND2_320(.VSS(VSS),.VDD(VDD),.Y(g13563),.A(g12711),.B(g3722));
  NAND2 NAND2_321(.VSS(VSS),.VDD(VDD),.Y(g13564),.A(g12711),.B(g3722));
  NAND2 NAND2_322(.VSS(VSS),.VDD(VDD),.Y(g13599),.A(g12886),.B(g3366));
  NAND2 NAND2_323(.VSS(VSS),.VDD(VDD),.Y(g13611),.A(g12926),.B(g3522));
  NAND2 NAND2_324(.VSS(VSS),.VDD(VDD),.Y(g13621),.A(g12955),.B(g3678));
  NAND2 NAND2_325(.VSS(VSS),.VDD(VDD),.Y(g13633),.A(g12984),.B(g3834));
  NAND2 NAND2_326(.VSS(VSS),.VDD(VDD),.Y(g13893),.A(g8580),.B(g12463));
  NAND3 NAND3_0(.VSS(VSS),.VDD(VDD),.Y(g13915),.A(g8822),.B(g12473),.C(g12463));
  NAND2 NAND2_327(.VSS(VSS),.VDD(VDD),.Y(g13934),.A(g8587),.B(g12478));
  NAND2 NAND2_328(.VSS(VSS),.VDD(VDD),.Y(g13957),.A(g10730),.B(g12473));
  NAND3 NAND3_1(.VSS(VSS),.VDD(VDD),.Y(g13971),.A(g8846),.B(g12490),.C(g12478));
  NAND2 NAND2_329(.VSS(VSS),.VDD(VDD),.Y(g13990),.A(g8594),.B(g12495));
  NAND2 NAND2_330(.VSS(VSS),.VDD(VDD),.Y(g14027),.A(g10749),.B(g12490));
  NAND3 NAND3_2(.VSS(VSS),.VDD(VDD),.Y(g14041),.A(g8873),.B(g12510),.C(g12495));
  NAND2 NAND2_331(.VSS(VSS),.VDD(VDD),.Y(g14060),.A(g8605),.B(g12515));
  NAND2 NAND2_332(.VSS(VSS),.VDD(VDD),.Y(g14118),.A(g10767),.B(g12510));
  NAND3 NAND3_3(.VSS(VSS),.VDD(VDD),.Y(g14132),.A(g8911),.B(g12527),.C(g12515));
  NAND2 NAND2_333(.VSS(VSS),.VDD(VDD),.Y(g14233),.A(g10773),.B(g12527));
  NAND3 NAND3_4(.VSS(VSS),.VDD(VDD),.Y(g15454),.A(g9232),.B(g9150),.C(g12780));
  NAND3 NAND3_5(.VSS(VSS),.VDD(VDD),.Y(g15540),.A(g9310),.B(g9174),.C(g12819));
  NAND3 NAND3_6(.VSS(VSS),.VDD(VDD),.Y(g15618),.A(g9391),.B(g9216),.C(g12857));
  NAND2 NAND2_334(.VSS(VSS),.VDD(VDD),.Y(g15660),.A(g13401),.B(g12354));
  NAND2 NAND2_335(.VSS(VSS),.VDD(VDD),.Y(g15664),.A(g12565),.B(g6314));
  NAND3 NAND3_7(.VSS(VSS),.VDD(VDD),.Y(g15694),.A(g9488),.B(g9277),.C(g12898));
  NAND2 NAND2_336(.VSS(VSS),.VDD(VDD),.Y(g15718),.A(g13286),.B(g12354));
  NAND2 NAND2_337(.VSS(VSS),.VDD(VDD),.Y(g15719),.A(g13401),.B(g12392));
  NAND2 NAND2_338(.VSS(VSS),.VDD(VDD),.Y(g15720),.A(g12565),.B(g6232));
  NAND2 NAND2_339(.VSS(VSS),.VDD(VDD),.Y(g15721),.A(g12565),.B(g6314));
  NAND2 NAND2_340(.VSS(VSS),.VDD(VDD),.Y(g15723),.A(g12611),.B(g6519));
  NAND2 NAND2_341(.VSS(VSS),.VDD(VDD),.Y(g15756),.A(g13313),.B(g12354));
  NAND2 NAND2_342(.VSS(VSS),.VDD(VDD),.Y(g15757),.A(g11622),.B(g12392));
  NAND2 NAND2_343(.VSS(VSS),.VDD(VDD),.Y(g15758),.A(g12565),.B(g6232));
  NAND2 NAND2_344(.VSS(VSS),.VDD(VDD),.Y(g15759),.A(g12565),.B(g6314));
  NAND2 NAND2_345(.VSS(VSS),.VDD(VDD),.Y(g15760),.A(g12611),.B(g6369));
  NAND2 NAND2_346(.VSS(VSS),.VDD(VDD),.Y(g15761),.A(g12611),.B(g6519));
  NAND2 NAND2_347(.VSS(VSS),.VDD(VDD),.Y(g15763),.A(g12657),.B(g6783));
  NAND2 NAND2_348(.VSS(VSS),.VDD(VDD),.Y(g15782),.A(g13332),.B(g12354));
  NAND2 NAND2_349(.VSS(VSS),.VDD(VDD),.Y(g15783),.A(g11643),.B(g12392));
  NAND2 NAND2_350(.VSS(VSS),.VDD(VDD),.Y(g15784),.A(g12565),.B(g6232));
  NAND2 NAND2_351(.VSS(VSS),.VDD(VDD),.Y(g15785),.A(g12565),.B(g6314));
  NAND2 NAND2_352(.VSS(VSS),.VDD(VDD),.Y(g15786),.A(g12611),.B(g6369));
  NAND2 NAND2_353(.VSS(VSS),.VDD(VDD),.Y(g15787),.A(g12611),.B(g6519));
  NAND2 NAND2_354(.VSS(VSS),.VDD(VDD),.Y(g15788),.A(g12657),.B(g6574));
  NAND2 NAND2_355(.VSS(VSS),.VDD(VDD),.Y(g15789),.A(g12657),.B(g6783));
  NAND2 NAND2_356(.VSS(VSS),.VDD(VDD),.Y(g15791),.A(g12711),.B(g7085));
  NAND2 NAND2_357(.VSS(VSS),.VDD(VDD),.Y(g15803),.A(g13375),.B(g12354));
  NAND2 NAND2_358(.VSS(VSS),.VDD(VDD),.Y(g15804),.A(g11660),.B(g12392));
  NAND2 NAND2_359(.VSS(VSS),.VDD(VDD),.Y(g15805),.A(g12565),.B(g6232));
  NAND2 NAND2_360(.VSS(VSS),.VDD(VDD),.Y(g15806),.A(g12565),.B(g6314));
  NAND2 NAND2_361(.VSS(VSS),.VDD(VDD),.Y(g15807),.A(g12611),.B(g6369));
  NAND2 NAND2_362(.VSS(VSS),.VDD(VDD),.Y(g15808),.A(g12611),.B(g6519));
  NAND2 NAND2_363(.VSS(VSS),.VDD(VDD),.Y(g15809),.A(g12657),.B(g6574));
  NAND2 NAND2_364(.VSS(VSS),.VDD(VDD),.Y(g15810),.A(g12657),.B(g6783));
  NAND2 NAND2_365(.VSS(VSS),.VDD(VDD),.Y(g15811),.A(g12711),.B(g6838));
  NAND2 NAND2_366(.VSS(VSS),.VDD(VDD),.Y(g15812),.A(g12711),.B(g7085));
  NAND2 NAND2_367(.VSS(VSS),.VDD(VDD),.Y(I22062),.A(g12999),.B(g12988));
  NAND2 NAND2_368(.VSS(VSS),.VDD(VDD),.Y(I22063),.A(g12999),.B(I22062));
  NAND2 NAND2_369(.VSS(VSS),.VDD(VDD),.Y(I22064),.A(g12988),.B(I22062));
  NAND2 NAND2_370(.VSS(VSS),.VDD(VDD),.Y(g15814),.A(I22063),.B(I22064));
  NAND2 NAND2_371(.VSS(VSS),.VDD(VDD),.Y(g15818),.A(g13024),.B(g12354));
  NAND2 NAND2_372(.VSS(VSS),.VDD(VDD),.Y(g15819),.A(g13286),.B(g12392));
  NAND2 NAND2_373(.VSS(VSS),.VDD(VDD),.Y(g15820),.A(g12565),.B(g6232));
  NAND2 NAND2_374(.VSS(VSS),.VDD(VDD),.Y(g15821),.A(g12565),.B(g6314));
  NAND2 NAND2_375(.VSS(VSS),.VDD(VDD),.Y(g15822),.A(g12611),.B(g6369));
  NAND2 NAND2_376(.VSS(VSS),.VDD(VDD),.Y(g15823),.A(g12611),.B(g6519));
  NAND2 NAND2_377(.VSS(VSS),.VDD(VDD),.Y(g15824),.A(g12657),.B(g6574));
  NAND2 NAND2_378(.VSS(VSS),.VDD(VDD),.Y(g15825),.A(g12657),.B(g6783));
  NAND2 NAND2_379(.VSS(VSS),.VDD(VDD),.Y(g15826),.A(g12711),.B(g6838));
  NAND2 NAND2_380(.VSS(VSS),.VDD(VDD),.Y(g15827),.A(g12711),.B(g7085));
  NAND2 NAND2_381(.VSS(VSS),.VDD(VDD),.Y(g15830),.A(g13310),.B(g12392));
  NAND2 NAND2_382(.VSS(VSS),.VDD(VDD),.Y(g15831),.A(g13313),.B(g12392));
  NAND2 NAND2_383(.VSS(VSS),.VDD(VDD),.Y(g15832),.A(g12565),.B(g6232));
  NAND2 NAND2_384(.VSS(VSS),.VDD(VDD),.Y(g15833),.A(g12565),.B(g6314));
  NAND2 NAND2_385(.VSS(VSS),.VDD(VDD),.Y(g15834),.A(g12611),.B(g6369));
  NAND2 NAND2_386(.VSS(VSS),.VDD(VDD),.Y(g15835),.A(g12611),.B(g6519));
  NAND2 NAND2_387(.VSS(VSS),.VDD(VDD),.Y(g15836),.A(g12657),.B(g6574));
  NAND2 NAND2_388(.VSS(VSS),.VDD(VDD),.Y(g15837),.A(g12657),.B(g6783));
  NAND2 NAND2_389(.VSS(VSS),.VDD(VDD),.Y(g15838),.A(g12711),.B(g6838));
  NAND2 NAND2_390(.VSS(VSS),.VDD(VDD),.Y(g15839),.A(g12711),.B(g7085));
  NAND2 NAND2_391(.VSS(VSS),.VDD(VDD),.Y(g15841),.A(g13331),.B(g12392));
  NAND2 NAND2_392(.VSS(VSS),.VDD(VDD),.Y(g15842),.A(g13332),.B(g12392));
  NAND2 NAND2_393(.VSS(VSS),.VDD(VDD),.Y(g15843),.A(g12565),.B(g6314));
  NAND2 NAND2_394(.VSS(VSS),.VDD(VDD),.Y(g15844),.A(g12565),.B(g6232));
  NAND2 NAND2_395(.VSS(VSS),.VDD(VDD),.Y(g15845),.A(g12565),.B(g6314));
  NAND2 NAND2_396(.VSS(VSS),.VDD(VDD),.Y(g15846),.A(g12611),.B(g6369));
  NAND2 NAND2_397(.VSS(VSS),.VDD(VDD),.Y(g15847),.A(g12611),.B(g6519));
  NAND2 NAND2_398(.VSS(VSS),.VDD(VDD),.Y(g15848),.A(g12657),.B(g6574));
  NAND2 NAND2_399(.VSS(VSS),.VDD(VDD),.Y(g15849),.A(g12657),.B(g6783));
  NAND2 NAND2_400(.VSS(VSS),.VDD(VDD),.Y(g15850),.A(g12711),.B(g6838));
  NAND2 NAND2_401(.VSS(VSS),.VDD(VDD),.Y(g15851),.A(g12711),.B(g7085));
  NAND2 NAND2_402(.VSS(VSS),.VDD(VDD),.Y(g15853),.A(g13310),.B(g12354));
  NAND2 NAND2_403(.VSS(VSS),.VDD(VDD),.Y(g15854),.A(g13353),.B(g12392));
  NAND2 NAND2_404(.VSS(VSS),.VDD(VDD),.Y(g15855),.A(g13354),.B(g12392));
  NAND2 NAND2_405(.VSS(VSS),.VDD(VDD),.Y(g15856),.A(g12565),.B(g6232));
  NAND2 NAND2_406(.VSS(VSS),.VDD(VDD),.Y(g15857),.A(g12565),.B(g6314));
  NAND2 NAND2_407(.VSS(VSS),.VDD(VDD),.Y(g15858),.A(g12565),.B(g6232));
  NAND2 NAND2_408(.VSS(VSS),.VDD(VDD),.Y(g15866),.A(g12611),.B(g6519));
  NAND2 NAND2_409(.VSS(VSS),.VDD(VDD),.Y(g15867),.A(g12611),.B(g6369));
  NAND2 NAND2_410(.VSS(VSS),.VDD(VDD),.Y(g15868),.A(g12611),.B(g6519));
  NAND2 NAND2_411(.VSS(VSS),.VDD(VDD),.Y(g15869),.A(g12657),.B(g6574));
  NAND2 NAND2_412(.VSS(VSS),.VDD(VDD),.Y(g15870),.A(g12657),.B(g6783));
  NAND2 NAND2_413(.VSS(VSS),.VDD(VDD),.Y(g15871),.A(g12711),.B(g6838));
  NAND2 NAND2_414(.VSS(VSS),.VDD(VDD),.Y(g15872),.A(g12711),.B(g7085));
  NAND2 NAND2_415(.VSS(VSS),.VDD(VDD),.Y(g15877),.A(g13374),.B(g12392));
  NAND2 NAND2_416(.VSS(VSS),.VDD(VDD),.Y(g15878),.A(g13375),.B(g12392));
  NAND2 NAND2_417(.VSS(VSS),.VDD(VDD),.Y(g15879),.A(g12565),.B(g6232));
  NAND2 NAND2_418(.VSS(VSS),.VDD(VDD),.Y(g15887),.A(g12611),.B(g6369));
  NAND2 NAND2_419(.VSS(VSS),.VDD(VDD),.Y(g15888),.A(g12611),.B(g6519));
  NAND2 NAND2_420(.VSS(VSS),.VDD(VDD),.Y(g15889),.A(g12611),.B(g6369));
  NAND2 NAND2_421(.VSS(VSS),.VDD(VDD),.Y(g15897),.A(g12657),.B(g6783));
  NAND2 NAND2_422(.VSS(VSS),.VDD(VDD),.Y(g15898),.A(g12657),.B(g6574));
  NAND2 NAND2_423(.VSS(VSS),.VDD(VDD),.Y(g15899),.A(g12657),.B(g6783));
  NAND2 NAND2_424(.VSS(VSS),.VDD(VDD),.Y(g15900),.A(g12711),.B(g6838));
  NAND2 NAND2_425(.VSS(VSS),.VDD(VDD),.Y(g15901),.A(g12711),.B(g7085));
  NAND2 NAND2_426(.VSS(VSS),.VDD(VDD),.Y(g15903),.A(g13404),.B(g12392));
  NAND2 NAND2_427(.VSS(VSS),.VDD(VDD),.Y(g15912),.A(g12611),.B(g6369));
  NAND2 NAND2_428(.VSS(VSS),.VDD(VDD),.Y(g15920),.A(g12657),.B(g6574));
  NAND2 NAND2_429(.VSS(VSS),.VDD(VDD),.Y(g15921),.A(g12657),.B(g6783));
  NAND2 NAND2_430(.VSS(VSS),.VDD(VDD),.Y(g15922),.A(g12657),.B(g6574));
  NAND2 NAND2_431(.VSS(VSS),.VDD(VDD),.Y(g15930),.A(g12711),.B(g7085));
  NAND2 NAND2_432(.VSS(VSS),.VDD(VDD),.Y(g15931),.A(g12711),.B(g6838));
  NAND2 NAND2_433(.VSS(VSS),.VDD(VDD),.Y(g15932),.A(g12711),.B(g7085));
  NAND2 NAND2_434(.VSS(VSS),.VDD(VDD),.Y(g15941),.A(g12657),.B(g6574));
  NAND2 NAND2_435(.VSS(VSS),.VDD(VDD),.Y(g15949),.A(g12711),.B(g6838));
  NAND2 NAND2_436(.VSS(VSS),.VDD(VDD),.Y(g15950),.A(g12711),.B(g7085));
  NAND2 NAND2_437(.VSS(VSS),.VDD(VDD),.Y(g15951),.A(g12711),.B(g6838));
  NAND2 NAND2_438(.VSS(VSS),.VDD(VDD),.Y(g15970),.A(g12711),.B(g6838));
  NAND2 NAND2_439(.VSS(VSS),.VDD(VDD),.Y(g15990),.A(g12886),.B(g6912));
  NAND2 NAND2_440(.VSS(VSS),.VDD(VDD),.Y(g15992),.A(g12886),.B(g6678));
  NAND2 NAND2_441(.VSS(VSS),.VDD(VDD),.Y(g15993),.A(g12926),.B(g7162));
  NAND2 NAND2_442(.VSS(VSS),.VDD(VDD),.Y(g15995),.A(g12926),.B(g6980));
  NAND2 NAND2_443(.VSS(VSS),.VDD(VDD),.Y(g15996),.A(g12955),.B(g7358));
  NAND2 NAND2_444(.VSS(VSS),.VDD(VDD),.Y(g15999),.A(g12955),.B(g7230));
  NAND2 NAND2_445(.VSS(VSS),.VDD(VDD),.Y(g16000),.A(g12984),.B(g7488));
  NAND2 NAND2_446(.VSS(VSS),.VDD(VDD),.Y(g16006),.A(g12984),.B(g7426));
  NAND2 NAND2_447(.VSS(VSS),.VDD(VDD),.Y(g16085),.A(g12883),.B(g633));
  NAND2 NAND2_448(.VSS(VSS),.VDD(VDD),.Y(g16123),.A(g12923),.B(g1319));
  NAND2 NAND2_449(.VSS(VSS),.VDD(VDD),.Y(I22282),.A(g2962),.B(g13348));
  NAND2 NAND2_450(.VSS(VSS),.VDD(VDD),.Y(I22283),.A(g2962),.B(I22282));
  NAND2 NAND2_451(.VSS(VSS),.VDD(VDD),.Y(I22284),.A(g13348),.B(I22282));
  NAND2 NAND2_452(.VSS(VSS),.VDD(VDD),.Y(g16132),.A(I22283),.B(I22284));
  NAND2 NAND2_453(.VSS(VSS),.VDD(VDD),.Y(g16174),.A(g12952),.B(g2013));
  NAND2 NAND2_454(.VSS(VSS),.VDD(VDD),.Y(I22316),.A(g2934),.B(g13370));
  NAND2 NAND2_455(.VSS(VSS),.VDD(VDD),.Y(I22317),.A(g2934),.B(I22316));
  NAND2 NAND2_456(.VSS(VSS),.VDD(VDD),.Y(I22318),.A(g13370),.B(I22316));
  NAND2 NAND2_457(.VSS(VSS),.VDD(VDD),.Y(g16181),.A(I22317),.B(I22318));
  NAND2 NAND2_458(.VSS(VSS),.VDD(VDD),.Y(g16233),.A(g12981),.B(g2707));
  NAND2 NAND2_459(.VSS(VSS),.VDD(VDD),.Y(g16341),.A(g12377),.B(g12407));
  NAND2 NAND2_460(.VSS(VSS),.VDD(VDD),.Y(g16412),.A(g12565),.B(g3254));
  NAND2 NAND2_461(.VSS(VSS),.VDD(VDD),.Y(g16439),.A(g13082),.B(g2912));
  NAND2 NAND2_462(.VSS(VSS),.VDD(VDD),.Y(g16442),.A(g12565),.B(g3254));
  NAND2 NAND2_463(.VSS(VSS),.VDD(VDD),.Y(g16446),.A(g12611),.B(g3410));
  NAND2 NAND2_464(.VSS(VSS),.VDD(VDD),.Y(g16463),.A(g13004),.B(g3018));
  NAND2 NAND2_465(.VSS(VSS),.VDD(VDD),.Y(g16536),.A(g15873),.B(g2896));
  NAND2 NAND2_466(.VSS(VSS),.VDD(VDD),.Y(I22630),.A(g13507),.B(g15978));
  NAND2 NAND2_467(.VSS(VSS),.VDD(VDD),.Y(I22631),.A(g13507),.B(I22630));
  NAND2 NAND2_468(.VSS(VSS),.VDD(VDD),.Y(I22632),.A(g15978),.B(I22630));
  NAND2 NAND2_469(.VSS(VSS),.VDD(VDD),.Y(g16566),.A(I22631),.B(I22632));
  NAND2 NAND2_470(.VSS(VSS),.VDD(VDD),.Y(I22705),.A(g13348),.B(g15661));
  NAND2 NAND2_471(.VSS(VSS),.VDD(VDD),.Y(I22706),.A(g13348),.B(I22705));
  NAND2 NAND2_472(.VSS(VSS),.VDD(VDD),.Y(I22707),.A(g15661),.B(I22705));
  NAND2 NAND2_473(.VSS(VSS),.VDD(VDD),.Y(g16662),.A(I22706),.B(I22707));
  NAND2 NAND2_474(.VSS(VSS),.VDD(VDD),.Y(I22884),.A(g13370),.B(g15661));
  NAND2 NAND2_475(.VSS(VSS),.VDD(VDD),.Y(I22885),.A(g13370),.B(I22884));
  NAND2 NAND2_476(.VSS(VSS),.VDD(VDD),.Y(I22886),.A(g15661),.B(I22884));
  NAND2 NAND2_477(.VSS(VSS),.VDD(VDD),.Y(g16935),.A(I22885),.B(I22886));
  NAND2 NAND2_478(.VSS(VSS),.VDD(VDD),.Y(I22900),.A(g15022),.B(g14000));
  NAND2 NAND2_479(.VSS(VSS),.VDD(VDD),.Y(I22901),.A(g15022),.B(I22900));
  NAND2 NAND2_480(.VSS(VSS),.VDD(VDD),.Y(I22902),.A(g14000),.B(I22900));
  NAND2 NAND2_481(.VSS(VSS),.VDD(VDD),.Y(g16965),.A(I22901),.B(I22902));
  NAND2 NAND2_482(.VSS(VSS),.VDD(VDD),.Y(I22917),.A(g15096),.B(g13945));
  NAND2 NAND2_483(.VSS(VSS),.VDD(VDD),.Y(I22918),.A(g15096),.B(I22917));
  NAND2 NAND2_484(.VSS(VSS),.VDD(VDD),.Y(I22919),.A(g13945),.B(I22917));
  NAND2 NAND2_485(.VSS(VSS),.VDD(VDD),.Y(g16985),.A(I22918),.B(I22919));
  NAND2 NAND2_486(.VSS(VSS),.VDD(VDD),.Y(I22924),.A(g15118),.B(g14091));
  NAND2 NAND2_487(.VSS(VSS),.VDD(VDD),.Y(I22925),.A(g15118),.B(I22924));
  NAND2 NAND2_488(.VSS(VSS),.VDD(VDD),.Y(I22926),.A(g14091),.B(I22924));
  NAND2 NAND2_489(.VSS(VSS),.VDD(VDD),.Y(g16986),.A(I22925),.B(I22926));
  NAND2 NAND2_490(.VSS(VSS),.VDD(VDD),.Y(I22936),.A(g9150),.B(g13906));
  NAND2 NAND2_491(.VSS(VSS),.VDD(VDD),.Y(I22937),.A(g9150),.B(I22936));
  NAND2 NAND2_492(.VSS(VSS),.VDD(VDD),.Y(I22938),.A(g13906),.B(I22936));
  NAND2 NAND2_493(.VSS(VSS),.VDD(VDD),.Y(g16992),.A(I22937),.B(I22938));
  NAND2 NAND2_494(.VSS(VSS),.VDD(VDD),.Y(I22945),.A(g15188),.B(g14015));
  NAND2 NAND2_495(.VSS(VSS),.VDD(VDD),.Y(I22946),.A(g15188),.B(I22945));
  NAND2 NAND2_496(.VSS(VSS),.VDD(VDD),.Y(I22947),.A(g14015),.B(I22945));
  NAND2 NAND2_497(.VSS(VSS),.VDD(VDD),.Y(g16995),.A(I22946),.B(I22947));
  NAND2 NAND2_498(.VSS(VSS),.VDD(VDD),.Y(I22952),.A(g15210),.B(g14206));
  NAND2 NAND2_499(.VSS(VSS),.VDD(VDD),.Y(I22953),.A(g15210),.B(I22952));
  NAND2 NAND2_500(.VSS(VSS),.VDD(VDD),.Y(I22954),.A(g14206),.B(I22952));
  NAND2 NAND2_501(.VSS(VSS),.VDD(VDD),.Y(g16996),.A(I22953),.B(I22954));
  NAND2 NAND2_502(.VSS(VSS),.VDD(VDD),.Y(I22962),.A(g9161),.B(g13885));
  NAND2 NAND2_503(.VSS(VSS),.VDD(VDD),.Y(I22963),.A(g9161),.B(I22962));
  NAND2 NAND2_504(.VSS(VSS),.VDD(VDD),.Y(I22964),.A(g13885),.B(I22962));
  NAND2 NAND2_505(.VSS(VSS),.VDD(VDD),.Y(g17000),.A(I22963),.B(I22964));
  NAND2 NAND2_506(.VSS(VSS),.VDD(VDD),.Y(I22972),.A(g9174),.B(g13962));
  NAND2 NAND2_507(.VSS(VSS),.VDD(VDD),.Y(I22973),.A(g9174),.B(I22972));
  NAND2 NAND2_508(.VSS(VSS),.VDD(VDD),.Y(I22974),.A(g13962),.B(I22972));
  NAND2 NAND2_509(.VSS(VSS),.VDD(VDD),.Y(g17016),.A(I22973),.B(I22974));
  NAND2 NAND2_510(.VSS(VSS),.VDD(VDD),.Y(I22981),.A(g15274),.B(g14106));
  NAND2 NAND2_511(.VSS(VSS),.VDD(VDD),.Y(I22982),.A(g15274),.B(I22981));
  NAND2 NAND2_512(.VSS(VSS),.VDD(VDD),.Y(I22983),.A(g14106),.B(I22981));
  NAND2 NAND2_513(.VSS(VSS),.VDD(VDD),.Y(g17019),.A(I22982),.B(I22983));
  NAND2 NAND2_514(.VSS(VSS),.VDD(VDD),.Y(I22988),.A(g15296),.B(g14321));
  NAND2 NAND2_515(.VSS(VSS),.VDD(VDD),.Y(I22989),.A(g15296),.B(I22988));
  NAND2 NAND2_516(.VSS(VSS),.VDD(VDD),.Y(I22990),.A(g14321),.B(I22988));
  NAND2 NAND2_517(.VSS(VSS),.VDD(VDD),.Y(g17020),.A(I22989),.B(I22990));
  NAND2 NAND2_518(.VSS(VSS),.VDD(VDD),.Y(I22998),.A(g9187),.B(g13872));
  NAND2 NAND2_519(.VSS(VSS),.VDD(VDD),.Y(I22999),.A(g9187),.B(I22998));
  NAND2 NAND2_520(.VSS(VSS),.VDD(VDD),.Y(I23000),.A(g13872),.B(I22998));
  NAND2 NAND2_521(.VSS(VSS),.VDD(VDD),.Y(g17024),.A(I22999),.B(I23000));
  NAND2 NAND2_522(.VSS(VSS),.VDD(VDD),.Y(I23008),.A(g9203),.B(g13926));
  NAND2 NAND2_523(.VSS(VSS),.VDD(VDD),.Y(I23009),.A(g9203),.B(I23008));
  NAND2 NAND2_524(.VSS(VSS),.VDD(VDD),.Y(I23010),.A(g13926),.B(I23008));
  NAND2 NAND2_525(.VSS(VSS),.VDD(VDD),.Y(g17030),.A(I23009),.B(I23010));
  NAND2 NAND2_526(.VSS(VSS),.VDD(VDD),.Y(I23018),.A(g9216),.B(g14032));
  NAND2 NAND2_527(.VSS(VSS),.VDD(VDD),.Y(I23019),.A(g9216),.B(I23018));
  NAND2 NAND2_528(.VSS(VSS),.VDD(VDD),.Y(I23020),.A(g14032),.B(I23018));
  NAND2 NAND2_529(.VSS(VSS),.VDD(VDD),.Y(g17046),.A(I23019),.B(I23020));
  NAND2 NAND2_530(.VSS(VSS),.VDD(VDD),.Y(I23027),.A(g15366),.B(g14221));
  NAND2 NAND2_531(.VSS(VSS),.VDD(VDD),.Y(I23028),.A(g15366),.B(I23027));
  NAND2 NAND2_532(.VSS(VSS),.VDD(VDD),.Y(I23029),.A(g14221),.B(I23027));
  NAND2 NAND2_533(.VSS(VSS),.VDD(VDD),.Y(g17049),.A(I23028),.B(I23029));
  NAND2 NAND2_534(.VSS(VSS),.VDD(VDD),.Y(I23034),.A(g9232),.B(g13864));
  NAND2 NAND2_535(.VSS(VSS),.VDD(VDD),.Y(I23035),.A(g9232),.B(I23034));
  NAND2 NAND2_536(.VSS(VSS),.VDD(VDD),.Y(I23036),.A(g13864),.B(I23034));
  NAND2 NAND2_537(.VSS(VSS),.VDD(VDD),.Y(g17050),.A(I23035),.B(I23036));
  NAND2 NAND2_538(.VSS(VSS),.VDD(VDD),.Y(I23045),.A(g9248),.B(g13894));
  NAND2 NAND2_539(.VSS(VSS),.VDD(VDD),.Y(I23046),.A(g9248),.B(I23045));
  NAND2 NAND2_540(.VSS(VSS),.VDD(VDD),.Y(I23047),.A(g13894),.B(I23045));
  NAND2 NAND2_541(.VSS(VSS),.VDD(VDD),.Y(g17058),.A(I23046),.B(I23047));
  NAND2 NAND2_542(.VSS(VSS),.VDD(VDD),.Y(I23055),.A(g9264),.B(g13982));
  NAND2 NAND2_543(.VSS(VSS),.VDD(VDD),.Y(I23056),.A(g9264),.B(I23055));
  NAND2 NAND2_544(.VSS(VSS),.VDD(VDD),.Y(I23057),.A(g13982),.B(I23055));
  NAND2 NAND2_545(.VSS(VSS),.VDD(VDD),.Y(g17064),.A(I23056),.B(I23057));
  NAND2 NAND2_546(.VSS(VSS),.VDD(VDD),.Y(I23065),.A(g9277),.B(g14123));
  NAND2 NAND2_547(.VSS(VSS),.VDD(VDD),.Y(I23066),.A(g9277),.B(I23065));
  NAND2 NAND2_548(.VSS(VSS),.VDD(VDD),.Y(I23067),.A(g14123),.B(I23065));
  NAND2 NAND2_549(.VSS(VSS),.VDD(VDD),.Y(g17080),.A(I23066),.B(I23067));
  NAND2 NAND2_550(.VSS(VSS),.VDD(VDD),.Y(I23074),.A(g9293),.B(g13856));
  NAND2 NAND2_551(.VSS(VSS),.VDD(VDD),.Y(I23075),.A(g9293),.B(I23074));
  NAND2 NAND2_552(.VSS(VSS),.VDD(VDD),.Y(I23076),.A(g13856),.B(I23074));
  NAND2 NAND2_553(.VSS(VSS),.VDD(VDD),.Y(g17083),.A(I23075),.B(I23076));
  NAND2 NAND2_554(.VSS(VSS),.VDD(VDD),.Y(I23082),.A(g9310),.B(g13879));
  NAND2 NAND2_555(.VSS(VSS),.VDD(VDD),.Y(I23083),.A(g9310),.B(I23082));
  NAND2 NAND2_556(.VSS(VSS),.VDD(VDD),.Y(I23084),.A(g13879),.B(I23082));
  NAND2 NAND2_557(.VSS(VSS),.VDD(VDD),.Y(g17085),.A(I23083),.B(I23084));
  NAND2 NAND2_558(.VSS(VSS),.VDD(VDD),.Y(I23093),.A(g9326),.B(g13935));
  NAND2 NAND2_559(.VSS(VSS),.VDD(VDD),.Y(I23094),.A(g9326),.B(I23093));
  NAND2 NAND2_560(.VSS(VSS),.VDD(VDD),.Y(I23095),.A(g13935),.B(I23093));
  NAND2 NAND2_561(.VSS(VSS),.VDD(VDD),.Y(g17093),.A(I23094),.B(I23095));
  NAND2 NAND2_562(.VSS(VSS),.VDD(VDD),.Y(I23103),.A(g9342),.B(g14052));
  NAND2 NAND2_563(.VSS(VSS),.VDD(VDD),.Y(I23104),.A(g9342),.B(I23103));
  NAND2 NAND2_564(.VSS(VSS),.VDD(VDD),.Y(I23105),.A(g14052),.B(I23103));
  NAND2 NAND2_565(.VSS(VSS),.VDD(VDD),.Y(g17099),.A(I23104),.B(I23105));
  NAND2 NAND2_566(.VSS(VSS),.VDD(VDD),.Y(I23113),.A(g9356),.B(g13848));
  NAND2 NAND2_567(.VSS(VSS),.VDD(VDD),.Y(I23114),.A(g9356),.B(I23113));
  NAND2 NAND2_568(.VSS(VSS),.VDD(VDD),.Y(I23115),.A(g13848),.B(I23113));
  NAND2 NAND2_569(.VSS(VSS),.VDD(VDD),.Y(g17115),.A(I23114),.B(I23115));
  NAND2 NAND2_570(.VSS(VSS),.VDD(VDD),.Y(g17118),.A(g13915),.B(g13893));
  NAND2 NAND2_571(.VSS(VSS),.VDD(VDD),.Y(I23123),.A(g9374),.B(g13866));
  NAND2 NAND2_572(.VSS(VSS),.VDD(VDD),.Y(I23124),.A(g9374),.B(I23123));
  NAND2 NAND2_573(.VSS(VSS),.VDD(VDD),.Y(I23125),.A(g13866),.B(I23123));
  NAND2 NAND2_574(.VSS(VSS),.VDD(VDD),.Y(g17121),.A(I23124),.B(I23125));
  NAND2 NAND2_575(.VSS(VSS),.VDD(VDD),.Y(I23131),.A(g9391),.B(g13901));
  NAND2 NAND2_576(.VSS(VSS),.VDD(VDD),.Y(I23132),.A(g9391),.B(I23131));
  NAND2 NAND2_577(.VSS(VSS),.VDD(VDD),.Y(I23133),.A(g13901),.B(I23131));
  NAND2 NAND2_578(.VSS(VSS),.VDD(VDD),.Y(g17123),.A(I23132),.B(I23133));
  NAND2 NAND2_579(.VSS(VSS),.VDD(VDD),.Y(I23142),.A(g9407),.B(g13991));
  NAND2 NAND2_580(.VSS(VSS),.VDD(VDD),.Y(I23143),.A(g9407),.B(I23142));
  NAND2 NAND2_581(.VSS(VSS),.VDD(VDD),.Y(I23144),.A(g13991),.B(I23142));
  NAND2 NAND2_582(.VSS(VSS),.VDD(VDD),.Y(g17131),.A(I23143),.B(I23144));
  NAND2 NAND2_583(.VSS(VSS),.VDD(VDD),.Y(I23152),.A(g9427),.B(g14061));
  NAND2 NAND2_584(.VSS(VSS),.VDD(VDD),.Y(I23153),.A(g9427),.B(I23152));
  NAND2 NAND2_585(.VSS(VSS),.VDD(VDD),.Y(I23154),.A(g14061),.B(I23152));
  NAND2 NAND2_586(.VSS(VSS),.VDD(VDD),.Y(g17137),.A(I23153),.B(I23154));
  NAND2 NAND2_587(.VSS(VSS),.VDD(VDD),.Y(g17139),.A(g13957),.B(g13915));
  NAND2 NAND2_588(.VSS(VSS),.VDD(VDD),.Y(I23161),.A(g9453),.B(g13857));
  NAND2 NAND2_589(.VSS(VSS),.VDD(VDD),.Y(I23162),.A(g9453),.B(I23161));
  NAND2 NAND2_590(.VSS(VSS),.VDD(VDD),.Y(I23163),.A(g13857),.B(I23161));
  NAND2 NAND2_591(.VSS(VSS),.VDD(VDD),.Y(g17142),.A(I23162),.B(I23163));
  NAND2 NAND2_592(.VSS(VSS),.VDD(VDD),.Y(g17145),.A(g13971),.B(g13934));
  NAND2 NAND2_593(.VSS(VSS),.VDD(VDD),.Y(I23171),.A(g9471),.B(g13881));
  NAND2 NAND2_594(.VSS(VSS),.VDD(VDD),.Y(I23172),.A(g9471),.B(I23171));
  NAND2 NAND2_595(.VSS(VSS),.VDD(VDD),.Y(I23173),.A(g13881),.B(I23171));
  NAND2 NAND2_596(.VSS(VSS),.VDD(VDD),.Y(g17148),.A(I23172),.B(I23173));
  NAND2 NAND2_597(.VSS(VSS),.VDD(VDD),.Y(I23179),.A(g9488),.B(g13942));
  NAND2 NAND2_598(.VSS(VSS),.VDD(VDD),.Y(I23180),.A(g9488),.B(I23179));
  NAND2 NAND2_599(.VSS(VSS),.VDD(VDD),.Y(I23181),.A(g13942),.B(I23179));
  NAND2 NAND2_600(.VSS(VSS),.VDD(VDD),.Y(g17150),.A(I23180),.B(I23181));
  NAND2 NAND2_601(.VSS(VSS),.VDD(VDD),.Y(I23190),.A(g9507),.B(g13999));
  NAND2 NAND2_602(.VSS(VSS),.VDD(VDD),.Y(I23191),.A(g9507),.B(I23190));
  NAND2 NAND2_603(.VSS(VSS),.VDD(VDD),.Y(I23192),.A(g13999),.B(I23190));
  NAND2 NAND2_604(.VSS(VSS),.VDD(VDD),.Y(g17158),.A(I23191),.B(I23192));
  NAND2 NAND2_605(.VSS(VSS),.VDD(VDD),.Y(g17159),.A(g14642),.B(g14657));
  NAND2 NAND2_606(.VSS(VSS),.VDD(VDD),.Y(I23198),.A(g9569),.B(g14176));
  NAND2 NAND2_607(.VSS(VSS),.VDD(VDD),.Y(I23199),.A(g9569),.B(I23198));
  NAND2 NAND2_608(.VSS(VSS),.VDD(VDD),.Y(I23200),.A(g14176),.B(I23198));
  NAND2 NAND2_609(.VSS(VSS),.VDD(VDD),.Y(g17160),.A(I23199),.B(I23200));
  NAND2 NAND2_610(.VSS(VSS),.VDD(VDD),.Y(g17162),.A(g14027),.B(g13971));
  NAND2 NAND2_611(.VSS(VSS),.VDD(VDD),.Y(I23207),.A(g9595),.B(g13867));
  NAND2 NAND2_612(.VSS(VSS),.VDD(VDD),.Y(I23208),.A(g9595),.B(I23207));
  NAND2 NAND2_613(.VSS(VSS),.VDD(VDD),.Y(I23209),.A(g13867),.B(I23207));
  NAND2 NAND2_614(.VSS(VSS),.VDD(VDD),.Y(g17165),.A(I23208),.B(I23209));
  NAND2 NAND2_615(.VSS(VSS),.VDD(VDD),.Y(g17168),.A(g14041),.B(g13990));
  NAND2 NAND2_616(.VSS(VSS),.VDD(VDD),.Y(I23217),.A(g9613),.B(g13903));
  NAND2 NAND2_617(.VSS(VSS),.VDD(VDD),.Y(I23218),.A(g9613),.B(I23217));
  NAND2 NAND2_618(.VSS(VSS),.VDD(VDD),.Y(I23219),.A(g13903),.B(I23217));
  NAND2 NAND2_619(.VSS(VSS),.VDD(VDD),.Y(g17171),.A(I23218),.B(I23219));
  NAND2 NAND2_620(.VSS(VSS),.VDD(VDD),.Y(I23225),.A(g9649),.B(g14090));
  NAND2 NAND2_621(.VSS(VSS),.VDD(VDD),.Y(I23226),.A(g9649),.B(I23225));
  NAND2 NAND2_622(.VSS(VSS),.VDD(VDD),.Y(I23227),.A(g14090),.B(I23225));
  NAND2 NAND2_623(.VSS(VSS),.VDD(VDD),.Y(g17173),.A(I23226),.B(I23227));
  NAND2 NAND2_624(.VSS(VSS),.VDD(VDD),.Y(g17174),.A(g14669),.B(g14691));
  NAND2 NAND2_625(.VSS(VSS),.VDD(VDD),.Y(I23233),.A(g9711),.B(g14291));
  NAND2 NAND2_626(.VSS(VSS),.VDD(VDD),.Y(I23234),.A(g9711),.B(I23233));
  NAND2 NAND2_627(.VSS(VSS),.VDD(VDD),.Y(I23235),.A(g14291),.B(I23233));
  NAND2 NAND2_628(.VSS(VSS),.VDD(VDD),.Y(g17175),.A(I23234),.B(I23235));
  NAND2 NAND2_629(.VSS(VSS),.VDD(VDD),.Y(g17177),.A(g14118),.B(g14041));
  NAND2 NAND2_630(.VSS(VSS),.VDD(VDD),.Y(I23242),.A(g9737),.B(g13882));
  NAND2 NAND2_631(.VSS(VSS),.VDD(VDD),.Y(I23243),.A(g9737),.B(I23242));
  NAND2 NAND2_632(.VSS(VSS),.VDD(VDD),.Y(I23244),.A(g13882),.B(I23242));
  NAND2 NAND2_633(.VSS(VSS),.VDD(VDD),.Y(g17180),.A(I23243),.B(I23244));
  NAND2 NAND2_634(.VSS(VSS),.VDD(VDD),.Y(g17183),.A(g14132),.B(g14060));
  NAND2 NAND2_635(.VSS(VSS),.VDD(VDD),.Y(I23256),.A(g9795),.B(g14205));
  NAND2 NAND2_636(.VSS(VSS),.VDD(VDD),.Y(I23257),.A(g9795),.B(I23256));
  NAND2 NAND2_637(.VSS(VSS),.VDD(VDD),.Y(I23258),.A(g14205),.B(I23256));
  NAND2 NAND2_638(.VSS(VSS),.VDD(VDD),.Y(g17190),.A(I23257),.B(I23258));
  NAND2 NAND2_639(.VSS(VSS),.VDD(VDD),.Y(g17191),.A(g14703),.B(g14725));
  NAND2 NAND2_640(.VSS(VSS),.VDD(VDD),.Y(I23264),.A(g9857),.B(g14413));
  NAND2 NAND2_641(.VSS(VSS),.VDD(VDD),.Y(I23265),.A(g9857),.B(I23264));
  NAND2 NAND2_642(.VSS(VSS),.VDD(VDD),.Y(I23266),.A(g14413),.B(I23264));
  NAND2 NAND2_643(.VSS(VSS),.VDD(VDD),.Y(g17192),.A(I23265),.B(I23266));
  NAND2 NAND2_644(.VSS(VSS),.VDD(VDD),.Y(g17194),.A(g14233),.B(g14132));
  NAND2 NAND2_645(.VSS(VSS),.VDD(VDD),.Y(I23277),.A(g9941),.B(g14320));
  NAND2 NAND2_646(.VSS(VSS),.VDD(VDD),.Y(I23278),.A(g9941),.B(I23277));
  NAND2 NAND2_647(.VSS(VSS),.VDD(VDD),.Y(I23279),.A(g14320),.B(I23277));
  NAND2 NAND2_648(.VSS(VSS),.VDD(VDD),.Y(g17201),.A(I23278),.B(I23279));
  NAND2 NAND2_649(.VSS(VSS),.VDD(VDD),.Y(g17202),.A(g14737),.B(g14753));
  NAND2 NAND2_650(.VSS(VSS),.VDD(VDD),.Y(I23806),.A(g14062),.B(g9150));
  NAND2 NAND2_651(.VSS(VSS),.VDD(VDD),.Y(I23807),.A(g14062),.B(I23806));
  NAND2 NAND2_652(.VSS(VSS),.VDD(VDD),.Y(I23808),.A(g9150),.B(I23806));
  NAND2 NAND2_653(.VSS(VSS),.VDD(VDD),.Y(g17729),.A(I23807),.B(I23808));
  NAND2 NAND2_654(.VSS(VSS),.VDD(VDD),.Y(I23878),.A(g14001),.B(g9187));
  NAND2 NAND2_655(.VSS(VSS),.VDD(VDD),.Y(I23879),.A(g14001),.B(I23878));
  NAND2 NAND2_656(.VSS(VSS),.VDD(VDD),.Y(I23880),.A(g9187),.B(I23878));
  NAND2 NAND2_657(.VSS(VSS),.VDD(VDD),.Y(g17807),.A(I23879),.B(I23880));
  NAND2 NAND2_658(.VSS(VSS),.VDD(VDD),.Y(I23893),.A(g14177),.B(g9174));
  NAND2 NAND2_659(.VSS(VSS),.VDD(VDD),.Y(I23894),.A(g14177),.B(I23893));
  NAND2 NAND2_660(.VSS(VSS),.VDD(VDD),.Y(I23895),.A(g9174),.B(I23893));
  NAND2 NAND2_661(.VSS(VSS),.VDD(VDD),.Y(g17830),.A(I23894),.B(I23895));
  NAND2 NAND2_662(.VSS(VSS),.VDD(VDD),.Y(I23941),.A(g13946),.B(g9293));
  NAND2 NAND2_663(.VSS(VSS),.VDD(VDD),.Y(I23942),.A(g13946),.B(I23941));
  NAND2 NAND2_664(.VSS(VSS),.VDD(VDD),.Y(I23943),.A(g9293),.B(I23941));
  NAND2 NAND2_665(.VSS(VSS),.VDD(VDD),.Y(g17887),.A(I23942),.B(I23943));
  NAND2 NAND2_666(.VSS(VSS),.VDD(VDD),.Y(I23958),.A(g6513),.B(g14171));
  NAND2 NAND2_667(.VSS(VSS),.VDD(VDD),.Y(I23959),.A(g6513),.B(I23958));
  NAND2 NAND2_668(.VSS(VSS),.VDD(VDD),.Y(I23960),.A(g14171),.B(I23958));
  NAND2 NAND2_669(.VSS(VSS),.VDD(VDD),.Y(g17913),.A(I23959),.B(I23960));
  NAND2 NAND2_670(.VSS(VSS),.VDD(VDD),.Y(I23966),.A(g14092),.B(g9248));
  NAND2 NAND2_671(.VSS(VSS),.VDD(VDD),.Y(I23967),.A(g14092),.B(I23966));
  NAND2 NAND2_672(.VSS(VSS),.VDD(VDD),.Y(I23968),.A(g9248),.B(I23966));
  NAND2 NAND2_673(.VSS(VSS),.VDD(VDD),.Y(g17919),.A(I23967),.B(I23968));
  NAND2 NAND2_674(.VSS(VSS),.VDD(VDD),.Y(I23981),.A(g14292),.B(g9216));
  NAND2 NAND2_675(.VSS(VSS),.VDD(VDD),.Y(I23982),.A(g14292),.B(I23981));
  NAND2 NAND2_676(.VSS(VSS),.VDD(VDD),.Y(I23983),.A(g9216),.B(I23981));
  NAND2 NAND2_677(.VSS(VSS),.VDD(VDD),.Y(g17942),.A(I23982),.B(I23983));
  NAND2 NAND2_678(.VSS(VSS),.VDD(VDD),.Y(I24005),.A(g7548),.B(g15814));
  NAND2 NAND2_679(.VSS(VSS),.VDD(VDD),.Y(I24006),.A(g7548),.B(I24005));
  NAND2 NAND2_680(.VSS(VSS),.VDD(VDD),.Y(I24007),.A(g15814),.B(I24005));
  NAND2 NAND2_681(.VSS(VSS),.VDD(VDD),.Y(g17968),.A(I24006),.B(I24007));
  NAND2 NAND2_682(.VSS(VSS),.VDD(VDD),.Y(I24015),.A(g13907),.B(g9427));
  NAND2 NAND2_683(.VSS(VSS),.VDD(VDD),.Y(I24016),.A(g13907),.B(I24015));
  NAND2 NAND2_684(.VSS(VSS),.VDD(VDD),.Y(I24017),.A(g9427),.B(I24015));
  NAND2 NAND2_685(.VSS(VSS),.VDD(VDD),.Y(g17979),.A(I24016),.B(I24017));
  NAND2 NAND2_686(.VSS(VSS),.VDD(VDD),.Y(g17985),.A(g14641),.B(g9636));
  NAND2 NAND2_687(.VSS(VSS),.VDD(VDD),.Y(I24028),.A(g6201),.B(g14086));
  NAND2 NAND2_688(.VSS(VSS),.VDD(VDD),.Y(I24029),.A(g6201),.B(I24028));
  NAND2 NAND2_689(.VSS(VSS),.VDD(VDD),.Y(I24030),.A(g14086),.B(I24028));
  NAND2 NAND2_690(.VSS(VSS),.VDD(VDD),.Y(g17992),.A(I24029),.B(I24030));
  NAND2 NAND2_691(.VSS(VSS),.VDD(VDD),.Y(I24036),.A(g14016),.B(g9374));
  NAND2 NAND2_692(.VSS(VSS),.VDD(VDD),.Y(I24037),.A(g14016),.B(I24036));
  NAND2 NAND2_693(.VSS(VSS),.VDD(VDD),.Y(I24038),.A(g9374),.B(I24036));
  NAND2 NAND2_694(.VSS(VSS),.VDD(VDD),.Y(g17998),.A(I24037),.B(I24038));
  NAND2 NAND2_695(.VSS(VSS),.VDD(VDD),.Y(I24053),.A(g6777),.B(g14286));
  NAND2 NAND2_696(.VSS(VSS),.VDD(VDD),.Y(I24054),.A(g6777),.B(I24053));
  NAND2 NAND2_697(.VSS(VSS),.VDD(VDD),.Y(I24055),.A(g14286),.B(I24053));
  NAND2 NAND2_698(.VSS(VSS),.VDD(VDD),.Y(g18024),.A(I24054),.B(I24055));
  NAND2 NAND2_699(.VSS(VSS),.VDD(VDD),.Y(I24061),.A(g14207),.B(g9326));
  NAND2 NAND2_700(.VSS(VSS),.VDD(VDD),.Y(I24062),.A(g14207),.B(I24061));
  NAND2 NAND2_701(.VSS(VSS),.VDD(VDD),.Y(I24063),.A(g9326),.B(I24061));
  NAND2 NAND2_702(.VSS(VSS),.VDD(VDD),.Y(g18030),.A(I24062),.B(I24063));
  NAND2 NAND2_703(.VSS(VSS),.VDD(VDD),.Y(I24076),.A(g14414),.B(g9277));
  NAND2 NAND2_704(.VSS(VSS),.VDD(VDD),.Y(I24077),.A(g14414),.B(I24076));
  NAND2 NAND2_705(.VSS(VSS),.VDD(VDD),.Y(I24078),.A(g9277),.B(I24076));
  NAND2 NAND2_706(.VSS(VSS),.VDD(VDD),.Y(g18053),.A(I24077),.B(I24078));
  NAND2 NAND2_707(.VSS(VSS),.VDD(VDD),.Y(I24091),.A(g13886),.B(g15096));
  NAND2 NAND2_708(.VSS(VSS),.VDD(VDD),.Y(I24092),.A(g13886),.B(I24091));
  NAND2 NAND2_709(.VSS(VSS),.VDD(VDD),.Y(I24093),.A(g15096),.B(I24091));
  NAND2 NAND2_710(.VSS(VSS),.VDD(VDD),.Y(g18079),.A(I24092),.B(I24093));
  NAND2 NAND2_711(.VSS(VSS),.VDD(VDD),.Y(I24102),.A(g6363),.B(g14011));
  NAND2 NAND2_712(.VSS(VSS),.VDD(VDD),.Y(I24103),.A(g6363),.B(I24102));
  NAND2 NAND2_713(.VSS(VSS),.VDD(VDD),.Y(I24104),.A(g14011),.B(I24102));
  NAND2 NAND2_714(.VSS(VSS),.VDD(VDD),.Y(g18090),.A(I24103),.B(I24104));
  NAND2 NAND2_715(.VSS(VSS),.VDD(VDD),.Y(I24110),.A(g13963),.B(g9569));
  NAND2 NAND2_716(.VSS(VSS),.VDD(VDD),.Y(I24111),.A(g13963),.B(I24110));
  NAND2 NAND2_717(.VSS(VSS),.VDD(VDD),.Y(I24112),.A(g9569),.B(I24110));
  NAND2 NAND2_718(.VSS(VSS),.VDD(VDD),.Y(g18096),.A(I24111),.B(I24112));
  NAND2 NAND2_719(.VSS(VSS),.VDD(VDD),.Y(g18102),.A(g14668),.B(g9782));
  NAND2 NAND2_720(.VSS(VSS),.VDD(VDD),.Y(I24123),.A(g6290),.B(g14201));
  NAND2 NAND2_721(.VSS(VSS),.VDD(VDD),.Y(I24124),.A(g6290),.B(I24123));
  NAND2 NAND2_722(.VSS(VSS),.VDD(VDD),.Y(I24125),.A(g14201),.B(I24123));
  NAND2 NAND2_723(.VSS(VSS),.VDD(VDD),.Y(g18109),.A(I24124),.B(I24125));
  NAND2 NAND2_724(.VSS(VSS),.VDD(VDD),.Y(I24131),.A(g14107),.B(g9471));
  NAND2 NAND2_725(.VSS(VSS),.VDD(VDD),.Y(I24132),.A(g14107),.B(I24131));
  NAND2 NAND2_726(.VSS(VSS),.VDD(VDD),.Y(I24133),.A(g9471),.B(I24131));
  NAND2 NAND2_727(.VSS(VSS),.VDD(VDD),.Y(g18115),.A(I24132),.B(I24133));
  NAND2 NAND2_728(.VSS(VSS),.VDD(VDD),.Y(I24148),.A(g7079),.B(g14408));
  NAND2 NAND2_729(.VSS(VSS),.VDD(VDD),.Y(I24149),.A(g7079),.B(I24148));
  NAND2 NAND2_730(.VSS(VSS),.VDD(VDD),.Y(I24150),.A(g14408),.B(I24148));
  NAND2 NAND2_731(.VSS(VSS),.VDD(VDD),.Y(g18141),.A(I24149),.B(I24150));
  NAND2 NAND2_732(.VSS(VSS),.VDD(VDD),.Y(I24156),.A(g14322),.B(g9407));
  NAND2 NAND2_733(.VSS(VSS),.VDD(VDD),.Y(I24157),.A(g14322),.B(I24156));
  NAND2 NAND2_734(.VSS(VSS),.VDD(VDD),.Y(I24158),.A(g9407),.B(I24156));
  NAND2 NAND2_735(.VSS(VSS),.VDD(VDD),.Y(g18147),.A(I24157),.B(I24158));
  NAND2 NAND2_736(.VSS(VSS),.VDD(VDD),.Y(I24178),.A(g13873),.B(g9161));
  NAND2 NAND2_737(.VSS(VSS),.VDD(VDD),.Y(I24179),.A(g13873),.B(I24178));
  NAND2 NAND2_738(.VSS(VSS),.VDD(VDD),.Y(I24180),.A(g9161),.B(I24178));
  NAND2 NAND2_739(.VSS(VSS),.VDD(VDD),.Y(g18183),.A(I24179),.B(I24180));
  NAND2 NAND2_740(.VSS(VSS),.VDD(VDD),.Y(I24186),.A(g6177),.B(g13958));
  NAND2 NAND2_741(.VSS(VSS),.VDD(VDD),.Y(I24187),.A(g6177),.B(I24186));
  NAND2 NAND2_742(.VSS(VSS),.VDD(VDD),.Y(I24188),.A(g13958),.B(I24186));
  NAND2 NAND2_743(.VSS(VSS),.VDD(VDD),.Y(g18189),.A(I24187),.B(I24188));
  NAND2 NAND2_744(.VSS(VSS),.VDD(VDD),.Y(I24194),.A(g13927),.B(g15188));
  NAND2 NAND2_745(.VSS(VSS),.VDD(VDD),.Y(I24195),.A(g13927),.B(I24194));
  NAND2 NAND2_746(.VSS(VSS),.VDD(VDD),.Y(I24196),.A(g15188),.B(I24194));
  NAND2 NAND2_747(.VSS(VSS),.VDD(VDD),.Y(g18195),.A(I24195),.B(I24196));
  NAND2 NAND2_748(.VSS(VSS),.VDD(VDD),.Y(I24205),.A(g6568),.B(g14102));
  NAND2 NAND2_749(.VSS(VSS),.VDD(VDD),.Y(I24206),.A(g6568),.B(I24205));
  NAND2 NAND2_750(.VSS(VSS),.VDD(VDD),.Y(I24207),.A(g14102),.B(I24205));
  NAND2 NAND2_751(.VSS(VSS),.VDD(VDD),.Y(g18206),.A(I24206),.B(I24207));
  NAND2 NAND2_752(.VSS(VSS),.VDD(VDD),.Y(I24213),.A(g14033),.B(g9711));
  NAND2 NAND2_753(.VSS(VSS),.VDD(VDD),.Y(I24214),.A(g14033),.B(I24213));
  NAND2 NAND2_754(.VSS(VSS),.VDD(VDD),.Y(I24215),.A(g9711),.B(I24213));
  NAND2 NAND2_755(.VSS(VSS),.VDD(VDD),.Y(g18212),.A(I24214),.B(I24215));
  NAND2 NAND2_756(.VSS(VSS),.VDD(VDD),.Y(g18218),.A(g14702),.B(g9928));
  NAND2 NAND2_757(.VSS(VSS),.VDD(VDD),.Y(I24226),.A(g6427),.B(g14316));
  NAND2 NAND2_758(.VSS(VSS),.VDD(VDD),.Y(I24227),.A(g6427),.B(I24226));
  NAND2 NAND2_759(.VSS(VSS),.VDD(VDD),.Y(I24228),.A(g14316),.B(I24226));
  NAND2 NAND2_760(.VSS(VSS),.VDD(VDD),.Y(g18225),.A(I24227),.B(I24228));
  NAND2 NAND2_761(.VSS(VSS),.VDD(VDD),.Y(I24234),.A(g14222),.B(g9613));
  NAND2 NAND2_762(.VSS(VSS),.VDD(VDD),.Y(I24235),.A(g14222),.B(I24234));
  NAND2 NAND2_763(.VSS(VSS),.VDD(VDD),.Y(I24236),.A(g9613),.B(I24234));
  NAND2 NAND2_764(.VSS(VSS),.VDD(VDD),.Y(g18231),.A(I24235),.B(I24236));
  NAND2 NAND2_765(.VSS(VSS),.VDD(VDD),.Y(I24251),.A(g7329),.B(g14520));
  NAND2 NAND2_766(.VSS(VSS),.VDD(VDD),.Y(I24252),.A(g7329),.B(I24251));
  NAND2 NAND2_767(.VSS(VSS),.VDD(VDD),.Y(I24253),.A(g14520),.B(I24251));
  NAND2 NAND2_768(.VSS(VSS),.VDD(VDD),.Y(g18257),.A(I24252),.B(I24253));
  NAND2 NAND2_769(.VSS(VSS),.VDD(VDD),.Y(I24263),.A(g14342),.B(g9232));
  NAND2 NAND2_770(.VSS(VSS),.VDD(VDD),.Y(I24264),.A(g14342),.B(I24263));
  NAND2 NAND2_771(.VSS(VSS),.VDD(VDD),.Y(I24265),.A(g9232),.B(I24263));
  NAND2 NAND2_772(.VSS(VSS),.VDD(VDD),.Y(g18270),.A(I24264),.B(I24265));
  NAND2 NAND2_773(.VSS(VSS),.VDD(VDD),.Y(I24271),.A(g6180),.B(g13922));
  NAND2 NAND2_774(.VSS(VSS),.VDD(VDD),.Y(I24272),.A(g6180),.B(I24271));
  NAND2 NAND2_775(.VSS(VSS),.VDD(VDD),.Y(I24273),.A(g13922),.B(I24271));
  NAND2 NAND2_776(.VSS(VSS),.VDD(VDD),.Y(g18276),.A(I24272),.B(I24273));
  NAND2 NAND2_777(.VSS(VSS),.VDD(VDD),.Y(I24278),.A(g6284),.B(g13918));
  NAND2 NAND2_778(.VSS(VSS),.VDD(VDD),.Y(I24279),.A(g6284),.B(I24278));
  NAND2 NAND2_779(.VSS(VSS),.VDD(VDD),.Y(I24280),.A(g13918),.B(I24278));
  NAND2 NAND2_780(.VSS(VSS),.VDD(VDD),.Y(g18277),.A(I24279),.B(I24280));
  NAND2 NAND2_781(.VSS(VSS),.VDD(VDD),.Y(I24290),.A(g13895),.B(g9203));
  NAND2 NAND2_782(.VSS(VSS),.VDD(VDD),.Y(I24291),.A(g13895),.B(I24290));
  NAND2 NAND2_783(.VSS(VSS),.VDD(VDD),.Y(I24292),.A(g9203),.B(I24290));
  NAND2 NAND2_784(.VSS(VSS),.VDD(VDD),.Y(g18290),.A(I24291),.B(I24292));
  NAND2 NAND2_785(.VSS(VSS),.VDD(VDD),.Y(I24298),.A(g6209),.B(g14028));
  NAND2 NAND2_786(.VSS(VSS),.VDD(VDD),.Y(I24299),.A(g6209),.B(I24298));
  NAND2 NAND2_787(.VSS(VSS),.VDD(VDD),.Y(I24300),.A(g14028),.B(I24298));
  NAND2 NAND2_788(.VSS(VSS),.VDD(VDD),.Y(g18296),.A(I24299),.B(I24300));
  NAND2 NAND2_789(.VSS(VSS),.VDD(VDD),.Y(I24306),.A(g13983),.B(g15274));
  NAND2 NAND2_790(.VSS(VSS),.VDD(VDD),.Y(I24307),.A(g13983),.B(I24306));
  NAND2 NAND2_791(.VSS(VSS),.VDD(VDD),.Y(I24308),.A(g15274),.B(I24306));
  NAND2 NAND2_792(.VSS(VSS),.VDD(VDD),.Y(g18302),.A(I24307),.B(I24308));
  NAND2 NAND2_793(.VSS(VSS),.VDD(VDD),.Y(I24317),.A(g6832),.B(g14217));
  NAND2 NAND2_794(.VSS(VSS),.VDD(VDD),.Y(I24318),.A(g6832),.B(I24317));
  NAND2 NAND2_795(.VSS(VSS),.VDD(VDD),.Y(I24319),.A(g14217),.B(I24317));
  NAND2 NAND2_796(.VSS(VSS),.VDD(VDD),.Y(g18313),.A(I24318),.B(I24319));
  NAND2 NAND2_797(.VSS(VSS),.VDD(VDD),.Y(I24325),.A(g14124),.B(g9857));
  NAND2 NAND2_798(.VSS(VSS),.VDD(VDD),.Y(I24326),.A(g14124),.B(I24325));
  NAND2 NAND2_799(.VSS(VSS),.VDD(VDD),.Y(I24327),.A(g9857),.B(I24325));
  NAND2 NAND2_800(.VSS(VSS),.VDD(VDD),.Y(g18319),.A(I24326),.B(I24327));
  NAND2 NAND2_801(.VSS(VSS),.VDD(VDD),.Y(g18325),.A(g14736),.B(g10082));
  NAND2 NAND2_802(.VSS(VSS),.VDD(VDD),.Y(I24338),.A(g6632),.B(g14438));
  NAND2 NAND2_803(.VSS(VSS),.VDD(VDD),.Y(I24339),.A(g6632),.B(I24338));
  NAND2 NAND2_804(.VSS(VSS),.VDD(VDD),.Y(I24340),.A(g14438),.B(I24338));
  NAND2 NAND2_805(.VSS(VSS),.VDD(VDD),.Y(g18332),.A(I24339),.B(I24340));
  NAND2 NAND2_806(.VSS(VSS),.VDD(VDD),.Y(I24351),.A(g14238),.B(g9356));
  NAND2 NAND2_807(.VSS(VSS),.VDD(VDD),.Y(I24352),.A(g14238),.B(I24351));
  NAND2 NAND2_808(.VSS(VSS),.VDD(VDD),.Y(I24353),.A(g9356),.B(I24351));
  NAND2 NAND2_809(.VSS(VSS),.VDD(VDD),.Y(g18346),.A(I24352),.B(I24353));
  NAND2 NAND2_810(.VSS(VSS),.VDD(VDD),.Y(I24361),.A(g6157),.B(g14525));
  NAND2 NAND2_811(.VSS(VSS),.VDD(VDD),.Y(I24362),.A(g6157),.B(I24361));
  NAND2 NAND2_812(.VSS(VSS),.VDD(VDD),.Y(I24363),.A(g14525),.B(I24361));
  NAND2 NAND2_813(.VSS(VSS),.VDD(VDD),.Y(g18354),.A(I24362),.B(I24363));
  NAND2 NAND2_814(.VSS(VSS),.VDD(VDD),.Y(I24372),.A(g14454),.B(g9310));
  NAND2 NAND2_815(.VSS(VSS),.VDD(VDD),.Y(I24373),.A(g14454),.B(I24372));
  NAND2 NAND2_816(.VSS(VSS),.VDD(VDD),.Y(I24374),.A(g9310),.B(I24372));
  NAND2 NAND2_817(.VSS(VSS),.VDD(VDD),.Y(g18363),.A(I24373),.B(I24374));
  NAND2 NAND2_818(.VSS(VSS),.VDD(VDD),.Y(I24380),.A(g6212),.B(g13978));
  NAND2 NAND2_819(.VSS(VSS),.VDD(VDD),.Y(I24381),.A(g6212),.B(I24380));
  NAND2 NAND2_820(.VSS(VSS),.VDD(VDD),.Y(I24382),.A(g13978),.B(I24380));
  NAND2 NAND2_821(.VSS(VSS),.VDD(VDD),.Y(g18369),.A(I24381),.B(I24382));
  NAND2 NAND2_822(.VSS(VSS),.VDD(VDD),.Y(I24387),.A(g6421),.B(g13974));
  NAND2 NAND2_823(.VSS(VSS),.VDD(VDD),.Y(I24388),.A(g6421),.B(I24387));
  NAND2 NAND2_824(.VSS(VSS),.VDD(VDD),.Y(I24389),.A(g13974),.B(I24387));
  NAND2 NAND2_825(.VSS(VSS),.VDD(VDD),.Y(g18370),.A(I24388),.B(I24389));
  NAND2 NAND2_826(.VSS(VSS),.VDD(VDD),.Y(I24399),.A(g13936),.B(g9264));
  NAND2 NAND2_827(.VSS(VSS),.VDD(VDD),.Y(I24400),.A(g13936),.B(I24399));
  NAND2 NAND2_828(.VSS(VSS),.VDD(VDD),.Y(I24401),.A(g9264),.B(I24399));
  NAND2 NAND2_829(.VSS(VSS),.VDD(VDD),.Y(g18383),.A(I24400),.B(I24401));
  NAND2 NAND2_830(.VSS(VSS),.VDD(VDD),.Y(I24407),.A(g6298),.B(g14119));
  NAND2 NAND2_831(.VSS(VSS),.VDD(VDD),.Y(I24408),.A(g6298),.B(I24407));
  NAND2 NAND2_832(.VSS(VSS),.VDD(VDD),.Y(I24409),.A(g14119),.B(I24407));
  NAND2 NAND2_833(.VSS(VSS),.VDD(VDD),.Y(g18389),.A(I24408),.B(I24409));
  NAND2 NAND2_834(.VSS(VSS),.VDD(VDD),.Y(I24415),.A(g14053),.B(g15366));
  NAND2 NAND2_835(.VSS(VSS),.VDD(VDD),.Y(I24416),.A(g14053),.B(I24415));
  NAND2 NAND2_836(.VSS(VSS),.VDD(VDD),.Y(I24417),.A(g15366),.B(I24415));
  NAND2 NAND2_837(.VSS(VSS),.VDD(VDD),.Y(g18395),.A(I24416),.B(I24417));
  NAND2 NAND2_838(.VSS(VSS),.VDD(VDD),.Y(I24426),.A(g7134),.B(g14332));
  NAND2 NAND2_839(.VSS(VSS),.VDD(VDD),.Y(I24427),.A(g7134),.B(I24426));
  NAND2 NAND2_840(.VSS(VSS),.VDD(VDD),.Y(I24428),.A(g14332),.B(I24426));
  NAND2 NAND2_841(.VSS(VSS),.VDD(VDD),.Y(g18406),.A(I24427),.B(I24428));
  NAND2 NAND2_842(.VSS(VSS),.VDD(VDD),.Y(I24436),.A(g14153),.B(g15022));
  NAND2 NAND2_843(.VSS(VSS),.VDD(VDD),.Y(I24437),.A(g14153),.B(I24436));
  NAND2 NAND2_844(.VSS(VSS),.VDD(VDD),.Y(I24438),.A(g15022),.B(I24436));
  NAND2 NAND2_845(.VSS(VSS),.VDD(VDD),.Y(g18419),.A(I24437),.B(I24438));
  NAND2 NAND2_846(.VSS(VSS),.VDD(VDD),.Y(I24443),.A(g14148),.B(g9507));
  NAND2 NAND2_847(.VSS(VSS),.VDD(VDD),.Y(I24444),.A(g14148),.B(I24443));
  NAND2 NAND2_848(.VSS(VSS),.VDD(VDD),.Y(I24445),.A(g9507),.B(I24443));
  NAND2 NAND2_849(.VSS(VSS),.VDD(VDD),.Y(g18424),.A(I24444),.B(I24445));
  NAND2 NAND2_850(.VSS(VSS),.VDD(VDD),.Y(I24452),.A(g6142),.B(g14450));
  NAND2 NAND2_851(.VSS(VSS),.VDD(VDD),.Y(I24453),.A(g6142),.B(I24452));
  NAND2 NAND2_852(.VSS(VSS),.VDD(VDD),.Y(I24454),.A(g14450),.B(I24452));
  NAND2 NAND2_853(.VSS(VSS),.VDD(VDD),.Y(g18431),.A(I24453),.B(I24454));
  NAND2 NAND2_854(.VSS(VSS),.VDD(VDD),.Y(I24464),.A(g14360),.B(g9453));
  NAND2 NAND2_855(.VSS(VSS),.VDD(VDD),.Y(I24465),.A(g14360),.B(I24464));
  NAND2 NAND2_856(.VSS(VSS),.VDD(VDD),.Y(I24466),.A(g9453),.B(I24464));
  NAND2 NAND2_857(.VSS(VSS),.VDD(VDD),.Y(g18441),.A(I24465),.B(I24466));
  NAND2 NAND2_858(.VSS(VSS),.VDD(VDD),.Y(I24474),.A(g6184),.B(g14580));
  NAND2 NAND2_859(.VSS(VSS),.VDD(VDD),.Y(I24475),.A(g6184),.B(I24474));
  NAND2 NAND2_860(.VSS(VSS),.VDD(VDD),.Y(I24476),.A(g14580),.B(I24474));
  NAND2 NAND2_861(.VSS(VSS),.VDD(VDD),.Y(g18449),.A(I24475),.B(I24476));
  NAND2 NAND2_862(.VSS(VSS),.VDD(VDD),.Y(I24485),.A(g14541),.B(g9391));
  NAND2 NAND2_863(.VSS(VSS),.VDD(VDD),.Y(I24486),.A(g14541),.B(I24485));
  NAND2 NAND2_864(.VSS(VSS),.VDD(VDD),.Y(I24487),.A(g9391),.B(I24485));
  NAND2 NAND2_865(.VSS(VSS),.VDD(VDD),.Y(g18458),.A(I24486),.B(I24487));
  NAND2 NAND2_866(.VSS(VSS),.VDD(VDD),.Y(I24493),.A(g6301),.B(g14048));
  NAND2 NAND2_867(.VSS(VSS),.VDD(VDD),.Y(I24494),.A(g6301),.B(I24493));
  NAND2 NAND2_868(.VSS(VSS),.VDD(VDD),.Y(I24495),.A(g14048),.B(I24493));
  NAND2 NAND2_869(.VSS(VSS),.VDD(VDD),.Y(g18464),.A(I24494),.B(I24495));
  NAND2 NAND2_870(.VSS(VSS),.VDD(VDD),.Y(I24500),.A(g6626),.B(g14044));
  NAND2 NAND2_871(.VSS(VSS),.VDD(VDD),.Y(I24501),.A(g6626),.B(I24500));
  NAND2 NAND2_872(.VSS(VSS),.VDD(VDD),.Y(I24502),.A(g14044),.B(I24500));
  NAND2 NAND2_873(.VSS(VSS),.VDD(VDD),.Y(g18465),.A(I24501),.B(I24502));
  NAND2 NAND2_874(.VSS(VSS),.VDD(VDD),.Y(I24512),.A(g13992),.B(g9342));
  NAND2 NAND2_875(.VSS(VSS),.VDD(VDD),.Y(I24513),.A(g13992),.B(I24512));
  NAND2 NAND2_876(.VSS(VSS),.VDD(VDD),.Y(I24514),.A(g9342),.B(I24512));
  NAND2 NAND2_877(.VSS(VSS),.VDD(VDD),.Y(g18478),.A(I24513),.B(I24514));
  NAND2 NAND2_878(.VSS(VSS),.VDD(VDD),.Y(I24520),.A(g6435),.B(g14234));
  NAND2 NAND2_879(.VSS(VSS),.VDD(VDD),.Y(I24521),.A(g6435),.B(I24520));
  NAND2 NAND2_880(.VSS(VSS),.VDD(VDD),.Y(I24522),.A(g14234),.B(I24520));
  NAND2 NAND2_881(.VSS(VSS),.VDD(VDD),.Y(g18484),.A(I24521),.B(I24522));
  NAND2 NAND2_882(.VSS(VSS),.VDD(VDD),.Y(I24530),.A(g6707),.B(g14355));
  NAND2 NAND2_883(.VSS(VSS),.VDD(VDD),.Y(I24531),.A(g6707),.B(I24530));
  NAND2 NAND2_884(.VSS(VSS),.VDD(VDD),.Y(I24532),.A(g14355),.B(I24530));
  NAND2 NAND2_885(.VSS(VSS),.VDD(VDD),.Y(g18491),.A(I24531),.B(I24532));
  NAND2 NAND2_886(.VSS(VSS),.VDD(VDD),.Y(I24537),.A(g14268),.B(g15118));
  NAND2 NAND2_887(.VSS(VSS),.VDD(VDD),.Y(I24538),.A(g14268),.B(I24537));
  NAND2 NAND2_888(.VSS(VSS),.VDD(VDD),.Y(I24539),.A(g15118),.B(I24537));
  NAND2 NAND2_889(.VSS(VSS),.VDD(VDD),.Y(g18492),.A(I24538),.B(I24539));
  NAND2 NAND2_890(.VSS(VSS),.VDD(VDD),.Y(I24544),.A(g14263),.B(g9649));
  NAND2 NAND2_891(.VSS(VSS),.VDD(VDD),.Y(I24545),.A(g14263),.B(I24544));
  NAND2 NAND2_892(.VSS(VSS),.VDD(VDD),.Y(I24546),.A(g9649),.B(I24544));
  NAND2 NAND2_893(.VSS(VSS),.VDD(VDD),.Y(g18497),.A(I24545),.B(I24546));
  NAND2 NAND2_894(.VSS(VSS),.VDD(VDD),.Y(I24553),.A(g6163),.B(g14537));
  NAND2 NAND2_895(.VSS(VSS),.VDD(VDD),.Y(I24554),.A(g6163),.B(I24553));
  NAND2 NAND2_896(.VSS(VSS),.VDD(VDD),.Y(I24555),.A(g14537),.B(I24553));
  NAND2 NAND2_897(.VSS(VSS),.VDD(VDD),.Y(g18504),.A(I24554),.B(I24555));
  NAND2 NAND2_898(.VSS(VSS),.VDD(VDD),.Y(I24565),.A(g14472),.B(g9595));
  NAND2 NAND2_899(.VSS(VSS),.VDD(VDD),.Y(I24566),.A(g14472),.B(I24565));
  NAND2 NAND2_900(.VSS(VSS),.VDD(VDD),.Y(I24567),.A(g9595),.B(I24565));
  NAND2 NAND2_901(.VSS(VSS),.VDD(VDD),.Y(g18514),.A(I24566),.B(I24567));
  NAND2 NAND2_902(.VSS(VSS),.VDD(VDD),.Y(I24575),.A(g6216),.B(g14614));
  NAND2 NAND2_903(.VSS(VSS),.VDD(VDD),.Y(I24576),.A(g6216),.B(I24575));
  NAND2 NAND2_904(.VSS(VSS),.VDD(VDD),.Y(I24577),.A(g14614),.B(I24575));
  NAND2 NAND2_905(.VSS(VSS),.VDD(VDD),.Y(g18522),.A(I24576),.B(I24577));
  NAND2 NAND2_906(.VSS(VSS),.VDD(VDD),.Y(I24586),.A(g14596),.B(g9488));
  NAND2 NAND2_907(.VSS(VSS),.VDD(VDD),.Y(I24587),.A(g14596),.B(I24586));
  NAND2 NAND2_908(.VSS(VSS),.VDD(VDD),.Y(I24588),.A(g9488),.B(I24586));
  NAND2 NAND2_909(.VSS(VSS),.VDD(VDD),.Y(g18531),.A(I24587),.B(I24588));
  NAND2 NAND2_910(.VSS(VSS),.VDD(VDD),.Y(I24594),.A(g6438),.B(g14139));
  NAND2 NAND2_911(.VSS(VSS),.VDD(VDD),.Y(I24595),.A(g6438),.B(I24594));
  NAND2 NAND2_912(.VSS(VSS),.VDD(VDD),.Y(I24596),.A(g14139),.B(I24594));
  NAND2 NAND2_913(.VSS(VSS),.VDD(VDD),.Y(g18537),.A(I24595),.B(I24596));
  NAND2 NAND2_914(.VSS(VSS),.VDD(VDD),.Y(I24601),.A(g6890),.B(g14135));
  NAND2 NAND2_915(.VSS(VSS),.VDD(VDD),.Y(I24602),.A(g6890),.B(I24601));
  NAND2 NAND2_916(.VSS(VSS),.VDD(VDD),.Y(I24603),.A(g14135),.B(I24601));
  NAND2 NAND2_917(.VSS(VSS),.VDD(VDD),.Y(g18538),.A(I24602),.B(I24603));
  NAND2 NAND2_918(.VSS(VSS),.VDD(VDD),.Y(I24611),.A(g15814),.B(g15978));
  NAND2 NAND2_919(.VSS(VSS),.VDD(VDD),.Y(I24612),.A(g15814),.B(I24611));
  NAND2 NAND2_920(.VSS(VSS),.VDD(VDD),.Y(I24613),.A(g15978),.B(I24611));
  NAND2 NAND2_921(.VSS(VSS),.VDD(VDD),.Y(g18542),.A(I24612),.B(I24613));
  NAND2 NAND2_922(.VSS(VSS),.VDD(VDD),.Y(I24624),.A(g6136),.B(g14252));
  NAND2 NAND2_923(.VSS(VSS),.VDD(VDD),.Y(I24625),.A(g6136),.B(I24624));
  NAND2 NAND2_924(.VSS(VSS),.VDD(VDD),.Y(I24626),.A(g14252),.B(I24624));
  NAND2 NAND2_925(.VSS(VSS),.VDD(VDD),.Y(g18553),.A(I24625),.B(I24626));
  NAND2 NAND2_926(.VSS(VSS),.VDD(VDD),.Y(I24632),.A(g7009),.B(g14467));
  NAND2 NAND2_927(.VSS(VSS),.VDD(VDD),.Y(I24633),.A(g7009),.B(I24632));
  NAND2 NAND2_928(.VSS(VSS),.VDD(VDD),.Y(I24634),.A(g14467),.B(I24632));
  NAND2 NAND2_929(.VSS(VSS),.VDD(VDD),.Y(g18555),.A(I24633),.B(I24634));
  NAND2 NAND2_930(.VSS(VSS),.VDD(VDD),.Y(I24639),.A(g14390),.B(g15210));
  NAND2 NAND2_931(.VSS(VSS),.VDD(VDD),.Y(I24640),.A(g14390),.B(I24639));
  NAND2 NAND2_932(.VSS(VSS),.VDD(VDD),.Y(I24641),.A(g15210),.B(I24639));
  NAND2 NAND2_933(.VSS(VSS),.VDD(VDD),.Y(g18556),.A(I24640),.B(I24641));
  NAND2 NAND2_934(.VSS(VSS),.VDD(VDD),.Y(I24646),.A(g14385),.B(g9795));
  NAND2 NAND2_935(.VSS(VSS),.VDD(VDD),.Y(I24647),.A(g14385),.B(I24646));
  NAND2 NAND2_936(.VSS(VSS),.VDD(VDD),.Y(I24648),.A(g9795),.B(I24646));
  NAND2 NAND2_937(.VSS(VSS),.VDD(VDD),.Y(g18561),.A(I24647),.B(I24648));
  NAND2 NAND2_938(.VSS(VSS),.VDD(VDD),.Y(I24655),.A(g6190),.B(g14592));
  NAND2 NAND2_939(.VSS(VSS),.VDD(VDD),.Y(I24656),.A(g6190),.B(I24655));
  NAND2 NAND2_940(.VSS(VSS),.VDD(VDD),.Y(I24657),.A(g14592),.B(I24655));
  NAND2 NAND2_941(.VSS(VSS),.VDD(VDD),.Y(g18568),.A(I24656),.B(I24657));
  NAND2 NAND2_942(.VSS(VSS),.VDD(VDD),.Y(I24667),.A(g14559),.B(g9737));
  NAND2 NAND2_943(.VSS(VSS),.VDD(VDD),.Y(I24668),.A(g14559),.B(I24667));
  NAND2 NAND2_944(.VSS(VSS),.VDD(VDD),.Y(I24669),.A(g9737),.B(I24667));
  NAND2 NAND2_945(.VSS(VSS),.VDD(VDD),.Y(g18578),.A(I24668),.B(I24669));
  NAND2 NAND2_946(.VSS(VSS),.VDD(VDD),.Y(I24677),.A(g6305),.B(g14637));
  NAND2 NAND2_947(.VSS(VSS),.VDD(VDD),.Y(I24678),.A(g6305),.B(I24677));
  NAND2 NAND2_948(.VSS(VSS),.VDD(VDD),.Y(I24679),.A(g14637),.B(I24677));
  NAND2 NAND2_949(.VSS(VSS),.VDD(VDD),.Y(g18586),.A(I24678),.B(I24679));
  NAND2 NAND2_950(.VSS(VSS),.VDD(VDD),.Y(I24694),.A(g6146),.B(g14374));
  NAND2 NAND2_951(.VSS(VSS),.VDD(VDD),.Y(I24695),.A(g6146),.B(I24694));
  NAND2 NAND2_952(.VSS(VSS),.VDD(VDD),.Y(I24696),.A(g14374),.B(I24694));
  NAND2 NAND2_953(.VSS(VSS),.VDD(VDD),.Y(g18603),.A(I24695),.B(I24696));
  NAND2 NAND2_954(.VSS(VSS),.VDD(VDD),.Y(I24702),.A(g7259),.B(g14554));
  NAND2 NAND2_955(.VSS(VSS),.VDD(VDD),.Y(I24703),.A(g7259),.B(I24702));
  NAND2 NAND2_956(.VSS(VSS),.VDD(VDD),.Y(I24704),.A(g14554),.B(I24702));
  NAND2 NAND2_957(.VSS(VSS),.VDD(VDD),.Y(g18605),.A(I24703),.B(I24704));
  NAND2 NAND2_958(.VSS(VSS),.VDD(VDD),.Y(I24709),.A(g14502),.B(g15296));
  NAND2 NAND2_959(.VSS(VSS),.VDD(VDD),.Y(I24710),.A(g14502),.B(I24709));
  NAND2 NAND2_960(.VSS(VSS),.VDD(VDD),.Y(I24711),.A(g15296),.B(I24709));
  NAND2 NAND2_961(.VSS(VSS),.VDD(VDD),.Y(g18606),.A(I24710),.B(I24711));
  NAND2 NAND2_962(.VSS(VSS),.VDD(VDD),.Y(I24716),.A(g14497),.B(g9941));
  NAND2 NAND2_963(.VSS(VSS),.VDD(VDD),.Y(I24717),.A(g14497),.B(I24716));
  NAND2 NAND2_964(.VSS(VSS),.VDD(VDD),.Y(I24718),.A(g9941),.B(I24716));
  NAND2 NAND2_965(.VSS(VSS),.VDD(VDD),.Y(g18611),.A(I24717),.B(I24718));
  NAND2 NAND2_966(.VSS(VSS),.VDD(VDD),.Y(I24725),.A(g6222),.B(g14626));
  NAND2 NAND2_967(.VSS(VSS),.VDD(VDD),.Y(I24726),.A(g6222),.B(I24725));
  NAND2 NAND2_968(.VSS(VSS),.VDD(VDD),.Y(I24727),.A(g14626),.B(I24725));
  NAND2 NAND2_969(.VSS(VSS),.VDD(VDD),.Y(g18618),.A(I24726),.B(I24727));
  NAND2 NAND2_970(.VSS(VSS),.VDD(VDD),.Y(I24743),.A(g6167),.B(g14486));
  NAND2 NAND2_971(.VSS(VSS),.VDD(VDD),.Y(I24744),.A(g6167),.B(I24743));
  NAND2 NAND2_972(.VSS(VSS),.VDD(VDD),.Y(I24745),.A(g14486),.B(I24743));
  NAND2 NAND2_973(.VSS(VSS),.VDD(VDD),.Y(g18635),.A(I24744),.B(I24745));
  NAND2 NAND2_974(.VSS(VSS),.VDD(VDD),.Y(I24751),.A(g7455),.B(g14609));
  NAND2 NAND2_975(.VSS(VSS),.VDD(VDD),.Y(I24752),.A(g7455),.B(I24751));
  NAND2 NAND2_976(.VSS(VSS),.VDD(VDD),.Y(I24753),.A(g14609),.B(I24751));
  NAND2 NAND2_977(.VSS(VSS),.VDD(VDD),.Y(g18637),.A(I24752),.B(I24753));
  NAND2 NAND2_978(.VSS(VSS),.VDD(VDD),.Y(I24763),.A(g6194),.B(g14573));
  NAND2 NAND2_979(.VSS(VSS),.VDD(VDD),.Y(I24764),.A(g6194),.B(I24763));
  NAND2 NAND2_980(.VSS(VSS),.VDD(VDD),.Y(I24765),.A(g14573),.B(I24763));
  NAND2 NAND2_981(.VSS(VSS),.VDD(VDD),.Y(g18644),.A(I24764),.B(I24765));
  NAND2 NAND2_982(.VSS(VSS),.VDD(VDD),.Y(g18977),.A(g15797),.B(g3006));
  NAND2 NAND2_983(.VSS(VSS),.VDD(VDD),.Y(I25030),.A(g8029),.B(g13507));
  NAND2 NAND2_984(.VSS(VSS),.VDD(VDD),.Y(I25031),.A(g8029),.B(I25030));
  NAND2 NAND2_985(.VSS(VSS),.VDD(VDD),.Y(I25032),.A(g13507),.B(I25030));
  NAND2 NAND2_986(.VSS(VSS),.VDD(VDD),.Y(g18980),.A(I25031),.B(I25032));
  NAND2 NAND2_987(.VSS(VSS),.VDD(VDD),.Y(g19067),.A(g16554),.B(g16578));
  NAND2 NAND2_988(.VSS(VSS),.VDD(VDD),.Y(g19084),.A(g16586),.B(g16602));
  NAND2 NAND2_989(.VSS(VSS),.VDD(VDD),.Y(g19103),.A(g18590),.B(g2924));
  NAND2 NAND2_990(.VSS(VSS),.VDD(VDD),.Y(g19121),.A(g16682),.B(g16697));
  NAND2 NAND2_991(.VSS(VSS),.VDD(VDD),.Y(g19128),.A(g16708),.B(g16728));
  NAND2 NAND2_992(.VSS(VSS),.VDD(VDD),.Y(g19135),.A(g16739),.B(g16770));
  NAND2 NAND2_993(.VSS(VSS),.VDD(VDD),.Y(g19138),.A(g16781),.B(g16797));
  NAND2 NAND2_994(.VSS(VSS),.VDD(VDD),.Y(g19141),.A(g3088),.B(g16825));
  NAND2 NAND2_995(.VSS(VSS),.VDD(VDD),.Y(g19152),.A(g5378),.B(g18884));
  NAND2 NAND2_996(.VSS(VSS),.VDD(VDD),.Y(I25532),.A(g52),.B(g18179));
  NAND2 NAND2_997(.VSS(VSS),.VDD(VDD),.Y(I25533),.A(g52),.B(I25532));
  NAND2 NAND2_998(.VSS(VSS),.VDD(VDD),.Y(I25534),.A(g18179),.B(I25532));
  NAND2 NAND2_999(.VSS(VSS),.VDD(VDD),.Y(g19261),.A(I25533),.B(I25534));
  NAND2 NAND2_1000(.VSS(VSS),.VDD(VDD),.Y(I25539),.A(g92),.B(g18174));
  NAND2 NAND2_1001(.VSS(VSS),.VDD(VDD),.Y(I25540),.A(g92),.B(I25539));
  NAND2 NAND2_1002(.VSS(VSS),.VDD(VDD),.Y(I25541),.A(g18174),.B(I25539));
  NAND2 NAND2_1003(.VSS(VSS),.VDD(VDD),.Y(g19262),.A(I25540),.B(I25541));
  NAND2 NAND2_1004(.VSS(VSS),.VDD(VDD),.Y(I25560),.A(g56),.B(g17724));
  NAND2 NAND2_1005(.VSS(VSS),.VDD(VDD),.Y(I25561),.A(g56),.B(I25560));
  NAND2 NAND2_1006(.VSS(VSS),.VDD(VDD),.Y(I25562),.A(g17724),.B(I25560));
  NAND2 NAND2_1007(.VSS(VSS),.VDD(VDD),.Y(g19271),.A(I25561),.B(I25562));
  NAND2 NAND2_1008(.VSS(VSS),.VDD(VDD),.Y(I25571),.A(g740),.B(g18286));
  NAND2 NAND2_1009(.VSS(VSS),.VDD(VDD),.Y(I25572),.A(g740),.B(I25571));
  NAND2 NAND2_1010(.VSS(VSS),.VDD(VDD),.Y(I25573),.A(g18286),.B(I25571));
  NAND2 NAND2_1011(.VSS(VSS),.VDD(VDD),.Y(g19276),.A(I25572),.B(I25573));
  NAND2 NAND2_1012(.VSS(VSS),.VDD(VDD),.Y(I25578),.A(g780),.B(g18281));
  NAND2 NAND2_1013(.VSS(VSS),.VDD(VDD),.Y(I25579),.A(g780),.B(I25578));
  NAND2 NAND2_1014(.VSS(VSS),.VDD(VDD),.Y(I25580),.A(g18281),.B(I25578));
  NAND2 NAND2_1015(.VSS(VSS),.VDD(VDD),.Y(g19277),.A(I25579),.B(I25580));
  NAND2 NAND2_1016(.VSS(VSS),.VDD(VDD),.Y(I25595),.A(g61),.B(g18074));
  NAND2 NAND2_1017(.VSS(VSS),.VDD(VDD),.Y(I25596),.A(g61),.B(I25595));
  NAND2 NAND2_1018(.VSS(VSS),.VDD(VDD),.Y(I25597),.A(g18074),.B(I25595));
  NAND2 NAND2_1019(.VSS(VSS),.VDD(VDD),.Y(g19286),.A(I25596),.B(I25597));
  NAND3 NAND3_8(.VSS(VSS),.VDD(VDD),.Y(g19288),.A(g14685),.B(g8580),.C(g17057));
  NAND2 NAND2_1020(.VSS(VSS),.VDD(VDD),.Y(I25605),.A(g744),.B(g17825));
  NAND2 NAND2_1021(.VSS(VSS),.VDD(VDD),.Y(I25606),.A(g744),.B(I25605));
  NAND2 NAND2_1022(.VSS(VSS),.VDD(VDD),.Y(I25607),.A(g17825),.B(I25605));
  NAND2 NAND2_1023(.VSS(VSS),.VDD(VDD),.Y(g19290),.A(I25606),.B(I25607));
  NAND2 NAND2_1024(.VSS(VSS),.VDD(VDD),.Y(I25616),.A(g1426),.B(g18379));
  NAND2 NAND2_1025(.VSS(VSS),.VDD(VDD),.Y(I25617),.A(g1426),.B(I25616));
  NAND2 NAND2_1026(.VSS(VSS),.VDD(VDD),.Y(I25618),.A(g18379),.B(I25616));
  NAND2 NAND2_1027(.VSS(VSS),.VDD(VDD),.Y(g19295),.A(I25617),.B(I25618));
  NAND2 NAND2_1028(.VSS(VSS),.VDD(VDD),.Y(I25623),.A(g1466),.B(g18374));
  NAND2 NAND2_1029(.VSS(VSS),.VDD(VDD),.Y(I25624),.A(g1466),.B(I25623));
  NAND2 NAND2_1030(.VSS(VSS),.VDD(VDD),.Y(I25625),.A(g18374),.B(I25623));
  NAND2 NAND2_1031(.VSS(VSS),.VDD(VDD),.Y(g19296),.A(I25624),.B(I25625));
  NAND2 NAND2_1032(.VSS(VSS),.VDD(VDD),.Y(I25633),.A(g65),.B(g17640));
  NAND2 NAND2_1033(.VSS(VSS),.VDD(VDD),.Y(I25634),.A(g65),.B(I25633));
  NAND2 NAND2_1034(.VSS(VSS),.VDD(VDD),.Y(I25635),.A(g17640),.B(I25633));
  NAND2 NAND2_1035(.VSS(VSS),.VDD(VDD),.Y(g19300),.A(I25634),.B(I25635));
  NAND2 NAND2_1036(.VSS(VSS),.VDD(VDD),.Y(I25643),.A(g749),.B(g18190));
  NAND2 NAND2_1037(.VSS(VSS),.VDD(VDD),.Y(I25644),.A(g749),.B(I25643));
  NAND2 NAND2_1038(.VSS(VSS),.VDD(VDD),.Y(I25645),.A(g18190),.B(I25643));
  NAND2 NAND2_1039(.VSS(VSS),.VDD(VDD),.Y(g19304),.A(I25644),.B(I25645));
  NAND3 NAND3_9(.VSS(VSS),.VDD(VDD),.Y(g19306),.A(g14719),.B(g8587),.C(g17092));
  NAND2 NAND2_1040(.VSS(VSS),.VDD(VDD),.Y(I25653),.A(g1430),.B(g17937));
  NAND2 NAND2_1041(.VSS(VSS),.VDD(VDD),.Y(I25654),.A(g1430),.B(I25653));
  NAND2 NAND2_1042(.VSS(VSS),.VDD(VDD),.Y(I25655),.A(g17937),.B(I25653));
  NAND2 NAND2_1043(.VSS(VSS),.VDD(VDD),.Y(g19308),.A(I25654),.B(I25655));
  NAND2 NAND2_1044(.VSS(VSS),.VDD(VDD),.Y(I25664),.A(g2120),.B(g18474));
  NAND2 NAND2_1045(.VSS(VSS),.VDD(VDD),.Y(I25665),.A(g2120),.B(I25664));
  NAND2 NAND2_1046(.VSS(VSS),.VDD(VDD),.Y(I25666),.A(g18474),.B(I25664));
  NAND2 NAND2_1047(.VSS(VSS),.VDD(VDD),.Y(g19313),.A(I25665),.B(I25666));
  NAND2 NAND2_1048(.VSS(VSS),.VDD(VDD),.Y(I25671),.A(g2160),.B(g18469));
  NAND2 NAND2_1049(.VSS(VSS),.VDD(VDD),.Y(I25672),.A(g2160),.B(I25671));
  NAND2 NAND2_1050(.VSS(VSS),.VDD(VDD),.Y(I25673),.A(g18469),.B(I25671));
  NAND2 NAND2_1051(.VSS(VSS),.VDD(VDD),.Y(g19314),.A(I25672),.B(I25673));
  NAND2 NAND2_1052(.VSS(VSS),.VDD(VDD),.Y(I25681),.A(g70),.B(g17974));
  NAND2 NAND2_1053(.VSS(VSS),.VDD(VDD),.Y(I25682),.A(g70),.B(I25681));
  NAND2 NAND2_1054(.VSS(VSS),.VDD(VDD),.Y(I25683),.A(g17974),.B(I25681));
  NAND2 NAND2_1055(.VSS(VSS),.VDD(VDD),.Y(g19318),.A(I25682),.B(I25683));
  NAND2 NAND2_1056(.VSS(VSS),.VDD(VDD),.Y(I25690),.A(g753),.B(g17741));
  NAND2 NAND2_1057(.VSS(VSS),.VDD(VDD),.Y(I25691),.A(g753),.B(I25690));
  NAND2 NAND2_1058(.VSS(VSS),.VDD(VDD),.Y(I25692),.A(g17741),.B(I25690));
  NAND2 NAND2_1059(.VSS(VSS),.VDD(VDD),.Y(g19321),.A(I25691),.B(I25692));
  NAND2 NAND2_1060(.VSS(VSS),.VDD(VDD),.Y(I25700),.A(g1435),.B(g18297));
  NAND2 NAND2_1061(.VSS(VSS),.VDD(VDD),.Y(I25701),.A(g1435),.B(I25700));
  NAND2 NAND2_1062(.VSS(VSS),.VDD(VDD),.Y(I25702),.A(g18297),.B(I25700));
  NAND2 NAND2_1063(.VSS(VSS),.VDD(VDD),.Y(g19325),.A(I25701),.B(I25702));
  NAND3 NAND3_10(.VSS(VSS),.VDD(VDD),.Y(g19327),.A(g14747),.B(g8594),.C(g17130));
  NAND2 NAND2_1064(.VSS(VSS),.VDD(VDD),.Y(I25710),.A(g2124),.B(g18048));
  NAND2 NAND2_1065(.VSS(VSS),.VDD(VDD),.Y(I25711),.A(g2124),.B(I25710));
  NAND2 NAND2_1066(.VSS(VSS),.VDD(VDD),.Y(I25712),.A(g18048),.B(I25710));
  NAND2 NAND2_1067(.VSS(VSS),.VDD(VDD),.Y(g19329),.A(I25711),.B(I25712));
  NAND2 NAND2_1068(.VSS(VSS),.VDD(VDD),.Y(I25721),.A(g74),.B(g18341));
  NAND2 NAND2_1069(.VSS(VSS),.VDD(VDD),.Y(I25722),.A(g74),.B(I25721));
  NAND2 NAND2_1070(.VSS(VSS),.VDD(VDD),.Y(I25723),.A(g18341),.B(I25721));
  NAND2 NAND2_1071(.VSS(VSS),.VDD(VDD),.Y(g19334),.A(I25722),.B(I25723));
  NAND2 NAND2_1072(.VSS(VSS),.VDD(VDD),.Y(I25731),.A(g758),.B(g18091));
  NAND2 NAND2_1073(.VSS(VSS),.VDD(VDD),.Y(I25732),.A(g758),.B(I25731));
  NAND2 NAND2_1074(.VSS(VSS),.VDD(VDD),.Y(I25733),.A(g18091),.B(I25731));
  NAND2 NAND2_1075(.VSS(VSS),.VDD(VDD),.Y(g19345),.A(I25732),.B(I25733));
  NAND2 NAND2_1076(.VSS(VSS),.VDD(VDD),.Y(I25740),.A(g1439),.B(g17842));
  NAND2 NAND2_1077(.VSS(VSS),.VDD(VDD),.Y(I25741),.A(g1439),.B(I25740));
  NAND2 NAND2_1078(.VSS(VSS),.VDD(VDD),.Y(I25742),.A(g17842),.B(I25740));
  NAND2 NAND2_1079(.VSS(VSS),.VDD(VDD),.Y(g19348),.A(I25741),.B(I25742));
  NAND2 NAND2_1080(.VSS(VSS),.VDD(VDD),.Y(I25750),.A(g2129),.B(g18390));
  NAND2 NAND2_1081(.VSS(VSS),.VDD(VDD),.Y(I25751),.A(g2129),.B(I25750));
  NAND2 NAND2_1082(.VSS(VSS),.VDD(VDD),.Y(I25752),.A(g18390),.B(I25750));
  NAND2 NAND2_1083(.VSS(VSS),.VDD(VDD),.Y(g19352),.A(I25751),.B(I25752));
  NAND3 NAND3_11(.VSS(VSS),.VDD(VDD),.Y(g19354),.A(g14768),.B(g8605),.C(g17157));
  NAND2 NAND2_1084(.VSS(VSS),.VDD(VDD),.Y(I25761),.A(g79),.B(g17882));
  NAND2 NAND2_1085(.VSS(VSS),.VDD(VDD),.Y(I25762),.A(g79),.B(I25761));
  NAND2 NAND2_1086(.VSS(VSS),.VDD(VDD),.Y(I25763),.A(g17882),.B(I25761));
  NAND2 NAND2_1087(.VSS(VSS),.VDD(VDD),.Y(g19357),.A(I25762),.B(I25763));
  NAND2 NAND2_1088(.VSS(VSS),.VDD(VDD),.Y(I25771),.A(g762),.B(g18436));
  NAND2 NAND2_1089(.VSS(VSS),.VDD(VDD),.Y(I25772),.A(g762),.B(I25771));
  NAND2 NAND2_1090(.VSS(VSS),.VDD(VDD),.Y(I25773),.A(g18436),.B(I25771));
  NAND2 NAND2_1091(.VSS(VSS),.VDD(VDD),.Y(g19368),.A(I25772),.B(I25773));
  NAND2 NAND2_1092(.VSS(VSS),.VDD(VDD),.Y(I25781),.A(g1444),.B(g18207));
  NAND2 NAND2_1093(.VSS(VSS),.VDD(VDD),.Y(I25782),.A(g1444),.B(I25781));
  NAND2 NAND2_1094(.VSS(VSS),.VDD(VDD),.Y(I25783),.A(g18207),.B(I25781));
  NAND2 NAND2_1095(.VSS(VSS),.VDD(VDD),.Y(g19379),.A(I25782),.B(I25783));
  NAND2 NAND2_1096(.VSS(VSS),.VDD(VDD),.Y(I25790),.A(g2133),.B(g17954));
  NAND2 NAND2_1097(.VSS(VSS),.VDD(VDD),.Y(I25791),.A(g2133),.B(I25790));
  NAND2 NAND2_1098(.VSS(VSS),.VDD(VDD),.Y(I25792),.A(g17954),.B(I25790));
  NAND2 NAND2_1099(.VSS(VSS),.VDD(VDD),.Y(g19382),.A(I25791),.B(I25792));
  NAND2 NAND2_1100(.VSS(VSS),.VDD(VDD),.Y(I25800),.A(g83),.B(g18265));
  NAND2 NAND2_1101(.VSS(VSS),.VDD(VDD),.Y(I25801),.A(g83),.B(I25800));
  NAND2 NAND2_1102(.VSS(VSS),.VDD(VDD),.Y(I25802),.A(g18265),.B(I25800));
  NAND2 NAND2_1103(.VSS(VSS),.VDD(VDD),.Y(g19386),.A(I25801),.B(I25802));
  NAND2 NAND2_1104(.VSS(VSS),.VDD(VDD),.Y(I25809),.A(g767),.B(g17993));
  NAND2 NAND2_1105(.VSS(VSS),.VDD(VDD),.Y(I25810),.A(g767),.B(I25809));
  NAND2 NAND2_1106(.VSS(VSS),.VDD(VDD),.Y(I25811),.A(g17993),.B(I25809));
  NAND2 NAND2_1107(.VSS(VSS),.VDD(VDD),.Y(g19389),.A(I25810),.B(I25811));
  NAND2 NAND2_1108(.VSS(VSS),.VDD(VDD),.Y(I25819),.A(g1448),.B(g18509));
  NAND2 NAND2_1109(.VSS(VSS),.VDD(VDD),.Y(I25820),.A(g1448),.B(I25819));
  NAND2 NAND2_1110(.VSS(VSS),.VDD(VDD),.Y(I25821),.A(g18509),.B(I25819));
  NAND2 NAND2_1111(.VSS(VSS),.VDD(VDD),.Y(g19400),.A(I25820),.B(I25821));
  NAND2 NAND2_1112(.VSS(VSS),.VDD(VDD),.Y(I25829),.A(g2138),.B(g18314));
  NAND2 NAND2_1113(.VSS(VSS),.VDD(VDD),.Y(I25830),.A(g2138),.B(I25829));
  NAND2 NAND2_1114(.VSS(VSS),.VDD(VDD),.Y(I25831),.A(g18314),.B(I25829));
  NAND2 NAND2_1115(.VSS(VSS),.VDD(VDD),.Y(g19411),.A(I25830),.B(I25831));
  NAND2 NAND2_1116(.VSS(VSS),.VDD(VDD),.Y(I25838),.A(g88),.B(g17802));
  NAND2 NAND2_1117(.VSS(VSS),.VDD(VDD),.Y(I25839),.A(g88),.B(I25838));
  NAND2 NAND2_1118(.VSS(VSS),.VDD(VDD),.Y(I25840),.A(g17802),.B(I25838));
  NAND2 NAND2_1119(.VSS(VSS),.VDD(VDD),.Y(g19414),.A(I25839),.B(I25840));
  NAND2 NAND2_1120(.VSS(VSS),.VDD(VDD),.Y(I25846),.A(g771),.B(g18358));
  NAND2 NAND2_1121(.VSS(VSS),.VDD(VDD),.Y(I25847),.A(g771),.B(I25846));
  NAND2 NAND2_1122(.VSS(VSS),.VDD(VDD),.Y(I25848),.A(g18358),.B(I25846));
  NAND2 NAND2_1123(.VSS(VSS),.VDD(VDD),.Y(g19416),.A(I25847),.B(I25848));
  NAND2 NAND2_1124(.VSS(VSS),.VDD(VDD),.Y(I25855),.A(g1453),.B(g18110));
  NAND2 NAND2_1125(.VSS(VSS),.VDD(VDD),.Y(I25856),.A(g1453),.B(I25855));
  NAND2 NAND2_1126(.VSS(VSS),.VDD(VDD),.Y(I25857),.A(g18110),.B(I25855));
  NAND2 NAND2_1127(.VSS(VSS),.VDD(VDD),.Y(g19419),.A(I25856),.B(I25857));
  NAND2 NAND2_1128(.VSS(VSS),.VDD(VDD),.Y(I25865),.A(g2142),.B(g18573));
  NAND2 NAND2_1129(.VSS(VSS),.VDD(VDD),.Y(I25866),.A(g2142),.B(I25865));
  NAND2 NAND2_1130(.VSS(VSS),.VDD(VDD),.Y(I25867),.A(g18573),.B(I25865));
  NAND2 NAND2_1131(.VSS(VSS),.VDD(VDD),.Y(g19430),.A(I25866),.B(I25867));
  NAND2 NAND2_1132(.VSS(VSS),.VDD(VDD),.Y(I25880),.A(g776),.B(g17914));
  NAND2 NAND2_1133(.VSS(VSS),.VDD(VDD),.Y(I25881),.A(g776),.B(I25880));
  NAND2 NAND2_1134(.VSS(VSS),.VDD(VDD),.Y(I25882),.A(g17914),.B(I25880));
  NAND2 NAND2_1135(.VSS(VSS),.VDD(VDD),.Y(g19451),.A(I25881),.B(I25882));
  NAND2 NAND2_1136(.VSS(VSS),.VDD(VDD),.Y(I25888),.A(g1457),.B(g18453));
  NAND2 NAND2_1137(.VSS(VSS),.VDD(VDD),.Y(I25889),.A(g1457),.B(I25888));
  NAND2 NAND2_1138(.VSS(VSS),.VDD(VDD),.Y(I25890),.A(g18453),.B(I25888));
  NAND2 NAND2_1139(.VSS(VSS),.VDD(VDD),.Y(g19453),.A(I25889),.B(I25890));
  NAND2 NAND2_1140(.VSS(VSS),.VDD(VDD),.Y(I25897),.A(g2147),.B(g18226));
  NAND2 NAND2_1141(.VSS(VSS),.VDD(VDD),.Y(I25898),.A(g2147),.B(I25897));
  NAND2 NAND2_1142(.VSS(VSS),.VDD(VDD),.Y(I25899),.A(g18226),.B(I25897));
  NAND2 NAND2_1143(.VSS(VSS),.VDD(VDD),.Y(g19456),.A(I25898),.B(I25899));
  NAND2 NAND2_1144(.VSS(VSS),.VDD(VDD),.Y(I25913),.A(g1462),.B(g18025));
  NAND2 NAND2_1145(.VSS(VSS),.VDD(VDD),.Y(I25914),.A(g1462),.B(I25913));
  NAND2 NAND2_1146(.VSS(VSS),.VDD(VDD),.Y(I25915),.A(g18025),.B(I25913));
  NAND2 NAND2_1147(.VSS(VSS),.VDD(VDD),.Y(g19478),.A(I25914),.B(I25915));
  NAND2 NAND2_1148(.VSS(VSS),.VDD(VDD),.Y(I25921),.A(g2151),.B(g18526));
  NAND2 NAND2_1149(.VSS(VSS),.VDD(VDD),.Y(I25922),.A(g2151),.B(I25921));
  NAND2 NAND2_1150(.VSS(VSS),.VDD(VDD),.Y(I25923),.A(g18526),.B(I25921));
  NAND2 NAND2_1151(.VSS(VSS),.VDD(VDD),.Y(g19480),.A(I25922),.B(I25923));
  NAND2 NAND2_1152(.VSS(VSS),.VDD(VDD),.Y(I25938),.A(g2156),.B(g18142));
  NAND2 NAND2_1153(.VSS(VSS),.VDD(VDD),.Y(I25939),.A(g2156),.B(I25938));
  NAND2 NAND2_1154(.VSS(VSS),.VDD(VDD),.Y(I25940),.A(g18142),.B(I25938));
  NAND2 NAND2_1155(.VSS(VSS),.VDD(VDD),.Y(g19501),.A(I25939),.B(I25940));
  NAND2 NAND2_1156(.VSS(VSS),.VDD(VDD),.Y(g19865),.A(g16607),.B(g9636));
  NAND2 NAND2_1157(.VSS(VSS),.VDD(VDD),.Y(g19896),.A(g16625),.B(g9782));
  NAND2 NAND2_1158(.VSS(VSS),.VDD(VDD),.Y(g19921),.A(g16639),.B(g9928));
  NAND2 NAND2_1159(.VSS(VSS),.VDD(VDD),.Y(g19936),.A(g16650),.B(g10082));
  NAND2 NAND2_1160(.VSS(VSS),.VDD(VDD),.Y(g19954),.A(g17186),.B(g92));
  NAND2 NAND2_1161(.VSS(VSS),.VDD(VDD),.Y(g19984),.A(g17197),.B(g780));
  NAND2 NAND2_1162(.VSS(VSS),.VDD(VDD),.Y(g20022),.A(g17204),.B(g1466));
  NAND2 NAND2_1163(.VSS(VSS),.VDD(VDD),.Y(g20064),.A(g17209),.B(g2160));
  NAND2 NAND2_1164(.VSS(VSS),.VDD(VDD),.Y(g20473),.A(g18085),.B(g646));
  NAND2 NAND2_1165(.VSS(VSS),.VDD(VDD),.Y(g20481),.A(g18201),.B(g1332));
  NAND2 NAND2_1166(.VSS(VSS),.VDD(VDD),.Y(g20487),.A(g18308),.B(g2026));
  NAND2 NAND2_1167(.VSS(VSS),.VDD(VDD),.Y(g20493),.A(g18401),.B(g2720));
  NAND2 NAND2_1168(.VSS(VSS),.VDD(VDD),.Y(g20497),.A(g5410),.B(g18886));
  NAND2 NAND2_1169(.VSS(VSS),.VDD(VDD),.Y(g20522),.A(g16501),.B(g16515));
  NAND2 NAND2_1170(.VSS(VSS),.VDD(VDD),.Y(g20537),.A(g18626),.B(g3036));
  NAND2 NAND2_1171(.VSS(VSS),.VDD(VDD),.Y(g20542),.A(g16523),.B(g16546));
  NAND2 NAND2_1172(.VSS(VSS),.VDD(VDD),.Y(g20633),.A(g20164),.B(g3254));
  NAND2 NAND2_1173(.VSS(VSS),.VDD(VDD),.Y(g20648),.A(g20164),.B(g3254));
  NAND2 NAND2_1174(.VSS(VSS),.VDD(VDD),.Y(g20658),.A(g20198),.B(g3410));
  NAND2 NAND2_1175(.VSS(VSS),.VDD(VDD),.Y(g20672),.A(g20164),.B(g3254));
  NAND2 NAND2_1176(.VSS(VSS),.VDD(VDD),.Y(g20683),.A(g20198),.B(g3410));
  NAND2 NAND2_1177(.VSS(VSS),.VDD(VDD),.Y(g20693),.A(g20228),.B(g3566));
  NAND2 NAND2_1178(.VSS(VSS),.VDD(VDD),.Y(g20700),.A(g20153),.B(g2903));
  NAND2 NAND2_1179(.VSS(VSS),.VDD(VDD),.Y(g20703),.A(g20164),.B(g3254));
  NAND2 NAND2_1180(.VSS(VSS),.VDD(VDD),.Y(g20707),.A(g20198),.B(g3410));
  NAND2 NAND2_1181(.VSS(VSS),.VDD(VDD),.Y(g20718),.A(g20228),.B(g3566));
  NAND2 NAND2_1182(.VSS(VSS),.VDD(VDD),.Y(g20728),.A(g20255),.B(g3722));
  NAND2 NAND2_1183(.VSS(VSS),.VDD(VDD),.Y(g20738),.A(g20198),.B(g3410));
  NAND2 NAND2_1184(.VSS(VSS),.VDD(VDD),.Y(g20742),.A(g20228),.B(g3566));
  NAND2 NAND2_1185(.VSS(VSS),.VDD(VDD),.Y(g20753),.A(g20255),.B(g3722));
  NAND2 NAND2_1186(.VSS(VSS),.VDD(VDD),.Y(g20775),.A(g20228),.B(g3566));
  NAND2 NAND2_1187(.VSS(VSS),.VDD(VDD),.Y(g20779),.A(g20255),.B(g3722));
  NAND2 NAND2_1188(.VSS(VSS),.VDD(VDD),.Y(g20805),.A(g20255),.B(g3722));
  NAND2 NAND2_1189(.VSS(VSS),.VDD(VDD),.Y(g20825),.A(g19219),.B(g15959));
  NAND2 NAND2_1190(.VSS(VSS),.VDD(VDD),.Y(g21659),.A(g20164),.B(g6314));
  NAND2 NAND2_1191(.VSS(VSS),.VDD(VDD),.Y(I28189),.A(g14079),.B(g19444));
  NAND2 NAND2_1192(.VSS(VSS),.VDD(VDD),.Y(I28190),.A(g14079),.B(I28189));
  NAND2 NAND2_1193(.VSS(VSS),.VDD(VDD),.Y(I28191),.A(g19444),.B(I28189));
  NAND2 NAND2_1194(.VSS(VSS),.VDD(VDD),.Y(g21660),.A(I28190),.B(I28191));
  NAND2 NAND2_1195(.VSS(VSS),.VDD(VDD),.Y(g21685),.A(g20164),.B(g6232));
  NAND2 NAND2_1196(.VSS(VSS),.VDD(VDD),.Y(g21686),.A(g20164),.B(g6314));
  NAND2 NAND2_1197(.VSS(VSS),.VDD(VDD),.Y(g21688),.A(g20198),.B(g6519));
  NAND2 NAND2_1198(.VSS(VSS),.VDD(VDD),.Y(I28217),.A(g14194),.B(g19471));
  NAND2 NAND2_1199(.VSS(VSS),.VDD(VDD),.Y(I28218),.A(g14194),.B(I28217));
  NAND2 NAND2_1200(.VSS(VSS),.VDD(VDD),.Y(I28219),.A(g19471),.B(I28217));
  NAND2 NAND2_1201(.VSS(VSS),.VDD(VDD),.Y(g21689),.A(I28218),.B(I28219));
  NAND2 NAND2_1202(.VSS(VSS),.VDD(VDD),.Y(g21714),.A(g20164),.B(g6232));
  NAND2 NAND2_1203(.VSS(VSS),.VDD(VDD),.Y(g21715),.A(g20164),.B(g6314));
  NAND4 NAND4_1(.VSS(VSS),.VDD(VDD),.Y(g21720),.A(g14256),.B(g15177),.C(g19871),.D(g19842));
  NAND2 NAND2_1204(.VSS(VSS),.VDD(VDD),.Y(g21721),.A(g20198),.B(g6369));
  NAND2 NAND2_1205(.VSS(VSS),.VDD(VDD),.Y(g21722),.A(g20198),.B(g6519));
  NAND2 NAND2_1206(.VSS(VSS),.VDD(VDD),.Y(g21724),.A(g20228),.B(g6783));
  NAND2 NAND2_1207(.VSS(VSS),.VDD(VDD),.Y(I28247),.A(g14309),.B(g19494));
  NAND2 NAND2_1208(.VSS(VSS),.VDD(VDD),.Y(I28248),.A(g14309),.B(I28247));
  NAND2 NAND2_1209(.VSS(VSS),.VDD(VDD),.Y(I28249),.A(g19494),.B(I28247));
  NAND2 NAND2_1210(.VSS(VSS),.VDD(VDD),.Y(g21725),.A(I28248),.B(I28249));
  NAND2 NAND2_1211(.VSS(VSS),.VDD(VDD),.Y(g21736),.A(g20164),.B(g6232));
  NAND2 NAND2_1212(.VSS(VSS),.VDD(VDD),.Y(g21737),.A(g20164),.B(g6314));
  NAND2 NAND2_1213(.VSS(VSS),.VDD(VDD),.Y(g21740),.A(g20198),.B(g6369));
  NAND2 NAND2_1214(.VSS(VSS),.VDD(VDD),.Y(g21741),.A(g20198),.B(g6519));
  NAND4 NAND4_2(.VSS(VSS),.VDD(VDD),.Y(g21746),.A(g14378),.B(g15263),.C(g19902),.D(g19875));
  NAND2 NAND2_1215(.VSS(VSS),.VDD(VDD),.Y(g21747),.A(g20228),.B(g6574));
  NAND2 NAND2_1216(.VSS(VSS),.VDD(VDD),.Y(g21748),.A(g20228),.B(g6783));
  NAND2 NAND2_1217(.VSS(VSS),.VDD(VDD),.Y(g21750),.A(g20255),.B(g7085));
  NAND2 NAND2_1218(.VSS(VSS),.VDD(VDD),.Y(I28271),.A(g14431),.B(g19515));
  NAND2 NAND2_1219(.VSS(VSS),.VDD(VDD),.Y(I28272),.A(g14431),.B(I28271));
  NAND2 NAND2_1220(.VSS(VSS),.VDD(VDD),.Y(I28273),.A(g19515),.B(I28271));
  NAND2 NAND2_1221(.VSS(VSS),.VDD(VDD),.Y(g21751),.A(I28272),.B(I28273));
  NAND2 NAND2_1222(.VSS(VSS),.VDD(VDD),.Y(g21759),.A(g20164),.B(g6232));
  NAND2 NAND2_1223(.VSS(VSS),.VDD(VDD),.Y(g21760),.A(g20198),.B(g6369));
  NAND2 NAND2_1224(.VSS(VSS),.VDD(VDD),.Y(g21761),.A(g20198),.B(g6519));
  NAND2 NAND2_1225(.VSS(VSS),.VDD(VDD),.Y(g21764),.A(g20228),.B(g6574));
  NAND2 NAND2_1226(.VSS(VSS),.VDD(VDD),.Y(g21765),.A(g20228),.B(g6783));
  NAND4 NAND4_3(.VSS(VSS),.VDD(VDD),.Y(g21770),.A(g14490),.B(g15355),.C(g19927),.D(g19906));
  NAND2 NAND2_1227(.VSS(VSS),.VDD(VDD),.Y(g21771),.A(g20255),.B(g6838));
  NAND2 NAND2_1228(.VSS(VSS),.VDD(VDD),.Y(g21772),.A(g20255),.B(g7085));
  NAND2 NAND2_1229(.VSS(VSS),.VDD(VDD),.Y(g21775),.A(g20198),.B(g6369));
  NAND2 NAND2_1230(.VSS(VSS),.VDD(VDD),.Y(g21776),.A(g20228),.B(g6574));
  NAND2 NAND2_1231(.VSS(VSS),.VDD(VDD),.Y(g21777),.A(g20228),.B(g6783));
  NAND2 NAND2_1232(.VSS(VSS),.VDD(VDD),.Y(g21780),.A(g20255),.B(g6838));
  NAND2 NAND2_1233(.VSS(VSS),.VDD(VDD),.Y(g21781),.A(g20255),.B(g7085));
  NAND4 NAND4_4(.VSS(VSS),.VDD(VDD),.Y(g21786),.A(g14577),.B(g15441),.C(g19942),.D(g19931));
  NAND2 NAND2_1234(.VSS(VSS),.VDD(VDD),.Y(g21790),.A(g20228),.B(g6574));
  NAND2 NAND2_1235(.VSS(VSS),.VDD(VDD),.Y(g21791),.A(g20255),.B(g6838));
  NAND2 NAND2_1236(.VSS(VSS),.VDD(VDD),.Y(g21792),.A(g20255),.B(g7085));
  NAND2 NAND2_1237(.VSS(VSS),.VDD(VDD),.Y(g21804),.A(g20255),.B(g6838));
  NAND3 NAND3_12(.VSS(VSS),.VDD(VDD),.Y(g21848),.A(g17807),.B(g19181),.C(g19186));
  NAND3 NAND3_13(.VSS(VSS),.VDD(VDD),.Y(g21850),.A(g17979),.B(g19187),.C(g19191));
  NAND3 NAND3_14(.VSS(VSS),.VDD(VDD),.Y(g21855),.A(g17919),.B(g19188),.C(g19193));
  NAND3 NAND3_15(.VSS(VSS),.VDD(VDD),.Y(g21857),.A(g18079),.B(g19192),.C(g19200));
  NAND3 NAND3_16(.VSS(VSS),.VDD(VDD),.Y(g21858),.A(g18096),.B(g19194),.C(g19202));
  NAND3 NAND3_17(.VSS(VSS),.VDD(VDD),.Y(g21859),.A(g18030),.B(g19195),.C(g19204));
  NAND3 NAND3_18(.VSS(VSS),.VDD(VDD),.Y(g21860),.A(g18270),.B(g19201),.C(g19209));
  NAND3 NAND3_19(.VSS(VSS),.VDD(VDD),.Y(g21862),.A(g18195),.B(g19203),.C(g19211));
  NAND3 NAND3_20(.VSS(VSS),.VDD(VDD),.Y(g21863),.A(g18212),.B(g19205),.C(g19213));
  NAND3 NAND3_21(.VSS(VSS),.VDD(VDD),.Y(g21864),.A(g18147),.B(g19206),.C(g19215));
  NAND3 NAND3_22(.VSS(VSS),.VDD(VDD),.Y(g21865),.A(g18424),.B(g19210),.C(g19221));
  NAND3 NAND3_23(.VSS(VSS),.VDD(VDD),.Y(g21866),.A(g18363),.B(g19212),.C(g19222));
  NAND3 NAND3_24(.VSS(VSS),.VDD(VDD),.Y(g21868),.A(g18302),.B(g19214),.C(g19224));
  NAND3 NAND3_25(.VSS(VSS),.VDD(VDD),.Y(g21869),.A(g18319),.B(g19216),.C(g19226));
  NAND3 NAND3_26(.VSS(VSS),.VDD(VDD),.Y(g21870),.A(g18497),.B(g19223),.C(g19231));
  NAND3 NAND3_27(.VSS(VSS),.VDD(VDD),.Y(g21871),.A(g18458),.B(g19225),.C(g19232));
  NAND3 NAND3_28(.VSS(VSS),.VDD(VDD),.Y(g21873),.A(g18395),.B(g19227),.C(g19234));
  NAND3 NAND3_29(.VSS(VSS),.VDD(VDD),.Y(g21874),.A(g18561),.B(g19233),.C(g19244));
  NAND3 NAND3_30(.VSS(VSS),.VDD(VDD),.Y(g21875),.A(g18531),.B(g19235),.C(g19245));
  NAND3 NAND3_31(.VSS(VSS),.VDD(VDD),.Y(g21877),.A(g18611),.B(g19246),.C(g19257));
  NAND3 NAND3_32(.VSS(VSS),.VDD(VDD),.Y(g21879),.A(g18419),.B(g19250),.C(g19263));
  NAND3 NAND3_33(.VSS(VSS),.VDD(VDD),.Y(g21881),.A(g18492),.B(g19264),.C(g19278));
  NAND3 NAND3_34(.VSS(VSS),.VDD(VDD),.Y(g21885),.A(g18556),.B(g19279),.C(g19297));
  NAND3 NAND3_35(.VSS(VSS),.VDD(VDD),.Y(g21888),.A(g18606),.B(g19298),.C(g19315));
  NAND2 NAND2_1238(.VSS(VSS),.VDD(VDD),.Y(g21903),.A(g20008),.B(g3013));
  NAND3 NAND3_36(.VSS(VSS),.VDD(VDD),.Y(g21976),.A(g19242),.B(g21120),.C(g19275));
  NAND3 NAND3_37(.VSS(VSS),.VDD(VDD),.Y(g21983),.A(g19255),.B(g21139),.C(g19294));
  NAND2 NAND2_1239(.VSS(VSS),.VDD(VDD),.Y(g21989),.A(g21048),.B(g18623));
  NAND2 NAND2_1240(.VSS(VSS),.VDD(VDD),.Y(g21991),.A(g21501),.B(g21536));
  NAND3 NAND3_38(.VSS(VSS),.VDD(VDD),.Y(g21996),.A(g19268),.B(g21159),.C(g19312));
  NAND2 NAND2_1241(.VSS(VSS),.VDD(VDD),.Y(g22002),.A(g21065),.B(g21711));
  NAND2 NAND2_1242(.VSS(VSS),.VDD(VDD),.Y(g22005),.A(g21540),.B(g21572));
  NAND3 NAND3_39(.VSS(VSS),.VDD(VDD),.Y(g22009),.A(g19283),.B(g21179),.C(g19333));
  NAND2 NAND2_1243(.VSS(VSS),.VDD(VDD),.Y(g22016),.A(g21576),.B(g21605));
  NAND2 NAND2_1244(.VSS(VSS),.VDD(VDD),.Y(g22021),.A(g21609),.B(g21634));
  NAND3 NAND3_40(.VSS(VSS),.VDD(VDD),.Y(g22050),.A(g19450),.B(g21244),.C(g19503));
  NAND3 NAND3_41(.VSS(VSS),.VDD(VDD),.Y(g22069),.A(g19477),.B(g21253),.C(g19522));
  NAND2 NAND2_1245(.VSS(VSS),.VDD(VDD),.Y(g22083),.A(g21774),.B(g21787));
  NAND3 NAND3_42(.VSS(VSS),.VDD(VDD),.Y(g22093),.A(g19500),.B(g21261),.C(g19532));
  NAND2 NAND2_1246(.VSS(VSS),.VDD(VDD),.Y(g22108),.A(g21789),.B(g21801));
  NAND3 NAND3_43(.VSS(VSS),.VDD(VDD),.Y(g22118),.A(g19521),.B(g21269),.C(g19542));
  NAND2 NAND2_1247(.VSS(VSS),.VDD(VDD),.Y(g22134),.A(g21803),.B(g21809));
  NAND2 NAND2_1248(.VSS(VSS),.VDD(VDD),.Y(g22157),.A(g21811),.B(g21816));
  NAND2 NAND2_1249(.VSS(VSS),.VDD(VDD),.Y(I28726),.A(g21887),.B(g13519));
  NAND2 NAND2_1250(.VSS(VSS),.VDD(VDD),.Y(I28727),.A(g21887),.B(I28726));
  NAND2 NAND2_1251(.VSS(VSS),.VDD(VDD),.Y(I28728),.A(g13519),.B(I28726));
  NAND2 NAND2_1252(.VSS(VSS),.VDD(VDD),.Y(g22188),.A(I28727),.B(I28728));
  NAND2 NAND2_1253(.VSS(VSS),.VDD(VDD),.Y(I28741),.A(g21890),.B(g13530));
  NAND2 NAND2_1254(.VSS(VSS),.VDD(VDD),.Y(I28742),.A(g21890),.B(I28741));
  NAND2 NAND2_1255(.VSS(VSS),.VDD(VDD),.Y(I28743),.A(g13530),.B(I28741));
  NAND2 NAND2_1256(.VSS(VSS),.VDD(VDD),.Y(g22197),.A(I28742),.B(I28743));
  NAND2 NAND2_1257(.VSS(VSS),.VDD(VDD),.Y(I28753),.A(g21893),.B(g13541));
  NAND2 NAND2_1258(.VSS(VSS),.VDD(VDD),.Y(I28754),.A(g21893),.B(I28753));
  NAND2 NAND2_1259(.VSS(VSS),.VDD(VDD),.Y(I28755),.A(g13541),.B(I28753));
  NAND2 NAND2_1260(.VSS(VSS),.VDD(VDD),.Y(g22203),.A(I28754),.B(I28755));
  NAND2 NAND2_1261(.VSS(VSS),.VDD(VDD),.Y(I28765),.A(g21901),.B(g13552));
  NAND2 NAND2_1262(.VSS(VSS),.VDD(VDD),.Y(I28766),.A(g21901),.B(I28765));
  NAND2 NAND2_1263(.VSS(VSS),.VDD(VDD),.Y(I28767),.A(g13552),.B(I28765));
  NAND2 NAND2_1264(.VSS(VSS),.VDD(VDD),.Y(g22209),.A(I28766),.B(I28767));
  NAND3 NAND3_44(.VSS(VSS),.VDD(VDD),.Y(g22317),.A(g21152),.B(g21241),.C(g21136));
  NAND3 NAND3_45(.VSS(VSS),.VDD(VDD),.Y(g22339),.A(g14442),.B(g21149),.C(g10694));
  NAND3 NAND3_46(.VSS(VSS),.VDD(VDD),.Y(g22342),.A(g21172),.B(g21249),.C(g21156));
  NAND3 NAND3_47(.VSS(VSS),.VDD(VDD),.Y(g22362),.A(g14529),.B(g21169),.C(g10714));
  NAND3 NAND3_48(.VSS(VSS),.VDD(VDD),.Y(g22365),.A(g21192),.B(g21258),.C(g21176));
  NAND3 NAND3_49(.VSS(VSS),.VDD(VDD),.Y(g22381),.A(g21211),.B(g14442),.C(g10694));
  NAND3 NAND3_50(.VSS(VSS),.VDD(VDD),.Y(g22382),.A(g14584),.B(g21189),.C(g10735));
  NAND3 NAND3_51(.VSS(VSS),.VDD(VDD),.Y(g22385),.A(g21207),.B(g21266),.C(g21196));
  NAND3 NAND3_52(.VSS(VSS),.VDD(VDD),.Y(g22396),.A(g21219),.B(g14529),.C(g10714));
  NAND3 NAND3_53(.VSS(VSS),.VDD(VDD),.Y(g22397),.A(g14618),.B(g21204),.C(g10754));
  NAND3 NAND3_54(.VSS(VSS),.VDD(VDD),.Y(g22399),.A(g21230),.B(g14584),.C(g10735));
  NAND3 NAND3_55(.VSS(VSS),.VDD(VDD),.Y(g22400),.A(g21235),.B(g14618),.C(g10754));
  NAND2 NAND2_1265(.VSS(VSS),.VDD(VDD),.Y(g22608),.A(g20842),.B(g20885));
  NAND2 NAND2_1266(.VSS(VSS),.VDD(VDD),.Y(g22644),.A(g20850),.B(g20904));
  NAND2 NAND2_1267(.VSS(VSS),.VDD(VDD),.Y(g22668),.A(g16075),.B(g21271));
  NAND2 NAND2_1268(.VSS(VSS),.VDD(VDD),.Y(g22680),.A(g20858),.B(g20928));
  NAND2 NAND2_1269(.VSS(VSS),.VDD(VDD),.Y(g22708),.A(g16113),.B(g21278));
  NAND2 NAND2_1270(.VSS(VSS),.VDD(VDD),.Y(g22720),.A(g20866),.B(g20956));
  NAND2 NAND2_1271(.VSS(VSS),.VDD(VDD),.Y(g22739),.A(g16164),.B(g21285));
  NAND2 NAND2_1272(.VSS(VSS),.VDD(VDD),.Y(g22771),.A(g16223),.B(g21293));
  NAND3 NAND3_56(.VSS(VSS),.VDD(VDD),.Y(g22809),.A(g21850),.B(g21848),.C(g21879));
  NAND3 NAND3_57(.VSS(VSS),.VDD(VDD),.Y(g22844),.A(g21865),.B(g21860),.C(g21857));
  NAND2 NAND2_1273(.VSS(VSS),.VDD(VDD),.Y(g22845),.A(g19441),.B(g20885));
  NAND2 NAND2_1274(.VSS(VSS),.VDD(VDD),.Y(g22846),.A(g8278),.B(g21660));
  NAND3 NAND3_58(.VSS(VSS),.VDD(VDD),.Y(g22850),.A(g21858),.B(g21855),.C(g21881));
  NAND2 NAND2_1275(.VSS(VSS),.VDD(VDD),.Y(g22876),.A(g21238),.B(g83));
  NAND3 NAND3_59(.VSS(VSS),.VDD(VDD),.Y(g22879),.A(g21870),.B(g21866),.C(g21862));
  NAND2 NAND2_1276(.VSS(VSS),.VDD(VDD),.Y(g22880),.A(g19468),.B(g20904));
  NAND2 NAND2_1277(.VSS(VSS),.VDD(VDD),.Y(g22881),.A(g8287),.B(g21689));
  NAND3 NAND3_60(.VSS(VSS),.VDD(VDD),.Y(g22885),.A(g21863),.B(g21859),.C(g21885));
  NAND2 NAND2_1278(.VSS(VSS),.VDD(VDD),.Y(g22911),.A(g21246),.B(g771));
  NAND3 NAND3_61(.VSS(VSS),.VDD(VDD),.Y(g22914),.A(g21874),.B(g21871),.C(g21868));
  NAND2 NAND2_1279(.VSS(VSS),.VDD(VDD),.Y(g22915),.A(g19491),.B(g20928));
  NAND2 NAND2_1280(.VSS(VSS),.VDD(VDD),.Y(g22916),.A(g8296),.B(g21725));
  NAND3 NAND3_62(.VSS(VSS),.VDD(VDD),.Y(g22920),.A(g21869),.B(g21864),.C(g21888));
  NAND2 NAND2_1281(.VSS(VSS),.VDD(VDD),.Y(g22936),.A(g21255),.B(g1457));
  NAND3 NAND3_63(.VSS(VSS),.VDD(VDD),.Y(g22939),.A(g21877),.B(g21875),.C(g21873));
  NAND2 NAND2_1282(.VSS(VSS),.VDD(VDD),.Y(g22940),.A(g19512),.B(g20956));
  NAND2 NAND2_1283(.VSS(VSS),.VDD(VDD),.Y(g22941),.A(g8305),.B(g21751));
  NAND2 NAND2_1284(.VSS(VSS),.VDD(VDD),.Y(g22942),.A(g21263),.B(g2151));
  NAND2 NAND2_1285(.VSS(VSS),.VDD(VDD),.Y(g22992),.A(g21636),.B(g672));
  NAND2 NAND2_1286(.VSS(VSS),.VDD(VDD),.Y(g23003),.A(g21667),.B(g1358));
  NAND2 NAND2_1287(.VSS(VSS),.VDD(VDD),.Y(g23017),.A(g21696),.B(g2052));
  NAND2 NAND2_1288(.VSS(VSS),.VDD(VDD),.Y(g23033),.A(g21732),.B(g2746));
  NAND2 NAND2_1289(.VSS(VSS),.VDD(VDD),.Y(g23320),.A(g23066),.B(g23051));
  NAND2 NAND2_1290(.VSS(VSS),.VDD(VDD),.Y(g23325),.A(g23080),.B(g23070));
  NAND2 NAND2_1291(.VSS(VSS),.VDD(VDD),.Y(g23331),.A(g22999),.B(g22174));
  NAND2 NAND2_1292(.VSS(VSS),.VDD(VDD),.Y(g23335),.A(g23096),.B(g23083));
  NAND2 NAND2_1293(.VSS(VSS),.VDD(VDD),.Y(g23340),.A(g23013),.B(g22189));
  NAND2 NAND2_1294(.VSS(VSS),.VDD(VDD),.Y(g23344),.A(g23113),.B(g23099));
  NAND2 NAND2_1295(.VSS(VSS),.VDD(VDD),.Y(g23349),.A(g23029),.B(g22198));
  NAND2 NAND2_1296(.VSS(VSS),.VDD(VDD),.Y(g23353),.A(g23046),.B(g22204));
  NAND2 NAND2_1297(.VSS(VSS),.VDD(VDD),.Y(g23360),.A(g21980),.B(g21975));
  NAND2 NAND2_1298(.VSS(VSS),.VDD(VDD),.Y(g23364),.A(g21987),.B(g21981));
  NAND2 NAND2_1299(.VSS(VSS),.VDD(VDD),.Y(g23368),.A(g23135),.B(g22288));
  NAND2 NAND2_1300(.VSS(VSS),.VDD(VDD),.Y(g23372),.A(g22000),.B(g21988));
  NAND2 NAND2_1301(.VSS(VSS),.VDD(VDD),.Y(g23376),.A(g18435),.B(g22812));
  NAND2 NAND2_1302(.VSS(VSS),.VDD(VDD),.Y(g23377),.A(g21968),.B(g22308));
  NAND2 NAND2_1303(.VSS(VSS),.VDD(VDD),.Y(g23381),.A(g22013),.B(g22001));
  NAND2 NAND2_1304(.VSS(VSS),.VDD(VDD),.Y(g23387),.A(g18508),.B(g22852));
  NAND2 NAND2_1305(.VSS(VSS),.VDD(VDD),.Y(g23388),.A(g21971),.B(g22336));
  NAND2 NAND2_1306(.VSS(VSS),.VDD(VDD),.Y(g23394),.A(g18572),.B(g22887));
  NAND2 NAND2_1307(.VSS(VSS),.VDD(VDD),.Y(g23395),.A(g21973),.B(g22361));
  NAND2 NAND2_1308(.VSS(VSS),.VDD(VDD),.Y(g23402),.A(g18622),.B(g22922));
  NAND3 NAND3_64(.VSS(VSS),.VDD(VDD),.Y(g23478),.A(g22809),.B(g14442),.C(g10694));
  NAND3 NAND3_65(.VSS(VSS),.VDD(VDD),.Y(g23486),.A(g22844),.B(g14442),.C(g10694));
  NAND3 NAND3_66(.VSS(VSS),.VDD(VDD),.Y(g23489),.A(g22850),.B(g14529),.C(g10714));
  NAND3 NAND3_67(.VSS(VSS),.VDD(VDD),.Y(g23495),.A(g10694),.B(g14442),.C(g22316));
  NAND3 NAND3_68(.VSS(VSS),.VDD(VDD),.Y(g23502),.A(g22879),.B(g14529),.C(g10714));
  NAND3 NAND3_69(.VSS(VSS),.VDD(VDD),.Y(g23505),.A(g22885),.B(g14584),.C(g10735));
  NAND3 NAND3_70(.VSS(VSS),.VDD(VDD),.Y(g23511),.A(g10714),.B(g14529),.C(g22341));
  NAND3 NAND3_71(.VSS(VSS),.VDD(VDD),.Y(g23518),.A(g22914),.B(g14584),.C(g10735));
  NAND3 NAND3_72(.VSS(VSS),.VDD(VDD),.Y(g23521),.A(g22920),.B(g14618),.C(g10754));
  NAND3 NAND3_73(.VSS(VSS),.VDD(VDD),.Y(g23526),.A(g10735),.B(g14584),.C(g22364));
  NAND3 NAND3_74(.VSS(VSS),.VDD(VDD),.Y(g23533),.A(g22939),.B(g14618),.C(g10754));
  NAND3 NAND3_75(.VSS(VSS),.VDD(VDD),.Y(g23537),.A(g10754),.B(g14618),.C(g22384));
  NAND2 NAND2_1309(.VSS(VSS),.VDD(VDD),.Y(I30790),.A(g22846),.B(g14079));
  NAND2 NAND2_1310(.VSS(VSS),.VDD(VDD),.Y(I30791),.A(g22846),.B(I30790));
  NAND2 NAND2_1311(.VSS(VSS),.VDD(VDD),.Y(I30792),.A(g14079),.B(I30790));
  NAND2 NAND2_1312(.VSS(VSS),.VDD(VDD),.Y(g23660),.A(I30791),.B(I30792));
  NAND2 NAND2_1313(.VSS(VSS),.VDD(VDD),.Y(I30868),.A(g22881),.B(g14194));
  NAND2 NAND2_1314(.VSS(VSS),.VDD(VDD),.Y(I30869),.A(g22881),.B(I30868));
  NAND2 NAND2_1315(.VSS(VSS),.VDD(VDD),.Y(I30870),.A(g14194),.B(I30868));
  NAND2 NAND2_1316(.VSS(VSS),.VDD(VDD),.Y(g23710),.A(I30869),.B(I30870));
  NAND2 NAND2_1317(.VSS(VSS),.VDD(VDD),.Y(I30952),.A(g22916),.B(g14309));
  NAND2 NAND2_1318(.VSS(VSS),.VDD(VDD),.Y(I30953),.A(g22916),.B(I30952));
  NAND2 NAND2_1319(.VSS(VSS),.VDD(VDD),.Y(I30954),.A(g14309),.B(I30952));
  NAND2 NAND2_1320(.VSS(VSS),.VDD(VDD),.Y(g23764),.A(I30953),.B(I30954));
  NAND2 NAND2_1321(.VSS(VSS),.VDD(VDD),.Y(I31035),.A(g22941),.B(g14431));
  NAND2 NAND2_1322(.VSS(VSS),.VDD(VDD),.Y(I31036),.A(g22941),.B(I31035));
  NAND2 NAND2_1323(.VSS(VSS),.VDD(VDD),.Y(I31037),.A(g14431),.B(I31035));
  NAND2 NAND2_1324(.VSS(VSS),.VDD(VDD),.Y(g23819),.A(I31036),.B(I31037));
  NAND2 NAND2_1325(.VSS(VSS),.VDD(VDD),.Y(g23906),.A(g22812),.B(g13958));
  NAND2 NAND2_1326(.VSS(VSS),.VDD(VDD),.Y(g23936),.A(g22812),.B(g13922));
  NAND2 NAND2_1327(.VSS(VSS),.VDD(VDD),.Y(g23937),.A(g22812),.B(g13918));
  NAND2 NAND2_1328(.VSS(VSS),.VDD(VDD),.Y(g23938),.A(g22852),.B(g14028));
  NAND2 NAND2_1329(.VSS(VSS),.VDD(VDD),.Y(g23953),.A(g22812),.B(g14525));
  NAND2 NAND2_1330(.VSS(VSS),.VDD(VDD),.Y(g23968),.A(g22852),.B(g13978));
  NAND2 NAND2_1331(.VSS(VSS),.VDD(VDD),.Y(g23969),.A(g22852),.B(g13974));
  NAND2 NAND2_1332(.VSS(VSS),.VDD(VDD),.Y(g23970),.A(g22887),.B(g14119));
  NAND2 NAND2_1333(.VSS(VSS),.VDD(VDD),.Y(g23973),.A(g22812),.B(g14450));
  NAND2 NAND2_1334(.VSS(VSS),.VDD(VDD),.Y(g23982),.A(g22852),.B(g14580));
  NAND2 NAND2_1335(.VSS(VSS),.VDD(VDD),.Y(g23997),.A(g22887),.B(g14048));
  NAND2 NAND2_1336(.VSS(VSS),.VDD(VDD),.Y(g23998),.A(g22887),.B(g14044));
  NAND2 NAND2_1337(.VSS(VSS),.VDD(VDD),.Y(g23999),.A(g22922),.B(g14234));
  NAND2 NAND2_1338(.VSS(VSS),.VDD(VDD),.Y(g24002),.A(g22812),.B(g14355));
  NAND2 NAND2_1339(.VSS(VSS),.VDD(VDD),.Y(g24003),.A(g22852),.B(g14537));
  NAND2 NAND2_1340(.VSS(VSS),.VDD(VDD),.Y(g24012),.A(g22887),.B(g14614));
  NAND2 NAND2_1341(.VSS(VSS),.VDD(VDD),.Y(g24027),.A(g22922),.B(g14139));
  NAND2 NAND2_1342(.VSS(VSS),.VDD(VDD),.Y(g24028),.A(g22922),.B(g14135));
  NAND2 NAND2_1343(.VSS(VSS),.VDD(VDD),.Y(g24034),.A(g22812),.B(g14252));
  NAND2 NAND2_1344(.VSS(VSS),.VDD(VDD),.Y(g24036),.A(g22852),.B(g14467));
  NAND2 NAND2_1345(.VSS(VSS),.VDD(VDD),.Y(g24037),.A(g22887),.B(g14592));
  NAND2 NAND2_1346(.VSS(VSS),.VDD(VDD),.Y(g24046),.A(g22922),.B(g14637));
  NAND2 NAND2_1347(.VSS(VSS),.VDD(VDD),.Y(g24052),.A(g22812),.B(g14171));
  NAND2 NAND2_1348(.VSS(VSS),.VDD(VDD),.Y(g24054),.A(g22852),.B(g14374));
  NAND2 NAND2_1349(.VSS(VSS),.VDD(VDD),.Y(g24056),.A(g22887),.B(g14554));
  NAND2 NAND2_1350(.VSS(VSS),.VDD(VDD),.Y(g24057),.A(g22922),.B(g14626));
  NAND2 NAND2_1351(.VSS(VSS),.VDD(VDD),.Y(g24058),.A(g22812),.B(g14086));
  NAND2 NAND2_1352(.VSS(VSS),.VDD(VDD),.Y(g24065),.A(g22852),.B(g14286));
  NAND2 NAND2_1353(.VSS(VSS),.VDD(VDD),.Y(g24067),.A(g22887),.B(g14486));
  NAND2 NAND2_1354(.VSS(VSS),.VDD(VDD),.Y(g24069),.A(g22922),.B(g14609));
  NAND2 NAND2_1355(.VSS(VSS),.VDD(VDD),.Y(g24070),.A(g22812),.B(g14011));
  NAND2 NAND2_1356(.VSS(VSS),.VDD(VDD),.Y(g24071),.A(g22852),.B(g14201));
  NAND2 NAND2_1357(.VSS(VSS),.VDD(VDD),.Y(g24078),.A(g22887),.B(g14408));
  NAND2 NAND2_1358(.VSS(VSS),.VDD(VDD),.Y(g24080),.A(g22922),.B(g14573));
  NAND2 NAND2_1359(.VSS(VSS),.VDD(VDD),.Y(g24081),.A(g22852),.B(g14102));
  NAND2 NAND2_1360(.VSS(VSS),.VDD(VDD),.Y(g24082),.A(g22887),.B(g14316));
  NAND2 NAND2_1361(.VSS(VSS),.VDD(VDD),.Y(g24089),.A(g22922),.B(g14520));
  NAND2 NAND2_1362(.VSS(VSS),.VDD(VDD),.Y(g24090),.A(g22887),.B(g14217));
  NAND2 NAND2_1363(.VSS(VSS),.VDD(VDD),.Y(g24091),.A(g22922),.B(g14438));
  NAND2 NAND2_1364(.VSS(VSS),.VDD(VDD),.Y(g24093),.A(g22922),.B(g14332));
  NAND2 NAND2_1365(.VSS(VSS),.VDD(VDD),.Y(g24100),.A(g20885),.B(g22175));
  NAND2 NAND2_1366(.VSS(VSS),.VDD(VDD),.Y(g24109),.A(g20904),.B(g22190));
  NAND2 NAND2_1367(.VSS(VSS),.VDD(VDD),.Y(g24126),.A(g20928),.B(g22199));
  NAND2 NAND2_1368(.VSS(VSS),.VDD(VDD),.Y(g24145),.A(g20956),.B(g22205));
  NAND2 NAND2_1369(.VSS(VSS),.VDD(VDD),.Y(g24442),.A(g23644),.B(g3306));
  NAND2 NAND2_1370(.VSS(VSS),.VDD(VDD),.Y(g24443),.A(g23644),.B(g3306));
  NAND2 NAND2_1371(.VSS(VSS),.VDD(VDD),.Y(g24444),.A(g23694),.B(g3462));
  NAND2 NAND2_1372(.VSS(VSS),.VDD(VDD),.Y(g24447),.A(g23644),.B(g3306));
  NAND2 NAND2_1373(.VSS(VSS),.VDD(VDD),.Y(g24448),.A(g23923),.B(g3338));
  NAND2 NAND2_1374(.VSS(VSS),.VDD(VDD),.Y(g24449),.A(g23694),.B(g3462));
  NAND2 NAND2_1375(.VSS(VSS),.VDD(VDD),.Y(g24450),.A(g23748),.B(g3618));
  NAND2 NAND2_1376(.VSS(VSS),.VDD(VDD),.Y(g24451),.A(g23644),.B(g3306));
  NAND2 NAND2_1377(.VSS(VSS),.VDD(VDD),.Y(g24452),.A(g23923),.B(g3338));
  NAND2 NAND2_1378(.VSS(VSS),.VDD(VDD),.Y(g24453),.A(g23694),.B(g3462));
  NAND2 NAND2_1379(.VSS(VSS),.VDD(VDD),.Y(g24454),.A(g23955),.B(g3494));
  NAND2 NAND2_1380(.VSS(VSS),.VDD(VDD),.Y(g24455),.A(g23748),.B(g3618));
  NAND2 NAND2_1381(.VSS(VSS),.VDD(VDD),.Y(g24456),.A(g23803),.B(g3774));
  NAND2 NAND2_1382(.VSS(VSS),.VDD(VDD),.Y(g24457),.A(g23923),.B(g3338));
  NAND2 NAND2_1383(.VSS(VSS),.VDD(VDD),.Y(g24458),.A(g23694),.B(g3462));
  NAND2 NAND2_1384(.VSS(VSS),.VDD(VDD),.Y(g24459),.A(g23955),.B(g3494));
  NAND2 NAND2_1385(.VSS(VSS),.VDD(VDD),.Y(g24460),.A(g23748),.B(g3618));
  NAND2 NAND2_1386(.VSS(VSS),.VDD(VDD),.Y(g24461),.A(g23984),.B(g3650));
  NAND2 NAND2_1387(.VSS(VSS),.VDD(VDD),.Y(g24462),.A(g23803),.B(g3774));
  NAND2 NAND2_1388(.VSS(VSS),.VDD(VDD),.Y(g24463),.A(g23923),.B(g3338));
  NAND2 NAND2_1389(.VSS(VSS),.VDD(VDD),.Y(g24464),.A(g23955),.B(g3494));
  NAND2 NAND2_1390(.VSS(VSS),.VDD(VDD),.Y(g24465),.A(g23748),.B(g3618));
  NAND2 NAND2_1391(.VSS(VSS),.VDD(VDD),.Y(g24466),.A(g23984),.B(g3650));
  NAND2 NAND2_1392(.VSS(VSS),.VDD(VDD),.Y(g24467),.A(g23803),.B(g3774));
  NAND2 NAND2_1393(.VSS(VSS),.VDD(VDD),.Y(g24468),.A(g24014),.B(g3806));
  NAND2 NAND2_1394(.VSS(VSS),.VDD(VDD),.Y(g24469),.A(g23955),.B(g3494));
  NAND2 NAND2_1395(.VSS(VSS),.VDD(VDD),.Y(g24470),.A(g23984),.B(g3650));
  NAND2 NAND2_1396(.VSS(VSS),.VDD(VDD),.Y(g24471),.A(g23803),.B(g3774));
  NAND2 NAND2_1397(.VSS(VSS),.VDD(VDD),.Y(g24472),.A(g24014),.B(g3806));
  NAND2 NAND2_1398(.VSS(VSS),.VDD(VDD),.Y(g24474),.A(g23984),.B(g3650));
  NAND2 NAND2_1399(.VSS(VSS),.VDD(VDD),.Y(g24475),.A(g24014),.B(g3806));
  NAND2 NAND2_1400(.VSS(VSS),.VDD(VDD),.Y(g24477),.A(g24014),.B(g3806));
  NAND2 NAND2_1401(.VSS(VSS),.VDD(VDD),.Y(g24616),.A(g499),.B(g23376));
  NAND2 NAND2_1402(.VSS(VSS),.VDD(VDD),.Y(g24627),.A(g1186),.B(g23387));
  NAND2 NAND2_1403(.VSS(VSS),.VDD(VDD),.Y(g24641),.A(g1880),.B(g23394));
  NAND2 NAND2_1404(.VSS(VSS),.VDD(VDD),.Y(g24660),.A(g2574),.B(g23402));
  NAND2 NAND2_1405(.VSS(VSS),.VDD(VDD),.Y(I32265),.A(g17903),.B(g23936));
  NAND2 NAND2_1406(.VSS(VSS),.VDD(VDD),.Y(I32266),.A(g17903),.B(I32265));
  NAND2 NAND2_1407(.VSS(VSS),.VDD(VDD),.Y(I32267),.A(g23936),.B(I32265));
  NAND2 NAND2_1408(.VSS(VSS),.VDD(VDD),.Y(g24753),.A(I32266),.B(I32267));
  NAND2 NAND2_1409(.VSS(VSS),.VDD(VDD),.Y(I32284),.A(g17815),.B(g23953));
  NAND2 NAND2_1410(.VSS(VSS),.VDD(VDD),.Y(I32285),.A(g17815),.B(I32284));
  NAND2 NAND2_1411(.VSS(VSS),.VDD(VDD),.Y(I32286),.A(g23953),.B(I32284));
  NAND2 NAND2_1412(.VSS(VSS),.VDD(VDD),.Y(g24766),.A(I32285),.B(I32286));
  NAND2 NAND2_1413(.VSS(VSS),.VDD(VDD),.Y(I32295),.A(g18014),.B(g23968));
  NAND2 NAND2_1414(.VSS(VSS),.VDD(VDD),.Y(I32296),.A(g18014),.B(I32295));
  NAND2 NAND2_1415(.VSS(VSS),.VDD(VDD),.Y(I32297),.A(g23968),.B(I32295));
  NAND2 NAND2_1416(.VSS(VSS),.VDD(VDD),.Y(g24771),.A(I32296),.B(I32297));
  NAND2 NAND2_1417(.VSS(VSS),.VDD(VDD),.Y(I32308),.A(g17903),.B(g23973));
  NAND2 NAND2_1418(.VSS(VSS),.VDD(VDD),.Y(I32309),.A(g17903),.B(I32308));
  NAND2 NAND2_1419(.VSS(VSS),.VDD(VDD),.Y(I32310),.A(g23973),.B(I32308));
  NAND2 NAND2_1420(.VSS(VSS),.VDD(VDD),.Y(g24778),.A(I32309),.B(I32310));
  NAND2 NAND2_1421(.VSS(VSS),.VDD(VDD),.Y(I32323),.A(g17927),.B(g23982));
  NAND2 NAND2_1422(.VSS(VSS),.VDD(VDD),.Y(I32324),.A(g17927),.B(I32323));
  NAND2 NAND2_1423(.VSS(VSS),.VDD(VDD),.Y(I32325),.A(g23982),.B(I32323));
  NAND2 NAND2_1424(.VSS(VSS),.VDD(VDD),.Y(g24787),.A(I32324),.B(I32325));
  NAND2 NAND2_1425(.VSS(VSS),.VDD(VDD),.Y(I32333),.A(g18131),.B(g23997));
  NAND2 NAND2_1426(.VSS(VSS),.VDD(VDD),.Y(I32334),.A(g18131),.B(I32333));
  NAND2 NAND2_1427(.VSS(VSS),.VDD(VDD),.Y(I32335),.A(g23997),.B(I32333));
  NAND2 NAND2_1428(.VSS(VSS),.VDD(VDD),.Y(g24791),.A(I32334),.B(I32335));
  NAND2 NAND2_1429(.VSS(VSS),.VDD(VDD),.Y(I32345),.A(g17815),.B(g24002));
  NAND2 NAND2_1430(.VSS(VSS),.VDD(VDD),.Y(I32346),.A(g17815),.B(I32345));
  NAND2 NAND2_1431(.VSS(VSS),.VDD(VDD),.Y(I32347),.A(g24002),.B(I32345));
  NAND2 NAND2_1432(.VSS(VSS),.VDD(VDD),.Y(g24797),.A(I32346),.B(I32347));
  NAND2 NAND2_1433(.VSS(VSS),.VDD(VDD),.Y(I32355),.A(g18014),.B(g24003));
  NAND2 NAND2_1434(.VSS(VSS),.VDD(VDD),.Y(I32356),.A(g18014),.B(I32355));
  NAND2 NAND2_1435(.VSS(VSS),.VDD(VDD),.Y(I32357),.A(g24003),.B(I32355));
  NAND2 NAND2_1436(.VSS(VSS),.VDD(VDD),.Y(g24801),.A(I32356),.B(I32357));
  NAND2 NAND2_1437(.VSS(VSS),.VDD(VDD),.Y(I32368),.A(g18038),.B(g24012));
  NAND2 NAND2_1438(.VSS(VSS),.VDD(VDD),.Y(I32369),.A(g18038),.B(I32368));
  NAND2 NAND2_1439(.VSS(VSS),.VDD(VDD),.Y(I32370),.A(g24012),.B(I32368));
  NAND2 NAND2_1440(.VSS(VSS),.VDD(VDD),.Y(g24808),.A(I32369),.B(I32370));
  NAND2 NAND2_1441(.VSS(VSS),.VDD(VDD),.Y(I32378),.A(g18247),.B(g24027));
  NAND2 NAND2_1442(.VSS(VSS),.VDD(VDD),.Y(I32379),.A(g18247),.B(I32378));
  NAND2 NAND2_1443(.VSS(VSS),.VDD(VDD),.Y(I32380),.A(g24027),.B(I32378));
  NAND2 NAND2_1444(.VSS(VSS),.VDD(VDD),.Y(g24812),.A(I32379),.B(I32380));
  NAND2 NAND2_1445(.VSS(VSS),.VDD(VDD),.Y(g24814),.A(g24239),.B(g24244));
  NAND2 NAND2_1446(.VSS(VSS),.VDD(VDD),.Y(I32391),.A(g17903),.B(g24034));
  NAND2 NAND2_1447(.VSS(VSS),.VDD(VDD),.Y(I32392),.A(g17903),.B(I32391));
  NAND2 NAND2_1448(.VSS(VSS),.VDD(VDD),.Y(I32393),.A(g24034),.B(I32391));
  NAND2 NAND2_1449(.VSS(VSS),.VDD(VDD),.Y(g24817),.A(I32392),.B(I32393));
  NAND2 NAND2_1450(.VSS(VSS),.VDD(VDD),.Y(I32400),.A(g17927),.B(g24036));
  NAND2 NAND2_1451(.VSS(VSS),.VDD(VDD),.Y(I32401),.A(g17927),.B(I32400));
  NAND2 NAND2_1452(.VSS(VSS),.VDD(VDD),.Y(I32402),.A(g24036),.B(I32400));
  NAND2 NAND2_1453(.VSS(VSS),.VDD(VDD),.Y(g24820),.A(I32401),.B(I32402));
  NAND2 NAND2_1454(.VSS(VSS),.VDD(VDD),.Y(I32409),.A(g18131),.B(g24037));
  NAND2 NAND2_1455(.VSS(VSS),.VDD(VDD),.Y(I32410),.A(g18131),.B(I32409));
  NAND2 NAND2_1456(.VSS(VSS),.VDD(VDD),.Y(I32411),.A(g24037),.B(I32409));
  NAND2 NAND2_1457(.VSS(VSS),.VDD(VDD),.Y(g24823),.A(I32410),.B(I32411));
  NAND2 NAND2_1458(.VSS(VSS),.VDD(VDD),.Y(I32422),.A(g18155),.B(g24046));
  NAND2 NAND2_1459(.VSS(VSS),.VDD(VDD),.Y(I32423),.A(g18155),.B(I32422));
  NAND2 NAND2_1460(.VSS(VSS),.VDD(VDD),.Y(I32424),.A(g24046),.B(I32422));
  NAND2 NAND2_1461(.VSS(VSS),.VDD(VDD),.Y(g24830),.A(I32423),.B(I32424));
  NAND2 NAND2_1462(.VSS(VSS),.VDD(VDD),.Y(I32430),.A(g17815),.B(g24052));
  NAND2 NAND2_1463(.VSS(VSS),.VDD(VDD),.Y(I32431),.A(g17815),.B(I32430));
  NAND2 NAND2_1464(.VSS(VSS),.VDD(VDD),.Y(I32432),.A(g24052),.B(I32430));
  NAND2 NAND2_1465(.VSS(VSS),.VDD(VDD),.Y(g24832),.A(I32431),.B(I32432));
  NAND2 NAND2_1466(.VSS(VSS),.VDD(VDD),.Y(g24833),.A(g24245),.B(g24252));
  NAND2 NAND2_1467(.VSS(VSS),.VDD(VDD),.Y(I32443),.A(g18014),.B(g24054));
  NAND2 NAND2_1468(.VSS(VSS),.VDD(VDD),.Y(I32444),.A(g18014),.B(I32443));
  NAND2 NAND2_1469(.VSS(VSS),.VDD(VDD),.Y(I32445),.A(g24054),.B(I32443));
  NAND2 NAND2_1470(.VSS(VSS),.VDD(VDD),.Y(g24837),.A(I32444),.B(I32445));
  NAND2 NAND2_1471(.VSS(VSS),.VDD(VDD),.Y(I32451),.A(g18038),.B(g24056));
  NAND2 NAND2_1472(.VSS(VSS),.VDD(VDD),.Y(I32452),.A(g18038),.B(I32451));
  NAND2 NAND2_1473(.VSS(VSS),.VDD(VDD),.Y(I32453),.A(g24056),.B(I32451));
  NAND2 NAND2_1474(.VSS(VSS),.VDD(VDD),.Y(g24839),.A(I32452),.B(I32453));
  NAND2 NAND2_1475(.VSS(VSS),.VDD(VDD),.Y(I32460),.A(g18247),.B(g24057));
  NAND2 NAND2_1476(.VSS(VSS),.VDD(VDD),.Y(I32461),.A(g18247),.B(I32460));
  NAND2 NAND2_1477(.VSS(VSS),.VDD(VDD),.Y(I32462),.A(g24057),.B(I32460));
  NAND2 NAND2_1478(.VSS(VSS),.VDD(VDD),.Y(g24842),.A(I32461),.B(I32462));
  NAND2 NAND2_1479(.VSS(VSS),.VDD(VDD),.Y(I32468),.A(g17903),.B(g24058));
  NAND2 NAND2_1480(.VSS(VSS),.VDD(VDD),.Y(I32469),.A(g17903),.B(I32468));
  NAND2 NAND2_1481(.VSS(VSS),.VDD(VDD),.Y(I32470),.A(g24058),.B(I32468));
  NAND2 NAND2_1482(.VSS(VSS),.VDD(VDD),.Y(g24844),.A(I32469),.B(I32470));
  NAND2 NAND2_1483(.VSS(VSS),.VDD(VDD),.Y(I32478),.A(g17927),.B(g24065));
  NAND2 NAND2_1484(.VSS(VSS),.VDD(VDD),.Y(I32479),.A(g17927),.B(I32478));
  NAND2 NAND2_1485(.VSS(VSS),.VDD(VDD),.Y(I32480),.A(g24065),.B(I32478));
  NAND2 NAND2_1486(.VSS(VSS),.VDD(VDD),.Y(g24848),.A(I32479),.B(I32480));
  NAND2 NAND2_1487(.VSS(VSS),.VDD(VDD),.Y(g24849),.A(g24254),.B(g24257));
  NAND2 NAND2_1488(.VSS(VSS),.VDD(VDD),.Y(I32490),.A(g18131),.B(g24067));
  NAND2 NAND2_1489(.VSS(VSS),.VDD(VDD),.Y(I32491),.A(g18131),.B(I32490));
  NAND2 NAND2_1490(.VSS(VSS),.VDD(VDD),.Y(I32492),.A(g24067),.B(I32490));
  NAND2 NAND2_1491(.VSS(VSS),.VDD(VDD),.Y(g24852),.A(I32491),.B(I32492));
  NAND2 NAND2_1492(.VSS(VSS),.VDD(VDD),.Y(I32498),.A(g18155),.B(g24069));
  NAND2 NAND2_1493(.VSS(VSS),.VDD(VDD),.Y(I32499),.A(g18155),.B(I32498));
  NAND2 NAND2_1494(.VSS(VSS),.VDD(VDD),.Y(I32500),.A(g24069),.B(I32498));
  NAND2 NAND2_1495(.VSS(VSS),.VDD(VDD),.Y(g24854),.A(I32499),.B(I32500));
  NAND2 NAND2_1496(.VSS(VSS),.VDD(VDD),.Y(I32509),.A(g17815),.B(g24070));
  NAND2 NAND2_1497(.VSS(VSS),.VDD(VDD),.Y(I32510),.A(g17815),.B(I32509));
  NAND2 NAND2_1498(.VSS(VSS),.VDD(VDD),.Y(I32511),.A(g24070),.B(I32509));
  NAND2 NAND2_1499(.VSS(VSS),.VDD(VDD),.Y(g24857),.A(I32510),.B(I32511));
  NAND2 NAND2_1500(.VSS(VSS),.VDD(VDD),.Y(I32518),.A(g18014),.B(g24071));
  NAND2 NAND2_1501(.VSS(VSS),.VDD(VDD),.Y(I32519),.A(g18014),.B(I32518));
  NAND2 NAND2_1502(.VSS(VSS),.VDD(VDD),.Y(I32520),.A(g24071),.B(I32518));
  NAND2 NAND2_1503(.VSS(VSS),.VDD(VDD),.Y(g24860),.A(I32519),.B(I32520));
  NAND2 NAND2_1504(.VSS(VSS),.VDD(VDD),.Y(I32526),.A(g18038),.B(g24078));
  NAND2 NAND2_1505(.VSS(VSS),.VDD(VDD),.Y(I32527),.A(g18038),.B(I32526));
  NAND2 NAND2_1506(.VSS(VSS),.VDD(VDD),.Y(I32528),.A(g24078),.B(I32526));
  NAND2 NAND2_1507(.VSS(VSS),.VDD(VDD),.Y(g24862),.A(I32527),.B(I32528));
  NAND2 NAND2_1508(.VSS(VSS),.VDD(VDD),.Y(g24863),.A(g24258),.B(g23319));
  NAND2 NAND2_1509(.VSS(VSS),.VDD(VDD),.Y(I32538),.A(g18247),.B(g24080));
  NAND2 NAND2_1510(.VSS(VSS),.VDD(VDD),.Y(I32539),.A(g18247),.B(I32538));
  NAND2 NAND2_1511(.VSS(VSS),.VDD(VDD),.Y(I32540),.A(g24080),.B(I32538));
  NAND2 NAND2_1512(.VSS(VSS),.VDD(VDD),.Y(g24866),.A(I32539),.B(I32540));
  NAND2 NAND2_1513(.VSS(VSS),.VDD(VDD),.Y(I32546),.A(g17903),.B(g23906));
  NAND2 NAND2_1514(.VSS(VSS),.VDD(VDD),.Y(I32547),.A(g17903),.B(I32546));
  NAND2 NAND2_1515(.VSS(VSS),.VDD(VDD),.Y(I32548),.A(g23906),.B(I32546));
  NAND2 NAND2_1516(.VSS(VSS),.VDD(VDD),.Y(g24868),.A(I32547),.B(I32548));
  NAND2 NAND2_1517(.VSS(VSS),.VDD(VDD),.Y(I32559),.A(g17927),.B(g24081));
  NAND2 NAND2_1518(.VSS(VSS),.VDD(VDD),.Y(I32560),.A(g17927),.B(I32559));
  NAND2 NAND2_1519(.VSS(VSS),.VDD(VDD),.Y(I32561),.A(g24081),.B(I32559));
  NAND2 NAND2_1520(.VSS(VSS),.VDD(VDD),.Y(g24873),.A(I32560),.B(I32561));
  NAND2 NAND2_1521(.VSS(VSS),.VDD(VDD),.Y(I32567),.A(g18131),.B(g24082));
  NAND2 NAND2_1522(.VSS(VSS),.VDD(VDD),.Y(I32568),.A(g18131),.B(I32567));
  NAND2 NAND2_1523(.VSS(VSS),.VDD(VDD),.Y(I32569),.A(g24082),.B(I32567));
  NAND2 NAND2_1524(.VSS(VSS),.VDD(VDD),.Y(g24875),.A(I32568),.B(I32569));
  NAND2 NAND2_1525(.VSS(VSS),.VDD(VDD),.Y(I32575),.A(g18155),.B(g24089));
  NAND2 NAND2_1526(.VSS(VSS),.VDD(VDD),.Y(I32576),.A(g18155),.B(I32575));
  NAND2 NAND2_1527(.VSS(VSS),.VDD(VDD),.Y(I32577),.A(g24089),.B(I32575));
  NAND2 NAND2_1528(.VSS(VSS),.VDD(VDD),.Y(g24877),.A(I32576),.B(I32577));
  NAND2 NAND2_1529(.VSS(VSS),.VDD(VDD),.Y(I32586),.A(g17815),.B(g23937));
  NAND2 NAND2_1530(.VSS(VSS),.VDD(VDD),.Y(I32587),.A(g17815),.B(I32586));
  NAND2 NAND2_1531(.VSS(VSS),.VDD(VDD),.Y(I32588),.A(g23937),.B(I32586));
  NAND2 NAND2_1532(.VSS(VSS),.VDD(VDD),.Y(g24880),.A(I32587),.B(I32588));
  NAND2 NAND2_1533(.VSS(VSS),.VDD(VDD),.Y(I32595),.A(g18014),.B(g23938));
  NAND2 NAND2_1534(.VSS(VSS),.VDD(VDD),.Y(I32596),.A(g18014),.B(I32595));
  NAND2 NAND2_1535(.VSS(VSS),.VDD(VDD),.Y(I32597),.A(g23938),.B(I32595));
  NAND2 NAND2_1536(.VSS(VSS),.VDD(VDD),.Y(g24883),.A(I32596),.B(I32597));
  NAND2 NAND2_1537(.VSS(VSS),.VDD(VDD),.Y(I32607),.A(g18038),.B(g24090));
  NAND2 NAND2_1538(.VSS(VSS),.VDD(VDD),.Y(I32608),.A(g18038),.B(I32607));
  NAND2 NAND2_1539(.VSS(VSS),.VDD(VDD),.Y(I32609),.A(g24090),.B(I32607));
  NAND2 NAND2_1540(.VSS(VSS),.VDD(VDD),.Y(g24887),.A(I32608),.B(I32609));
  NAND2 NAND2_1541(.VSS(VSS),.VDD(VDD),.Y(I32615),.A(g18247),.B(g24091));
  NAND2 NAND2_1542(.VSS(VSS),.VDD(VDD),.Y(I32616),.A(g18247),.B(I32615));
  NAND2 NAND2_1543(.VSS(VSS),.VDD(VDD),.Y(I32617),.A(g24091),.B(I32615));
  NAND2 NAND2_1544(.VSS(VSS),.VDD(VDD),.Y(g24889),.A(I32616),.B(I32617));
  NAND2 NAND2_1545(.VSS(VSS),.VDD(VDD),.Y(I32624),.A(g17927),.B(g23969));
  NAND2 NAND2_1546(.VSS(VSS),.VDD(VDD),.Y(I32625),.A(g17927),.B(I32624));
  NAND2 NAND2_1547(.VSS(VSS),.VDD(VDD),.Y(I32626),.A(g23969),.B(I32624));
  NAND2 NAND2_1548(.VSS(VSS),.VDD(VDD),.Y(g24897),.A(I32625),.B(I32626));
  NAND2 NAND2_1549(.VSS(VSS),.VDD(VDD),.Y(I32633),.A(g18131),.B(g23970));
  NAND2 NAND2_1550(.VSS(VSS),.VDD(VDD),.Y(I32634),.A(g18131),.B(I32633));
  NAND2 NAND2_1551(.VSS(VSS),.VDD(VDD),.Y(I32635),.A(g23970),.B(I32633));
  NAND2 NAND2_1552(.VSS(VSS),.VDD(VDD),.Y(g24900),.A(I32634),.B(I32635));
  NAND2 NAND2_1553(.VSS(VSS),.VDD(VDD),.Y(I32645),.A(g18155),.B(g24093));
  NAND2 NAND2_1554(.VSS(VSS),.VDD(VDD),.Y(I32646),.A(g18155),.B(I32645));
  NAND2 NAND2_1555(.VSS(VSS),.VDD(VDD),.Y(I32647),.A(g24093),.B(I32645));
  NAND2 NAND2_1556(.VSS(VSS),.VDD(VDD),.Y(g24904),.A(I32646),.B(I32647));
  NAND2 NAND2_1557(.VSS(VSS),.VDD(VDD),.Y(I32659),.A(g18038),.B(g23998));
  NAND2 NAND2_1558(.VSS(VSS),.VDD(VDD),.Y(I32660),.A(g18038),.B(I32659));
  NAND2 NAND2_1559(.VSS(VSS),.VDD(VDD),.Y(I32661),.A(g23998),.B(I32659));
  NAND2 NAND2_1560(.VSS(VSS),.VDD(VDD),.Y(g24920),.A(I32660),.B(I32661));
  NAND2 NAND2_1561(.VSS(VSS),.VDD(VDD),.Y(I32668),.A(g18247),.B(g23999));
  NAND2 NAND2_1562(.VSS(VSS),.VDD(VDD),.Y(I32669),.A(g18247),.B(I32668));
  NAND2 NAND2_1563(.VSS(VSS),.VDD(VDD),.Y(I32670),.A(g23999),.B(I32668));
  NAND2 NAND2_1564(.VSS(VSS),.VDD(VDD),.Y(g24923),.A(I32669),.B(I32670));
  NAND2 NAND2_1565(.VSS(VSS),.VDD(VDD),.Y(I32677),.A(g23823),.B(g14165));
  NAND2 NAND2_1566(.VSS(VSS),.VDD(VDD),.Y(I32678),.A(g23823),.B(I32677));
  NAND2 NAND2_1567(.VSS(VSS),.VDD(VDD),.Y(I32679),.A(g14165),.B(I32677));
  NAND2 NAND2_1568(.VSS(VSS),.VDD(VDD),.Y(g24928),.A(I32678),.B(I32679));
  NAND2 NAND2_1569(.VSS(VSS),.VDD(VDD),.Y(I32686),.A(g18155),.B(g24028));
  NAND2 NAND2_1570(.VSS(VSS),.VDD(VDD),.Y(I32687),.A(g18155),.B(I32686));
  NAND2 NAND2_1571(.VSS(VSS),.VDD(VDD),.Y(I32688),.A(g24028),.B(I32686));
  NAND2 NAND2_1572(.VSS(VSS),.VDD(VDD),.Y(g24937),.A(I32687),.B(I32688));
  NAND2 NAND2_1573(.VSS(VSS),.VDD(VDD),.Y(I32695),.A(g23858),.B(g14280));
  NAND2 NAND2_1574(.VSS(VSS),.VDD(VDD),.Y(I32696),.A(g23858),.B(I32695));
  NAND2 NAND2_1575(.VSS(VSS),.VDD(VDD),.Y(I32697),.A(g14280),.B(I32695));
  NAND2 NAND2_1576(.VSS(VSS),.VDD(VDD),.Y(g24940),.A(I32696),.B(I32697));
  NAND2 NAND2_1577(.VSS(VSS),.VDD(VDD),.Y(I32708),.A(g23892),.B(g14402));
  NAND2 NAND2_1578(.VSS(VSS),.VDD(VDD),.Y(I32709),.A(g23892),.B(I32708));
  NAND2 NAND2_1579(.VSS(VSS),.VDD(VDD),.Y(I32710),.A(g14402),.B(I32708));
  NAND2 NAND2_1580(.VSS(VSS),.VDD(VDD),.Y(g24951),.A(I32709),.B(I32710));
  NAND2 NAND2_1581(.VSS(VSS),.VDD(VDD),.Y(I32724),.A(g23913),.B(g14514));
  NAND2 NAND2_1582(.VSS(VSS),.VDD(VDD),.Y(I32725),.A(g23913),.B(I32724));
  NAND2 NAND2_1583(.VSS(VSS),.VDD(VDD),.Y(I32726),.A(g14514),.B(I32724));
  NAND2 NAND2_1584(.VSS(VSS),.VDD(VDD),.Y(g24963),.A(I32725),.B(I32726));
  NAND2 NAND2_1585(.VSS(VSS),.VDD(VDD),.Y(g24975),.A(g23497),.B(g74));
  NAND2 NAND2_1586(.VSS(VSS),.VDD(VDD),.Y(g24986),.A(g23513),.B(g762));
  NAND2 NAND2_1587(.VSS(VSS),.VDD(VDD),.Y(g24997),.A(g23528),.B(g1448));
  NAND2 NAND2_1588(.VSS(VSS),.VDD(VDD),.Y(g25004),.A(g23644),.B(g6448));
  NAND2 NAND2_1589(.VSS(VSS),.VDD(VDD),.Y(g25005),.A(g23539),.B(g2142));
  NAND2 NAND2_1590(.VSS(VSS),.VDD(VDD),.Y(g25008),.A(g23644),.B(g5438));
  NAND2 NAND2_1591(.VSS(VSS),.VDD(VDD),.Y(g25009),.A(g23644),.B(g6448));
  NAND2 NAND2_1592(.VSS(VSS),.VDD(VDD),.Y(g25010),.A(g23694),.B(g6713));
  NAND2 NAND2_1593(.VSS(VSS),.VDD(VDD),.Y(g25011),.A(g23644),.B(g5438));
  NAND2 NAND2_1594(.VSS(VSS),.VDD(VDD),.Y(g25012),.A(g23644),.B(g6448));
  NAND2 NAND2_1595(.VSS(VSS),.VDD(VDD),.Y(g25013),.A(g23923),.B(g6643));
  NAND2 NAND2_1596(.VSS(VSS),.VDD(VDD),.Y(g25014),.A(g23694),.B(g5473));
  NAND2 NAND2_1597(.VSS(VSS),.VDD(VDD),.Y(g25015),.A(g23694),.B(g6713));
  NAND2 NAND2_1598(.VSS(VSS),.VDD(VDD),.Y(g25016),.A(g23748),.B(g7015));
  NAND2 NAND2_1599(.VSS(VSS),.VDD(VDD),.Y(g25017),.A(g23644),.B(g5438));
  NAND2 NAND2_1600(.VSS(VSS),.VDD(VDD),.Y(g25018),.A(g23644),.B(g6448));
  NAND2 NAND2_1601(.VSS(VSS),.VDD(VDD),.Y(g25019),.A(g23923),.B(g6486));
  NAND2 NAND2_1602(.VSS(VSS),.VDD(VDD),.Y(g25020),.A(g23923),.B(g6643));
  NAND2 NAND2_1603(.VSS(VSS),.VDD(VDD),.Y(g25021),.A(g23694),.B(g5473));
  NAND2 NAND2_1604(.VSS(VSS),.VDD(VDD),.Y(g25022),.A(g23694),.B(g6713));
  NAND2 NAND2_1605(.VSS(VSS),.VDD(VDD),.Y(g25023),.A(g23955),.B(g6945));
  NAND2 NAND2_1606(.VSS(VSS),.VDD(VDD),.Y(g25024),.A(g23748),.B(g5512));
  NAND2 NAND2_1607(.VSS(VSS),.VDD(VDD),.Y(g25025),.A(g23748),.B(g7015));
  NAND2 NAND2_1608(.VSS(VSS),.VDD(VDD),.Y(g25026),.A(g23803),.B(g7265));
  NAND2 NAND2_1609(.VSS(VSS),.VDD(VDD),.Y(g25028),.A(g23644),.B(g5438));
  NAND2 NAND2_1610(.VSS(VSS),.VDD(VDD),.Y(g25029),.A(g23923),.B(g6486));
  NAND2 NAND2_1611(.VSS(VSS),.VDD(VDD),.Y(g25030),.A(g23923),.B(g6643));
  NAND2 NAND2_1612(.VSS(VSS),.VDD(VDD),.Y(g25031),.A(g23694),.B(g5473));
  NAND2 NAND2_1613(.VSS(VSS),.VDD(VDD),.Y(g25032),.A(g23694),.B(g6713));
  NAND2 NAND2_1614(.VSS(VSS),.VDD(VDD),.Y(g25033),.A(g23955),.B(g6751));
  NAND2 NAND2_1615(.VSS(VSS),.VDD(VDD),.Y(g25034),.A(g23955),.B(g6945));
  NAND2 NAND2_1616(.VSS(VSS),.VDD(VDD),.Y(g25035),.A(g23748),.B(g5512));
  NAND2 NAND2_1617(.VSS(VSS),.VDD(VDD),.Y(g25036),.A(g23748),.B(g7015));
  NAND2 NAND2_1618(.VSS(VSS),.VDD(VDD),.Y(g25037),.A(g23984),.B(g7195));
  NAND2 NAND2_1619(.VSS(VSS),.VDD(VDD),.Y(g25038),.A(g23803),.B(g5556));
  NAND2 NAND2_1620(.VSS(VSS),.VDD(VDD),.Y(g25039),.A(g23803),.B(g7265));
  NAND2 NAND2_1621(.VSS(VSS),.VDD(VDD),.Y(g25040),.A(g23923),.B(g6486));
  NAND2 NAND2_1622(.VSS(VSS),.VDD(VDD),.Y(g25041),.A(g23923),.B(g6643));
  NAND2 NAND2_1623(.VSS(VSS),.VDD(VDD),.Y(g25043),.A(g23694),.B(g5473));
  NAND2 NAND2_1624(.VSS(VSS),.VDD(VDD),.Y(g25044),.A(g23955),.B(g6751));
  NAND2 NAND2_1625(.VSS(VSS),.VDD(VDD),.Y(g25045),.A(g23955),.B(g6945));
  NAND2 NAND2_1626(.VSS(VSS),.VDD(VDD),.Y(g25046),.A(g23748),.B(g5512));
  NAND2 NAND2_1627(.VSS(VSS),.VDD(VDD),.Y(g25047),.A(g23748),.B(g7015));
  NAND2 NAND2_1628(.VSS(VSS),.VDD(VDD),.Y(g25048),.A(g23984),.B(g7053));
  NAND2 NAND2_1629(.VSS(VSS),.VDD(VDD),.Y(g25049),.A(g23984),.B(g7195));
  NAND2 NAND2_1630(.VSS(VSS),.VDD(VDD),.Y(g25050),.A(g23803),.B(g5556));
  NAND2 NAND2_1631(.VSS(VSS),.VDD(VDD),.Y(g25051),.A(g23803),.B(g7265));
  NAND2 NAND2_1632(.VSS(VSS),.VDD(VDD),.Y(g25052),.A(g24014),.B(g7391));
  NAND2 NAND2_1633(.VSS(VSS),.VDD(VDD),.Y(g25053),.A(g23923),.B(g6486));
  NAND2 NAND2_1634(.VSS(VSS),.VDD(VDD),.Y(g25054),.A(g23955),.B(g6751));
  NAND2 NAND2_1635(.VSS(VSS),.VDD(VDD),.Y(g25055),.A(g23955),.B(g6945));
  NAND2 NAND2_1636(.VSS(VSS),.VDD(VDD),.Y(g25057),.A(g23748),.B(g5512));
  NAND2 NAND2_1637(.VSS(VSS),.VDD(VDD),.Y(g25058),.A(g23984),.B(g7053));
  NAND2 NAND2_1638(.VSS(VSS),.VDD(VDD),.Y(g25059),.A(g23984),.B(g7195));
  NAND2 NAND2_1639(.VSS(VSS),.VDD(VDD),.Y(g25060),.A(g23803),.B(g5556));
  NAND2 NAND2_1640(.VSS(VSS),.VDD(VDD),.Y(g25061),.A(g23803),.B(g7265));
  NAND2 NAND2_1641(.VSS(VSS),.VDD(VDD),.Y(g25062),.A(g24014),.B(g7303));
  NAND2 NAND2_1642(.VSS(VSS),.VDD(VDD),.Y(g25063),.A(g24014),.B(g7391));
  NAND2 NAND2_1643(.VSS(VSS),.VDD(VDD),.Y(g25064),.A(g23955),.B(g6751));
  NAND2 NAND2_1644(.VSS(VSS),.VDD(VDD),.Y(g25065),.A(g23984),.B(g7053));
  NAND2 NAND2_1645(.VSS(VSS),.VDD(VDD),.Y(g25066),.A(g23984),.B(g7195));
  NAND2 NAND2_1646(.VSS(VSS),.VDD(VDD),.Y(g25068),.A(g23803),.B(g5556));
  NAND2 NAND2_1647(.VSS(VSS),.VDD(VDD),.Y(g25069),.A(g24014),.B(g7303));
  NAND2 NAND2_1648(.VSS(VSS),.VDD(VDD),.Y(g25070),.A(g24014),.B(g7391));
  NAND2 NAND2_1649(.VSS(VSS),.VDD(VDD),.Y(g25071),.A(g23984),.B(g7053));
  NAND2 NAND2_1650(.VSS(VSS),.VDD(VDD),.Y(g25072),.A(g24014),.B(g7303));
  NAND2 NAND2_1651(.VSS(VSS),.VDD(VDD),.Y(g25073),.A(g24014),.B(g7391));
  NAND2 NAND2_1652(.VSS(VSS),.VDD(VDD),.Y(g25074),.A(g24014),.B(g7303));
  NAND2 NAND2_1653(.VSS(VSS),.VDD(VDD),.Y(g25088),.A(g23950),.B(g679));
  NAND2 NAND2_1654(.VSS(VSS),.VDD(VDD),.Y(g25096),.A(g23979),.B(g1365));
  NAND2 NAND2_1655(.VSS(VSS),.VDD(VDD),.Y(g25106),.A(g24009),.B(g2059));
  NAND2 NAND2_1656(.VSS(VSS),.VDD(VDD),.Y(g25112),.A(g24043),.B(g2753));
  NAND2 NAND2_1657(.VSS(VSS),.VDD(VDD),.Y(g25200),.A(g24965),.B(g3306));
  NAND2 NAND2_1658(.VSS(VSS),.VDD(VDD),.Y(g25203),.A(g24978),.B(g3462));
  NAND2 NAND2_1659(.VSS(VSS),.VDD(VDD),.Y(g25205),.A(g24989),.B(g3618));
  NAND2 NAND2_1660(.VSS(VSS),.VDD(VDD),.Y(g25210),.A(g25000),.B(g3774));
  NAND4 NAND4_5(.VSS(VSS),.VDD(VDD),.Y(g25312),.A(g21211),.B(g14442),.C(g10694),.D(g24590));
  NAND4 NAND4_6(.VSS(VSS),.VDD(VDD),.Y(g25320),.A(g21219),.B(g14529),.C(g10714),.D(g24595));
  NAND4 NAND4_7(.VSS(VSS),.VDD(VDD),.Y(g25331),.A(g21230),.B(g14584),.C(g10735),.D(g24603));
  NAND4 NAND4_8(.VSS(VSS),.VDD(VDD),.Y(g25340),.A(g21235),.B(g14618),.C(g10754),.D(g24610));
  NAND2 NAND2_1661(.VSS(VSS),.VDD(VDD),.Y(g25927),.A(g24965),.B(g6448));
  NAND2 NAND2_1662(.VSS(VSS),.VDD(VDD),.Y(g25928),.A(g24965),.B(g5438));
  NAND2 NAND2_1663(.VSS(VSS),.VDD(VDD),.Y(g25929),.A(g24978),.B(g6713));
  NAND2 NAND2_1664(.VSS(VSS),.VDD(VDD),.Y(g25930),.A(g24978),.B(g5473));
  NAND2 NAND2_1665(.VSS(VSS),.VDD(VDD),.Y(g25931),.A(g24989),.B(g7015));
  NAND2 NAND2_1666(.VSS(VSS),.VDD(VDD),.Y(g25933),.A(g24989),.B(g5512));
  NAND2 NAND2_1667(.VSS(VSS),.VDD(VDD),.Y(g25934),.A(g25000),.B(g7265));
  NAND2 NAND2_1668(.VSS(VSS),.VDD(VDD),.Y(g25936),.A(g25000),.B(g5556));
  NAND2 NAND2_1669(.VSS(VSS),.VDD(VDD),.Y(g25954),.A(g22806),.B(g24517));
  NAND2 NAND2_1670(.VSS(VSS),.VDD(VDD),.Y(g25958),.A(g22847),.B(g24530));
  NAND2 NAND2_1671(.VSS(VSS),.VDD(VDD),.Y(g25964),.A(g22882),.B(g24543));
  NAND2 NAND2_1672(.VSS(VSS),.VDD(VDD),.Y(g25969),.A(g22917),.B(g24555));
  NAND3 NAND3_76(.VSS(VSS),.VDD(VDD),.Y(g26059),.A(g25422),.B(g25379),.C(g25274));
  NAND3 NAND3_77(.VSS(VSS),.VDD(VDD),.Y(g26066),.A(g25431),.B(g25395),.C(g25283));
  NAND3 NAND3_78(.VSS(VSS),.VDD(VDD),.Y(g26073),.A(g25438),.B(g25405),.C(g25291));
  NAND3 NAND3_79(.VSS(VSS),.VDD(VDD),.Y(g26079),.A(g25445),.B(g25413),.C(g25301));
  NAND2 NAND2_1673(.VSS(VSS),.VDD(VDD),.Y(g26106),.A(g23644),.B(g25354));
  NAND4 NAND4_9(.VSS(VSS),.VDD(VDD),.Y(g26119),.A(g8278),.B(g14657),.C(g25422),.D(g25379));
  NAND2 NAND2_1674(.VSS(VSS),.VDD(VDD),.Y(g26120),.A(g23694),.B(g25369));
  NAND4 NAND4_10(.VSS(VSS),.VDD(VDD),.Y(g26129),.A(g8287),.B(g14691),.C(g25431),.D(g25395));
  NAND2 NAND2_1675(.VSS(VSS),.VDD(VDD),.Y(g26130),.A(g23748),.B(g25386));
  NAND4 NAND4_11(.VSS(VSS),.VDD(VDD),.Y(g26143),.A(g8296),.B(g14725),.C(g25438),.D(g25405));
  NAND2 NAND2_1676(.VSS(VSS),.VDD(VDD),.Y(g26144),.A(g23803),.B(g25402));
  NAND4 NAND4_12(.VSS(VSS),.VDD(VDD),.Y(g26148),.A(g8305),.B(g14753),.C(g25445),.D(g25413));
  NAND2 NAND2_1677(.VSS(VSS),.VDD(VDD),.Y(g26356),.A(g16539),.B(g25183));
  NAND2 NAND2_1678(.VSS(VSS),.VDD(VDD),.Y(g26399),.A(g16571),.B(g25186));
  NAND2 NAND2_1679(.VSS(VSS),.VDD(VDD),.Y(g26440),.A(g16595),.B(g25190));
  NAND2 NAND2_1680(.VSS(VSS),.VDD(VDD),.Y(g26458),.A(g25343),.B(g65));
  NAND2 NAND2_1681(.VSS(VSS),.VDD(VDD),.Y(g26472),.A(g16615),.B(g25195));
  NAND2 NAND2_1682(.VSS(VSS),.VDD(VDD),.Y(g26482),.A(g25357),.B(g753));
  NAND2 NAND2_1683(.VSS(VSS),.VDD(VDD),.Y(g26498),.A(g25372),.B(g1439));
  NAND2 NAND2_1684(.VSS(VSS),.VDD(VDD),.Y(g26513),.A(g25389),.B(g2133));
  NAND2 NAND2_1685(.VSS(VSS),.VDD(VDD),.Y(g26772),.A(g26320),.B(g3306));
  NAND2 NAND2_1686(.VSS(VSS),.VDD(VDD),.Y(g26779),.A(g26367),.B(g3462));
  NAND2 NAND2_1687(.VSS(VSS),.VDD(VDD),.Y(g26785),.A(g26410),.B(g3618));
  NAND2 NAND2_1688(.VSS(VSS),.VDD(VDD),.Y(g26792),.A(g26451),.B(g3774));
  NAND2 NAND2_1689(.VSS(VSS),.VDD(VDD),.Y(I35020),.A(g26110),.B(g26099));
  NAND2 NAND2_1690(.VSS(VSS),.VDD(VDD),.Y(I35021),.A(g26110),.B(I35020));
  NAND2 NAND2_1691(.VSS(VSS),.VDD(VDD),.Y(I35022),.A(g26099),.B(I35020));
  NAND2 NAND2_1692(.VSS(VSS),.VDD(VDD),.Y(g26859),.A(I35021),.B(I35022));
  NAND2 NAND2_1693(.VSS(VSS),.VDD(VDD),.Y(I35034),.A(g26087),.B(g26154));
  NAND2 NAND2_1694(.VSS(VSS),.VDD(VDD),.Y(I35035),.A(g26087),.B(I35034));
  NAND2 NAND2_1695(.VSS(VSS),.VDD(VDD),.Y(I35036),.A(g26154),.B(I35034));
  NAND2 NAND2_1696(.VSS(VSS),.VDD(VDD),.Y(g26865),.A(I35035),.B(I35036));
  NAND2 NAND2_1697(.VSS(VSS),.VDD(VDD),.Y(I35042),.A(g26151),.B(g26145));
  NAND2 NAND2_1698(.VSS(VSS),.VDD(VDD),.Y(I35043),.A(g26151),.B(I35042));
  NAND2 NAND2_1699(.VSS(VSS),.VDD(VDD),.Y(I35044),.A(g26145),.B(I35042));
  NAND2 NAND2_1700(.VSS(VSS),.VDD(VDD),.Y(g26867),.A(I35043),.B(I35044));
  NAND2 NAND2_1701(.VSS(VSS),.VDD(VDD),.Y(I35057),.A(g26137),.B(g26126));
  NAND2 NAND2_1702(.VSS(VSS),.VDD(VDD),.Y(I35058),.A(g26137),.B(I35057));
  NAND2 NAND2_1703(.VSS(VSS),.VDD(VDD),.Y(I35059),.A(g26126),.B(I35057));
  NAND2 NAND2_1704(.VSS(VSS),.VDD(VDD),.Y(g26874),.A(I35058),.B(I35059));
  NAND4 NAND4_13(.VSS(VSS),.VDD(VDD),.Y(g26892),.A(g25699),.B(g26283),.C(g25569),.D(g25631));
  NAND3 NAND3_80(.VSS(VSS),.VDD(VDD),.Y(g26902),.A(g25631),.B(g26283),.C(g25569));
  NAND4 NAND4_14(.VSS(VSS),.VDD(VDD),.Y(g26906),.A(g25772),.B(g26327),.C(g25648),.D(g25708));
  NAND2 NAND2_1705(.VSS(VSS),.VDD(VDD),.Y(g26911),.A(g25569),.B(g26283));
  NAND3 NAND3_81(.VSS(VSS),.VDD(VDD),.Y(g26915),.A(g25708),.B(g26327),.C(g25648));
  NAND4 NAND4_15(.VSS(VSS),.VDD(VDD),.Y(g26918),.A(g25826),.B(g26374),.C(g25725),.D(g25781));
  NAND2 NAND2_1706(.VSS(VSS),.VDD(VDD),.Y(g26925),.A(g25648),.B(g26327));
  NAND3 NAND3_82(.VSS(VSS),.VDD(VDD),.Y(g26928),.A(g25781),.B(g26374),.C(g25725));
  NAND4 NAND4_16(.VSS(VSS),.VDD(VDD),.Y(g26931),.A(g25861),.B(g26417),.C(g25798),.D(g25835));
  NAND2 NAND2_1707(.VSS(VSS),.VDD(VDD),.Y(I35123),.A(g26107),.B(g26096));
  NAND2 NAND2_1708(.VSS(VSS),.VDD(VDD),.Y(I35124),.A(g26107),.B(I35123));
  NAND2 NAND2_1709(.VSS(VSS),.VDD(VDD),.Y(I35125),.A(g26096),.B(I35123));
  NAND2 NAND2_1710(.VSS(VSS),.VDD(VDD),.Y(g26934),.A(I35124),.B(I35125));
  NAND2 NAND2_1711(.VSS(VSS),.VDD(VDD),.Y(g26938),.A(g25725),.B(g26374));
  NAND3 NAND3_83(.VSS(VSS),.VDD(VDD),.Y(g26941),.A(g25835),.B(g26417),.C(g25798));
  NAND2 NAND2_1712(.VSS(VSS),.VDD(VDD),.Y(g26947),.A(g25798),.B(g26417));
  NAND2 NAND2_1713(.VSS(VSS),.VDD(VDD),.Y(g27117),.A(g26320),.B(g6448));
  NAND2 NAND2_1714(.VSS(VSS),.VDD(VDD),.Y(g27118),.A(g26320),.B(g5438));
  NAND2 NAND2_1715(.VSS(VSS),.VDD(VDD),.Y(g27119),.A(g26367),.B(g6713));
  NAND2 NAND2_1716(.VSS(VSS),.VDD(VDD),.Y(g27121),.A(g26367),.B(g5473));
  NAND2 NAND2_1717(.VSS(VSS),.VDD(VDD),.Y(g27122),.A(g26410),.B(g7015));
  NAND2 NAND2_1718(.VSS(VSS),.VDD(VDD),.Y(g27124),.A(g26410),.B(g5512));
  NAND2 NAND2_1719(.VSS(VSS),.VDD(VDD),.Y(g27125),.A(g26451),.B(g7265));
  NAND2 NAND2_1720(.VSS(VSS),.VDD(VDD),.Y(g27130),.A(g26451),.B(g5556));
  NAND2 NAND2_1721(.VSS(VSS),.VDD(VDD),.Y(I35701),.A(g26867),.B(g26874));
  NAND2 NAND2_1722(.VSS(VSS),.VDD(VDD),.Y(I35702),.A(g26867),.B(I35701));
  NAND2 NAND2_1723(.VSS(VSS),.VDD(VDD),.Y(I35703),.A(g26874),.B(I35701));
  NAND2 NAND2_1724(.VSS(VSS),.VDD(VDD),.Y(g27379),.A(I35702),.B(I35703));
  NAND2 NAND2_1725(.VSS(VSS),.VDD(VDD),.Y(I35714),.A(g26859),.B(g26865));
  NAND2 NAND2_1726(.VSS(VSS),.VDD(VDD),.Y(I35715),.A(g26859),.B(I35714));
  NAND2 NAND2_1727(.VSS(VSS),.VDD(VDD),.Y(I35716),.A(g26865),.B(I35714));
  NAND2 NAND2_1728(.VSS(VSS),.VDD(VDD),.Y(g27382),.A(I35715),.B(I35716));
  NAND2 NAND2_1729(.VSS(VSS),.VDD(VDD),.Y(g27390),.A(g26989),.B(g6448));
  NAND2 NAND2_1730(.VSS(VSS),.VDD(VDD),.Y(g27395),.A(g26989),.B(g5438));
  NAND2 NAND2_1731(.VSS(VSS),.VDD(VDD),.Y(g27400),.A(g27012),.B(g6713));
  NAND2 NAND2_1732(.VSS(VSS),.VDD(VDD),.Y(g27408),.A(g27012),.B(g5473));
  NAND2 NAND2_1733(.VSS(VSS),.VDD(VDD),.Y(g27413),.A(g27038),.B(g7015));
  NAND2 NAND2_1734(.VSS(VSS),.VDD(VDD),.Y(g27426),.A(g27038),.B(g5512));
  NAND2 NAND2_1735(.VSS(VSS),.VDD(VDD),.Y(g27431),.A(g27066),.B(g7265));
  NAND2 NAND2_1736(.VSS(VSS),.VDD(VDD),.Y(g27447),.A(g27066),.B(g5556));
  NAND2 NAND2_1737(.VSS(VSS),.VDD(VDD),.Y(I35904),.A(g27051),.B(g14831));
  NAND2 NAND2_1738(.VSS(VSS),.VDD(VDD),.Y(I35905),.A(g27051),.B(I35904));
  NAND2 NAND2_1739(.VSS(VSS),.VDD(VDD),.Y(I35906),.A(g14831),.B(I35904));
  NAND2 NAND2_1740(.VSS(VSS),.VDD(VDD),.Y(g27528),.A(I35905),.B(I35906));
  NAND2 NAND2_1741(.VSS(VSS),.VDD(VDD),.Y(I35944),.A(g27078),.B(g14904));
  NAND2 NAND2_1742(.VSS(VSS),.VDD(VDD),.Y(I35945),.A(g27078),.B(I35944));
  NAND2 NAND2_1743(.VSS(VSS),.VDD(VDD),.Y(I35946),.A(g14904),.B(I35944));
  NAND2 NAND2_1744(.VSS(VSS),.VDD(VDD),.Y(g27550),.A(I35945),.B(I35946));
  NAND2 NAND2_1745(.VSS(VSS),.VDD(VDD),.Y(I35974),.A(g27094),.B(g14985));
  NAND2 NAND2_1746(.VSS(VSS),.VDD(VDD),.Y(I35975),.A(g27094),.B(I35974));
  NAND2 NAND2_1747(.VSS(VSS),.VDD(VDD),.Y(I35976),.A(g14985),.B(I35974));
  NAND2 NAND2_1748(.VSS(VSS),.VDD(VDD),.Y(g27566),.A(I35975),.B(I35976));
  NAND2 NAND2_1749(.VSS(VSS),.VDD(VDD),.Y(g27571),.A(g26869),.B(g56));
  NAND2 NAND2_1750(.VSS(VSS),.VDD(VDD),.Y(I35992),.A(g27106),.B(g15074));
  NAND2 NAND2_1751(.VSS(VSS),.VDD(VDD),.Y(I35993),.A(g27106),.B(I35992));
  NAND2 NAND2_1752(.VSS(VSS),.VDD(VDD),.Y(I35994),.A(g15074),.B(I35992));
  NAND2 NAND2_1753(.VSS(VSS),.VDD(VDD),.Y(g27576),.A(I35993),.B(I35994));
  NAND2 NAND2_1754(.VSS(VSS),.VDD(VDD),.Y(g27580),.A(g26878),.B(g744));
  NAND2 NAND2_1755(.VSS(VSS),.VDD(VDD),.Y(g27583),.A(g26887),.B(g1430));
  NAND2 NAND2_1756(.VSS(VSS),.VDD(VDD),.Y(g27587),.A(g26897),.B(g2124));
  NAND2 NAND2_1757(.VSS(VSS),.VDD(VDD),.Y(g27626),.A(g26989),.B(g3306));
  NAND2 NAND2_1758(.VSS(VSS),.VDD(VDD),.Y(g27627),.A(g27012),.B(g3462));
  NAND2 NAND2_1759(.VSS(VSS),.VDD(VDD),.Y(g27628),.A(g27038),.B(g3618));
  NAND2 NAND2_1760(.VSS(VSS),.VDD(VDD),.Y(g27630),.A(g27066),.B(g3774));
  NAND2 NAND2_1761(.VSS(VSS),.VDD(VDD),.Y(g27738),.A(g25367),.B(g27415));
  NAND2 NAND2_1762(.VSS(VSS),.VDD(VDD),.Y(g27743),.A(g25384),.B(g27436));
  NAND2 NAND2_1763(.VSS(VSS),.VDD(VDD),.Y(g27751),.A(g25400),.B(g27455));
  NAND2 NAND2_1764(.VSS(VSS),.VDD(VDD),.Y(g27756),.A(g25410),.B(g27471));
  NAND2 NAND2_1765(.VSS(VSS),.VDD(VDD),.Y(I36256),.A(g27527),.B(g15859));
  NAND2 NAND2_1766(.VSS(VSS),.VDD(VDD),.Y(I36257),.A(g27527),.B(I36256));
  NAND2 NAND2_1767(.VSS(VSS),.VDD(VDD),.Y(I36258),.A(g15859),.B(I36256));
  NAND2 NAND2_1768(.VSS(VSS),.VDD(VDD),.Y(g27801),.A(I36257),.B(I36258));
  NAND2 NAND2_1769(.VSS(VSS),.VDD(VDD),.Y(I36270),.A(g27549),.B(g15890));
  NAND2 NAND2_1770(.VSS(VSS),.VDD(VDD),.Y(I36271),.A(g27549),.B(I36270));
  NAND2 NAND2_1771(.VSS(VSS),.VDD(VDD),.Y(I36272),.A(g15890),.B(I36270));
  NAND2 NAND2_1772(.VSS(VSS),.VDD(VDD),.Y(g27809),.A(I36271),.B(I36272));
  NAND2 NAND2_1773(.VSS(VSS),.VDD(VDD),.Y(I36289),.A(g27565),.B(g15923));
  NAND2 NAND2_1774(.VSS(VSS),.VDD(VDD),.Y(I36290),.A(g27565),.B(I36289));
  NAND2 NAND2_1775(.VSS(VSS),.VDD(VDD),.Y(I36291),.A(g15923),.B(I36289));
  NAND2 NAND2_1776(.VSS(VSS),.VDD(VDD),.Y(g27830),.A(I36290),.B(I36291));
  NAND2 NAND2_1777(.VSS(VSS),.VDD(VDD),.Y(I36300),.A(g27382),.B(g27379));
  NAND2 NAND2_1778(.VSS(VSS),.VDD(VDD),.Y(I36301),.A(g27382),.B(I36300));
  NAND2 NAND2_1779(.VSS(VSS),.VDD(VDD),.Y(I36302),.A(g27379),.B(I36300));
  NAND2 NAND2_1780(.VSS(VSS),.VDD(VDD),.Y(g27838),.A(I36301),.B(I36302));
  NAND2 NAND2_1781(.VSS(VSS),.VDD(VDD),.Y(I36314),.A(g27575),.B(g15952));
  NAND2 NAND2_1782(.VSS(VSS),.VDD(VDD),.Y(I36315),.A(g27575),.B(I36314));
  NAND2 NAND2_1783(.VSS(VSS),.VDD(VDD),.Y(I36316),.A(g15952),.B(I36314));
  NAND2 NAND2_1784(.VSS(VSS),.VDD(VDD),.Y(g27846),.A(I36315),.B(I36316));
  NAND2 NAND2_1785(.VSS(VSS),.VDD(VDD),.Y(I36591),.A(g27529),.B(g14885));
  NAND2 NAND2_1786(.VSS(VSS),.VDD(VDD),.Y(I36592),.A(g27529),.B(I36591));
  NAND2 NAND2_1787(.VSS(VSS),.VDD(VDD),.Y(I36593),.A(g14885),.B(I36591));
  NAND2 NAND2_1788(.VSS(VSS),.VDD(VDD),.Y(g28046),.A(I36592),.B(I36593));
  NAND2 NAND2_1789(.VSS(VSS),.VDD(VDD),.Y(I36666),.A(g27551),.B(g14966));
  NAND2 NAND2_1790(.VSS(VSS),.VDD(VDD),.Y(I36667),.A(g27551),.B(I36666));
  NAND2 NAND2_1791(.VSS(VSS),.VDD(VDD),.Y(I36668),.A(g14966),.B(I36666));
  NAND2 NAND2_1792(.VSS(VSS),.VDD(VDD),.Y(g28075),.A(I36667),.B(I36668));
  NAND2 NAND2_1793(.VSS(VSS),.VDD(VDD),.Y(I36731),.A(g27567),.B(g15055));
  NAND2 NAND2_1794(.VSS(VSS),.VDD(VDD),.Y(I36732),.A(g27567),.B(I36731));
  NAND2 NAND2_1795(.VSS(VSS),.VDD(VDD),.Y(I36733),.A(g15055),.B(I36731));
  NAND2 NAND2_1796(.VSS(VSS),.VDD(VDD),.Y(g28100),.A(I36732),.B(I36733));
  NAND2 NAND2_1797(.VSS(VSS),.VDD(VDD),.Y(I36779),.A(g27577),.B(g15151));
  NAND2 NAND2_1798(.VSS(VSS),.VDD(VDD),.Y(I36780),.A(g27577),.B(I36779));
  NAND2 NAND2_1799(.VSS(VSS),.VDD(VDD),.Y(I36781),.A(g15151),.B(I36779));
  NAND2 NAND2_1800(.VSS(VSS),.VDD(VDD),.Y(g28118),.A(I36780),.B(I36781));
  NAND2 NAND2_1801(.VSS(VSS),.VDD(VDD),.Y(I37295),.A(g27827),.B(g27814));
  NAND2 NAND2_1802(.VSS(VSS),.VDD(VDD),.Y(I37296),.A(g27827),.B(I37295));
  NAND2 NAND2_1803(.VSS(VSS),.VDD(VDD),.Y(I37297),.A(g27814),.B(I37295));
  NAND2 NAND2_1804(.VSS(VSS),.VDD(VDD),.Y(g28384),.A(I37296),.B(I37297));
  NAND2 NAND2_1805(.VSS(VSS),.VDD(VDD),.Y(I37303),.A(g27802),.B(g27900));
  NAND2 NAND2_1806(.VSS(VSS),.VDD(VDD),.Y(I37304),.A(g27802),.B(I37303));
  NAND2 NAND2_1807(.VSS(VSS),.VDD(VDD),.Y(I37305),.A(g27900),.B(I37303));
  NAND2 NAND2_1808(.VSS(VSS),.VDD(VDD),.Y(g28386),.A(I37304),.B(I37305));
  NAND2 NAND2_1809(.VSS(VSS),.VDD(VDD),.Y(I37311),.A(g27897),.B(g27883));
  NAND2 NAND2_1810(.VSS(VSS),.VDD(VDD),.Y(I37312),.A(g27897),.B(I37311));
  NAND2 NAND2_1811(.VSS(VSS),.VDD(VDD),.Y(I37313),.A(g27883),.B(I37311));
  NAND2 NAND2_1812(.VSS(VSS),.VDD(VDD),.Y(g28388),.A(I37312),.B(I37313));
  NAND2 NAND2_1813(.VSS(VSS),.VDD(VDD),.Y(I37322),.A(g27865),.B(g27855));
  NAND2 NAND2_1814(.VSS(VSS),.VDD(VDD),.Y(I37323),.A(g27865),.B(I37322));
  NAND2 NAND2_1815(.VSS(VSS),.VDD(VDD),.Y(I37324),.A(g27855),.B(I37322));
  NAND2 NAND2_1816(.VSS(VSS),.VDD(VDD),.Y(g28391),.A(I37323),.B(I37324));
  NAND2 NAND2_1817(.VSS(VSS),.VDD(VDD),.Y(I37356),.A(g27824),.B(g27811));
  NAND2 NAND2_1818(.VSS(VSS),.VDD(VDD),.Y(I37357),.A(g27824),.B(I37356));
  NAND2 NAND2_1819(.VSS(VSS),.VDD(VDD),.Y(I37358),.A(g27811),.B(I37356));
  NAND2 NAND2_1820(.VSS(VSS),.VDD(VDD),.Y(g28415),.A(I37357),.B(I37358));
  NAND2 NAND2_1821(.VSS(VSS),.VDD(VDD),.Y(I37813),.A(g28388),.B(g28391));
  NAND2 NAND2_1822(.VSS(VSS),.VDD(VDD),.Y(I37814),.A(g28388),.B(I37813));
  NAND2 NAND2_1823(.VSS(VSS),.VDD(VDD),.Y(I37815),.A(g28391),.B(I37813));
  NAND2 NAND2_1824(.VSS(VSS),.VDD(VDD),.Y(g28842),.A(I37814),.B(I37815));
  NAND2 NAND2_1825(.VSS(VSS),.VDD(VDD),.Y(I37822),.A(g28384),.B(g28386));
  NAND2 NAND2_1826(.VSS(VSS),.VDD(VDD),.Y(I37823),.A(g28384),.B(I37822));
  NAND2 NAND2_1827(.VSS(VSS),.VDD(VDD),.Y(I37824),.A(g28386),.B(I37822));
  NAND2 NAND2_1828(.VSS(VSS),.VDD(VDD),.Y(g28845),.A(I37823),.B(I37824));
  NAND2 NAND2_1829(.VSS(VSS),.VDD(VDD),.Y(g28978),.A(g9150),.B(g28512));
  NAND2 NAND2_1830(.VSS(VSS),.VDD(VDD),.Y(g29001),.A(g9161),.B(g28512));
  NAND2 NAND2_1831(.VSS(VSS),.VDD(VDD),.Y(g29008),.A(g9174),.B(g28540));
  NAND2 NAND2_1832(.VSS(VSS),.VDD(VDD),.Y(g29026),.A(g9187),.B(g28512));
  NAND2 NAND2_1833(.VSS(VSS),.VDD(VDD),.Y(g29030),.A(g9203),.B(g28540));
  NAND2 NAND2_1834(.VSS(VSS),.VDD(VDD),.Y(g29038),.A(g9216),.B(g28567));
  NAND2 NAND2_1835(.VSS(VSS),.VDD(VDD),.Y(g29045),.A(g9232),.B(g28512));
  NAND2 NAND2_1836(.VSS(VSS),.VDD(VDD),.Y(g29049),.A(g9248),.B(g28540));
  NAND2 NAND2_1837(.VSS(VSS),.VDD(VDD),.Y(g29053),.A(g9264),.B(g28567));
  NAND2 NAND2_1838(.VSS(VSS),.VDD(VDD),.Y(g29060),.A(g9277),.B(g28595));
  NAND2 NAND2_1839(.VSS(VSS),.VDD(VDD),.Y(g29062),.A(g9310),.B(g28540));
  NAND2 NAND2_1840(.VSS(VSS),.VDD(VDD),.Y(g29068),.A(g9326),.B(g28567));
  NAND2 NAND2_1841(.VSS(VSS),.VDD(VDD),.Y(g29072),.A(g9342),.B(g28595));
  NAND2 NAND2_1842(.VSS(VSS),.VDD(VDD),.Y(g29076),.A(g9391),.B(g28567));
  NAND2 NAND2_1843(.VSS(VSS),.VDD(VDD),.Y(g29080),.A(g9407),.B(g28595));
  NAND2 NAND2_1844(.VSS(VSS),.VDD(VDD),.Y(g29087),.A(g9488),.B(g28595));
  NAND2 NAND2_1845(.VSS(VSS),.VDD(VDD),.Y(g29088),.A(g9507),.B(g28512));
  NAND2 NAND2_1846(.VSS(VSS),.VDD(VDD),.Y(g29096),.A(g9649),.B(g28540));
  NAND2 NAND2_1847(.VSS(VSS),.VDD(VDD),.Y(g29103),.A(g9795),.B(g28567));
  NAND2 NAND2_1848(.VSS(VSS),.VDD(VDD),.Y(g29107),.A(g9941),.B(g28595));
  NAND2 NAND2_1849(.VSS(VSS),.VDD(VDD),.Y(I38378),.A(g28845),.B(g28842));
  NAND2 NAND2_1850(.VSS(VSS),.VDD(VDD),.Y(I38379),.A(g28845),.B(I38378));
  NAND2 NAND2_1851(.VSS(VSS),.VDD(VDD),.Y(I38380),.A(g28842),.B(I38378));
  NAND2 NAND2_1852(.VSS(VSS),.VDD(VDD),.Y(g29265),.A(I38379),.B(I38380));
  NAND2 NAND2_1853(.VSS(VSS),.VDD(VDD),.Y(I38810),.A(g29303),.B(g15904));
  NAND2 NAND2_1854(.VSS(VSS),.VDD(VDD),.Y(I38811),.A(g29303),.B(I38810));
  NAND2 NAND2_1855(.VSS(VSS),.VDD(VDD),.Y(I38812),.A(g15904),.B(I38810));
  NAND2 NAND2_1856(.VSS(VSS),.VDD(VDD),.Y(g29498),.A(I38811),.B(I38812));
  NAND2 NAND2_1857(.VSS(VSS),.VDD(VDD),.Y(I38820),.A(g29313),.B(g15933));
  NAND2 NAND2_1858(.VSS(VSS),.VDD(VDD),.Y(I38821),.A(g29313),.B(I38820));
  NAND2 NAND2_1859(.VSS(VSS),.VDD(VDD),.Y(I38822),.A(g15933),.B(I38820));
  NAND2 NAND2_1860(.VSS(VSS),.VDD(VDD),.Y(g29500),.A(I38821),.B(I38822));
  NAND2 NAND2_1861(.VSS(VSS),.VDD(VDD),.Y(I38831),.A(g29324),.B(g15962));
  NAND2 NAND2_1862(.VSS(VSS),.VDD(VDD),.Y(I38832),.A(g29324),.B(I38831));
  NAND2 NAND2_1863(.VSS(VSS),.VDD(VDD),.Y(I38833),.A(g15962),.B(I38831));
  NAND2 NAND2_1864(.VSS(VSS),.VDD(VDD),.Y(g29503),.A(I38832),.B(I38833));
  NAND2 NAND2_1865(.VSS(VSS),.VDD(VDD),.Y(I38841),.A(g29333),.B(g15981));
  NAND2 NAND2_1866(.VSS(VSS),.VDD(VDD),.Y(I38842),.A(g29333),.B(I38841));
  NAND2 NAND2_1867(.VSS(VSS),.VDD(VDD),.Y(I38843),.A(g15981),.B(I38841));
  NAND2 NAND2_1868(.VSS(VSS),.VDD(VDD),.Y(g29505),.A(I38842),.B(I38843));
  NAND2 NAND2_1869(.VSS(VSS),.VDD(VDD),.Y(I39323),.A(g29721),.B(g29713));
  NAND2 NAND2_1870(.VSS(VSS),.VDD(VDD),.Y(I39324),.A(g29721),.B(I39323));
  NAND2 NAND2_1871(.VSS(VSS),.VDD(VDD),.Y(I39325),.A(g29713),.B(I39323));
  NAND2 NAND2_1872(.VSS(VSS),.VDD(VDD),.Y(g29911),.A(I39324),.B(I39325));
  NAND2 NAND2_1873(.VSS(VSS),.VDD(VDD),.Y(I39331),.A(g29705),.B(g29751));
  NAND2 NAND2_1874(.VSS(VSS),.VDD(VDD),.Y(I39332),.A(g29705),.B(I39331));
  NAND2 NAND2_1875(.VSS(VSS),.VDD(VDD),.Y(I39333),.A(g29751),.B(I39331));
  NAND2 NAND2_1876(.VSS(VSS),.VDD(VDD),.Y(g29913),.A(I39332),.B(I39333));
  NAND2 NAND2_1877(.VSS(VSS),.VDD(VDD),.Y(I39339),.A(g29748),.B(g29741));
  NAND2 NAND2_1878(.VSS(VSS),.VDD(VDD),.Y(I39340),.A(g29748),.B(I39339));
  NAND2 NAND2_1879(.VSS(VSS),.VDD(VDD),.Y(I39341),.A(g29741),.B(I39339));
  NAND2 NAND2_1880(.VSS(VSS),.VDD(VDD),.Y(g29915),.A(I39340),.B(I39341));
  NAND2 NAND2_1881(.VSS(VSS),.VDD(VDD),.Y(I39347),.A(g29732),.B(g29728));
  NAND2 NAND2_1882(.VSS(VSS),.VDD(VDD),.Y(I39348),.A(g29732),.B(I39347));
  NAND2 NAND2_1883(.VSS(VSS),.VDD(VDD),.Y(I39349),.A(g29728),.B(I39347));
  NAND2 NAND2_1884(.VSS(VSS),.VDD(VDD),.Y(g29917),.A(I39348),.B(I39349));
  NAND2 NAND2_1885(.VSS(VSS),.VDD(VDD),.Y(I39359),.A(g29766),.B(g15880));
  NAND2 NAND2_1886(.VSS(VSS),.VDD(VDD),.Y(I39360),.A(g29766),.B(I39359));
  NAND2 NAND2_1887(.VSS(VSS),.VDD(VDD),.Y(I39361),.A(g15880),.B(I39359));
  NAND2 NAND2_1888(.VSS(VSS),.VDD(VDD),.Y(g29923),.A(I39360),.B(I39361));
  NAND2 NAND2_1889(.VSS(VSS),.VDD(VDD),.Y(I39367),.A(g29767),.B(g15913));
  NAND2 NAND2_1890(.VSS(VSS),.VDD(VDD),.Y(I39368),.A(g29767),.B(I39367));
  NAND2 NAND2_1891(.VSS(VSS),.VDD(VDD),.Y(I39369),.A(g15913),.B(I39367));
  NAND2 NAND2_1892(.VSS(VSS),.VDD(VDD),.Y(g29925),.A(I39368),.B(I39369));
  NAND2 NAND2_1893(.VSS(VSS),.VDD(VDD),.Y(I39375),.A(g29768),.B(g15942));
  NAND2 NAND2_1894(.VSS(VSS),.VDD(VDD),.Y(I39376),.A(g29768),.B(I39375));
  NAND2 NAND2_1895(.VSS(VSS),.VDD(VDD),.Y(I39377),.A(g15942),.B(I39375));
  NAND2 NAND2_1896(.VSS(VSS),.VDD(VDD),.Y(g29927),.A(I39376),.B(I39377));
  NAND2 NAND2_1897(.VSS(VSS),.VDD(VDD),.Y(I39384),.A(g29718),.B(g29710));
  NAND2 NAND2_1898(.VSS(VSS),.VDD(VDD),.Y(I39385),.A(g29718),.B(I39384));
  NAND2 NAND2_1899(.VSS(VSS),.VDD(VDD),.Y(I39386),.A(g29710),.B(I39384));
  NAND2 NAND2_1900(.VSS(VSS),.VDD(VDD),.Y(g29930),.A(I39385),.B(I39386));
  NAND2 NAND2_1901(.VSS(VSS),.VDD(VDD),.Y(I39391),.A(g29769),.B(g15971));
  NAND2 NAND2_1902(.VSS(VSS),.VDD(VDD),.Y(I39392),.A(g29769),.B(I39391));
  NAND2 NAND2_1903(.VSS(VSS),.VDD(VDD),.Y(I39393),.A(g15971),.B(I39391));
  NAND2 NAND2_1904(.VSS(VSS),.VDD(VDD),.Y(g29931),.A(I39392),.B(I39393));
  NAND2 NAND2_1905(.VSS(VSS),.VDD(VDD),.Y(I39532),.A(g29915),.B(g29917));
  NAND2 NAND2_1906(.VSS(VSS),.VDD(VDD),.Y(I39533),.A(g29915),.B(I39532));
  NAND2 NAND2_1907(.VSS(VSS),.VDD(VDD),.Y(I39534),.A(g29917),.B(I39532));
  NAND2 NAND2_1908(.VSS(VSS),.VDD(VDD),.Y(g30034),.A(I39533),.B(I39534));
  NAND2 NAND2_1909(.VSS(VSS),.VDD(VDD),.Y(I39539),.A(g29911),.B(g29913));
  NAND2 NAND2_1910(.VSS(VSS),.VDD(VDD),.Y(I39540),.A(g29911),.B(I39539));
  NAND2 NAND2_1911(.VSS(VSS),.VDD(VDD),.Y(I39541),.A(g29913),.B(I39539));
  NAND2 NAND2_1912(.VSS(VSS),.VDD(VDD),.Y(g30035),.A(I39540),.B(I39541));
  NAND2 NAND2_1913(.VSS(VSS),.VDD(VDD),.Y(I39689),.A(g30035),.B(g30034));
  NAND2 NAND2_1914(.VSS(VSS),.VDD(VDD),.Y(I39690),.A(g30035),.B(I39689));
  NAND2 NAND2_1915(.VSS(VSS),.VDD(VDD),.Y(I39691),.A(g30034),.B(I39689));
  NAND2 NAND2_1916(.VSS(VSS),.VDD(VDD),.Y(g30228),.A(I39690),.B(I39691));
  NAND2 NAND2_1917(.VSS(VSS),.VDD(VDD),.Y(I40558),.A(g30605),.B(g30597));
  NAND2 NAND2_1918(.VSS(VSS),.VDD(VDD),.Y(I40559),.A(g30605),.B(I40558));
  NAND2 NAND2_1919(.VSS(VSS),.VDD(VDD),.Y(I40560),.A(g30597),.B(I40558));
  NAND2 NAND2_1920(.VSS(VSS),.VDD(VDD),.Y(g30768),.A(I40559),.B(I40560));
  NAND2 NAND2_1921(.VSS(VSS),.VDD(VDD),.Y(I40571),.A(g30588),.B(g30632));
  NAND2 NAND2_1922(.VSS(VSS),.VDD(VDD),.Y(I40572),.A(g30588),.B(I40571));
  NAND2 NAND2_1923(.VSS(VSS),.VDD(VDD),.Y(I40573),.A(g30632),.B(I40571));
  NAND2 NAND2_1924(.VSS(VSS),.VDD(VDD),.Y(g30771),.A(I40572),.B(I40573));
  NAND2 NAND2_1925(.VSS(VSS),.VDD(VDD),.Y(I40587),.A(g30629),.B(g30622));
  NAND2 NAND2_1926(.VSS(VSS),.VDD(VDD),.Y(I40588),.A(g30629),.B(I40587));
  NAND2 NAND2_1927(.VSS(VSS),.VDD(VDD),.Y(I40589),.A(g30622),.B(I40587));
  NAND2 NAND2_1928(.VSS(VSS),.VDD(VDD),.Y(g30775),.A(I40588),.B(I40589));
  NAND2 NAND2_1929(.VSS(VSS),.VDD(VDD),.Y(I40603),.A(g30614),.B(g30610));
  NAND2 NAND2_1930(.VSS(VSS),.VDD(VDD),.Y(I40604),.A(g30614),.B(I40603));
  NAND2 NAND2_1931(.VSS(VSS),.VDD(VDD),.Y(I40605),.A(g30610),.B(I40603));
  NAND2 NAND2_1932(.VSS(VSS),.VDD(VDD),.Y(g30779),.A(I40604),.B(I40605));
  NAND2 NAND2_1933(.VSS(VSS),.VDD(VDD),.Y(I40627),.A(g30602),.B(g30594));
  NAND2 NAND2_1934(.VSS(VSS),.VDD(VDD),.Y(I40628),.A(g30602),.B(I40627));
  NAND2 NAND2_1935(.VSS(VSS),.VDD(VDD),.Y(I40629),.A(g30594),.B(I40627));
  NAND2 NAND2_1936(.VSS(VSS),.VDD(VDD),.Y(g30791),.A(I40628),.B(I40629));
  NAND2 NAND2_1937(.VSS(VSS),.VDD(VDD),.Y(I41010),.A(g30775),.B(g30779));
  NAND2 NAND2_1938(.VSS(VSS),.VDD(VDD),.Y(I41011),.A(g30775),.B(I41010));
  NAND2 NAND2_1939(.VSS(VSS),.VDD(VDD),.Y(I41012),.A(g30779),.B(I41010));
  NAND2 NAND2_1940(.VSS(VSS),.VDD(VDD),.Y(g30926),.A(I41011),.B(I41012));
  NAND2 NAND2_1941(.VSS(VSS),.VDD(VDD),.Y(I41017),.A(g30768),.B(g30771));
  NAND2 NAND2_1942(.VSS(VSS),.VDD(VDD),.Y(I41018),.A(g30768),.B(I41017));
  NAND2 NAND2_1943(.VSS(VSS),.VDD(VDD),.Y(I41019),.A(g30771),.B(I41017));
  NAND2 NAND2_1944(.VSS(VSS),.VDD(VDD),.Y(g30927),.A(I41018),.B(I41019));
  NAND2 NAND2_1945(.VSS(VSS),.VDD(VDD),.Y(I41064),.A(g30927),.B(g30926));
  NAND2 NAND2_1946(.VSS(VSS),.VDD(VDD),.Y(I41065),.A(g30927),.B(I41064));
  NAND2 NAND2_1947(.VSS(VSS),.VDD(VDD),.Y(I41066),.A(g30926),.B(I41064));
  NAND2 NAND2_1948(.VSS(VSS),.VDD(VDD),.Y(g30952),.A(I41065),.B(I41066));
//
  NOR3 NOR3_0(.VSS(VSS),.VDD(VDD),.Y(g7528),.A(g3151),.B(g3142),.C(g3147));
  NOR2 NOR2_0(.VSS(VSS),.VDD(VDD),.Y(g7575),.A(g2984),.B(g2985));
  NOR2 NOR2_1(.VSS(VSS),.VDD(VDD),.Y(g7795),.A(g2992),.B(g2991));
  NOR4 NOR4_0(.VSS(VSS),.VDD(VDD),.Y(g8430),.A(g3198),.B(g8120),.C(g3194),.D(g3191));
  NOR3 NOR3_1(.VSS(VSS),.VDD(VDD),.Y(g10784),.A(g5630),.B(g5649),.C(g5676));
  NOR3 NOR3_2(.VSS(VSS),.VDD(VDD),.Y(g10789),.A(g5650),.B(g5677),.C(g5709));
  NOR3 NOR3_3(.VSS(VSS),.VDD(VDD),.Y(g10793),.A(g5658),.B(g5687),.C(g5728));
  NOR3 NOR3_4(.VSS(VSS),.VDD(VDD),.Y(g10797),.A(g5678),.B(g5710),.C(g5757));
  NOR3 NOR3_5(.VSS(VSS),.VDD(VDD),.Y(g10801),.A(g5688),.B(g5729),.C(g5767));
  NOR3 NOR3_6(.VSS(VSS),.VDD(VDD),.Y(g10805),.A(g5696),.B(g5739),.C(g5786));
  NOR3 NOR3_7(.VSS(VSS),.VDD(VDD),.Y(g10810),.A(g5711),.B(g5758),.C(g5807));
  NOR3 NOR3_8(.VSS(VSS),.VDD(VDD),.Y(g10814),.A(g5730),.B(g5768),.C(g5816));
  NOR3 NOR3_9(.VSS(VSS),.VDD(VDD),.Y(g10818),.A(g5740),.B(g5787),.C(g5826));
  NOR3 NOR3_10(.VSS(VSS),.VDD(VDD),.Y(g10822),.A(g5748),.B(g5797),.C(g5845));
  NOR3 NOR3_11(.VSS(VSS),.VDD(VDD),.Y(g10831),.A(g5769),.B(g5817),.C(g5863));
  NOR3 NOR3_12(.VSS(VSS),.VDD(VDD),.Y(g10835),.A(g5788),.B(g5827),.C(g5872));
  NOR3 NOR3_13(.VSS(VSS),.VDD(VDD),.Y(g10839),.A(g5798),.B(g5846),.C(g5882));
  NOR3 NOR3_14(.VSS(VSS),.VDD(VDD),.Y(g10851),.A(g5828),.B(g5873),.C(g5910));
  NOR3 NOR3_15(.VSS(VSS),.VDD(VDD),.Y(g10855),.A(g5847),.B(g5883),.C(g5919));
  NOR3 NOR3_16(.VSS(VSS),.VDD(VDD),.Y(g10872),.A(g5884),.B(g5920),.C(g5949));
  NOR3 NOR3_17(.VSS(VSS),.VDD(VDD),.Y(g11600),.A(g9049),.B(g9064),.C(g9078));
  NOR4 NOR4_1(.VSS(VSS),.VDD(VDD),.Y(g11622),.A(g8183),.B(g11332),.C(g7928),.D(g11069));
  NOR3 NOR3_18(.VSS(VSS),.VDD(VDD),.Y(g11624),.A(g9062),.B(g9075),.C(g9091));
  NOR3 NOR3_19(.VSS(VSS),.VDD(VDD),.Y(g11627),.A(g9063),.B(g9077),.C(g9093));
  NOR3 NOR3_20(.VSS(VSS),.VDD(VDD),.Y(g11630),.A(g9066),.B(g9081),.C(g9097));
  NOR4 NOR4_2(.VSS(VSS),.VDD(VDD),.Y(g11643),.A(g11481),.B(g8045),.C(g7928),.D(g11069));
  NOR3 NOR3_21(.VSS(VSS),.VDD(VDD),.Y(g11644),.A(g9076),.B(g9092),.C(g9102));
  NOR3 NOR3_22(.VSS(VSS),.VDD(VDD),.Y(g11647),.A(g9079),.B(g9094),.C(g9103));
  NOR3 NOR3_23(.VSS(VSS),.VDD(VDD),.Y(g11650),.A(g9080),.B(g9096),.C(g9105));
  NOR3 NOR3_24(.VSS(VSS),.VDD(VDD),.Y(g11653),.A(g9083),.B(g9100),.C(g9109));
  NOR4 NOR4_3(.VSS(VSS),.VDD(VDD),.Y(g11660),.A(g8183),.B(g8045),.C(g7928),.D(g11069));
  NOR3 NOR3_25(.VSS(VSS),.VDD(VDD),.Y(g11663),.A(g9095),.B(g9104),.C(g9112));
  NOR3 NOR3_26(.VSS(VSS),.VDD(VDD),.Y(g11666),.A(g9098),.B(g9106),.C(g9113));
  NOR3 NOR3_27(.VSS(VSS),.VDD(VDD),.Y(g11669),.A(g9099),.B(g9108),.C(g9115));
  NOR3 NOR3_28(.VSS(VSS),.VDD(VDD),.Y(g11675),.A(g9107),.B(g9114),.C(g9120));
  NOR3 NOR3_29(.VSS(VSS),.VDD(VDD),.Y(g11678),.A(g9110),.B(g9116),.C(g9121));
  NOR3 NOR3_30(.VSS(VSS),.VDD(VDD),.Y(g11681),.A(g9111),.B(g9118),.C(g9123));
  NOR3 NOR3_31(.VSS(VSS),.VDD(VDD),.Y(g11687),.A(g9117),.B(g9122),.C(g9126));
  NOR3 NOR3_32(.VSS(VSS),.VDD(VDD),.Y(g11690),.A(g9119),.B(g9124),.C(g9127));
  NOR3 NOR3_33(.VSS(VSS),.VDD(VDD),.Y(g11697),.A(g9125),.B(g9131),.C(g9133));
  NOR3 NOR3_34(.VSS(VSS),.VDD(VDD),.Y(g11703),.A(g9132),.B(g9137),.C(g9139));
  NOR3 NOR3_35(.VSS(VSS),.VDD(VDD),.Y(g11711),.A(g9138),.B(g9143),.C(g9145));
  NOR3 NOR3_36(.VSS(VSS),.VDD(VDD),.Y(g11744),.A(g9241),.B(g9301),.C(g9364));
  NOR3 NOR3_37(.VSS(VSS),.VDD(VDD),.Y(g11759),.A(g9302),.B(g9365),.C(g9438));
  NOR3 NOR3_38(.VSS(VSS),.VDD(VDD),.Y(g11760),.A(g9319),.B(g9382),.C(g9461));
  NOR3 NOR3_39(.VSS(VSS),.VDD(VDD),.Y(g11767),.A(g9366),.B(g9439),.C(g9518));
  NOR3 NOR3_40(.VSS(VSS),.VDD(VDD),.Y(g11768),.A(g9367),.B(g9441),.C(g9521));
  NOR3 NOR3_41(.VSS(VSS),.VDD(VDD),.Y(g11772),.A(g9383),.B(g9462),.C(g9580));
  NOR3 NOR3_42(.VSS(VSS),.VDD(VDD),.Y(g11773),.A(g9400),.B(g9479),.C(g9603));
  NOR3 NOR3_43(.VSS(VSS),.VDD(VDD),.Y(g11780),.A(g9440),.B(g9519),.C(g9630));
  NOR3 NOR3_44(.VSS(VSS),.VDD(VDD),.Y(g11781),.A(g9442),.B(g9522),.C(g9633));
  NOR3 NOR3_45(.VSS(VSS),.VDD(VDD),.Y(g11784),.A(g9463),.B(g9581),.C(g9660));
  NOR3 NOR3_46(.VSS(VSS),.VDD(VDD),.Y(g11785),.A(g9464),.B(g9583),.C(g9663));
  NOR3 NOR3_47(.VSS(VSS),.VDD(VDD),.Y(g11789),.A(g9480),.B(g9604),.C(g9722));
  NOR3 NOR3_48(.VSS(VSS),.VDD(VDD),.Y(g11790),.A(g9497),.B(g9621),.C(g9745));
  NOR3 NOR3_49(.VSS(VSS),.VDD(VDD),.Y(g11799),.A(g9520),.B(g9631),.C(g9759));
  NOR3 NOR3_50(.VSS(VSS),.VDD(VDD),.Y(g11800),.A(g9523),.B(g9634),.C(g9762));
  NOR3 NOR3_51(.VSS(VSS),.VDD(VDD),.Y(g11806),.A(g9582),.B(g9661),.C(g9776));
  NOR3 NOR3_52(.VSS(VSS),.VDD(VDD),.Y(g11807),.A(g9584),.B(g9664),.C(g9779));
  NOR3 NOR3_53(.VSS(VSS),.VDD(VDD),.Y(g11810),.A(g9605),.B(g9723),.C(g9806));
  NOR3 NOR3_54(.VSS(VSS),.VDD(VDD),.Y(g11811),.A(g9606),.B(g9725),.C(g9809));
  NOR3 NOR3_55(.VSS(VSS),.VDD(VDD),.Y(g11815),.A(g9622),.B(g9746),.C(g9868));
  NOR3 NOR3_56(.VSS(VSS),.VDD(VDD),.Y(g11822),.A(g9632),.B(g9760),.C(g9888));
  NOR3 NOR3_57(.VSS(VSS),.VDD(VDD),.Y(g11823),.A(g9635),.B(g9763),.C(g9891));
  NOR3 NOR3_58(.VSS(VSS),.VDD(VDD),.Y(g11828),.A(g9639),.B(g9764),.C(g9892));
  NOR3 NOR3_59(.VSS(VSS),.VDD(VDD),.Y(g11830),.A(g9647),.B(g9773),.C(g9901));
  NOR3 NOR3_60(.VSS(VSS),.VDD(VDD),.Y(g11831),.A(g9648),.B(g9775),.C(g9904));
  NOR3 NOR3_61(.VSS(VSS),.VDD(VDD),.Y(g11832),.A(g9662),.B(g9777),.C(g9905));
  NOR3 NOR3_62(.VSS(VSS),.VDD(VDD),.Y(g11833),.A(g9665),.B(g9780),.C(g9908));
  NOR3 NOR3_63(.VSS(VSS),.VDD(VDD),.Y(g11839),.A(g9724),.B(g9807),.C(g9922));
  NOR3 NOR3_64(.VSS(VSS),.VDD(VDD),.Y(g11840),.A(g9726),.B(g9810),.C(g9925));
  NOR3 NOR3_65(.VSS(VSS),.VDD(VDD),.Y(g11843),.A(g9747),.B(g9869),.C(g9952));
  NOR3 NOR3_66(.VSS(VSS),.VDD(VDD),.Y(g11844),.A(g9748),.B(g9871),.C(g9955));
  NOR3 NOR3_67(.VSS(VSS),.VDD(VDD),.Y(g11855),.A(g9761),.B(g9889),.C(g10009));
  NOR3 NOR3_68(.VSS(VSS),.VDD(VDD),.Y(g11860),.A(g9765),.B(g9893),.C(g10012));
  NOR3 NOR3_69(.VSS(VSS),.VDD(VDD),.Y(g11861),.A(g9766),.B(g9894),.C(g10013));
  NOR3 NOR3_70(.VSS(VSS),.VDD(VDD),.Y(g11863),.A(g9774),.B(g9902),.C(g10035));
  NOR3 NOR3_71(.VSS(VSS),.VDD(VDD),.Y(g11864),.A(g9778),.B(g9906),.C(g10042));
  NOR3 NOR3_72(.VSS(VSS),.VDD(VDD),.Y(g11865),.A(g9781),.B(g9909),.C(g10045));
  NOR3 NOR3_73(.VSS(VSS),.VDD(VDD),.Y(g11870),.A(g9785),.B(g9910),.C(g10046));
  NOR3 NOR3_74(.VSS(VSS),.VDD(VDD),.Y(g11872),.A(g9793),.B(g9919),.C(g10055));
  NOR3 NOR3_75(.VSS(VSS),.VDD(VDD),.Y(g11873),.A(g9794),.B(g9921),.C(g10058));
  NOR3 NOR3_76(.VSS(VSS),.VDD(VDD),.Y(g11874),.A(g9808),.B(g9923),.C(g10059));
  NOR3 NOR3_77(.VSS(VSS),.VDD(VDD),.Y(g11875),.A(g9811),.B(g9926),.C(g10062));
  NOR3 NOR3_78(.VSS(VSS),.VDD(VDD),.Y(g11881),.A(g9870),.B(g9953),.C(g10076));
  NOR3 NOR3_79(.VSS(VSS),.VDD(VDD),.Y(g11882),.A(g9872),.B(g9956),.C(g10079));
  NOR3 NOR3_80(.VSS(VSS),.VDD(VDD),.Y(g11889),.A(g9887),.B(g10007),.C(g10101));
  NOR3 NOR3_81(.VSS(VSS),.VDD(VDD),.Y(g11890),.A(g9890),.B(g10010),.C(g10103));
  NOR3 NOR3_82(.VSS(VSS),.VDD(VDD),.Y(g11896),.A(g9903),.B(g10036),.C(g10112));
  NOR3 NOR3_83(.VSS(VSS),.VDD(VDD),.Y(g11897),.A(g9907),.B(g10043),.C(g10118));
  NOR3 NOR3_84(.VSS(VSS),.VDD(VDD),.Y(g11902),.A(g9911),.B(g10047),.C(g10121));
  NOR3 NOR3_85(.VSS(VSS),.VDD(VDD),.Y(g11903),.A(g9912),.B(g10048),.C(g10122));
  NOR3 NOR3_86(.VSS(VSS),.VDD(VDD),.Y(g11905),.A(g9920),.B(g10056),.C(g10144));
  NOR3 NOR3_87(.VSS(VSS),.VDD(VDD),.Y(g11906),.A(g9924),.B(g10060),.C(g10151));
  NOR3 NOR3_88(.VSS(VSS),.VDD(VDD),.Y(g11907),.A(g9927),.B(g10063),.C(g10154));
  NOR3 NOR3_89(.VSS(VSS),.VDD(VDD),.Y(g11912),.A(g9931),.B(g10064),.C(g10155));
  NOR3 NOR3_90(.VSS(VSS),.VDD(VDD),.Y(g11914),.A(g9939),.B(g10073),.C(g10164));
  NOR3 NOR3_91(.VSS(VSS),.VDD(VDD),.Y(g11915),.A(g9940),.B(g10075),.C(g10167));
  NOR3 NOR3_92(.VSS(VSS),.VDD(VDD),.Y(g11916),.A(g9954),.B(g10077),.C(g10168));
  NOR3 NOR3_93(.VSS(VSS),.VDD(VDD),.Y(g11917),.A(g9957),.B(g10080),.C(g10171));
  NOR3 NOR3_94(.VSS(VSS),.VDD(VDD),.Y(g11928),.A(g10008),.B(g10102),.C(g10192));
  NOR3 NOR3_95(.VSS(VSS),.VDD(VDD),.Y(g11934),.A(g10011),.B(g10104),.C(g10193));
  NOR3 NOR3_96(.VSS(VSS),.VDD(VDD),.Y(g11935),.A(g10014),.B(g10106),.C(g10196));
  NOR3 NOR3_97(.VSS(VSS),.VDD(VDD),.Y(g11938),.A(g10037),.B(g10113),.C(g10201));
  NOR3 NOR3_98(.VSS(VSS),.VDD(VDD),.Y(g11939),.A(g10041),.B(g10116),.C(g10206));
  NOR3 NOR3_99(.VSS(VSS),.VDD(VDD),.Y(g11940),.A(g10044),.B(g10119),.C(g10208));
  NOR3 NOR3_100(.VSS(VSS),.VDD(VDD),.Y(g11946),.A(g10057),.B(g10145),.C(g10217));
  NOR3 NOR3_101(.VSS(VSS),.VDD(VDD),.Y(g11947),.A(g10061),.B(g10152),.C(g10223));
  NOR3 NOR3_102(.VSS(VSS),.VDD(VDD),.Y(g11952),.A(g10065),.B(g10156),.C(g10226));
  NOR3 NOR3_103(.VSS(VSS),.VDD(VDD),.Y(g11953),.A(g10066),.B(g10157),.C(g10227));
  NOR3 NOR3_104(.VSS(VSS),.VDD(VDD),.Y(g11955),.A(g10074),.B(g10165),.C(g10249));
  NOR3 NOR3_105(.VSS(VSS),.VDD(VDD),.Y(g11956),.A(g10078),.B(g10169),.C(g10256));
  NOR3 NOR3_106(.VSS(VSS),.VDD(VDD),.Y(g11957),.A(g10081),.B(g10172),.C(g10259));
  NOR3 NOR3_107(.VSS(VSS),.VDD(VDD),.Y(g11962),.A(g10085),.B(g10173),.C(g10260));
  NOR3 NOR3_108(.VSS(VSS),.VDD(VDD),.Y(g11964),.A(g10093),.B(g10182),.C(g10269));
  NOR3 NOR3_109(.VSS(VSS),.VDD(VDD),.Y(g11965),.A(g10094),.B(g10184),.C(g10272));
  NOR3 NOR3_110(.VSS(VSS),.VDD(VDD),.Y(g11974),.A(g10105),.B(g10194),.C(g10279));
  NOR3 NOR3_111(.VSS(VSS),.VDD(VDD),.Y(g11975),.A(g10107),.B(g10197),.C(g10282));
  NOR3 NOR3_112(.VSS(VSS),.VDD(VDD),.Y(g11979),.A(g10114),.B(g10202),.C(g10288));
  NOR3 NOR3_113(.VSS(VSS),.VDD(VDD),.Y(g11980),.A(g10115),.B(g10204),.C(g10291));
  NOR3 NOR3_114(.VSS(VSS),.VDD(VDD),.Y(g11981),.A(g10117),.B(g10207),.C(g10294));
  NOR3 NOR3_115(.VSS(VSS),.VDD(VDD),.Y(g11987),.A(g10120),.B(g10209),.C(g10295));
  NOR3 NOR3_116(.VSS(VSS),.VDD(VDD),.Y(g11988),.A(g10123),.B(g10211),.C(g10298));
  NOR3 NOR3_117(.VSS(VSS),.VDD(VDD),.Y(g11991),.A(g10146),.B(g10218),.C(g10303));
  NOR3 NOR3_118(.VSS(VSS),.VDD(VDD),.Y(g11992),.A(g10150),.B(g10221),.C(g10308));
  NOR3 NOR3_119(.VSS(VSS),.VDD(VDD),.Y(g11993),.A(g10153),.B(g10224),.C(g10310));
  NOR3 NOR3_120(.VSS(VSS),.VDD(VDD),.Y(g11999),.A(g10166),.B(g10250),.C(g10319));
  NOR3 NOR3_121(.VSS(VSS),.VDD(VDD),.Y(g12000),.A(g10170),.B(g10257),.C(g10325));
  NOR3 NOR3_122(.VSS(VSS),.VDD(VDD),.Y(g12005),.A(g10174),.B(g10261),.C(g10328));
  NOR3 NOR3_123(.VSS(VSS),.VDD(VDD),.Y(g12006),.A(g10175),.B(g10262),.C(g10329));
  NOR3 NOR3_124(.VSS(VSS),.VDD(VDD),.Y(g12008),.A(g10183),.B(g10270),.C(g10351));
  NOR3 NOR3_125(.VSS(VSS),.VDD(VDD),.Y(g12026),.A(g10195),.B(g10280),.C(g10360));
  NOR3 NOR3_126(.VSS(VSS),.VDD(VDD),.Y(g12033),.A(g10199),.B(g10284),.C(g10362));
  NOR3 NOR3_127(.VSS(VSS),.VDD(VDD),.Y(g12034),.A(g10200),.B(g10286),.C(g10365));
  NOR3 NOR3_128(.VSS(VSS),.VDD(VDD),.Y(g12035),.A(g10203),.B(g10289),.C(g10367));
  NOR3 NOR3_129(.VSS(VSS),.VDD(VDD),.Y(g12036),.A(g10205),.B(g10292),.C(g10370));
  NOR3 NOR3_130(.VSS(VSS),.VDD(VDD),.Y(g12043),.A(g10210),.B(g10296),.C(g10372));
  NOR3 NOR3_131(.VSS(VSS),.VDD(VDD),.Y(g12044),.A(g10212),.B(g10299),.C(g10375));
  NOR3 NOR3_132(.VSS(VSS),.VDD(VDD),.Y(g12048),.A(g10219),.B(g10304),.C(g10381));
  NOR3 NOR3_133(.VSS(VSS),.VDD(VDD),.Y(g12049),.A(g10220),.B(g10306),.C(g10384));
  NOR3 NOR3_134(.VSS(VSS),.VDD(VDD),.Y(g12050),.A(g10222),.B(g10309),.C(g10387));
  NOR3 NOR3_135(.VSS(VSS),.VDD(VDD),.Y(g12056),.A(g10225),.B(g10311),.C(g10388));
  NOR3 NOR3_136(.VSS(VSS),.VDD(VDD),.Y(g12057),.A(g10228),.B(g10313),.C(g10391));
  NOR3 NOR3_137(.VSS(VSS),.VDD(VDD),.Y(g12060),.A(g10251),.B(g10320),.C(g10396));
  NOR3 NOR3_138(.VSS(VSS),.VDD(VDD),.Y(g12061),.A(g10255),.B(g10323),.C(g10401));
  NOR3 NOR3_139(.VSS(VSS),.VDD(VDD),.Y(g12062),.A(g10258),.B(g10326),.C(g10403));
  NOR3 NOR3_140(.VSS(VSS),.VDD(VDD),.Y(g12068),.A(g10271),.B(g10352),.C(g10412));
  NOR3 NOR3_141(.VSS(VSS),.VDD(VDD),.Y(g12079),.A(g10281),.B(g10361),.C(g10422));
  NOR3 NOR3_142(.VSS(VSS),.VDD(VDD),.Y(g12080),.A(g10285),.B(g10363),.C(g10430));
  NOR3 NOR3_143(.VSS(VSS),.VDD(VDD),.Y(g12081),.A(g10287),.B(g10366),.C(g10433));
  NOR3 NOR3_144(.VSS(VSS),.VDD(VDD),.Y(g12082),.A(g10290),.B(g10368),.C(g10435));
  NOR3 NOR3_145(.VSS(VSS),.VDD(VDD),.Y(g12083),.A(g10293),.B(g10371),.C(g10438));
  NOR3 NOR3_146(.VSS(VSS),.VDD(VDD),.Y(g12090),.A(g10297),.B(g10373),.C(g10439));
  NOR3 NOR3_147(.VSS(VSS),.VDD(VDD),.Y(g12097),.A(g10301),.B(g10377),.C(g10441));
  NOR3 NOR3_148(.VSS(VSS),.VDD(VDD),.Y(g12098),.A(g10302),.B(g10379),.C(g10444));
  NOR3 NOR3_149(.VSS(VSS),.VDD(VDD),.Y(g12099),.A(g10305),.B(g10382),.C(g10446));
  NOR3 NOR3_150(.VSS(VSS),.VDD(VDD),.Y(g12100),.A(g10307),.B(g10385),.C(g10449));
  NOR3 NOR3_151(.VSS(VSS),.VDD(VDD),.Y(g12107),.A(g10312),.B(g10389),.C(g10451));
  NOR3 NOR3_152(.VSS(VSS),.VDD(VDD),.Y(g12108),.A(g10314),.B(g10392),.C(g10454));
  NOR3 NOR3_153(.VSS(VSS),.VDD(VDD),.Y(g12112),.A(g10321),.B(g10397),.C(g10460));
  NOR3 NOR3_154(.VSS(VSS),.VDD(VDD),.Y(g12113),.A(g10322),.B(g10399),.C(g10463));
  NOR3 NOR3_155(.VSS(VSS),.VDD(VDD),.Y(g12114),.A(g10324),.B(g10402),.C(g10466));
  NOR3 NOR3_156(.VSS(VSS),.VDD(VDD),.Y(g12120),.A(g10327),.B(g10404),.C(g10467));
  NOR3 NOR3_157(.VSS(VSS),.VDD(VDD),.Y(g12121),.A(g10330),.B(g10406),.C(g10470));
  NOR3 NOR3_158(.VSS(VSS),.VDD(VDD),.Y(g12124),.A(g10353),.B(g10413),.C(g10475));
  NOR3 NOR3_159(.VSS(VSS),.VDD(VDD),.Y(g12145),.A(g10364),.B(g10431),.C(g10492));
  NOR3 NOR3_160(.VSS(VSS),.VDD(VDD),.Y(g12146),.A(g10369),.B(g10436),.C(g10496));
  NOR3 NOR3_161(.VSS(VSS),.VDD(VDD),.Y(g12151),.A(g10374),.B(g10440),.C(g10498));
  NOR3 NOR3_162(.VSS(VSS),.VDD(VDD),.Y(g12152),.A(g10378),.B(g10442),.C(g10506));
  NOR3 NOR3_163(.VSS(VSS),.VDD(VDD),.Y(g12153),.A(g10380),.B(g10445),.C(g10509));
  NOR3 NOR3_164(.VSS(VSS),.VDD(VDD),.Y(g12154),.A(g10383),.B(g10447),.C(g10511));
  NOR3 NOR3_165(.VSS(VSS),.VDD(VDD),.Y(g12155),.A(g10386),.B(g10450),.C(g10514));
  NOR3 NOR3_166(.VSS(VSS),.VDD(VDD),.Y(g12162),.A(g10390),.B(g10452),.C(g10515));
  NOR3 NOR3_167(.VSS(VSS),.VDD(VDD),.Y(g12169),.A(g10394),.B(g10456),.C(g10517));
  NOR3 NOR3_168(.VSS(VSS),.VDD(VDD),.Y(g12170),.A(g10395),.B(g10458),.C(g10520));
  NOR3 NOR3_169(.VSS(VSS),.VDD(VDD),.Y(g12171),.A(g10398),.B(g10461),.C(g10522));
  NOR3 NOR3_170(.VSS(VSS),.VDD(VDD),.Y(g12172),.A(g10400),.B(g10464),.C(g10525));
  NOR3 NOR3_171(.VSS(VSS),.VDD(VDD),.Y(g12179),.A(g10405),.B(g10468),.C(g10527));
  NOR3 NOR3_172(.VSS(VSS),.VDD(VDD),.Y(g12180),.A(g10407),.B(g10471),.C(g10530));
  NOR3 NOR3_173(.VSS(VSS),.VDD(VDD),.Y(g12184),.A(g10414),.B(g10476),.C(g10536));
  NOR3 NOR3_174(.VSS(VSS),.VDD(VDD),.Y(g12185),.A(g10415),.B(g10478),.C(g10539));
  NOR3 NOR3_175(.VSS(VSS),.VDD(VDD),.Y(g12192),.A(g10423),.B(g10485),.C(g10548));
  NOR3 NOR3_176(.VSS(VSS),.VDD(VDD),.Y(g12193),.A(g10432),.B(g10493),.C(g10555));
  NOR3 NOR3_177(.VSS(VSS),.VDD(VDD),.Y(g12194),.A(g10434),.B(g10494),.C(g10556));
  NOR3 NOR3_178(.VSS(VSS),.VDD(VDD),.Y(g12195),.A(g10437),.B(g10497),.C(g10558));
  NOR3 NOR3_179(.VSS(VSS),.VDD(VDD),.Y(g12207),.A(g10443),.B(g10507),.C(g10566));
  NOR3 NOR3_180(.VSS(VSS),.VDD(VDD),.Y(g12208),.A(g10448),.B(g10512),.C(g10570));
  NOR3 NOR3_181(.VSS(VSS),.VDD(VDD),.Y(g12213),.A(g10453),.B(g10516),.C(g10572));
  NOR3 NOR3_182(.VSS(VSS),.VDD(VDD),.Y(g12214),.A(g10457),.B(g10518),.C(g10580));
  NOR3 NOR3_183(.VSS(VSS),.VDD(VDD),.Y(g12215),.A(g10459),.B(g10521),.C(g10583));
  NOR3 NOR3_184(.VSS(VSS),.VDD(VDD),.Y(g12216),.A(g10462),.B(g10523),.C(g10585));
  NOR3 NOR3_185(.VSS(VSS),.VDD(VDD),.Y(g12217),.A(g10465),.B(g10526),.C(g10588));
  NOR3 NOR3_186(.VSS(VSS),.VDD(VDD),.Y(g12224),.A(g10469),.B(g10528),.C(g10589));
  NOR3 NOR3_187(.VSS(VSS),.VDD(VDD),.Y(g12231),.A(g10473),.B(g10532),.C(g10591));
  NOR3 NOR3_188(.VSS(VSS),.VDD(VDD),.Y(g12232),.A(g10474),.B(g10534),.C(g10594));
  NOR3 NOR3_189(.VSS(VSS),.VDD(VDD),.Y(g12233),.A(g10477),.B(g10537),.C(g10596));
  NOR3 NOR3_190(.VSS(VSS),.VDD(VDD),.Y(g12234),.A(g10479),.B(g10540),.C(g10599));
  NOR3 NOR3_191(.VSS(VSS),.VDD(VDD),.Y(g12245),.A(g10495),.B(g10557),.C(g10604));
  NOR3 NOR3_192(.VSS(VSS),.VDD(VDD),.Y(g12247),.A(g10499),.B(g10559),.C(g10605));
  NOR3 NOR3_193(.VSS(VSS),.VDD(VDD),.Y(g12248),.A(g10508),.B(g10567),.C(g10612));
  NOR3 NOR3_194(.VSS(VSS),.VDD(VDD),.Y(g12249),.A(g10510),.B(g10568),.C(g10613));
  NOR3 NOR3_195(.VSS(VSS),.VDD(VDD),.Y(g12250),.A(g10513),.B(g10571),.C(g10615));
  NOR3 NOR3_196(.VSS(VSS),.VDD(VDD),.Y(g12262),.A(g10519),.B(g10581),.C(g10623));
  NOR3 NOR3_197(.VSS(VSS),.VDD(VDD),.Y(g12263),.A(g10524),.B(g10586),.C(g10627));
  NOR3 NOR3_198(.VSS(VSS),.VDD(VDD),.Y(g12268),.A(g10529),.B(g10590),.C(g10629));
  NOR3 NOR3_199(.VSS(VSS),.VDD(VDD),.Y(g12269),.A(g10533),.B(g10592),.C(g10637));
  NOR3 NOR3_200(.VSS(VSS),.VDD(VDD),.Y(g12270),.A(g10535),.B(g10595),.C(g10640));
  NOR3 NOR3_201(.VSS(VSS),.VDD(VDD),.Y(g12271),.A(g10538),.B(g10597),.C(g10642));
  NOR3 NOR3_202(.VSS(VSS),.VDD(VDD),.Y(g12272),.A(g10541),.B(g10600),.C(g10645));
  NOR3 NOR3_203(.VSS(VSS),.VDD(VDD),.Y(g12288),.A(g10569),.B(g10614),.C(g10651));
  NOR3 NOR3_204(.VSS(VSS),.VDD(VDD),.Y(g12290),.A(g10573),.B(g10616),.C(g10652));
  NOR3 NOR3_205(.VSS(VSS),.VDD(VDD),.Y(g12291),.A(g10582),.B(g10624),.C(g10659));
  NOR3 NOR3_206(.VSS(VSS),.VDD(VDD),.Y(g12292),.A(g10584),.B(g10625),.C(g10660));
  NOR3 NOR3_207(.VSS(VSS),.VDD(VDD),.Y(g12293),.A(g10587),.B(g10628),.C(g10662));
  NOR3 NOR3_208(.VSS(VSS),.VDD(VDD),.Y(g12305),.A(g10593),.B(g10638),.C(g10670));
  NOR3 NOR3_209(.VSS(VSS),.VDD(VDD),.Y(g12306),.A(g10598),.B(g10643),.C(g10674));
  NOR3 NOR3_210(.VSS(VSS),.VDD(VDD),.Y(g12324),.A(g10626),.B(g10661),.C(g10681));
  NOR3 NOR3_211(.VSS(VSS),.VDD(VDD),.Y(g12326),.A(g10630),.B(g10663),.C(g10682));
  NOR3 NOR3_212(.VSS(VSS),.VDD(VDD),.Y(g12327),.A(g10639),.B(g10671),.C(g10689));
  NOR3 NOR3_213(.VSS(VSS),.VDD(VDD),.Y(g12328),.A(g10641),.B(g10672),.C(g10690));
  NOR3 NOR3_214(.VSS(VSS),.VDD(VDD),.Y(g12329),.A(g10644),.B(g10675),.C(g10692));
  NOR3 NOR3_215(.VSS(VSS),.VDD(VDD),.Y(g12339),.A(g10650),.B(g10678),.C(g10704));
  NOR3 NOR3_216(.VSS(VSS),.VDD(VDD),.Y(g12352),.A(g10673),.B(g10691),.C(g10710));
  NOR3 NOR3_217(.VSS(VSS),.VDD(VDD),.Y(g12369),.A(g10680),.B(g10707),.C(g10724));
  NOR3 NOR3_218(.VSS(VSS),.VDD(VDD),.Y(g12388),.A(g10709),.B(g10727),.C(g10745));
  NOR3 NOR3_219(.VSS(VSS),.VDD(VDD),.Y(g12418),.A(g10729),.B(g10748),.C(g10764));
  NOR2 NOR2_2(.VSS(VSS),.VDD(VDD),.Y(g12431),.A(g8580),.B(g10730));
  NOR2 NOR2_3(.VSS(VSS),.VDD(VDD),.Y(g12436),.A(g8587),.B(g10749));
  NOR2 NOR2_4(.VSS(VSS),.VDD(VDD),.Y(g12441),.A(g8594),.B(g10767));
  NOR2 NOR2_5(.VSS(VSS),.VDD(VDD),.Y(g12446),.A(g8605),.B(g10773));
  NOR2 NOR2_6(.VSS(VSS),.VDD(VDD),.Y(g12451),.A(g499),.B(g8983));
  NOR3 NOR3_220(.VSS(VSS),.VDD(VDD),.Y(g12457),.A(g9009),.B(g9033),.C(g9048));
  NOR3 NOR3_221(.VSS(VSS),.VDD(VDD),.Y(g12467),.A(g9034),.B(g9056),.C(g9065));
  NOR3 NOR3_222(.VSS(VSS),.VDD(VDD),.Y(g12482),.A(g9057),.B(g9073),.C(g9082));
  NOR3 NOR3_223(.VSS(VSS),.VDD(VDD),.Y(g12487),.A(g10108),.B(g10198),.C(g10283));
  NOR3 NOR3_224(.VSS(VSS),.VDD(VDD),.Y(g12499),.A(g9074),.B(g9090),.C(g9101));
  NOR3 NOR3_225(.VSS(VSS),.VDD(VDD),.Y(g12507),.A(g10213),.B(g10300),.C(g10376));
  NOR3 NOR3_226(.VSS(VSS),.VDD(VDD),.Y(g12524),.A(g10315),.B(g10393),.C(g10455));
  NOR3 NOR3_227(.VSS(VSS),.VDD(VDD),.Y(g12539),.A(g10408),.B(g10472),.C(g10531));
  NOR3 NOR3_228(.VSS(VSS),.VDD(VDD),.Y(g12698),.A(g11347),.B(g11420),.C(g8327));
  NOR3 NOR3_229(.VSS(VSS),.VDD(VDD),.Y(g12747),.A(g11421),.B(g8328),.C(g8385));
  NOR3 NOR3_230(.VSS(VSS),.VDD(VDD),.Y(g12755),.A(g11431),.B(g8339),.C(g8394));
  NOR2 NOR2_7(.VSS(VSS),.VDD(VDD),.Y(g12780),.A(g9187),.B(g9161));
  NOR3 NOR3_231(.VSS(VSS),.VDD(VDD),.Y(g12781),.A(g8329),.B(g8386),.C(g8431));
  NOR3 NOR3_232(.VSS(VSS),.VDD(VDD),.Y(g12789),.A(g8340),.B(g8395),.C(g8437));
  NOR3 NOR3_233(.VSS(VSS),.VDD(VDD),.Y(g12797),.A(g8350),.B(g8406),.C(g8446));
  NOR3 NOR3_234(.VSS(VSS),.VDD(VDD),.Y(g12814),.A(g8387),.B(g8432),.C(g8463));
  NOR2 NOR2_8(.VSS(VSS),.VDD(VDD),.Y(g12819),.A(g9248),.B(g9203));
  NOR3 NOR3_235(.VSS(VSS),.VDD(VDD),.Y(g12820),.A(g8396),.B(g8438),.C(g8466));
  NOR3 NOR3_236(.VSS(VSS),.VDD(VDD),.Y(g12828),.A(g8407),.B(g8447),.C(g8472));
  NOR3 NOR3_237(.VSS(VSS),.VDD(VDD),.Y(g12836),.A(g8417),.B(g8458),.C(g8481));
  NOR3 NOR3_238(.VSS(VSS),.VDD(VDD),.Y(g12849),.A(g8433),.B(g8464),.C(g8485));
  NOR3 NOR3_239(.VSS(VSS),.VDD(VDD),.Y(g12852),.A(g8439),.B(g8467),.C(g8488));
  NOR2 NOR2_9(.VSS(VSS),.VDD(VDD),.Y(g12857),.A(g9326),.B(g9264));
  NOR3 NOR3_240(.VSS(VSS),.VDD(VDD),.Y(g12858),.A(g8448),.B(g8473),.C(g8491));
  NOR3 NOR3_241(.VSS(VSS),.VDD(VDD),.Y(g12866),.A(g8459),.B(g8482),.C(g8497));
  NOR3 NOR3_242(.VSS(VSS),.VDD(VDD),.Y(g12880),.A(g8465),.B(g8486),.C(g8502));
  NOR2 NOR2_10(.VSS(VSS),.VDD(VDD),.Y(g12883),.A(g10038),.B(g6284));
  NOR3 NOR3_243(.VSS(VSS),.VDD(VDD),.Y(g12890),.A(g8468),.B(g8489),.C(g8505));
  NOR3 NOR3_244(.VSS(VSS),.VDD(VDD),.Y(g12893),.A(g8474),.B(g8492),.C(g8508));
  NOR2 NOR2_11(.VSS(VSS),.VDD(VDD),.Y(g12898),.A(g9407),.B(g9342));
  NOR3 NOR3_245(.VSS(VSS),.VDD(VDD),.Y(g12899),.A(g8483),.B(g8498),.C(g8511));
  NOR3 NOR3_246(.VSS(VSS),.VDD(VDD),.Y(g12912),.A(g8484),.B(g8500),.C(g8515));
  NOR3 NOR3_247(.VSS(VSS),.VDD(VDD),.Y(g12913),.A(g8487),.B(g8503),.C(g8518));
  NOR3 NOR3_248(.VSS(VSS),.VDD(VDD),.Y(g12920),.A(g8490),.B(g8506),.C(g8521));
  NOR2 NOR2_12(.VSS(VSS),.VDD(VDD),.Y(g12923),.A(g10147),.B(g6421));
  NOR3 NOR3_249(.VSS(VSS),.VDD(VDD),.Y(g12930),.A(g8493),.B(g8509),.C(g8524));
  NOR3 NOR3_250(.VSS(VSS),.VDD(VDD),.Y(g12933),.A(g8499),.B(g8512),.C(g8527));
  NOR3 NOR3_251(.VSS(VSS),.VDD(VDD),.Y(g12939),.A(g8501),.B(g8516),.C(g8531));
  NOR3 NOR3_252(.VSS(VSS),.VDD(VDD),.Y(g12941),.A(g8504),.B(g8519),.C(g8534));
  NOR3 NOR3_253(.VSS(VSS),.VDD(VDD),.Y(g12942),.A(g8507),.B(g8522),.C(g8537));
  NOR3 NOR3_254(.VSS(VSS),.VDD(VDD),.Y(g12949),.A(g8510),.B(g8525),.C(g8540));
  NOR2 NOR2_13(.VSS(VSS),.VDD(VDD),.Y(g12952),.A(g10252),.B(g6626));
  NOR3 NOR3_255(.VSS(VSS),.VDD(VDD),.Y(g12959),.A(g8513),.B(g8528),.C(g8543));
  NOR3 NOR3_256(.VSS(VSS),.VDD(VDD),.Y(g12967),.A(g8517),.B(g8532),.C(g8546));
  NOR3 NOR3_257(.VSS(VSS),.VDD(VDD),.Y(g12968),.A(g8520),.B(g8535),.C(g8548));
  NOR3 NOR3_258(.VSS(VSS),.VDD(VDD),.Y(g12970),.A(g8523),.B(g8538),.C(g8551));
  NOR3 NOR3_259(.VSS(VSS),.VDD(VDD),.Y(g12971),.A(g8526),.B(g8541),.C(g8554));
  NOR3 NOR3_260(.VSS(VSS),.VDD(VDD),.Y(g12978),.A(g8529),.B(g8544),.C(g8557));
  NOR2 NOR2_14(.VSS(VSS),.VDD(VDD),.Y(g12981),.A(g10354),.B(g6890));
  NOR3 NOR3_261(.VSS(VSS),.VDD(VDD),.Y(g12991),.A(g8536),.B(g8549),.C(g8559));
  NOR3 NOR3_262(.VSS(VSS),.VDD(VDD),.Y(g12992),.A(g8539),.B(g8552),.C(g8561));
  NOR3 NOR3_263(.VSS(VSS),.VDD(VDD),.Y(g12994),.A(g8542),.B(g8555),.C(g8564));
  NOR3 NOR3_264(.VSS(VSS),.VDD(VDD),.Y(g12995),.A(g8545),.B(g8558),.C(g8567));
  NOR3 NOR3_265(.VSS(VSS),.VDD(VDD),.Y(g13001),.A(g8553),.B(g8562),.C(g8570));
  NOR3 NOR3_266(.VSS(VSS),.VDD(VDD),.Y(g13002),.A(g8556),.B(g8565),.C(g8572));
  NOR3 NOR3_267(.VSS(VSS),.VDD(VDD),.Y(g13022),.A(g8566),.B(g8573),.C(g8576));
  NOR4 NOR4_4(.VSS(VSS),.VDD(VDD),.Y(g13024),.A(g11481),.B(g8045),.C(g7928),.D(g7880));
  NOR3 NOR3_268(.VSS(VSS),.VDD(VDD),.Y(g13111),.A(g8601),.B(g8612),.C(g8621));
  NOR3 NOR3_269(.VSS(VSS),.VDD(VDD),.Y(g13124),.A(g8613),.B(g8625),.C(g8631));
  NOR3 NOR3_270(.VSS(VSS),.VDD(VDD),.Y(g13135),.A(g8626),.B(g8635),.C(g8650));
  NOR3 NOR3_271(.VSS(VSS),.VDD(VDD),.Y(g13143),.A(g8636),.B(g8654),.C(g8666));
  NOR3 NOR3_272(.VSS(VSS),.VDD(VDD),.Y(g13149),.A(g8676),.B(g8687),.C(g8703));
  NOR3 NOR3_273(.VSS(VSS),.VDD(VDD),.Y(g13155),.A(g8688),.B(g8705),.C(g8722));
  NOR3 NOR3_274(.VSS(VSS),.VDD(VDD),.Y(g13160),.A(g8704),.B(g8717),.C(g8751));
  NOR3 NOR3_275(.VSS(VSS),.VDD(VDD),.Y(g13164),.A(g8706),.B(g8724),.C(g8760));
  NOR3 NOR3_276(.VSS(VSS),.VDD(VDD),.Y(g13171),.A(g8723),.B(g8755),.C(g8774));
  NOR3 NOR3_277(.VSS(VSS),.VDD(VDD),.Y(g13175),.A(g8725),.B(g8762),.C(g8783));
  NOR3 NOR3_278(.VSS(VSS),.VDD(VDD),.Y(g13182),.A(g8761),.B(g8778),.C(g8797));
  NOR3 NOR3_279(.VSS(VSS),.VDD(VDD),.Y(g13194),.A(g8784),.B(g8801),.C(g8816));
  NOR3 NOR3_280(.VSS(VSS),.VDD(VDD),.Y(g13228),.A(g8841),.B(g8861),.C(g8892));
  NOR3 NOR3_281(.VSS(VSS),.VDD(VDD),.Y(g13251),.A(g8868),.B(g8899),.C(g8932));
  NOR3 NOR3_282(.VSS(VSS),.VDD(VDD),.Y(g13274),.A(g8906),.B(g8939),.C(g8972));
  NOR4 NOR4_5(.VSS(VSS),.VDD(VDD),.Y(g13286),.A(g11481),.B(g11332),.C(g11190),.D(g7880));
  NOR3 NOR3_283(.VSS(VSS),.VDD(VDD),.Y(g13299),.A(g8946),.B(g8979),.C(g9004));
  NOR4 NOR4_6(.VSS(VSS),.VDD(VDD),.Y(g13310),.A(g11481),.B(g11332),.C(g11190),.D(g11069));
  NOR4 NOR4_7(.VSS(VSS),.VDD(VDD),.Y(g13313),.A(g8183),.B(g11332),.C(g11190),.D(g7880));
  NOR4 NOR4_8(.VSS(VSS),.VDD(VDD),.Y(g13331),.A(g8183),.B(g11332),.C(g11190),.D(g11069));
  NOR4 NOR4_9(.VSS(VSS),.VDD(VDD),.Y(g13332),.A(g11481),.B(g8045),.C(g11190),.D(g7880));
  NOR4 NOR4_10(.VSS(VSS),.VDD(VDD),.Y(g13353),.A(g11481),.B(g8045),.C(g11190),.D(g11069));
  NOR4 NOR4_11(.VSS(VSS),.VDD(VDD),.Y(g13354),.A(g8183),.B(g8045),.C(g11190),.D(g7880));
  NOR4 NOR4_12(.VSS(VSS),.VDD(VDD),.Y(g13374),.A(g8183),.B(g8045),.C(g11190),.D(g11069));
  NOR4 NOR4_13(.VSS(VSS),.VDD(VDD),.Y(g13375),.A(g11481),.B(g11332),.C(g7928),.D(g7880));
  NOR3 NOR3_284(.VSS(VSS),.VDD(VDD),.Y(g13378),.A(g9026),.B(g9047),.C(g9061));
  NOR4 NOR4_14(.VSS(VSS),.VDD(VDD),.Y(g13401),.A(g11481),.B(g11332),.C(g7928),.D(g11069));
  NOR4 NOR4_15(.VSS(VSS),.VDD(VDD),.Y(g13404),.A(g8183),.B(g11332),.C(g7928),.D(g7880));
  NOR2 NOR2_15(.VSS(VSS),.VDD(VDD),.Y(g15661),.A(g11737),.B(g7345));
  NOR2 NOR2_16(.VSS(VSS),.VDD(VDD),.Y(g15797),.A(g13305),.B(g7143));
  NOR2 NOR2_17(.VSS(VSS),.VDD(VDD),.Y(g15873),.A(g11617),.B(g7562));
  NOR2 NOR2_18(.VSS(VSS),.VDD(VDD),.Y(g15959),.A(g2814),.B(g13082));
  NOR2 NOR2_19(.VSS(VSS),.VDD(VDD),.Y(g15978),.A(g11737),.B(g7152));
  NOR3 NOR3_285(.VSS(VSS),.VDD(VDD),.Y(g16020),.A(g6200),.B(g12457),.C(g10952));
  NOR3 NOR3_286(.VSS(VSS),.VDD(VDD),.Y(g16036),.A(g6289),.B(g12467),.C(g10952));
  NOR3 NOR3_287(.VSS(VSS),.VDD(VDD),.Y(g16058),.A(g6426),.B(g12482),.C(g10952));
  NOR3 NOR3_288(.VSS(VSS),.VDD(VDD),.Y(g16082),.A(g10952),.B(g6140),.C(g12487));
  NOR3 NOR3_289(.VSS(VSS),.VDD(VDD),.Y(g16094),.A(g6631),.B(g12499),.C(g10952));
  NOR3 NOR3_290(.VSS(VSS),.VDD(VDD),.Y(g16120),.A(g10952),.B(g6161),.C(g12507));
  NOR3 NOR3_291(.VSS(VSS),.VDD(VDD),.Y(g16171),.A(g10952),.B(g6188),.C(g12524));
  NOR3 NOR3_292(.VSS(VSS),.VDD(VDD),.Y(g16230),.A(g10952),.B(g6220),.C(g12539));
  NOR2 NOR2_20(.VSS(VSS),.VDD(VDD),.Y(g16498),.A(g14158),.B(g14347));
  NOR2 NOR2_21(.VSS(VSS),.VDD(VDD),.Y(g16520),.A(g14273),.B(g14459));
  NOR2 NOR2_22(.VSS(VSS),.VDD(VDD),.Y(g16551),.A(g14395),.B(g14546));
  NOR3 NOR3_293(.VSS(VSS),.VDD(VDD),.Y(g16567),.A(g15904),.B(g15880),.C(g15859));
  NOR3 NOR3_294(.VSS(VSS),.VDD(VDD),.Y(g16570),.A(g15904),.B(g15880),.C(g14630));
  NOR2 NOR2_23(.VSS(VSS),.VDD(VDD),.Y(g16583),.A(g14507),.B(g14601));
  NOR3 NOR3_295(.VSS(VSS),.VDD(VDD),.Y(g16591),.A(g15933),.B(g15913),.C(g15890));
  NOR3 NOR3_296(.VSS(VSS),.VDD(VDD),.Y(g16594),.A(g15933),.B(g15913),.C(g14650));
  NOR3 NOR3_297(.VSS(VSS),.VDD(VDD),.Y(g16611),.A(g15962),.B(g15942),.C(g15923));
  NOR3 NOR3_298(.VSS(VSS),.VDD(VDD),.Y(g16614),.A(g15962),.B(g15942),.C(g14677));
  NOR3 NOR3_299(.VSS(VSS),.VDD(VDD),.Y(g16629),.A(g15981),.B(g15971),.C(g15952));
  NOR3 NOR3_300(.VSS(VSS),.VDD(VDD),.Y(g16632),.A(g15981),.B(g15971),.C(g14711));
  NOR3 NOR3_301(.VSS(VSS),.VDD(VDD),.Y(g16643),.A(g15904),.B(g14642),.C(g15859));
  NOR2 NOR2_24(.VSS(VSS),.VDD(VDD),.Y(g16654),.A(g14690),.B(g12477));
  NOR3 NOR3_302(.VSS(VSS),.VDD(VDD),.Y(g16655),.A(g15933),.B(g14669),.C(g15890));
  NOR2 NOR2_25(.VSS(VSS),.VDD(VDD),.Y(g16671),.A(g14724),.B(g12494));
  NOR3 NOR3_303(.VSS(VSS),.VDD(VDD),.Y(g16672),.A(g15962),.B(g14703),.C(g15923));
  NOR2 NOR2_26(.VSS(VSS),.VDD(VDD),.Y(g16679),.A(g14797),.B(g14895));
  NOR2 NOR2_27(.VSS(VSS),.VDD(VDD),.Y(g16692),.A(g14752),.B(g12514));
  NOR3 NOR3_304(.VSS(VSS),.VDD(VDD),.Y(g16693),.A(g15981),.B(g14737),.C(g15952));
  NOR2 NOR2_28(.VSS(VSS),.VDD(VDD),.Y(g16705),.A(g14849),.B(g14976));
  NOR2 NOR2_29(.VSS(VSS),.VDD(VDD),.Y(g16718),.A(g14773),.B(g12531));
  NOR2 NOR2_30(.VSS(VSS),.VDD(VDD),.Y(g16736),.A(g14922),.B(g15065));
  NOR2 NOR2_31(.VSS(VSS),.VDD(VDD),.Y(g16778),.A(g15003),.B(g15161));
  NOR2 NOR2_32(.VSS(VSS),.VDD(VDD),.Y(g16802),.A(g13469),.B(g3897));
  NOR2 NOR2_33(.VSS(VSS),.VDD(VDD),.Y(g16803),.A(g15593),.B(g12908));
  NOR2 NOR2_34(.VSS(VSS),.VDD(VDD),.Y(g16823),.A(g5362),.B(g13469));
  NOR2 NOR2_35(.VSS(VSS),.VDD(VDD),.Y(g16824),.A(g15658),.B(g12938));
  NOR2 NOR2_36(.VSS(VSS),.VDD(VDD),.Y(g16829),.A(g14956),.B(g12564));
  NOR2 NOR2_37(.VSS(VSS),.VDD(VDD),.Y(g16835),.A(g15717),.B(g12966));
  NOR2 NOR2_38(.VSS(VSS),.VDD(VDD),.Y(g16841),.A(g15021),.B(g12607));
  NOR2 NOR2_39(.VSS(VSS),.VDD(VDD),.Y(g16844),.A(g15754),.B(g12989));
  NOR2 NOR2_40(.VSS(VSS),.VDD(VDD),.Y(g16845),.A(g15755),.B(g12990));
  NOR2 NOR2_41(.VSS(VSS),.VDD(VDD),.Y(g16847),.A(g15095),.B(g12650));
  NOR2 NOR2_42(.VSS(VSS),.VDD(VDD),.Y(g16851),.A(g15781),.B(g13000));
  NOR2 NOR2_43(.VSS(VSS),.VDD(VDD),.Y(g16853),.A(g15801),.B(g13009));
  NOR2 NOR2_44(.VSS(VSS),.VDD(VDD),.Y(g16854),.A(g15802),.B(g13010));
  NOR2 NOR2_45(.VSS(VSS),.VDD(VDD),.Y(g16857),.A(g15817),.B(g13023));
  NOR2 NOR2_46(.VSS(VSS),.VDD(VDD),.Y(g16860),.A(g15828),.B(g13031));
  NOR2 NOR2_47(.VSS(VSS),.VDD(VDD),.Y(g16861),.A(g15829),.B(g13032));
  NOR2 NOR2_48(.VSS(VSS),.VDD(VDD),.Y(g16866),.A(g15840),.B(g13042));
  NOR2 NOR2_49(.VSS(VSS),.VDD(VDD),.Y(g16880),.A(g15852),.B(g13056));
  NOR3 NOR3_305(.VSS(VSS),.VDD(VDD),.Y(g17012),.A(g14657),.B(g14642),.C(g15859));
  NOR3 NOR3_306(.VSS(VSS),.VDD(VDD),.Y(g17025),.A(g15904),.B(g15880),.C(g15859));
  NOR3 NOR3_307(.VSS(VSS),.VDD(VDD),.Y(g17042),.A(g14691),.B(g14669),.C(g15890));
  NOR3 NOR3_308(.VSS(VSS),.VDD(VDD),.Y(g17051),.A(g14657),.B(g15880),.C(g14630));
  NOR3 NOR3_309(.VSS(VSS),.VDD(VDD),.Y(g17059),.A(g15933),.B(g15913),.C(g15890));
  NOR3 NOR3_310(.VSS(VSS),.VDD(VDD),.Y(g17076),.A(g14725),.B(g14703),.C(g15923));
  NOR3 NOR3_311(.VSS(VSS),.VDD(VDD),.Y(g17086),.A(g14691),.B(g15913),.C(g14650));
  NOR3 NOR3_312(.VSS(VSS),.VDD(VDD),.Y(g17094),.A(g15962),.B(g15942),.C(g15923));
  NOR3 NOR3_313(.VSS(VSS),.VDD(VDD),.Y(g17111),.A(g14753),.B(g14737),.C(g15952));
  NOR3 NOR3_314(.VSS(VSS),.VDD(VDD),.Y(g17124),.A(g14725),.B(g15942),.C(g14677));
  NOR3 NOR3_315(.VSS(VSS),.VDD(VDD),.Y(g17132),.A(g15981),.B(g15971),.C(g15952));
  NOR3 NOR3_316(.VSS(VSS),.VDD(VDD),.Y(g17151),.A(g14753),.B(g15971),.C(g14711));
  NOR2 NOR2_50(.VSS(VSS),.VDD(VDD),.Y(g17186),.A(g7949),.B(g14144));
  NOR2 NOR2_51(.VSS(VSS),.VDD(VDD),.Y(g17197),.A(g8000),.B(g14259));
  NOR2 NOR2_52(.VSS(VSS),.VDD(VDD),.Y(g17204),.A(g8075),.B(g14381));
  NOR2 NOR2_53(.VSS(VSS),.VDD(VDD),.Y(g17209),.A(g8160),.B(g14493));
  NOR2 NOR2_54(.VSS(VSS),.VDD(VDD),.Y(g17213),.A(g4326),.B(g14442));
  NOR2 NOR2_55(.VSS(VSS),.VDD(VDD),.Y(g17215),.A(g15904),.B(g14642));
  NOR2 NOR2_56(.VSS(VSS),.VDD(VDD),.Y(g17216),.A(g4495),.B(g14529));
  NOR2 NOR2_57(.VSS(VSS),.VDD(VDD),.Y(g17218),.A(g15933),.B(g14669));
  NOR2 NOR2_58(.VSS(VSS),.VDD(VDD),.Y(g17219),.A(g4671),.B(g14584));
  NOR2 NOR2_59(.VSS(VSS),.VDD(VDD),.Y(g17220),.A(g15962),.B(g14703));
  NOR2 NOR2_60(.VSS(VSS),.VDD(VDD),.Y(g17221),.A(g4848),.B(g14618));
  NOR2 NOR2_61(.VSS(VSS),.VDD(VDD),.Y(g17222),.A(g15998),.B(g16003));
  NOR2 NOR2_62(.VSS(VSS),.VDD(VDD),.Y(g17223),.A(g15981),.B(g14737));
  NOR2 NOR2_63(.VSS(VSS),.VDD(VDD),.Y(g17224),.A(g16004),.B(g16009));
  NOR2 NOR2_64(.VSS(VSS),.VDD(VDD),.Y(g17225),.A(g16008),.B(g16015));
  NOR2 NOR2_65(.VSS(VSS),.VDD(VDD),.Y(g17226),.A(g16010),.B(g16017));
  NOR2 NOR2_66(.VSS(VSS),.VDD(VDD),.Y(g17228),.A(g16016),.B(g16029));
  NOR2 NOR2_67(.VSS(VSS),.VDD(VDD),.Y(g17229),.A(g16019),.B(g16032));
  NOR2 NOR2_68(.VSS(VSS),.VDD(VDD),.Y(g17234),.A(g16028),.B(g16045));
  NOR2 NOR2_69(.VSS(VSS),.VDD(VDD),.Y(g17235),.A(g16030),.B(g16047));
  NOR2 NOR2_70(.VSS(VSS),.VDD(VDD),.Y(g17236),.A(g16033),.B(g16051));
  NOR2 NOR2_71(.VSS(VSS),.VDD(VDD),.Y(g17246),.A(g16046),.B(g16066));
  NOR2 NOR2_72(.VSS(VSS),.VDD(VDD),.Y(g17247),.A(g16050),.B(g16070));
  NOR2 NOR2_73(.VSS(VSS),.VDD(VDD),.Y(g17248),.A(g16052),.B(g16072));
  NOR2 NOR2_74(.VSS(VSS),.VDD(VDD),.Y(g17269),.A(g16067),.B(g16100));
  NOR2 NOR2_75(.VSS(VSS),.VDD(VDD),.Y(g17270),.A(g16071),.B(g16104));
  NOR2 NOR2_76(.VSS(VSS),.VDD(VDD),.Y(g17271),.A(g16073),.B(g16106));
  NOR2 NOR2_77(.VSS(VSS),.VDD(VDD),.Y(g17302),.A(g16103),.B(g16135));
  NOR2 NOR2_78(.VSS(VSS),.VDD(VDD),.Y(g17303),.A(g16105),.B(g16137));
  NOR2 NOR2_79(.VSS(VSS),.VDD(VDD),.Y(g17340),.A(g16136),.B(g16183));
  NOR2 NOR2_80(.VSS(VSS),.VDD(VDD),.Y(g17341),.A(g16138),.B(g16185));
  NOR2 NOR2_81(.VSS(VSS),.VDD(VDD),.Y(g17383),.A(g16184),.B(g16238));
  NOR2 NOR2_82(.VSS(VSS),.VDD(VDD),.Y(g17429),.A(g16239),.B(g16288));
  NOR2 NOR2_83(.VSS(VSS),.VDD(VDD),.Y(g17507),.A(g16298),.B(g13318));
  NOR2 NOR2_84(.VSS(VSS),.VDD(VDD),.Y(g17896),.A(g14352),.B(g16020));
  NOR2 NOR2_85(.VSS(VSS),.VDD(VDD),.Y(g18007),.A(g14464),.B(g16036));
  NOR2 NOR2_86(.VSS(VSS),.VDD(VDD),.Y(g18085),.A(g16085),.B(g6363));
  NOR2 NOR2_87(.VSS(VSS),.VDD(VDD),.Y(g18124),.A(g14551),.B(g16058));
  NOR2 NOR2_88(.VSS(VSS),.VDD(VDD),.Y(g18201),.A(g16123),.B(g6568));
  NOR2 NOR2_89(.VSS(VSS),.VDD(VDD),.Y(g18240),.A(g14606),.B(g16094));
  NOR2 NOR2_90(.VSS(VSS),.VDD(VDD),.Y(g18308),.A(g16174),.B(g6832));
  NOR2 NOR2_91(.VSS(VSS),.VDD(VDD),.Y(g18352),.A(g16082),.B(g14249));
  NOR2 NOR2_92(.VSS(VSS),.VDD(VDD),.Y(g18401),.A(g16233),.B(g7134));
  NOR2 NOR2_93(.VSS(VSS),.VDD(VDD),.Y(g18430),.A(g16020),.B(g14352));
  NOR2 NOR2_94(.VSS(VSS),.VDD(VDD),.Y(g18447),.A(g16120),.B(g14371));
  NOR2 NOR2_95(.VSS(VSS),.VDD(VDD),.Y(g18503),.A(g16036),.B(g14464));
  NOR2 NOR2_96(.VSS(VSS),.VDD(VDD),.Y(g18520),.A(g16171),.B(g14483));
  NOR2 NOR2_97(.VSS(VSS),.VDD(VDD),.Y(g18548),.A(g14249),.B(g16082));
  NOR2 NOR2_98(.VSS(VSS),.VDD(VDD),.Y(g18567),.A(g16058),.B(g14551));
  NOR2 NOR2_99(.VSS(VSS),.VDD(VDD),.Y(g18584),.A(g16230),.B(g14570));
  NOR2 NOR2_100(.VSS(VSS),.VDD(VDD),.Y(g18590),.A(g16439),.B(g7522));
  NOR2 NOR2_101(.VSS(VSS),.VDD(VDD),.Y(g18598),.A(g14371),.B(g16120));
  NOR2 NOR2_102(.VSS(VSS),.VDD(VDD),.Y(g18617),.A(g16094),.B(g14606));
  NOR2 NOR2_103(.VSS(VSS),.VDD(VDD),.Y(g18623),.A(g15902),.B(g2814));
  NOR2 NOR2_104(.VSS(VSS),.VDD(VDD),.Y(g18626),.A(g16463),.B(g7549));
  NOR2 NOR2_105(.VSS(VSS),.VDD(VDD),.Y(g18630),.A(g14483),.B(g16171));
  NOR2 NOR2_106(.VSS(VSS),.VDD(VDD),.Y(g18639),.A(g14570),.B(g16230));
  NOR2 NOR2_107(.VSS(VSS),.VDD(VDD),.Y(g18669),.A(g13623),.B(g13634));
  NOR2 NOR2_108(.VSS(VSS),.VDD(VDD),.Y(g18678),.A(g13625),.B(g11771));
  NOR2 NOR2_109(.VSS(VSS),.VDD(VDD),.Y(g18707),.A(g13636),.B(g11788));
  NOR2 NOR2_110(.VSS(VSS),.VDD(VDD),.Y(g18719),.A(g13643),.B(g13656));
  NOR2 NOR2_111(.VSS(VSS),.VDD(VDD),.Y(g18726),.A(g13645),.B(g11805));
  NOR2 NOR2_112(.VSS(VSS),.VDD(VDD),.Y(g18743),.A(g13648),.B(g11814));
  NOR2 NOR2_113(.VSS(VSS),.VDD(VDD),.Y(g18754),.A(g13655),.B(g11816));
  NOR2 NOR2_114(.VSS(VSS),.VDD(VDD),.Y(g18755),.A(g13871),.B(g12274));
  NOR2 NOR2_115(.VSS(VSS),.VDD(VDD),.Y(g18763),.A(g13671),.B(g11838));
  NOR2 NOR2_116(.VSS(VSS),.VDD(VDD),.Y(g18780),.A(g13674),.B(g11847));
  NOR2 NOR2_117(.VSS(VSS),.VDD(VDD),.Y(g18781),.A(g13675),.B(g11851));
  NOR2 NOR2_118(.VSS(VSS),.VDD(VDD),.Y(g18782),.A(g13676),.B(g13705));
  NOR2 NOR2_119(.VSS(VSS),.VDD(VDD),.Y(g18794),.A(g13701),.B(g11880));
  NOR2 NOR2_120(.VSS(VSS),.VDD(VDD),.Y(g18803),.A(g13704),.B(g11885));
  NOR2 NOR2_121(.VSS(VSS),.VDD(VDD),.Y(g18804),.A(g13905),.B(g12331));
  NOR2 NOR2_122(.VSS(VSS),.VDD(VDD),.Y(g18820),.A(g13738),.B(g11922));
  NOR2 NOR2_123(.VSS(VSS),.VDD(VDD),.Y(g18821),.A(g13740),.B(g11926));
  NOR2 NOR2_124(.VSS(VSS),.VDD(VDD),.Y(g18835),.A(g13788),.B(g11966));
  NOR2 NOR2_125(.VSS(VSS),.VDD(VDD),.Y(g18836),.A(g13789),.B(g11967));
  NOR2 NOR2_126(.VSS(VSS),.VDD(VDD),.Y(g18837),.A(g13998),.B(g12376));
  NOR2 NOR2_127(.VSS(VSS),.VDD(VDD),.Y(g18852),.A(g13815),.B(g12012));
  NOR2 NOR2_128(.VSS(VSS),.VDD(VDD),.Y(g18866),.A(g13834),.B(g12069));
  NOR2 NOR2_129(.VSS(VSS),.VDD(VDD),.Y(g18867),.A(g13835),.B(g12070));
  NOR2 NOR2_130(.VSS(VSS),.VDD(VDD),.Y(g18868),.A(g14143),.B(g12419));
  NOR2 NOR2_131(.VSS(VSS),.VDD(VDD),.Y(g18883),.A(g13846),.B(g12128));
  NOR2 NOR2_132(.VSS(VSS),.VDD(VDD),.Y(g18885),.A(g13847),.B(g12129));
  NOR2 NOR2_133(.VSS(VSS),.VDD(VDD),.Y(g18906),.A(g13855),.B(g12186));
  NOR2 NOR2_134(.VSS(VSS),.VDD(VDD),.Y(g18907),.A(g14336),.B(g12429));
  NOR2 NOR2_135(.VSS(VSS),.VDD(VDD),.Y(g18942),.A(g13870),.B(g12273));
  NOR2 NOR2_136(.VSS(VSS),.VDD(VDD),.Y(g18957),.A(g13884),.B(g12307));
  NOR2 NOR2_137(.VSS(VSS),.VDD(VDD),.Y(g18968),.A(g13904),.B(g12330));
  NOR2 NOR2_138(.VSS(VSS),.VDD(VDD),.Y(g18975),.A(g13944),.B(g12353));
  NOR2 NOR2_139(.VSS(VSS),.VDD(VDD),.Y(g19144),.A(g17268),.B(g14884));
  NOR2 NOR2_140(.VSS(VSS),.VDD(VDD),.Y(g19149),.A(g17339),.B(g15020));
  NOR2 NOR2_141(.VSS(VSS),.VDD(VDD),.Y(g19153),.A(g17381),.B(g15093));
  NOR2 NOR2_142(.VSS(VSS),.VDD(VDD),.Y(g19154),.A(g17382),.B(g15094));
  NOR2 NOR2_143(.VSS(VSS),.VDD(VDD),.Y(g19157),.A(g17428),.B(g15171));
  NOR2 NOR2_144(.VSS(VSS),.VDD(VDD),.Y(g19160),.A(g17446),.B(g15178));
  NOR2 NOR2_145(.VSS(VSS),.VDD(VDD),.Y(g19162),.A(g17485),.B(g15243));
  NOR2 NOR2_146(.VSS(VSS),.VDD(VDD),.Y(g19163),.A(g17486),.B(g15244));
  NOR2 NOR2_147(.VSS(VSS),.VDD(VDD),.Y(g19165),.A(g17526),.B(g15264));
  NOR2 NOR2_148(.VSS(VSS),.VDD(VDD),.Y(g19167),.A(g17556),.B(g15320));
  NOR2 NOR2_149(.VSS(VSS),.VDD(VDD),.Y(g19171),.A(g17616),.B(g15356));
  NOR2 NOR2_150(.VSS(VSS),.VDD(VDD),.Y(g19172),.A(g17635),.B(g15388));
  NOR2 NOR2_151(.VSS(VSS),.VDD(VDD),.Y(g19173),.A(g17636),.B(g15389));
  NOR2 NOR2_152(.VSS(VSS),.VDD(VDD),.Y(g19177),.A(g17713),.B(g15442));
  NOR2 NOR2_153(.VSS(VSS),.VDD(VDD),.Y(g19178),.A(g17718),.B(g15452));
  NOR2 NOR2_154(.VSS(VSS),.VDD(VDD),.Y(g19179),.A(g17719),.B(g15453));
  NOR2 NOR2_155(.VSS(VSS),.VDD(VDD),.Y(g19184),.A(g17798),.B(g15520));
  NOR2 NOR2_156(.VSS(VSS),.VDD(VDD),.Y(g19219),.A(g18165),.B(g15753));
  NOR2 NOR2_157(.VSS(VSS),.VDD(VDD),.Y(g20008),.A(g18977),.B(g7338));
  NOR2 NOR2_158(.VSS(VSS),.VDD(VDD),.Y(g20054),.A(g19001),.B(g16867));
  NOR2 NOR2_159(.VSS(VSS),.VDD(VDD),.Y(g20095),.A(g16507),.B(g16895));
  NOR2 NOR2_160(.VSS(VSS),.VDD(VDD),.Y(g20120),.A(g16529),.B(g16924));
  NOR2 NOR2_161(.VSS(VSS),.VDD(VDD),.Y(g20150),.A(g16560),.B(g16954));
  NOR2 NOR2_162(.VSS(VSS),.VDD(VDD),.Y(g20153),.A(g16536),.B(g7583));
  NOR2 NOR2_163(.VSS(VSS),.VDD(VDD),.Y(g20299),.A(g16665),.B(g16884));
  NOR2 NOR2_164(.VSS(VSS),.VDD(VDD),.Y(g20310),.A(g16850),.B(g13654));
  NOR2 NOR2_165(.VSS(VSS),.VDD(VDD),.Y(g20314),.A(g13646),.B(g16855));
  NOR2 NOR2_166(.VSS(VSS),.VDD(VDD),.Y(g20318),.A(g16686),.B(g16913));
  NOR2 NOR2_167(.VSS(VSS),.VDD(VDD),.Y(g20333),.A(g13672),.B(g16859));
  NOR2 NOR2_168(.VSS(VSS),.VDD(VDD),.Y(g20337),.A(g16712),.B(g16943));
  NOR2 NOR2_169(.VSS(VSS),.VDD(VDD),.Y(g20343),.A(g16856),.B(g13703));
  NOR2 NOR2_170(.VSS(VSS),.VDD(VDD),.Y(g20353),.A(g13702),.B(g16864));
  NOR2 NOR2_171(.VSS(VSS),.VDD(VDD),.Y(g20357),.A(g16743),.B(g16974));
  NOR2 NOR2_172(.VSS(VSS),.VDD(VDD),.Y(g20375),.A(g13739),.B(g16879));
  NOR2 NOR2_173(.VSS(VSS),.VDD(VDD),.Y(g20376),.A(g16865),.B(g13787));
  NOR2 NOR2_174(.VSS(VSS),.VDD(VDD),.Y(g20417),.A(g16907),.B(g13833));
  NOR2 NOR2_175(.VSS(VSS),.VDD(VDD),.Y(g20682),.A(g19160),.B(g10024));
  NOR2 NOR2_176(.VSS(VSS),.VDD(VDD),.Y(g20717),.A(g19165),.B(g10133));
  NOR2 NOR2_177(.VSS(VSS),.VDD(VDD),.Y(g20752),.A(g19171),.B(g10238));
  NOR2 NOR2_178(.VSS(VSS),.VDD(VDD),.Y(g20789),.A(g19177),.B(g10340));
  NOR2 NOR2_179(.VSS(VSS),.VDD(VDD),.Y(g20841),.A(g14767),.B(g19552));
  NOR2 NOR2_180(.VSS(VSS),.VDD(VDD),.Y(g20874),.A(g17301),.B(g19594));
  NOR2 NOR2_181(.VSS(VSS),.VDD(VDD),.Y(g20875),.A(g19584),.B(g17352));
  NOR2 NOR2_182(.VSS(VSS),.VDD(VDD),.Y(g20876),.A(g19585),.B(g17353));
  NOR2 NOR2_183(.VSS(VSS),.VDD(VDD),.Y(g20877),.A(g3919),.B(g19830));
  NOR2 NOR2_184(.VSS(VSS),.VDD(VDD),.Y(g20878),.A(g19600),.B(g17395));
  NOR2 NOR2_185(.VSS(VSS),.VDD(VDD),.Y(g20879),.A(g19601),.B(g17396));
  NOR2 NOR2_186(.VSS(VSS),.VDD(VDD),.Y(g20880),.A(g19602),.B(g17397));
  NOR2 NOR2_187(.VSS(VSS),.VDD(VDD),.Y(g20881),.A(g19603),.B(g17398));
  NOR2 NOR2_188(.VSS(VSS),.VDD(VDD),.Y(g20882),.A(g19614),.B(g17408));
  NOR2 NOR2_189(.VSS(VSS),.VDD(VDD),.Y(g20883),.A(g19615),.B(g17409));
  NOR2 NOR2_190(.VSS(VSS),.VDD(VDD),.Y(g20884),.A(g5394),.B(g19830));
  NOR2 NOR2_191(.VSS(VSS),.VDD(VDD),.Y(g20891),.A(g19626),.B(g17447));
  NOR2 NOR2_192(.VSS(VSS),.VDD(VDD),.Y(g20892),.A(g19627),.B(g17448));
  NOR2 NOR2_193(.VSS(VSS),.VDD(VDD),.Y(g20893),.A(g19628),.B(g17449));
  NOR2 NOR2_194(.VSS(VSS),.VDD(VDD),.Y(g20894),.A(g19629),.B(g17450));
  NOR2 NOR2_195(.VSS(VSS),.VDD(VDD),.Y(g20895),.A(g19633),.B(g17461));
  NOR2 NOR2_196(.VSS(VSS),.VDD(VDD),.Y(g20896),.A(g19634),.B(g17462));
  NOR2 NOR2_197(.VSS(VSS),.VDD(VDD),.Y(g20897),.A(g19635),.B(g17463));
  NOR2 NOR2_198(.VSS(VSS),.VDD(VDD),.Y(g20898),.A(g19636),.B(g17464));
  NOR2 NOR2_199(.VSS(VSS),.VDD(VDD),.Y(g20899),.A(g19647),.B(g17474));
  NOR2 NOR2_200(.VSS(VSS),.VDD(VDD),.Y(g20900),.A(g19648),.B(g17475));
  NOR2 NOR2_201(.VSS(VSS),.VDD(VDD),.Y(g20901),.A(g19660),.B(g17508));
  NOR2 NOR2_202(.VSS(VSS),.VDD(VDD),.Y(g20902),.A(g19661),.B(g17509));
  NOR2 NOR2_203(.VSS(VSS),.VDD(VDD),.Y(g20903),.A(g19662),.B(g17510));
  NOR2 NOR2_204(.VSS(VSS),.VDD(VDD),.Y(g20910),.A(g19666),.B(g17527));
  NOR2 NOR2_205(.VSS(VSS),.VDD(VDD),.Y(g20911),.A(g19667),.B(g17528));
  NOR2 NOR2_206(.VSS(VSS),.VDD(VDD),.Y(g20912),.A(g19668),.B(g17529));
  NOR2 NOR2_207(.VSS(VSS),.VDD(VDD),.Y(g20913),.A(g19669),.B(g17530));
  NOR2 NOR2_208(.VSS(VSS),.VDD(VDD),.Y(g20914),.A(g19673),.B(g17541));
  NOR2 NOR2_209(.VSS(VSS),.VDD(VDD),.Y(g20915),.A(g19674),.B(g17542));
  NOR2 NOR2_210(.VSS(VSS),.VDD(VDD),.Y(g20916),.A(g19675),.B(g17543));
  NOR2 NOR2_211(.VSS(VSS),.VDD(VDD),.Y(g20917),.A(g19676),.B(g17544));
  NOR2 NOR2_212(.VSS(VSS),.VDD(VDD),.Y(g20918),.A(g19687),.B(g17554));
  NOR2 NOR2_213(.VSS(VSS),.VDD(VDD),.Y(g20919),.A(g19688),.B(g17555));
  NOR2 NOR2_214(.VSS(VSS),.VDD(VDD),.Y(g20920),.A(g19691),.B(g19726));
  NOR2 NOR2_215(.VSS(VSS),.VDD(VDD),.Y(g20921),.A(g19697),.B(g17576));
  NOR2 NOR2_216(.VSS(VSS),.VDD(VDD),.Y(g20922),.A(g19698),.B(g17577));
  NOR2 NOR2_217(.VSS(VSS),.VDD(VDD),.Y(g20923),.A(g19699),.B(g17578));
  NOR2 NOR2_218(.VSS(VSS),.VDD(VDD),.Y(g20924),.A(g19700),.B(g15257));
  NOR2 NOR2_219(.VSS(VSS),.VDD(VDD),.Y(g20925),.A(g19708),.B(g17598));
  NOR2 NOR2_220(.VSS(VSS),.VDD(VDD),.Y(g20926),.A(g19709),.B(g17599));
  NOR2 NOR2_221(.VSS(VSS),.VDD(VDD),.Y(g20927),.A(g19710),.B(g17600));
  NOR2 NOR2_222(.VSS(VSS),.VDD(VDD),.Y(g20934),.A(g19714),.B(g17617));
  NOR2 NOR2_223(.VSS(VSS),.VDD(VDD),.Y(g20935),.A(g19715),.B(g17618));
  NOR2 NOR2_224(.VSS(VSS),.VDD(VDD),.Y(g20936),.A(g19716),.B(g17619));
  NOR2 NOR2_225(.VSS(VSS),.VDD(VDD),.Y(g20937),.A(g19717),.B(g17620));
  NOR2 NOR2_226(.VSS(VSS),.VDD(VDD),.Y(g20938),.A(g19721),.B(g17631));
  NOR2 NOR2_227(.VSS(VSS),.VDD(VDD),.Y(g20939),.A(g19722),.B(g17632));
  NOR2 NOR2_228(.VSS(VSS),.VDD(VDD),.Y(g20940),.A(g19723),.B(g17633));
  NOR2 NOR2_229(.VSS(VSS),.VDD(VDD),.Y(g20941),.A(g19724),.B(g17634));
  NOR2 NOR2_230(.VSS(VSS),.VDD(VDD),.Y(g20944),.A(g19731),.B(g17652));
  NOR2 NOR2_231(.VSS(VSS),.VDD(VDD),.Y(g20945),.A(g19732),.B(g17653));
  NOR2 NOR2_232(.VSS(VSS),.VDD(VDD),.Y(g20946),.A(g19733),.B(g17654));
  NOR2 NOR2_233(.VSS(VSS),.VDD(VDD),.Y(g20947),.A(g19734),.B(g15335));
  NOR2 NOR2_234(.VSS(VSS),.VDD(VDD),.Y(g20948),.A(g19735),.B(g15336));
  NOR2 NOR2_235(.VSS(VSS),.VDD(VDD),.Y(g20949),.A(g19741),.B(g17673));
  NOR2 NOR2_236(.VSS(VSS),.VDD(VDD),.Y(g20950),.A(g19742),.B(g17674));
  NOR2 NOR2_237(.VSS(VSS),.VDD(VDD),.Y(g20951),.A(g19743),.B(g17675));
  NOR2 NOR2_238(.VSS(VSS),.VDD(VDD),.Y(g20952),.A(g19744),.B(g15349));
  NOR2 NOR2_239(.VSS(VSS),.VDD(VDD),.Y(g20953),.A(g19752),.B(g17695));
  NOR2 NOR2_240(.VSS(VSS),.VDD(VDD),.Y(g20954),.A(g19753),.B(g17696));
  NOR2 NOR2_241(.VSS(VSS),.VDD(VDD),.Y(g20955),.A(g19754),.B(g17697));
  NOR2 NOR2_242(.VSS(VSS),.VDD(VDD),.Y(g20962),.A(g19758),.B(g17714));
  NOR2 NOR2_243(.VSS(VSS),.VDD(VDD),.Y(g20963),.A(g19759),.B(g17715));
  NOR2 NOR2_244(.VSS(VSS),.VDD(VDD),.Y(g20964),.A(g19760),.B(g17716));
  NOR2 NOR2_245(.VSS(VSS),.VDD(VDD),.Y(g20965),.A(g19761),.B(g17717));
  NOR2 NOR2_246(.VSS(VSS),.VDD(VDD),.Y(g20966),.A(g19765),.B(g17734));
  NOR2 NOR2_247(.VSS(VSS),.VDD(VDD),.Y(g20967),.A(g19766),.B(g17735));
  NOR2 NOR2_248(.VSS(VSS),.VDD(VDD),.Y(g20968),.A(g19767),.B(g17736));
  NOR2 NOR2_249(.VSS(VSS),.VDD(VDD),.Y(g20969),.A(g19768),.B(g15402));
  NOR2 NOR2_250(.VSS(VSS),.VDD(VDD),.Y(g20970),.A(g19769),.B(g15403));
  NOR2 NOR2_251(.VSS(VSS),.VDD(VDD),.Y(g20972),.A(g19774),.B(g17752));
  NOR2 NOR2_252(.VSS(VSS),.VDD(VDD),.Y(g20973),.A(g19775),.B(g17753));
  NOR2 NOR2_253(.VSS(VSS),.VDD(VDD),.Y(g20974),.A(g19776),.B(g17754));
  NOR2 NOR2_254(.VSS(VSS),.VDD(VDD),.Y(g20975),.A(g19777),.B(g15421));
  NOR2 NOR2_255(.VSS(VSS),.VDD(VDD),.Y(g20976),.A(g19778),.B(g15422));
  NOR2 NOR2_256(.VSS(VSS),.VDD(VDD),.Y(g20977),.A(g19784),.B(g17773));
  NOR2 NOR2_257(.VSS(VSS),.VDD(VDD),.Y(g20978),.A(g19785),.B(g17774));
  NOR2 NOR2_258(.VSS(VSS),.VDD(VDD),.Y(g20979),.A(g19786),.B(g17775));
  NOR2 NOR2_259(.VSS(VSS),.VDD(VDD),.Y(g20980),.A(g19787),.B(g15435));
  NOR2 NOR2_260(.VSS(VSS),.VDD(VDD),.Y(g20981),.A(g19795),.B(g17795));
  NOR2 NOR2_261(.VSS(VSS),.VDD(VDD),.Y(g20982),.A(g19796),.B(g17796));
  NOR2 NOR2_262(.VSS(VSS),.VDD(VDD),.Y(g20983),.A(g19797),.B(g17797));
  NOR2 NOR2_263(.VSS(VSS),.VDD(VDD),.Y(g20989),.A(g19802),.B(g17812));
  NOR2 NOR2_264(.VSS(VSS),.VDD(VDD),.Y(g20990),.A(g19803),.B(g17813));
  NOR2 NOR2_265(.VSS(VSS),.VDD(VDD),.Y(g20991),.A(g19804),.B(g17814));
  NOR2 NOR2_266(.VSS(VSS),.VDD(VDD),.Y(g20992),.A(g19805),.B(g15470));
  NOR2 NOR2_267(.VSS(VSS),.VDD(VDD),.Y(g20993),.A(g19807),.B(g17835));
  NOR2 NOR2_268(.VSS(VSS),.VDD(VDD),.Y(g20994),.A(g19808),.B(g17836));
  NOR2 NOR2_269(.VSS(VSS),.VDD(VDD),.Y(g20995),.A(g19809),.B(g17837));
  NOR2 NOR2_270(.VSS(VSS),.VDD(VDD),.Y(g20996),.A(g19810),.B(g15486));
  NOR2 NOR2_271(.VSS(VSS),.VDD(VDD),.Y(g20997),.A(g19811),.B(g15487));
  NOR2 NOR2_272(.VSS(VSS),.VDD(VDD),.Y(g20999),.A(g19816),.B(g17853));
  NOR2 NOR2_273(.VSS(VSS),.VDD(VDD),.Y(g21000),.A(g19817),.B(g17854));
  NOR2 NOR2_274(.VSS(VSS),.VDD(VDD),.Y(g21001),.A(g19818),.B(g17855));
  NOR2 NOR2_275(.VSS(VSS),.VDD(VDD),.Y(g21002),.A(g19819),.B(g15505));
  NOR2 NOR2_276(.VSS(VSS),.VDD(VDD),.Y(g21003),.A(g19820),.B(g15506));
  NOR2 NOR2_277(.VSS(VSS),.VDD(VDD),.Y(g21004),.A(g19826),.B(g17874));
  NOR2 NOR2_278(.VSS(VSS),.VDD(VDD),.Y(g21005),.A(g19827),.B(g17875));
  NOR2 NOR2_279(.VSS(VSS),.VDD(VDD),.Y(g21006),.A(g19828),.B(g17876));
  NOR2 NOR2_280(.VSS(VSS),.VDD(VDD),.Y(g21007),.A(g19829),.B(g15519));
  NOR2 NOR2_281(.VSS(VSS),.VDD(VDD),.Y(g21008),.A(g19836),.B(g17877));
  NOR2 NOR2_282(.VSS(VSS),.VDD(VDD),.Y(g21009),.A(g19839),.B(g17900));
  NOR2 NOR2_283(.VSS(VSS),.VDD(VDD),.Y(g21010),.A(g19840),.B(g17901));
  NOR2 NOR2_284(.VSS(VSS),.VDD(VDD),.Y(g21011),.A(g19841),.B(g17902));
  NOR2 NOR2_285(.VSS(VSS),.VDD(VDD),.Y(g21015),.A(g19846),.B(g17924));
  NOR2 NOR2_286(.VSS(VSS),.VDD(VDD),.Y(g21016),.A(g19847),.B(g17925));
  NOR2 NOR2_287(.VSS(VSS),.VDD(VDD),.Y(g21017),.A(g19848),.B(g17926));
  NOR2 NOR2_288(.VSS(VSS),.VDD(VDD),.Y(g21018),.A(g19849),.B(g15556));
  NOR2 NOR2_289(.VSS(VSS),.VDD(VDD),.Y(g21019),.A(g19851),.B(g17947));
  NOR2 NOR2_290(.VSS(VSS),.VDD(VDD),.Y(g21020),.A(g19852),.B(g17948));
  NOR2 NOR2_291(.VSS(VSS),.VDD(VDD),.Y(g21021),.A(g19853),.B(g17949));
  NOR2 NOR2_292(.VSS(VSS),.VDD(VDD),.Y(g21022),.A(g19854),.B(g15572));
  NOR2 NOR2_293(.VSS(VSS),.VDD(VDD),.Y(g21023),.A(g19855),.B(g15573));
  NOR2 NOR2_294(.VSS(VSS),.VDD(VDD),.Y(g21025),.A(g19860),.B(g17965));
  NOR2 NOR2_295(.VSS(VSS),.VDD(VDD),.Y(g21026),.A(g19861),.B(g17966));
  NOR2 NOR2_296(.VSS(VSS),.VDD(VDD),.Y(g21027),.A(g19862),.B(g17967));
  NOR2 NOR2_297(.VSS(VSS),.VDD(VDD),.Y(g21028),.A(g19863),.B(g15591));
  NOR2 NOR2_298(.VSS(VSS),.VDD(VDD),.Y(g21029),.A(g19864),.B(g15592));
  NOR2 NOR2_299(.VSS(VSS),.VDD(VDD),.Y(g21031),.A(g19869),.B(g17989));
  NOR2 NOR2_300(.VSS(VSS),.VDD(VDD),.Y(g21032),.A(g19870),.B(g17990));
  NOR2 NOR2_301(.VSS(VSS),.VDD(VDD),.Y(g21033),.A(g19872),.B(g18011));
  NOR2 NOR2_302(.VSS(VSS),.VDD(VDD),.Y(g21034),.A(g19873),.B(g18012));
  NOR2 NOR2_303(.VSS(VSS),.VDD(VDD),.Y(g21035),.A(g19874),.B(g18013));
  NOR2 NOR2_304(.VSS(VSS),.VDD(VDD),.Y(g21039),.A(g19879),.B(g18035));
  NOR2 NOR2_305(.VSS(VSS),.VDD(VDD),.Y(g21040),.A(g19880),.B(g18036));
  NOR2 NOR2_306(.VSS(VSS),.VDD(VDD),.Y(g21041),.A(g19881),.B(g18037));
  NOR2 NOR2_307(.VSS(VSS),.VDD(VDD),.Y(g21042),.A(g19882),.B(g15634));
  NOR2 NOR2_308(.VSS(VSS),.VDD(VDD),.Y(g21043),.A(g19884),.B(g18058));
  NOR2 NOR2_309(.VSS(VSS),.VDD(VDD),.Y(g21044),.A(g19885),.B(g18059));
  NOR2 NOR2_310(.VSS(VSS),.VDD(VDD),.Y(g21045),.A(g19886),.B(g18060));
  NOR2 NOR2_311(.VSS(VSS),.VDD(VDD),.Y(g21046),.A(g19887),.B(g15650));
  NOR2 NOR2_312(.VSS(VSS),.VDD(VDD),.Y(g21047),.A(g19888),.B(g15651));
  NOR2 NOR2_313(.VSS(VSS),.VDD(VDD),.Y(g21048),.A(g19889),.B(g18062));
  NOR2 NOR2_314(.VSS(VSS),.VDD(VDD),.Y(g21051),.A(g19895),.B(g18088));
  NOR2 NOR2_315(.VSS(VSS),.VDD(VDD),.Y(g21052),.A(g19900),.B(g18106));
  NOR2 NOR2_316(.VSS(VSS),.VDD(VDD),.Y(g21053),.A(g19901),.B(g18107));
  NOR2 NOR2_317(.VSS(VSS),.VDD(VDD),.Y(g21054),.A(g19903),.B(g18128));
  NOR2 NOR2_318(.VSS(VSS),.VDD(VDD),.Y(g21055),.A(g19904),.B(g18129));
  NOR2 NOR2_319(.VSS(VSS),.VDD(VDD),.Y(g21056),.A(g19905),.B(g18130));
  NOR2 NOR2_320(.VSS(VSS),.VDD(VDD),.Y(g21060),.A(g19910),.B(g18152));
  NOR2 NOR2_321(.VSS(VSS),.VDD(VDD),.Y(g21061),.A(g19911),.B(g18153));
  NOR2 NOR2_322(.VSS(VSS),.VDD(VDD),.Y(g21062),.A(g19912),.B(g18154));
  NOR2 NOR2_323(.VSS(VSS),.VDD(VDD),.Y(g21063),.A(g19913),.B(g15710));
  NOR2 NOR2_324(.VSS(VSS),.VDD(VDD),.Y(g21065),.A(g19914),.B(g18169));
  NOR2 NOR2_325(.VSS(VSS),.VDD(VDD),.Y(g21070),.A(g19920),.B(g18204));
  NOR2 NOR2_326(.VSS(VSS),.VDD(VDD),.Y(g21071),.A(g19925),.B(g18222));
  NOR2 NOR2_327(.VSS(VSS),.VDD(VDD),.Y(g21072),.A(g19926),.B(g18223));
  NOR2 NOR2_328(.VSS(VSS),.VDD(VDD),.Y(g21073),.A(g19928),.B(g18244));
  NOR2 NOR2_329(.VSS(VSS),.VDD(VDD),.Y(g21074),.A(g19929),.B(g18245));
  NOR2 NOR2_330(.VSS(VSS),.VDD(VDD),.Y(g21075),.A(g19930),.B(g18246));
  NOR2 NOR2_331(.VSS(VSS),.VDD(VDD),.Y(g21080),.A(g19935),.B(g18311));
  NOR2 NOR2_332(.VSS(VSS),.VDD(VDD),.Y(g21081),.A(g19940),.B(g18329));
  NOR2 NOR2_333(.VSS(VSS),.VDD(VDD),.Y(g21082),.A(g19941),.B(g18330));
  NOR2 NOR2_334(.VSS(VSS),.VDD(VDD),.Y(g21083),.A(g19943),.B(g18333));
  NOR2 NOR2_335(.VSS(VSS),.VDD(VDD),.Y(g21084),.A(g20011),.B(g20048));
  NOR2 NOR2_336(.VSS(VSS),.VDD(VDD),.Y(g21094),.A(g19952),.B(g18404));
  NOR3 NOR3_317(.VSS(VSS),.VDD(VDD),.Y(g21095),.A(g20012),.B(g20049),.C(g20084));
  NOR3 NOR3_318(.VSS(VSS),.VDD(VDD),.Y(g21096),.A(g20013),.B(g20051),.C(g20087));
  NOR3 NOR3_319(.VSS(VSS),.VDD(VDD),.Y(g21104),.A(g20050),.B(g20085),.C(g20106));
  NOR3 NOR3_320(.VSS(VSS),.VDD(VDD),.Y(g21105),.A(g20052),.B(g20088),.C(g20109));
  NOR3 NOR3_321(.VSS(VSS),.VDD(VDD),.Y(g21106),.A(g20053),.B(g20090),.C(g20112));
  NOR3 NOR3_322(.VSS(VSS),.VDD(VDD),.Y(g21116),.A(g20086),.B(g20107),.C(g20131));
  NOR3 NOR3_323(.VSS(VSS),.VDD(VDD),.Y(g21117),.A(g20089),.B(g20110),.C(g20133));
  NOR3 NOR3_324(.VSS(VSS),.VDD(VDD),.Y(g21118),.A(g20091),.B(g20113),.C(g20136));
  NOR3 NOR3_325(.VSS(VSS),.VDD(VDD),.Y(g21119),.A(g20092),.B(g20115),.C(g20139));
  NOR3 NOR3_326(.VSS(VSS),.VDD(VDD),.Y(g21133),.A(g20108),.B(g20132),.C(g20156));
  NOR3 NOR3_327(.VSS(VSS),.VDD(VDD),.Y(g21134),.A(g20111),.B(g20134),.C(g20157));
  NOR3 NOR3_328(.VSS(VSS),.VDD(VDD),.Y(g21135),.A(g20114),.B(g20137),.C(g20160));
  NOR3 NOR3_329(.VSS(VSS),.VDD(VDD),.Y(g21147),.A(g20135),.B(g20158),.C(g20188));
  NOR3 NOR3_330(.VSS(VSS),.VDD(VDD),.Y(g21148),.A(g20138),.B(g20161),.C(g20190));
  NOR2 NOR2_337(.VSS(VSS),.VDD(VDD),.Y(g21149),.A(g20015),.B(g19981));
  NOR2 NOR2_338(.VSS(VSS),.VDD(VDD),.Y(g21167),.A(g20159),.B(g20189));
  NOR3 NOR3_331(.VSS(VSS),.VDD(VDD),.Y(g21168),.A(g20162),.B(g20191),.C(g20220));
  NOR2 NOR2_339(.VSS(VSS),.VDD(VDD),.Y(g21169),.A(g20057),.B(g20019));
  NOR2 NOR2_340(.VSS(VSS),.VDD(VDD),.Y(g21183),.A(g20192),.B(g20221));
  NOR2 NOR2_341(.VSS(VSS),.VDD(VDD),.Y(g21189),.A(g20098),.B(g20061));
  NOR2 NOR2_342(.VSS(VSS),.VDD(VDD),.Y(g21204),.A(g20123),.B(g20102));
  NOR2 NOR2_343(.VSS(VSS),.VDD(VDD),.Y(g21211),.A(g19240),.B(g19230));
  NOR2 NOR2_344(.VSS(VSS),.VDD(VDD),.Y(g21219),.A(g19253),.B(g19243));
  NOR3 NOR3_332(.VSS(VSS),.VDD(VDD),.Y(g21227),.A(g18414),.B(g18485),.C(g20295));
  NOR2 NOR2_345(.VSS(VSS),.VDD(VDD),.Y(g21228),.A(g19388),.B(g17118));
  NOR2 NOR2_346(.VSS(VSS),.VDD(VDD),.Y(g21230),.A(g19266),.B(g19256));
  NOR2 NOR2_347(.VSS(VSS),.VDD(VDD),.Y(g21233),.A(g19418),.B(g17145));
  NOR2 NOR2_348(.VSS(VSS),.VDD(VDD),.Y(g21235),.A(g19281),.B(g19269));
  NOR2 NOR2_349(.VSS(VSS),.VDD(VDD),.Y(g21238),.A(g19954),.B(g5890));
  NOR2 NOR2_350(.VSS(VSS),.VDD(VDD),.Y(g21242),.A(g19455),.B(g17168));
  NOR2 NOR2_351(.VSS(VSS),.VDD(VDD),.Y(g21246),.A(g19984),.B(g5929));
  NOR2 NOR2_352(.VSS(VSS),.VDD(VDD),.Y(g21250),.A(g19482),.B(g17183));
  NOR2 NOR2_353(.VSS(VSS),.VDD(VDD),.Y(g21255),.A(g20022),.B(g5963));
  NOR2 NOR2_354(.VSS(VSS),.VDD(VDD),.Y(g21263),.A(g20064),.B(g5992));
  NOR2 NOR2_355(.VSS(VSS),.VDD(VDD),.Y(g21316),.A(g20460),.B(g16111));
  NOR2 NOR2_356(.VSS(VSS),.VDD(VDD),.Y(g21331),.A(g20472),.B(g16153));
  NOR2 NOR2_357(.VSS(VSS),.VDD(VDD),.Y(g21346),.A(g20480),.B(g13247));
  NOR2 NOR2_358(.VSS(VSS),.VDD(VDD),.Y(g21364),.A(g20486),.B(g13266));
  NOR2 NOR2_359(.VSS(VSS),.VDD(VDD),.Y(g21385),.A(g20492),.B(g13289));
  NOR2 NOR2_360(.VSS(VSS),.VDD(VDD),.Y(g21407),.A(g20499),.B(g13316));
  NOR2 NOR2_361(.VSS(VSS),.VDD(VDD),.Y(g21432),.A(g20502),.B(g13335));
  NOR2 NOR2_362(.VSS(VSS),.VDD(VDD),.Y(g21435),.A(g20503),.B(g16385));
  NOR2 NOR2_363(.VSS(VSS),.VDD(VDD),.Y(g21467),.A(g20506),.B(g13355));
  NOR2 NOR2_364(.VSS(VSS),.VDD(VDD),.Y(g21470),.A(g20512),.B(g16417));
  NOR2 NOR2_365(.VSS(VSS),.VDD(VDD),.Y(g21502),.A(g20525),.B(g16445));
  NOR2 NOR2_366(.VSS(VSS),.VDD(VDD),.Y(g21615),.A(g16567),.B(g19957));
  NOR3 NOR3_333(.VSS(VSS),.VDD(VDD),.Y(g21618),.A(g20016),.B(g14079),.C(g14165));
  NOR2 NOR2_367(.VSS(VSS),.VDD(VDD),.Y(g21636),.A(g20473),.B(g6513));
  NOR2 NOR2_368(.VSS(VSS),.VDD(VDD),.Y(g21643),.A(g16591),.B(g19987));
  NOR3 NOR3_334(.VSS(VSS),.VDD(VDD),.Y(g21646),.A(g20058),.B(g14194),.C(g14280));
  NOR2 NOR2_369(.VSS(VSS),.VDD(VDD),.Y(g21665),.A(g20507),.B(g18352));
  NOR2 NOR2_370(.VSS(VSS),.VDD(VDD),.Y(g21667),.A(g20481),.B(g6777));
  NOR2 NOR2_371(.VSS(VSS),.VDD(VDD),.Y(g21674),.A(g16611),.B(g20025));
  NOR3 NOR3_335(.VSS(VSS),.VDD(VDD),.Y(g21677),.A(g20099),.B(g14309),.C(g14402));
  NOR2 NOR2_372(.VSS(VSS),.VDD(VDD),.Y(g21694),.A(g20526),.B(g18447));
  NOR2 NOR2_373(.VSS(VSS),.VDD(VDD),.Y(g21696),.A(g20487),.B(g7079));
  NOR2 NOR2_374(.VSS(VSS),.VDD(VDD),.Y(g21703),.A(g16629),.B(g20067));
  NOR3 NOR3_336(.VSS(VSS),.VDD(VDD),.Y(g21706),.A(g20124),.B(g14431),.C(g14514));
  NOR2 NOR2_375(.VSS(VSS),.VDD(VDD),.Y(g21711),.A(g19830),.B(g15780));
  NOR2 NOR2_376(.VSS(VSS),.VDD(VDD),.Y(g21730),.A(g20545),.B(g18520));
  NOR2 NOR2_377(.VSS(VSS),.VDD(VDD),.Y(g21732),.A(g20493),.B(g7329));
  NOR3 NOR3_337(.VSS(VSS),.VDD(VDD),.Y(g21738),.A(g19444),.B(g17893),.C(g14079));
  NOR2 NOR2_378(.VSS(VSS),.VDD(VDD),.Y(g21739),.A(g20507),.B(g18430));
  NOR2 NOR2_379(.VSS(VSS),.VDD(VDD),.Y(g21756),.A(g19070),.B(g18584));
  NOR3 NOR3_338(.VSS(VSS),.VDD(VDD),.Y(g21762),.A(g19471),.B(g18004),.C(g14194));
  NOR2 NOR2_380(.VSS(VSS),.VDD(VDD),.Y(g21763),.A(g20526),.B(g18503));
  NOR3 NOR3_339(.VSS(VSS),.VDD(VDD),.Y(g21778),.A(g19494),.B(g18121),.C(g14309));
  NOR2 NOR2_381(.VSS(VSS),.VDD(VDD),.Y(g21779),.A(g20545),.B(g18567));
  NOR3 NOR3_340(.VSS(VSS),.VDD(VDD),.Y(g21793),.A(g19515),.B(g18237),.C(g14431));
  NOR2 NOR2_382(.VSS(VSS),.VDD(VDD),.Y(g21794),.A(g19070),.B(g18617));
  NOR2 NOR2_383(.VSS(VSS),.VDD(VDD),.Y(g21796),.A(g19830),.B(g13004));
  NOR2 NOR2_384(.VSS(VSS),.VDD(VDD),.Y(g21842),.A(g13609),.B(g19150));
  NOR2 NOR2_385(.VSS(VSS),.VDD(VDD),.Y(g21843),.A(g13619),.B(g19155));
  NOR2 NOR2_386(.VSS(VSS),.VDD(VDD),.Y(g21845),.A(g13631),.B(g19161));
  NOR2 NOR2_387(.VSS(VSS),.VDD(VDD),.Y(g21847),.A(g13642),.B(g19166));
  NOR2 NOR2_388(.VSS(VSS),.VDD(VDD),.Y(g21851),.A(g19252),.B(g8842));
  NOR2 NOR2_389(.VSS(VSS),.VDD(VDD),.Y(g21878),.A(g16964),.B(g19228));
  NOR2 NOR2_390(.VSS(VSS),.VDD(VDD),.Y(g21880),.A(g13854),.B(g19236));
  NOR2 NOR2_391(.VSS(VSS),.VDD(VDD),.Y(g21882),.A(g13862),.B(g19248));
  NOR2 NOR2_392(.VSS(VSS),.VDD(VDD),.Y(g21884),.A(g19260),.B(g19284));
  NOR2 NOR2_393(.VSS(VSS),.VDD(VDD),.Y(g21887),.A(g13519),.B(g19289));
  NOR2 NOR2_394(.VSS(VSS),.VDD(VDD),.Y(g21889),.A(g19285),.B(g19316));
  NOR2 NOR2_395(.VSS(VSS),.VDD(VDD),.Y(g21890),.A(g13530),.B(g19307));
  NOR2 NOR2_396(.VSS(VSS),.VDD(VDD),.Y(g21893),.A(g13541),.B(g19328));
  NOR2 NOR2_397(.VSS(VSS),.VDD(VDD),.Y(g21894),.A(g19317),.B(g19356));
  NOR2 NOR2_398(.VSS(VSS),.VDD(VDD),.Y(g21901),.A(g13552),.B(g19355));
  NOR2 NOR2_399(.VSS(VSS),.VDD(VDD),.Y(g21968),.A(g21234),.B(g19476));
  NOR2 NOR2_400(.VSS(VSS),.VDD(VDD),.Y(g21969),.A(g20895),.B(g10133));
  NOR2 NOR2_401(.VSS(VSS),.VDD(VDD),.Y(g21970),.A(g17182),.B(g21226));
  NOR2 NOR2_402(.VSS(VSS),.VDD(VDD),.Y(g21971),.A(g21243),.B(g19499));
  NOR2 NOR2_403(.VSS(VSS),.VDD(VDD),.Y(g21972),.A(g20914),.B(g10238));
  NOR2 NOR2_404(.VSS(VSS),.VDD(VDD),.Y(g21973),.A(g21251),.B(g19520));
  NOR2 NOR2_405(.VSS(VSS),.VDD(VDD),.Y(g21974),.A(g20938),.B(g10340));
  NOR2 NOR2_406(.VSS(VSS),.VDD(VDD),.Y(g21975),.A(g21245),.B(g21259));
  NOR3 NOR3_341(.VSS(VSS),.VDD(VDD),.Y(g21980),.A(g21252),.B(g19531),.C(g19540));
  NOR2 NOR2_407(.VSS(VSS),.VDD(VDD),.Y(g21981),.A(g21254),.B(g21267));
  NOR3 NOR3_342(.VSS(VSS),.VDD(VDD),.Y(g21987),.A(g21260),.B(g19541),.C(g19544));
  NOR2 NOR2_408(.VSS(VSS),.VDD(VDD),.Y(g21988),.A(g21262),.B(g21276));
  NOR3 NOR3_343(.VSS(VSS),.VDD(VDD),.Y(g22000),.A(g21268),.B(g19545),.C(g19547));
  NOR2 NOR2_409(.VSS(VSS),.VDD(VDD),.Y(g22001),.A(g21270),.B(g21283));
  NOR3 NOR3_344(.VSS(VSS),.VDD(VDD),.Y(g22013),.A(g21277),.B(g19548),.C(g19551));
  NOR2 NOR2_410(.VSS(VSS),.VDD(VDD),.Y(g22025),.A(g21284),.B(g19549));
  NOR2 NOR2_411(.VSS(VSS),.VDD(VDD),.Y(g22026),.A(g21083),.B(g18407));
  NOR2 NOR2_412(.VSS(VSS),.VDD(VDD),.Y(g22027),.A(g21290),.B(g19553));
  NOR2 NOR2_413(.VSS(VSS),.VDD(VDD),.Y(g22028),.A(g21291),.B(g19554));
  NOR2 NOR2_414(.VSS(VSS),.VDD(VDD),.Y(g22029),.A(g21292),.B(g19555));
  NOR2 NOR2_415(.VSS(VSS),.VDD(VDD),.Y(g22030),.A(g21298),.B(g19557));
  NOR2 NOR2_416(.VSS(VSS),.VDD(VDD),.Y(g22031),.A(g21299),.B(g19558));
  NOR2 NOR2_417(.VSS(VSS),.VDD(VDD),.Y(g22032),.A(g21300),.B(g19559));
  NOR2 NOR2_418(.VSS(VSS),.VDD(VDD),.Y(g22033),.A(g21301),.B(g19560));
  NOR2 NOR2_419(.VSS(VSS),.VDD(VDD),.Y(g22034),.A(g21302),.B(g19561));
  NOR2 NOR2_420(.VSS(VSS),.VDD(VDD),.Y(g22035),.A(g21303),.B(g19562));
  NOR2 NOR2_421(.VSS(VSS),.VDD(VDD),.Y(g22037),.A(g21304),.B(g19564));
  NOR2 NOR2_422(.VSS(VSS),.VDD(VDD),.Y(g22038),.A(g21305),.B(g19565));
  NOR2 NOR2_423(.VSS(VSS),.VDD(VDD),.Y(g22039),.A(g21306),.B(g19566));
  NOR2 NOR2_424(.VSS(VSS),.VDD(VDD),.Y(g22040),.A(g21307),.B(g19567));
  NOR2 NOR2_425(.VSS(VSS),.VDD(VDD),.Y(g22041),.A(g21308),.B(g19568));
  NOR2 NOR2_426(.VSS(VSS),.VDD(VDD),.Y(g22042),.A(g21309),.B(g19569));
  NOR2 NOR2_427(.VSS(VSS),.VDD(VDD),.Y(g22043),.A(g21310),.B(g19570));
  NOR2 NOR2_428(.VSS(VSS),.VDD(VDD),.Y(g22044),.A(g21311),.B(g19571));
  NOR2 NOR2_429(.VSS(VSS),.VDD(VDD),.Y(g22045),.A(g21312),.B(g19572));
  NOR2 NOR2_430(.VSS(VSS),.VDD(VDD),.Y(g22047),.A(g21313),.B(g19574));
  NOR2 NOR2_431(.VSS(VSS),.VDD(VDD),.Y(g22048),.A(g21314),.B(g19575));
  NOR2 NOR2_432(.VSS(VSS),.VDD(VDD),.Y(g22049),.A(g21315),.B(g19576));
  NOR2 NOR2_433(.VSS(VSS),.VDD(VDD),.Y(g22054),.A(g21319),.B(g19586));
  NOR2 NOR2_434(.VSS(VSS),.VDD(VDD),.Y(g22055),.A(g21320),.B(g19587));
  NOR2 NOR2_435(.VSS(VSS),.VDD(VDD),.Y(g22056),.A(g21321),.B(g19588));
  NOR2 NOR2_436(.VSS(VSS),.VDD(VDD),.Y(g22057),.A(g21322),.B(g19589));
  NOR2 NOR2_437(.VSS(VSS),.VDD(VDD),.Y(g22058),.A(g21323),.B(g19590));
  NOR2 NOR2_438(.VSS(VSS),.VDD(VDD),.Y(g22059),.A(g21324),.B(g19591));
  NOR2 NOR2_439(.VSS(VSS),.VDD(VDD),.Y(g22060),.A(g21325),.B(g19592));
  NOR2 NOR2_440(.VSS(VSS),.VDD(VDD),.Y(g22061),.A(g21326),.B(g19593));
  NOR2 NOR2_441(.VSS(VSS),.VDD(VDD),.Y(g22063),.A(g21328),.B(g19597));
  NOR2 NOR2_442(.VSS(VSS),.VDD(VDD),.Y(g22064),.A(g21329),.B(g19598));
  NOR2 NOR2_443(.VSS(VSS),.VDD(VDD),.Y(g22065),.A(g21330),.B(g19599));
  NOR2 NOR2_444(.VSS(VSS),.VDD(VDD),.Y(g22066),.A(g21334),.B(g19604));
  NOR2 NOR2_445(.VSS(VSS),.VDD(VDD),.Y(g22067),.A(g21335),.B(g19605));
  NOR2 NOR2_446(.VSS(VSS),.VDD(VDD),.Y(g22068),.A(g21336),.B(g19606));
  NOR2 NOR2_447(.VSS(VSS),.VDD(VDD),.Y(g22073),.A(g21337),.B(g19616));
  NOR2 NOR2_448(.VSS(VSS),.VDD(VDD),.Y(g22074),.A(g21338),.B(g19617));
  NOR2 NOR2_449(.VSS(VSS),.VDD(VDD),.Y(g22075),.A(g21339),.B(g19618));
  NOR2 NOR2_450(.VSS(VSS),.VDD(VDD),.Y(g22076),.A(g21340),.B(g19619));
  NOR2 NOR2_451(.VSS(VSS),.VDD(VDD),.Y(g22077),.A(g21341),.B(g19620));
  NOR2 NOR2_452(.VSS(VSS),.VDD(VDD),.Y(g22078),.A(g21342),.B(g19621));
  NOR2 NOR2_453(.VSS(VSS),.VDD(VDD),.Y(g22079),.A(g21343),.B(g19623));
  NOR2 NOR2_454(.VSS(VSS),.VDD(VDD),.Y(g22080),.A(g21344),.B(g19624));
  NOR2 NOR2_455(.VSS(VSS),.VDD(VDD),.Y(g22081),.A(g21345),.B(g19625));
  NOR2 NOR2_456(.VSS(VSS),.VDD(VDD),.Y(g22087),.A(g21349),.B(g19630));
  NOR2 NOR2_457(.VSS(VSS),.VDD(VDD),.Y(g22088),.A(g21350),.B(g19631));
  NOR2 NOR2_458(.VSS(VSS),.VDD(VDD),.Y(g22089),.A(g21351),.B(g19632));
  NOR2 NOR2_459(.VSS(VSS),.VDD(VDD),.Y(g22090),.A(g21352),.B(g19637));
  NOR2 NOR2_460(.VSS(VSS),.VDD(VDD),.Y(g22091),.A(g21353),.B(g19638));
  NOR2 NOR2_461(.VSS(VSS),.VDD(VDD),.Y(g22092),.A(g21354),.B(g19639));
  NOR2 NOR2_462(.VSS(VSS),.VDD(VDD),.Y(g22097),.A(g21355),.B(g19649));
  NOR2 NOR2_463(.VSS(VSS),.VDD(VDD),.Y(g22098),.A(g21356),.B(g19650));
  NOR2 NOR2_464(.VSS(VSS),.VDD(VDD),.Y(g22099),.A(g21357),.B(g19651));
  NOR2 NOR2_465(.VSS(VSS),.VDD(VDD),.Y(g22100),.A(g21360),.B(g19653));
  NOR2 NOR2_466(.VSS(VSS),.VDD(VDD),.Y(g22101),.A(g21361),.B(g19654));
  NOR2 NOR2_467(.VSS(VSS),.VDD(VDD),.Y(g22102),.A(g21362),.B(g19655));
  NOR2 NOR2_468(.VSS(VSS),.VDD(VDD),.Y(g22103),.A(g21363),.B(g19656));
  NOR2 NOR2_469(.VSS(VSS),.VDD(VDD),.Y(g22104),.A(g21367),.B(g19663));
  NOR2 NOR2_470(.VSS(VSS),.VDD(VDD),.Y(g22105),.A(g21368),.B(g19664));
  NOR2 NOR2_471(.VSS(VSS),.VDD(VDD),.Y(g22106),.A(g21369),.B(g19665));
  NOR2 NOR2_472(.VSS(VSS),.VDD(VDD),.Y(g22112),.A(g21370),.B(g19670));
  NOR2 NOR2_473(.VSS(VSS),.VDD(VDD),.Y(g22113),.A(g21371),.B(g19671));
  NOR2 NOR2_474(.VSS(VSS),.VDD(VDD),.Y(g22114),.A(g21372),.B(g19672));
  NOR2 NOR2_475(.VSS(VSS),.VDD(VDD),.Y(g22115),.A(g21373),.B(g19677));
  NOR2 NOR2_476(.VSS(VSS),.VDD(VDD),.Y(g22116),.A(g21374),.B(g19678));
  NOR2 NOR2_477(.VSS(VSS),.VDD(VDD),.Y(g22117),.A(g21375),.B(g19679));
  NOR2 NOR2_478(.VSS(VSS),.VDD(VDD),.Y(g22122),.A(g21378),.B(g19692));
  NOR2 NOR2_479(.VSS(VSS),.VDD(VDD),.Y(g22123),.A(g21379),.B(g19693));
  NOR2 NOR2_480(.VSS(VSS),.VDD(VDD),.Y(g22124),.A(g21380),.B(g19694));
  NOR2 NOR2_481(.VSS(VSS),.VDD(VDD),.Y(g22125),.A(g21381),.B(g19695));
  NOR2 NOR2_482(.VSS(VSS),.VDD(VDD),.Y(g22126),.A(g21389),.B(g19701));
  NOR2 NOR2_483(.VSS(VSS),.VDD(VDD),.Y(g22127),.A(g21390),.B(g19702));
  NOR2 NOR2_484(.VSS(VSS),.VDD(VDD),.Y(g22128),.A(g21391),.B(g19703));
  NOR2 NOR2_485(.VSS(VSS),.VDD(VDD),.Y(g22129),.A(g21392),.B(g19704));
  NOR2 NOR2_486(.VSS(VSS),.VDD(VDD),.Y(g22130),.A(g21393),.B(g19711));
  NOR2 NOR2_487(.VSS(VSS),.VDD(VDD),.Y(g22131),.A(g21394),.B(g19712));
  NOR2 NOR2_488(.VSS(VSS),.VDD(VDD),.Y(g22132),.A(g21395),.B(g19713));
  NOR2 NOR2_489(.VSS(VSS),.VDD(VDD),.Y(g22138),.A(g21396),.B(g19718));
  NOR2 NOR2_490(.VSS(VSS),.VDD(VDD),.Y(g22139),.A(g21397),.B(g19719));
  NOR2 NOR2_491(.VSS(VSS),.VDD(VDD),.Y(g22140),.A(g21398),.B(g19720));
  NOR2 NOR2_492(.VSS(VSS),.VDD(VDD),.Y(g22141),.A(g21401),.B(g19727));
  NOR2 NOR2_493(.VSS(VSS),.VDD(VDD),.Y(g22142),.A(g21402),.B(g19728));
  NOR2 NOR2_494(.VSS(VSS),.VDD(VDD),.Y(g22143),.A(g21403),.B(g19729));
  NOR2 NOR2_495(.VSS(VSS),.VDD(VDD),.Y(g22144),.A(g21410),.B(g19730));
  NOR2 NOR2_496(.VSS(VSS),.VDD(VDD),.Y(g22145),.A(g21411),.B(g19736));
  NOR2 NOR2_497(.VSS(VSS),.VDD(VDD),.Y(g22146),.A(g21412),.B(g19737));
  NOR2 NOR2_498(.VSS(VSS),.VDD(VDD),.Y(g22147),.A(g21413),.B(g19738));
  NOR2 NOR2_499(.VSS(VSS),.VDD(VDD),.Y(g22148),.A(g21414),.B(g19739));
  NOR2 NOR2_500(.VSS(VSS),.VDD(VDD),.Y(g22149),.A(g21419),.B(g19745));
  NOR2 NOR2_501(.VSS(VSS),.VDD(VDD),.Y(g22150),.A(g21420),.B(g19746));
  NOR2 NOR2_502(.VSS(VSS),.VDD(VDD),.Y(g22151),.A(g21421),.B(g19747));
  NOR2 NOR2_503(.VSS(VSS),.VDD(VDD),.Y(g22152),.A(g21422),.B(g19748));
  NOR2 NOR2_504(.VSS(VSS),.VDD(VDD),.Y(g22153),.A(g21423),.B(g19755));
  NOR2 NOR2_505(.VSS(VSS),.VDD(VDD),.Y(g22154),.A(g21424),.B(g19756));
  NOR2 NOR2_506(.VSS(VSS),.VDD(VDD),.Y(g22155),.A(g21425),.B(g19757));
  NOR2 NOR2_507(.VSS(VSS),.VDD(VDD),.Y(g22161),.A(g21428),.B(g19764));
  NOR2 NOR2_508(.VSS(VSS),.VDD(VDD),.Y(g22162),.A(g21438),.B(g19770));
  NOR2 NOR2_509(.VSS(VSS),.VDD(VDD),.Y(g22163),.A(g21439),.B(g19771));
  NOR2 NOR2_510(.VSS(VSS),.VDD(VDD),.Y(g22164),.A(g21440),.B(g19772));
  NOR2 NOR2_511(.VSS(VSS),.VDD(VDD),.Y(g22165),.A(g21444),.B(g19773));
  NOR2 NOR2_512(.VSS(VSS),.VDD(VDD),.Y(g22166),.A(g21445),.B(g19779));
  NOR2 NOR2_513(.VSS(VSS),.VDD(VDD),.Y(g22167),.A(g21446),.B(g19780));
  NOR2 NOR2_514(.VSS(VSS),.VDD(VDD),.Y(g22168),.A(g21447),.B(g19781));
  NOR2 NOR2_515(.VSS(VSS),.VDD(VDD),.Y(g22169),.A(g21448),.B(g19782));
  NOR2 NOR2_516(.VSS(VSS),.VDD(VDD),.Y(g22170),.A(g21453),.B(g19788));
  NOR2 NOR2_517(.VSS(VSS),.VDD(VDD),.Y(g22171),.A(g21454),.B(g19789));
  NOR2 NOR2_518(.VSS(VSS),.VDD(VDD),.Y(g22172),.A(g21455),.B(g19790));
  NOR2 NOR2_519(.VSS(VSS),.VDD(VDD),.Y(g22173),.A(g21456),.B(g19791));
  NOR2 NOR2_520(.VSS(VSS),.VDD(VDD),.Y(g22174),.A(g19868),.B(g21593));
  NOR2 NOR2_521(.VSS(VSS),.VDD(VDD),.Y(g22177),.A(g21476),.B(g19806));
  NOR2 NOR2_522(.VSS(VSS),.VDD(VDD),.Y(g22178),.A(g21480),.B(g19812));
  NOR2 NOR2_523(.VSS(VSS),.VDD(VDD),.Y(g22179),.A(g21481),.B(g19813));
  NOR2 NOR2_524(.VSS(VSS),.VDD(VDD),.Y(g22180),.A(g21482),.B(g19814));
  NOR2 NOR2_525(.VSS(VSS),.VDD(VDD),.Y(g22181),.A(g21486),.B(g19815));
  NOR2 NOR2_526(.VSS(VSS),.VDD(VDD),.Y(g22182),.A(g21487),.B(g19821));
  NOR2 NOR2_527(.VSS(VSS),.VDD(VDD),.Y(g22183),.A(g21488),.B(g19822));
  NOR2 NOR2_528(.VSS(VSS),.VDD(VDD),.Y(g22184),.A(g21489),.B(g19823));
  NOR2 NOR2_529(.VSS(VSS),.VDD(VDD),.Y(g22185),.A(g21490),.B(g19824));
  NOR2 NOR2_530(.VSS(VSS),.VDD(VDD),.Y(g22186),.A(g21497),.B(g19837));
  NOR2 NOR2_531(.VSS(VSS),.VDD(VDD),.Y(g22189),.A(g19899),.B(g21622));
  NOR2 NOR2_532(.VSS(VSS),.VDD(VDD),.Y(g22191),.A(g21517),.B(g19850));
  NOR2 NOR2_533(.VSS(VSS),.VDD(VDD),.Y(g22192),.A(g21521),.B(g19856));
  NOR2 NOR2_534(.VSS(VSS),.VDD(VDD),.Y(g22193),.A(g21522),.B(g19857));
  NOR2 NOR2_535(.VSS(VSS),.VDD(VDD),.Y(g22194),.A(g21523),.B(g19858));
  NOR2 NOR2_536(.VSS(VSS),.VDD(VDD),.Y(g22195),.A(g21527),.B(g19859));
  NOR2 NOR2_537(.VSS(VSS),.VDD(VDD),.Y(g22198),.A(g19924),.B(g21650));
  NOR2 NOR2_538(.VSS(VSS),.VDD(VDD),.Y(g22200),.A(g21553),.B(g19883));
  NOR2 NOR2_539(.VSS(VSS),.VDD(VDD),.Y(g22204),.A(g19939),.B(g21681));
  NOR2 NOR2_540(.VSS(VSS),.VDD(VDD),.Y(g22210),.A(g21610),.B(g19932));
  NOR2 NOR2_541(.VSS(VSS),.VDD(VDD),.Y(g22216),.A(g21635),.B(g19944));
  NOR2 NOR2_542(.VSS(VSS),.VDD(VDD),.Y(g22218),.A(g21639),.B(g19949));
  NOR2 NOR2_543(.VSS(VSS),.VDD(VDD),.Y(g22227),.A(g21658),.B(g19953));
  NOR2 NOR2_544(.VSS(VSS),.VDD(VDD),.Y(g22231),.A(g21666),.B(g19971));
  NOR2 NOR2_545(.VSS(VSS),.VDD(VDD),.Y(g22234),.A(g21670),.B(g19976));
  NOR2 NOR2_546(.VSS(VSS),.VDD(VDD),.Y(g22242),.A(g21687),.B(g19983));
  NOR2 NOR2_547(.VSS(VSS),.VDD(VDD),.Y(g22247),.A(g21695),.B(g20001));
  NOR2 NOR2_548(.VSS(VSS),.VDD(VDD),.Y(g22249),.A(g21699),.B(g20006));
  NOR2 NOR2_549(.VSS(VSS),.VDD(VDD),.Y(g22263),.A(g21723),.B(g20021));
  NOR2 NOR2_550(.VSS(VSS),.VDD(VDD),.Y(g22267),.A(g21731),.B(g20039));
  NOR2 NOR2_551(.VSS(VSS),.VDD(VDD),.Y(g22269),.A(g21735),.B(g20044));
  NOR2 NOR2_552(.VSS(VSS),.VDD(VDD),.Y(g22280),.A(g21749),.B(g20063));
  NOR2 NOR2_553(.VSS(VSS),.VDD(VDD),.Y(g22284),.A(g21757),.B(g20081));
  NOR2 NOR2_554(.VSS(VSS),.VDD(VDD),.Y(g22288),.A(g20144),.B(g21805));
  NOR2 NOR2_555(.VSS(VSS),.VDD(VDD),.Y(g22299),.A(g21773),.B(g20104));
  NOR2 NOR2_556(.VSS(VSS),.VDD(VDD),.Y(g22308),.A(g20182),.B(g21812));
  NOR2 NOR2_557(.VSS(VSS),.VDD(VDD),.Y(g22336),.A(g20216),.B(g21818));
  NOR2 NOR2_558(.VSS(VSS),.VDD(VDD),.Y(g22361),.A(g20246),.B(g21822));
  NOR2 NOR2_559(.VSS(VSS),.VDD(VDD),.Y(g22454),.A(g17012),.B(g21891));
  NOR2 NOR2_560(.VSS(VSS),.VDD(VDD),.Y(g22493),.A(g17042),.B(g21899));
  NOR2 NOR2_561(.VSS(VSS),.VDD(VDD),.Y(g22536),.A(g17076),.B(g21911));
  NOR2 NOR2_562(.VSS(VSS),.VDD(VDD),.Y(g22576),.A(g17111),.B(g21925));
  NOR2 NOR2_563(.VSS(VSS),.VDD(VDD),.Y(g22578),.A(g21892),.B(g18982));
  NOR2 NOR2_564(.VSS(VSS),.VDD(VDD),.Y(g22615),.A(g21900),.B(g18990));
  NOR2 NOR2_565(.VSS(VSS),.VDD(VDD),.Y(g22651),.A(g21912),.B(g18997));
  NOR2 NOR2_566(.VSS(VSS),.VDD(VDD),.Y(g22687),.A(g21926),.B(g19010));
  NOR2 NOR2_567(.VSS(VSS),.VDD(VDD),.Y(g22755),.A(g21271),.B(g20842));
  NOR2 NOR2_568(.VSS(VSS),.VDD(VDD),.Y(g22784),.A(g16075),.B(g20885));
  NOR2 NOR2_569(.VSS(VSS),.VDD(VDD),.Y(g22789),.A(g21278),.B(g20850));
  NOR3 NOR3_345(.VSS(VSS),.VDD(VDD),.Y(g22810),.A(g16075),.B(g20842),.C(g21271));
  NOR2 NOR2_570(.VSS(VSS),.VDD(VDD),.Y(g22826),.A(g16113),.B(g20904));
  NOR2 NOR2_571(.VSS(VSS),.VDD(VDD),.Y(g22831),.A(g21285),.B(g20858));
  NOR3 NOR3_346(.VSS(VSS),.VDD(VDD),.Y(g22851),.A(g16113),.B(g20850),.C(g21278));
  NOR2 NOR2_572(.VSS(VSS),.VDD(VDD),.Y(g22865),.A(g16164),.B(g20928));
  NOR2 NOR2_573(.VSS(VSS),.VDD(VDD),.Y(g22870),.A(g21293),.B(g20866));
  NOR3 NOR3_347(.VSS(VSS),.VDD(VDD),.Y(g22886),.A(g16164),.B(g20858),.C(g21285));
  NOR2 NOR2_574(.VSS(VSS),.VDD(VDD),.Y(g22900),.A(g16223),.B(g20956));
  NOR3 NOR3_348(.VSS(VSS),.VDD(VDD),.Y(g22921),.A(g16223),.B(g20866),.C(g21293));
  NOR2 NOR2_575(.VSS(VSS),.VDD(VDD),.Y(g22935),.A(g21903),.B(g7466));
  NOR2 NOR2_576(.VSS(VSS),.VDD(VDD),.Y(g22953),.A(g20700),.B(g7595));
  NOR2 NOR2_577(.VSS(VSS),.VDD(VDD),.Y(g22985),.A(g21618),.B(g21049));
  NOR2 NOR2_578(.VSS(VSS),.VDD(VDD),.Y(g22987),.A(g21646),.B(g21068));
  NOR2 NOR2_579(.VSS(VSS),.VDD(VDD),.Y(g22990),.A(g21677),.B(g21078));
  NOR2 NOR2_580(.VSS(VSS),.VDD(VDD),.Y(g22997),.A(g21706),.B(g21092));
  NOR2 NOR2_581(.VSS(VSS),.VDD(VDD),.Y(g22999),.A(g21085),.B(g19241));
  NOR2 NOR2_582(.VSS(VSS),.VDD(VDD),.Y(g23000),.A(g16909),.B(g21067));
  NOR2 NOR2_583(.VSS(VSS),.VDD(VDD),.Y(g23009),.A(g21738),.B(g21107));
  NOR2 NOR2_584(.VSS(VSS),.VDD(VDD),.Y(g23013),.A(g21097),.B(g19254));
  NOR2 NOR2_585(.VSS(VSS),.VDD(VDD),.Y(g23014),.A(g16939),.B(g21077));
  NOR2 NOR2_586(.VSS(VSS),.VDD(VDD),.Y(g23022),.A(g16968),.B(g21086));
  NOR3 NOR3_349(.VSS(VSS),.VDD(VDD),.Y(g23023),.A(g14256),.B(g14175),.C(g21123));
  NOR2 NOR2_587(.VSS(VSS),.VDD(VDD),.Y(g23025),.A(g21762),.B(g21124));
  NOR2 NOR2_588(.VSS(VSS),.VDD(VDD),.Y(g23029),.A(g21111),.B(g19267));
  NOR2 NOR2_589(.VSS(VSS),.VDD(VDD),.Y(g23030),.A(g16970),.B(g21091));
  NOR2 NOR2_590(.VSS(VSS),.VDD(VDD),.Y(g23039),.A(g16989),.B(g21098));
  NOR3 NOR3_350(.VSS(VSS),.VDD(VDD),.Y(g23040),.A(g14378),.B(g14290),.C(g21142));
  NOR2 NOR2_591(.VSS(VSS),.VDD(VDD),.Y(g23042),.A(g21778),.B(g21143));
  NOR2 NOR2_592(.VSS(VSS),.VDD(VDD),.Y(g23046),.A(g21128),.B(g19282));
  NOR2 NOR2_593(.VSS(VSS),.VDD(VDD),.Y(g23047),.A(g16991),.B(g21103));
  NOR2 NOR2_594(.VSS(VSS),.VDD(VDD),.Y(g23051),.A(g21121),.B(g21153));
  NOR2 NOR2_595(.VSS(VSS),.VDD(VDD),.Y(g23058),.A(g16999),.B(g21112));
  NOR3 NOR3_351(.VSS(VSS),.VDD(VDD),.Y(g23059),.A(g14490),.B(g14412),.C(g21162));
  NOR2 NOR2_596(.VSS(VSS),.VDD(VDD),.Y(g23061),.A(g21793),.B(g21163));
  NOR3 NOR3_352(.VSS(VSS),.VDD(VDD),.Y(g23066),.A(g21138),.B(g19303),.C(g19320));
  NOR2 NOR2_597(.VSS(VSS),.VDD(VDD),.Y(g23067),.A(g17015),.B(g21122));
  NOR2 NOR2_598(.VSS(VSS),.VDD(VDD),.Y(g23070),.A(g21140),.B(g21173));
  NOR2 NOR2_599(.VSS(VSS),.VDD(VDD),.Y(g23076),.A(g17023),.B(g21129));
  NOR3 NOR3_353(.VSS(VSS),.VDD(VDD),.Y(g23077),.A(g14577),.B(g14524),.C(g21182));
  NOR3 NOR3_354(.VSS(VSS),.VDD(VDD),.Y(g23080),.A(g21158),.B(g19324),.C(g19347));
  NOR2 NOR2_600(.VSS(VSS),.VDD(VDD),.Y(g23081),.A(g17045),.B(g21141));
  NOR2 NOR2_601(.VSS(VSS),.VDD(VDD),.Y(g23083),.A(g21160),.B(g21193));
  NOR2 NOR2_602(.VSS(VSS),.VDD(VDD),.Y(g23092),.A(g17055),.B(g21154));
  NOR2 NOR2_603(.VSS(VSS),.VDD(VDD),.Y(g23093),.A(g17056),.B(g21155));
  NOR3 NOR3_355(.VSS(VSS),.VDD(VDD),.Y(g23096),.A(g21178),.B(g19351),.C(g19381));
  NOR2 NOR2_604(.VSS(VSS),.VDD(VDD),.Y(g23097),.A(g17079),.B(g21161));
  NOR2 NOR2_605(.VSS(VSS),.VDD(VDD),.Y(g23099),.A(g21180),.B(g21208));
  NOR2 NOR2_606(.VSS(VSS),.VDD(VDD),.Y(g23110),.A(g17090),.B(g21174));
  NOR2 NOR2_607(.VSS(VSS),.VDD(VDD),.Y(g23111),.A(g17091),.B(g21175));
  NOR3 NOR3_356(.VSS(VSS),.VDD(VDD),.Y(g23113),.A(g21198),.B(g19385),.C(g19413));
  NOR2 NOR2_608(.VSS(VSS),.VDD(VDD),.Y(g23114),.A(g17114),.B(g21181));
  NOR2 NOR2_609(.VSS(VSS),.VDD(VDD),.Y(g23117),.A(g17117),.B(g21188));
  NOR2 NOR2_610(.VSS(VSS),.VDD(VDD),.Y(g23123),.A(g17128),.B(g21194));
  NOR2 NOR2_611(.VSS(VSS),.VDD(VDD),.Y(g23124),.A(g17129),.B(g21195));
  NOR2 NOR2_612(.VSS(VSS),.VDD(VDD),.Y(g23126),.A(g17144),.B(g21203));
  NOR2 NOR2_613(.VSS(VSS),.VDD(VDD),.Y(g23132),.A(g17155),.B(g21209));
  NOR2 NOR2_614(.VSS(VSS),.VDD(VDD),.Y(g23133),.A(g17156),.B(g21210));
  NOR2 NOR2_615(.VSS(VSS),.VDD(VDD),.Y(g23135),.A(g21229),.B(g19449));
  NOR2 NOR2_616(.VSS(VSS),.VDD(VDD),.Y(g23136),.A(g20878),.B(g10024));
  NOR2 NOR2_617(.VSS(VSS),.VDD(VDD),.Y(g23137),.A(g17167),.B(g21218));
  NOR2 NOR2_618(.VSS(VSS),.VDD(VDD),.Y(g23324),.A(g22144),.B(g10024));
  NOR2 NOR2_619(.VSS(VSS),.VDD(VDD),.Y(g23329),.A(g22165),.B(g10133));
  NOR2 NOR2_620(.VSS(VSS),.VDD(VDD),.Y(g23330),.A(g22186),.B(g22777));
  NOR2 NOR2_621(.VSS(VSS),.VDD(VDD),.Y(g23339),.A(g22181),.B(g10238));
  NOR2 NOR2_622(.VSS(VSS),.VDD(VDD),.Y(g23348),.A(g22195),.B(g10340));
  NOR2 NOR2_623(.VSS(VSS),.VDD(VDD),.Y(g23357),.A(g22210),.B(g20127));
  NOR2 NOR2_624(.VSS(VSS),.VDD(VDD),.Y(g23358),.A(g22227),.B(g18407));
  NOR2 NOR2_625(.VSS(VSS),.VDD(VDD),.Y(g23359),.A(g22216),.B(g22907));
  NOR2 NOR2_626(.VSS(VSS),.VDD(VDD),.Y(g23385),.A(g17393),.B(g22517));
  NOR2 NOR2_627(.VSS(VSS),.VDD(VDD),.Y(g23386),.A(g22483),.B(g21388));
  NOR2 NOR2_628(.VSS(VSS),.VDD(VDD),.Y(g23392),.A(g17460),.B(g22557));
  NOR2 NOR2_629(.VSS(VSS),.VDD(VDD),.Y(g23393),.A(g22526),.B(g21418));
  NOR2 NOR2_630(.VSS(VSS),.VDD(VDD),.Y(g23399),.A(g17506),.B(g22581));
  NOR2 NOR2_631(.VSS(VSS),.VDD(VDD),.Y(g23400),.A(g17540),.B(g22597));
  NOR2 NOR2_632(.VSS(VSS),.VDD(VDD),.Y(g23401),.A(g22566),.B(g21452));
  NOR2 NOR2_633(.VSS(VSS),.VDD(VDD),.Y(g23406),.A(g17597),.B(g22618));
  NOR2 NOR2_634(.VSS(VSS),.VDD(VDD),.Y(g23407),.A(g17630),.B(g22634));
  NOR2 NOR2_635(.VSS(VSS),.VDD(VDD),.Y(g23408),.A(g22606),.B(g21494));
  NOR2 NOR2_636(.VSS(VSS),.VDD(VDD),.Y(g23413),.A(g17694),.B(g22654));
  NOR2 NOR2_637(.VSS(VSS),.VDD(VDD),.Y(g23418),.A(g17794),.B(g22690));
  NOR2 NOR2_638(.VSS(VSS),.VDD(VDD),.Y(g23427),.A(g22699),.B(g21589));
  NOR2 NOR2_639(.VSS(VSS),.VDD(VDD),.Y(g23433),.A(g22726),.B(g21611));
  NOR2 NOR2_640(.VSS(VSS),.VDD(VDD),.Y(g23461),.A(g22841),.B(g21707));
  NOR2 NOR2_641(.VSS(VSS),.VDD(VDD),.Y(g23477),.A(g22906),.B(g21758));
  NOR2 NOR2_642(.VSS(VSS),.VDD(VDD),.Y(g23497),.A(g22876),.B(g5606));
  NOR2 NOR2_643(.VSS(VSS),.VDD(VDD),.Y(g23513),.A(g22911),.B(g5631));
  NOR2 NOR2_644(.VSS(VSS),.VDD(VDD),.Y(g23528),.A(g22936),.B(g5659));
  NOR2 NOR2_645(.VSS(VSS),.VDD(VDD),.Y(g23539),.A(g22942),.B(g5697));
  NOR2 NOR2_646(.VSS(VSS),.VDD(VDD),.Y(g23545),.A(g22984),.B(g20285));
  NOR3 NOR3_357(.VSS(VSS),.VDD(VDD),.Y(g23823),.A(g23009),.B(g18490),.C(g4456));
  NOR3 NOR3_358(.VSS(VSS),.VDD(VDD),.Y(g23858),.A(g23025),.B(g18554),.C(g4632));
  NOR3 NOR3_359(.VSS(VSS),.VDD(VDD),.Y(g23892),.A(g23042),.B(g18604),.C(g4809));
  NOR3 NOR3_360(.VSS(VSS),.VDD(VDD),.Y(g23913),.A(g23061),.B(g18636),.C(g4985));
  NOR2 NOR2_647(.VSS(VSS),.VDD(VDD),.Y(g23922),.A(g4456),.B(g22985));
  NOR3 NOR3_361(.VSS(VSS),.VDD(VDD),.Y(g23945),.A(g4456),.B(g13565),.C(g23009));
  NOR2 NOR2_648(.VSS(VSS),.VDD(VDD),.Y(g23950),.A(g22992),.B(g6707));
  NOR2 NOR2_649(.VSS(VSS),.VDD(VDD),.Y(g23954),.A(g4632),.B(g22987));
  NOR3 NOR3_362(.VSS(VSS),.VDD(VDD),.Y(g23974),.A(g4632),.B(g13573),.C(g23025));
  NOR2 NOR2_650(.VSS(VSS),.VDD(VDD),.Y(g23979),.A(g23003),.B(g7009));
  NOR2 NOR2_651(.VSS(VSS),.VDD(VDD),.Y(g23983),.A(g4809),.B(g22990));
  NOR3 NOR3_363(.VSS(VSS),.VDD(VDD),.Y(g24004),.A(g4809),.B(g13582),.C(g23042));
  NOR2 NOR2_652(.VSS(VSS),.VDD(VDD),.Y(g24009),.A(g23017),.B(g7259));
  NOR2 NOR2_653(.VSS(VSS),.VDD(VDD),.Y(g24013),.A(g4985),.B(g22997));
  NOR3 NOR3_364(.VSS(VSS),.VDD(VDD),.Y(g24038),.A(g4985),.B(g13602),.C(g23061));
  NOR2 NOR2_654(.VSS(VSS),.VDD(VDD),.Y(g24043),.A(g23033),.B(g7455));
  NOR2 NOR2_655(.VSS(VSS),.VDD(VDD),.Y(g24059),.A(g21990),.B(g20809));
  NOR2 NOR2_656(.VSS(VSS),.VDD(VDD),.Y(g24072),.A(g22004),.B(g20826));
  NOR2 NOR2_657(.VSS(VSS),.VDD(VDD),.Y(g24083),.A(g22015),.B(g20836));
  NOR2 NOR2_658(.VSS(VSS),.VDD(VDD),.Y(g24092),.A(g22020),.B(g20840));
  NOR2 NOR2_659(.VSS(VSS),.VDD(VDD),.Y(g24174),.A(g16894),.B(g22206));
  NOR2 NOR2_660(.VSS(VSS),.VDD(VDD),.Y(g24178),.A(g16908),.B(g22211));
  NOR2 NOR2_661(.VSS(VSS),.VDD(VDD),.Y(g24179),.A(g16923),.B(g22214));
  NOR2 NOR2_662(.VSS(VSS),.VDD(VDD),.Y(g24181),.A(g16938),.B(g22220));
  NOR2 NOR2_663(.VSS(VSS),.VDD(VDD),.Y(g24182),.A(g16953),.B(g22223));
  NOR2 NOR2_664(.VSS(VSS),.VDD(VDD),.Y(g24206),.A(g16966),.B(g22228));
  NOR2 NOR2_665(.VSS(VSS),.VDD(VDD),.Y(g24207),.A(g16967),.B(g22229));
  NOR2 NOR2_666(.VSS(VSS),.VDD(VDD),.Y(g24208),.A(g16969),.B(g22235));
  NOR2 NOR2_667(.VSS(VSS),.VDD(VDD),.Y(g24209),.A(g16984),.B(g22238));
  NOR2 NOR2_668(.VSS(VSS),.VDD(VDD),.Y(g24212),.A(g16987),.B(g22244));
  NOR2 NOR2_669(.VSS(VSS),.VDD(VDD),.Y(g24213),.A(g16988),.B(g22245));
  NOR2 NOR2_670(.VSS(VSS),.VDD(VDD),.Y(g24214),.A(g16990),.B(g22250));
  NOR2 NOR2_671(.VSS(VSS),.VDD(VDD),.Y(g24215),.A(g16993),.B(g22254));
  NOR2 NOR2_672(.VSS(VSS),.VDD(VDD),.Y(g24216),.A(g16994),.B(g22255));
  NOR2 NOR2_673(.VSS(VSS),.VDD(VDD),.Y(g24218),.A(g16997),.B(g22264));
  NOR2 NOR2_674(.VSS(VSS),.VDD(VDD),.Y(g24219),.A(g16998),.B(g22265));
  NOR2 NOR2_675(.VSS(VSS),.VDD(VDD),.Y(g24222),.A(g17017),.B(g22272));
  NOR2 NOR2_676(.VSS(VSS),.VDD(VDD),.Y(g24223),.A(g17018),.B(g22273));
  NOR2 NOR2_677(.VSS(VSS),.VDD(VDD),.Y(g24225),.A(g17021),.B(g22281));
  NOR2 NOR2_678(.VSS(VSS),.VDD(VDD),.Y(g24226),.A(g17022),.B(g22282));
  NOR2 NOR2_679(.VSS(VSS),.VDD(VDD),.Y(g24227),.A(g22270),.B(g21137));
  NOR2 NOR2_680(.VSS(VSS),.VDD(VDD),.Y(g24228),.A(g17028),.B(g22285));
  NOR2 NOR2_681(.VSS(VSS),.VDD(VDD),.Y(g24230),.A(g17047),.B(g22291));
  NOR2 NOR2_682(.VSS(VSS),.VDD(VDD),.Y(g24231),.A(g17048),.B(g22292));
  NOR2 NOR2_683(.VSS(VSS),.VDD(VDD),.Y(g24232),.A(g22637),.B(g22665));
  NOR2 NOR2_684(.VSS(VSS),.VDD(VDD),.Y(g24234),.A(g22289),.B(g21157));
  NOR2 NOR2_685(.VSS(VSS),.VDD(VDD),.Y(g24235),.A(g17062),.B(g22305));
  NOR2 NOR2_686(.VSS(VSS),.VDD(VDD),.Y(g24237),.A(g17081),.B(g22311));
  NOR2 NOR2_687(.VSS(VSS),.VDD(VDD),.Y(g24238),.A(g17082),.B(g22312));
  NOR2 NOR2_688(.VSS(VSS),.VDD(VDD),.Y(g24242),.A(g22309),.B(g21177));
  NOR2 NOR2_689(.VSS(VSS),.VDD(VDD),.Y(g24243),.A(g17097),.B(g22333));
  NOR2 NOR2_690(.VSS(VSS),.VDD(VDD),.Y(g24249),.A(g22337),.B(g21197));
  NOR2 NOR2_691(.VSS(VSS),.VDD(VDD),.Y(g24250),.A(g17135),.B(g22358));
  NOR2 NOR2_692(.VSS(VSS),.VDD(VDD),.Y(g24426),.A(g23386),.B(g10024));
  NOR2 NOR2_693(.VSS(VSS),.VDD(VDD),.Y(g24428),.A(g23544),.B(g22398));
  NOR2 NOR2_694(.VSS(VSS),.VDD(VDD),.Y(g24430),.A(g23393),.B(g10133));
  NOR2 NOR2_695(.VSS(VSS),.VDD(VDD),.Y(g24434),.A(g23401),.B(g10238));
  NOR2 NOR2_696(.VSS(VSS),.VDD(VDD),.Y(g24438),.A(g23408),.B(g10340));
  NOR2 NOR2_697(.VSS(VSS),.VDD(VDD),.Y(g24445),.A(g23427),.B(g22777));
  NOR2 NOR2_698(.VSS(VSS),.VDD(VDD),.Y(g24446),.A(g23433),.B(g22907));
  NOR2 NOR2_699(.VSS(VSS),.VDD(VDD),.Y(g24473),.A(g23461),.B(g18407));
  NOR2 NOR2_700(.VSS(VSS),.VDD(VDD),.Y(g24476),.A(g23477),.B(g20127));
  NOR2 NOR2_701(.VSS(VSS),.VDD(VDD),.Y(g24479),.A(g23593),.B(g22516));
  NOR2 NOR2_702(.VSS(VSS),.VDD(VDD),.Y(g24480),.A(g23617),.B(g23659));
  NOR2 NOR2_703(.VSS(VSS),.VDD(VDD),.Y(g24481),.A(g23618),.B(g19696));
  NOR2 NOR2_704(.VSS(VSS),.VDD(VDD),.Y(g24485),.A(g23625),.B(g22556));
  NOR2 NOR2_705(.VSS(VSS),.VDD(VDD),.Y(g24486),.A(g23643),.B(g22577));
  NOR2 NOR2_706(.VSS(VSS),.VDD(VDD),.Y(g24487),.A(g23666),.B(g23709));
  NOR2 NOR2_707(.VSS(VSS),.VDD(VDD),.Y(g24488),.A(g23667),.B(g19740));
  NOR2 NOR2_708(.VSS(VSS),.VDD(VDD),.Y(g24489),.A(g23674),.B(g22596));
  NOR2 NOR2_709(.VSS(VSS),.VDD(VDD),.Y(g24490),.A(g23686),.B(g22607));
  NOR2 NOR2_710(.VSS(VSS),.VDD(VDD),.Y(g24491),.A(g15247),.B(g23735));
  NOR2 NOR2_711(.VSS(VSS),.VDD(VDD),.Y(g24492),.A(g23689),.B(g22610));
  NOR2 NOR2_712(.VSS(VSS),.VDD(VDD),.Y(g24493),.A(g23693),.B(g22614));
  NOR2 NOR2_713(.VSS(VSS),.VDD(VDD),.Y(g24494),.A(g23716),.B(g23763));
  NOR2 NOR2_714(.VSS(VSS),.VDD(VDD),.Y(g24495),.A(g23717),.B(g19783));
  NOR2 NOR2_715(.VSS(VSS),.VDD(VDD),.Y(g24496),.A(g23724),.B(g22633));
  NOR2 NOR2_716(.VSS(VSS),.VDD(VDD),.Y(g24497),.A(g23734),.B(g22638));
  NOR2 NOR2_717(.VSS(VSS),.VDD(VDD),.Y(g24498),.A(g15324),.B(g23777));
  NOR2 NOR2_718(.VSS(VSS),.VDD(VDD),.Y(g24499),.A(g15325),.B(g23778));
  NOR2 NOR2_719(.VSS(VSS),.VDD(VDD),.Y(g24500),.A(g23740),.B(g22643));
  NOR2 NOR2_720(.VSS(VSS),.VDD(VDD),.Y(g24501),.A(g15339),.B(g23790));
  NOR2 NOR2_721(.VSS(VSS),.VDD(VDD),.Y(g24502),.A(g23743),.B(g22646));
  NOR2 NOR2_722(.VSS(VSS),.VDD(VDD),.Y(g24503),.A(g23747),.B(g22650));
  NOR2 NOR2_723(.VSS(VSS),.VDD(VDD),.Y(g24504),.A(g23770),.B(g23818));
  NOR2 NOR2_724(.VSS(VSS),.VDD(VDD),.Y(g24505),.A(g23771),.B(g19825));
  NOR2 NOR2_725(.VSS(VSS),.VDD(VDD),.Y(g24506),.A(g23776),.B(g22667));
  NOR2 NOR2_726(.VSS(VSS),.VDD(VDD),.Y(g24507),.A(g15391),.B(g23824));
  NOR2 NOR2_727(.VSS(VSS),.VDD(VDD),.Y(g24508),.A(g15392),.B(g23825));
  NOR2 NOR2_728(.VSS(VSS),.VDD(VDD),.Y(g24509),.A(g23789),.B(g22674));
  NOR2 NOR2_729(.VSS(VSS),.VDD(VDD),.Y(g24510),.A(g15410),.B(g23830));
  NOR2 NOR2_730(.VSS(VSS),.VDD(VDD),.Y(g24511),.A(g15411),.B(g23831));
  NOR2 NOR2_731(.VSS(VSS),.VDD(VDD),.Y(g24512),.A(g23795),.B(g22679));
  NOR2 NOR2_732(.VSS(VSS),.VDD(VDD),.Y(g24513),.A(g15425),.B(g23843));
  NOR2 NOR2_733(.VSS(VSS),.VDD(VDD),.Y(g24514),.A(g23798),.B(g22682));
  NOR2 NOR2_734(.VSS(VSS),.VDD(VDD),.Y(g24515),.A(g23802),.B(g22686));
  NOR2 NOR2_735(.VSS(VSS),.VDD(VDD),.Y(g24516),.A(g23820),.B(g22700));
  NOR2 NOR2_736(.VSS(VSS),.VDD(VDD),.Y(g24517),.A(g23822),.B(g22701));
  NOR2 NOR2_737(.VSS(VSS),.VDD(VDD),.Y(g24519),.A(g15459),.B(g23855));
  NOR2 NOR2_738(.VSS(VSS),.VDD(VDD),.Y(g24520),.A(g23829),.B(g22707));
  NOR2 NOR2_739(.VSS(VSS),.VDD(VDD),.Y(g24521),.A(g15475),.B(g23859));
  NOR2 NOR2_740(.VSS(VSS),.VDD(VDD),.Y(g24522),.A(g15476),.B(g23860));
  NOR2 NOR2_741(.VSS(VSS),.VDD(VDD),.Y(g24523),.A(g23842),.B(g22714));
  NOR2 NOR2_742(.VSS(VSS),.VDD(VDD),.Y(g24524),.A(g15494),.B(g23865));
  NOR2 NOR2_743(.VSS(VSS),.VDD(VDD),.Y(g24525),.A(g15495),.B(g23866));
  NOR2 NOR2_744(.VSS(VSS),.VDD(VDD),.Y(g24526),.A(g23848),.B(g22719));
  NOR2 NOR2_745(.VSS(VSS),.VDD(VDD),.Y(g24527),.A(g15509),.B(g23878));
  NOR2 NOR2_746(.VSS(VSS),.VDD(VDD),.Y(g24528),.A(g23851),.B(g22722));
  NOR2 NOR2_747(.VSS(VSS),.VDD(VDD),.Y(g24530),.A(g23857),.B(g22732));
  NOR2 NOR2_748(.VSS(VSS),.VDD(VDD),.Y(g24532),.A(g15545),.B(g23889));
  NOR2 NOR2_749(.VSS(VSS),.VDD(VDD),.Y(g24533),.A(g23864),.B(g22738));
  NOR2 NOR2_750(.VSS(VSS),.VDD(VDD),.Y(g24534),.A(g15561),.B(g23893));
  NOR2 NOR2_751(.VSS(VSS),.VDD(VDD),.Y(g24535),.A(g15562),.B(g23894));
  NOR2 NOR2_752(.VSS(VSS),.VDD(VDD),.Y(g24536),.A(g23877),.B(g22745));
  NOR2 NOR2_753(.VSS(VSS),.VDD(VDD),.Y(g24537),.A(g15580),.B(g23899));
  NOR2 NOR2_754(.VSS(VSS),.VDD(VDD),.Y(g24538),.A(g15581),.B(g23900));
  NOR2 NOR2_755(.VSS(VSS),.VDD(VDD),.Y(g24543),.A(g23891),.B(g22764));
  NOR2 NOR2_756(.VSS(VSS),.VDD(VDD),.Y(g24545),.A(g15623),.B(g23910));
  NOR2 NOR2_757(.VSS(VSS),.VDD(VDD),.Y(g24546),.A(g23898),.B(g22770));
  NOR2 NOR2_758(.VSS(VSS),.VDD(VDD),.Y(g24547),.A(g15639),.B(g23914));
  NOR2 NOR2_759(.VSS(VSS),.VDD(VDD),.Y(g24548),.A(g15640),.B(g23915));
  NOR2 NOR2_760(.VSS(VSS),.VDD(VDD),.Y(g24555),.A(g23912),.B(g22798));
  NOR2 NOR2_761(.VSS(VSS),.VDD(VDD),.Y(g24557),.A(g15699),.B(g23942));
  NOR2 NOR2_762(.VSS(VSS),.VDD(VDD),.Y(g24558),.A(g23917),.B(g22804));
  NOR2 NOR2_763(.VSS(VSS),.VDD(VDD),.Y(g24566),.A(g23944),.B(g22842));
  NOR2 NOR2_764(.VSS(VSS),.VDD(VDD),.Y(g24575),.A(g23972),.B(g22874));
  NOR2 NOR2_765(.VSS(VSS),.VDD(VDD),.Y(g24606),.A(g24183),.B(g537));
  NOR2 NOR2_766(.VSS(VSS),.VDD(VDD),.Y(g24613),.A(g23592),.B(g22515));
  NOR2 NOR2_767(.VSS(VSS),.VDD(VDD),.Y(g24622),.A(g23616),.B(g22546));
  NOR2 NOR2_768(.VSS(VSS),.VDD(VDD),.Y(g24623),.A(g24183),.B(g529));
  NOR2 NOR2_769(.VSS(VSS),.VDD(VDD),.Y(g24624),.A(g23624),.B(g22555));
  NOR2 NOR2_770(.VSS(VSS),.VDD(VDD),.Y(g24636),.A(g24183),.B(g530));
  NOR2 NOR2_771(.VSS(VSS),.VDD(VDD),.Y(g24637),.A(g23665),.B(g22587));
  NOR2 NOR2_772(.VSS(VSS),.VDD(VDD),.Y(g24638),.A(g23673),.B(g22595));
  NOR2 NOR2_773(.VSS(VSS),.VDD(VDD),.Y(g24652),.A(g24183),.B(g531));
  NOR2 NOR2_774(.VSS(VSS),.VDD(VDD),.Y(g24656),.A(g23715),.B(g22624));
  NOR2 NOR2_775(.VSS(VSS),.VDD(VDD),.Y(g24657),.A(g23723),.B(g22632));
  NOR2 NOR2_776(.VSS(VSS),.VDD(VDD),.Y(g24663),.A(g24183),.B(g532));
  NOR2 NOR2_777(.VSS(VSS),.VDD(VDD),.Y(g24675),.A(g23769),.B(g22660));
  NOR2 NOR2_778(.VSS(VSS),.VDD(VDD),.Y(g24681),.A(g24183),.B(g533));
  NOR2 NOR2_779(.VSS(VSS),.VDD(VDD),.Y(g24682),.A(g23688),.B(g24183));
  NOR2 NOR2_780(.VSS(VSS),.VDD(VDD),.Y(g24694),.A(g24183),.B(g534));
  NOR2 NOR2_781(.VSS(VSS),.VDD(VDD),.Y(g24708),.A(g23854),.B(g22727));
  NOR2 NOR2_782(.VSS(VSS),.VDD(VDD),.Y(g24711),.A(g24183),.B(g536));
  NOR2 NOR2_783(.VSS(VSS),.VDD(VDD),.Y(g24717),.A(g23886),.B(g22754));
  NOR2 NOR2_784(.VSS(VSS),.VDD(VDD),.Y(g24720),.A(g23888),.B(g22759));
  NOR2 NOR2_785(.VSS(VSS),.VDD(VDD),.Y(g24728),.A(g23907),.B(g22788));
  NOR2 NOR2_786(.VSS(VSS),.VDD(VDD),.Y(g24731),.A(g23909),.B(g22793));
  NOR2 NOR2_787(.VSS(VSS),.VDD(VDD),.Y(g24736),.A(g23939),.B(g22830));
  NOR2 NOR2_788(.VSS(VSS),.VDD(VDD),.Y(g24739),.A(g23941),.B(g22835));
  NOR2 NOR2_789(.VSS(VSS),.VDD(VDD),.Y(g24742),.A(g23971),.B(g22869));
  NOR2 NOR2_790(.VSS(VSS),.VDD(VDD),.Y(g24756),.A(g16089),.B(g24211));
  NOR2 NOR2_791(.VSS(VSS),.VDD(VDD),.Y(g24770),.A(g16119),.B(g24217));
  NOR2 NOR2_792(.VSS(VSS),.VDD(VDD),.Y(g24782),.A(g16160),.B(g24221));
  NOR2 NOR2_793(.VSS(VSS),.VDD(VDD),.Y(g24783),.A(g16161),.B(g24224));
  NOR2 NOR2_794(.VSS(VSS),.VDD(VDD),.Y(g24800),.A(g16211),.B(g24229));
  NOR2 NOR2_795(.VSS(VSS),.VDD(VDD),.Y(g24819),.A(g16262),.B(g24236));
  NOR2 NOR2_796(.VSS(VSS),.VDD(VDD),.Y(g24836),.A(g16309),.B(g24241));
  NOR2 NOR2_797(.VSS(VSS),.VDD(VDD),.Y(g24845),.A(g16350),.B(g24246));
  NOR2 NOR2_798(.VSS(VSS),.VDD(VDD),.Y(g24847),.A(g16356),.B(g24247));
  NOR2 NOR2_799(.VSS(VSS),.VDD(VDD),.Y(g24859),.A(g16390),.B(g24253));
  NOR2 NOR2_800(.VSS(VSS),.VDD(VDD),.Y(g24871),.A(g16422),.B(g24256));
  NOR2 NOR2_801(.VSS(VSS),.VDD(VDD),.Y(g25027),.A(g24227),.B(g17001));
  NOR2 NOR2_802(.VSS(VSS),.VDD(VDD),.Y(g25042),.A(g24234),.B(g17031));
  NOR2 NOR2_803(.VSS(VSS),.VDD(VDD),.Y(g25056),.A(g24242),.B(g17065));
  NOR2 NOR2_804(.VSS(VSS),.VDD(VDD),.Y(g25067),.A(g24249),.B(g17100));
  NOR2 NOR2_805(.VSS(VSS),.VDD(VDD),.Y(g25075),.A(g13880),.B(g23483));
  NOR2 NOR2_806(.VSS(VSS),.VDD(VDD),.Y(g25076),.A(g23409),.B(g22187));
  NOR2 NOR2_807(.VSS(VSS),.VDD(VDD),.Y(g25077),.A(g23414),.B(g22196));
  NOR2 NOR2_808(.VSS(VSS),.VDD(VDD),.Y(g25078),.A(g23419),.B(g22201));
  NOR2 NOR2_809(.VSS(VSS),.VDD(VDD),.Y(g25081),.A(g23423),.B(g22202));
  NOR2 NOR2_810(.VSS(VSS),.VDD(VDD),.Y(g25082),.A(g23428),.B(g22207));
  NOR2 NOR2_811(.VSS(VSS),.VDD(VDD),.Y(g25085),.A(g23432),.B(g22208));
  NOR2 NOR2_812(.VSS(VSS),.VDD(VDD),.Y(g25091),.A(g23434),.B(g22215));
  NOR2 NOR2_813(.VSS(VSS),.VDD(VDD),.Y(g25099),.A(g23440),.B(g22224));
  NOR2 NOR2_814(.VSS(VSS),.VDD(VDD),.Y(g25125),.A(g23510),.B(g22340));
  NOR2 NOR2_815(.VSS(VSS),.VDD(VDD),.Y(g25127),.A(g23525),.B(g22363));
  NOR2 NOR2_816(.VSS(VSS),.VDD(VDD),.Y(g25129),.A(g23536),.B(g22383));
  NOR2 NOR2_817(.VSS(VSS),.VDD(VDD),.Y(g25185),.A(g24492),.B(g10024));
  NOR2 NOR2_818(.VSS(VSS),.VDD(VDD),.Y(g25189),.A(g24502),.B(g10133));
  NOR2 NOR2_819(.VSS(VSS),.VDD(VDD),.Y(g25191),.A(g24516),.B(g22777));
  NOR2 NOR2_820(.VSS(VSS),.VDD(VDD),.Y(g25194),.A(g24514),.B(g10238));
  NOR2 NOR2_821(.VSS(VSS),.VDD(VDD),.Y(g25197),.A(g24528),.B(g10340));
  NOR2 NOR2_822(.VSS(VSS),.VDD(VDD),.Y(g25199),.A(g24558),.B(g20127));
  NOR2 NOR2_823(.VSS(VSS),.VDD(VDD),.Y(g25201),.A(g24575),.B(g18407));
  NOR2 NOR2_824(.VSS(VSS),.VDD(VDD),.Y(g25202),.A(g24566),.B(g22907));
  NOR2 NOR2_825(.VSS(VSS),.VDD(VDD),.Y(g25204),.A(g24745),.B(g23547));
  NOR2 NOR2_826(.VSS(VSS),.VDD(VDD),.Y(g25206),.A(g24746),.B(g23550));
  NOR2 NOR2_827(.VSS(VSS),.VDD(VDD),.Y(g25207),.A(g24747),.B(g23551));
  NOR2 NOR2_828(.VSS(VSS),.VDD(VDD),.Y(g25208),.A(g24748),.B(g23552));
  NOR2 NOR2_829(.VSS(VSS),.VDD(VDD),.Y(g25209),.A(g24749),.B(g23554));
  NOR2 NOR2_830(.VSS(VSS),.VDD(VDD),.Y(g25211),.A(g24750),.B(g23558));
  NOR2 NOR2_831(.VSS(VSS),.VDD(VDD),.Y(g25212),.A(g24751),.B(g23559));
  NOR2 NOR2_832(.VSS(VSS),.VDD(VDD),.Y(g25213),.A(g24752),.B(g23560));
  NOR2 NOR2_833(.VSS(VSS),.VDD(VDD),.Y(g25214),.A(g24754),.B(g23563));
  NOR2 NOR2_834(.VSS(VSS),.VDD(VDD),.Y(g25215),.A(g24755),.B(g23564));
  NOR2 NOR2_835(.VSS(VSS),.VDD(VDD),.Y(g25216),.A(g24757),.B(g23565));
  NOR2 NOR2_836(.VSS(VSS),.VDD(VDD),.Y(g25217),.A(g24758),.B(g23567));
  NOR2 NOR2_837(.VSS(VSS),.VDD(VDD),.Y(g25218),.A(g24760),.B(g23571));
  NOR2 NOR2_838(.VSS(VSS),.VDD(VDD),.Y(g25219),.A(g24761),.B(g23572));
  NOR2 NOR2_839(.VSS(VSS),.VDD(VDD),.Y(g25220),.A(g24762),.B(g23573));
  NOR2 NOR2_840(.VSS(VSS),.VDD(VDD),.Y(g25221),.A(g24767),.B(g23577));
  NOR2 NOR2_841(.VSS(VSS),.VDD(VDD),.Y(g25222),.A(g24768),.B(g23578));
  NOR2 NOR2_842(.VSS(VSS),.VDD(VDD),.Y(g25223),.A(g24769),.B(g23579));
  NOR2 NOR2_843(.VSS(VSS),.VDD(VDD),.Y(g25224),.A(g24772),.B(g23582));
  NOR2 NOR2_844(.VSS(VSS),.VDD(VDD),.Y(g25225),.A(g24773),.B(g23583));
  NOR2 NOR2_845(.VSS(VSS),.VDD(VDD),.Y(g25226),.A(g24774),.B(g23584));
  NOR2 NOR2_846(.VSS(VSS),.VDD(VDD),.Y(g25227),.A(g24775),.B(g23586));
  NOR2 NOR2_847(.VSS(VSS),.VDD(VDD),.Y(g25228),.A(g24776),.B(g23590));
  NOR2 NOR2_848(.VSS(VSS),.VDD(VDD),.Y(g25229),.A(g24777),.B(g23591));
  NOR2 NOR2_849(.VSS(VSS),.VDD(VDD),.Y(g25230),.A(g24779),.B(g23598));
  NOR2 NOR2_850(.VSS(VSS),.VDD(VDD),.Y(g25231),.A(g24780),.B(g23599));
  NOR2 NOR2_851(.VSS(VSS),.VDD(VDD),.Y(g25232),.A(g24781),.B(g23600));
  NOR2 NOR2_852(.VSS(VSS),.VDD(VDD),.Y(g25233),.A(g24788),.B(g23604));
  NOR2 NOR2_853(.VSS(VSS),.VDD(VDD),.Y(g25234),.A(g24789),.B(g23605));
  NOR2 NOR2_854(.VSS(VSS),.VDD(VDD),.Y(g25235),.A(g24790),.B(g23606));
  NOR2 NOR2_855(.VSS(VSS),.VDD(VDD),.Y(g25236),.A(g24792),.B(g23609));
  NOR2 NOR2_856(.VSS(VSS),.VDD(VDD),.Y(g25237),.A(g24793),.B(g23610));
  NOR2 NOR2_857(.VSS(VSS),.VDD(VDD),.Y(g25238),.A(g24794),.B(g23611));
  NOR2 NOR2_858(.VSS(VSS),.VDD(VDD),.Y(g25239),.A(g24796),.B(g23615));
  NOR2 NOR2_859(.VSS(VSS),.VDD(VDD),.Y(g25240),.A(g24798),.B(g23622));
  NOR2 NOR2_860(.VSS(VSS),.VDD(VDD),.Y(g25241),.A(g24799),.B(g23623));
  NOR2 NOR2_861(.VSS(VSS),.VDD(VDD),.Y(g25242),.A(g24802),.B(g23630));
  NOR2 NOR2_862(.VSS(VSS),.VDD(VDD),.Y(g25243),.A(g24803),.B(g23631));
  NOR2 NOR2_863(.VSS(VSS),.VDD(VDD),.Y(g25244),.A(g24804),.B(g23632));
  NOR2 NOR2_864(.VSS(VSS),.VDD(VDD),.Y(g25245),.A(g24809),.B(g23636));
  NOR2 NOR2_865(.VSS(VSS),.VDD(VDD),.Y(g25246),.A(g24810),.B(g23637));
  NOR2 NOR2_866(.VSS(VSS),.VDD(VDD),.Y(g25247),.A(g24811),.B(g23638));
  NOR2 NOR2_867(.VSS(VSS),.VDD(VDD),.Y(g25248),.A(g24818),.B(g23664));
  NOR2 NOR2_868(.VSS(VSS),.VDD(VDD),.Y(g25249),.A(g24821),.B(g23671));
  NOR2 NOR2_869(.VSS(VSS),.VDD(VDD),.Y(g25250),.A(g24822),.B(g23672));
  NOR2 NOR2_870(.VSS(VSS),.VDD(VDD),.Y(g25251),.A(g24824),.B(g23679));
  NOR2 NOR2_871(.VSS(VSS),.VDD(VDD),.Y(g25252),.A(g24825),.B(g23680));
  NOR2 NOR2_872(.VSS(VSS),.VDD(VDD),.Y(g25253),.A(g24826),.B(g23681));
  NOR2 NOR2_873(.VSS(VSS),.VDD(VDD),.Y(g25254),.A(g24831),.B(g23687));
  NOR2 NOR2_874(.VSS(VSS),.VDD(VDD),.Y(g25255),.A(g24838),.B(g23714));
  NOR2 NOR2_875(.VSS(VSS),.VDD(VDD),.Y(g25256),.A(g24840),.B(g23721));
  NOR2 NOR2_876(.VSS(VSS),.VDD(VDD),.Y(g25257),.A(g24841),.B(g23722));
  NOR2 NOR2_877(.VSS(VSS),.VDD(VDD),.Y(g25258),.A(g24846),.B(g23741));
  NOR2 NOR2_878(.VSS(VSS),.VDD(VDD),.Y(g25259),.A(g24853),.B(g23768));
  NOR2 NOR2_879(.VSS(VSS),.VDD(VDD),.Y(g25260),.A(g24858),.B(g17737));
  NOR2 NOR2_880(.VSS(VSS),.VDD(VDD),.Y(g25261),.A(g24861),.B(g23796));
  NOR2 NOR2_881(.VSS(VSS),.VDD(VDD),.Y(g25262),.A(g24869),.B(g17824));
  NOR2 NOR2_882(.VSS(VSS),.VDD(VDD),.Y(g25263),.A(g24874),.B(g17838));
  NOR2 NOR2_883(.VSS(VSS),.VDD(VDD),.Y(g25264),.A(g24876),.B(g23849));
  NOR2 NOR2_884(.VSS(VSS),.VDD(VDD),.Y(g25265),.A(g24878),.B(g23852));
  NOR2 NOR2_885(.VSS(VSS),.VDD(VDD),.Y(g25266),.A(g24881),.B(g17912));
  NOR2 NOR2_886(.VSS(VSS),.VDD(VDD),.Y(g25267),.A(g24884),.B(g17936));
  NOR2 NOR2_887(.VSS(VSS),.VDD(VDD),.Y(g25268),.A(g24888),.B(g17950));
  NOR2 NOR2_888(.VSS(VSS),.VDD(VDD),.Y(g25270),.A(g24898),.B(g18023));
  NOR2 NOR2_889(.VSS(VSS),.VDD(VDD),.Y(g25271),.A(g24901),.B(g18047));
  NOR2 NOR2_890(.VSS(VSS),.VDD(VDD),.Y(g25272),.A(g24905),.B(g18061));
  NOR2 NOR2_891(.VSS(VSS),.VDD(VDD),.Y(g25273),.A(g24907),.B(g23904));
  NOR2 NOR2_892(.VSS(VSS),.VDD(VDD),.Y(g25279),.A(g24921),.B(g18140));
  NOR2 NOR2_893(.VSS(VSS),.VDD(VDD),.Y(g25280),.A(g24924),.B(g18164));
  NOR2 NOR2_894(.VSS(VSS),.VDD(VDD),.Y(g25288),.A(g24938),.B(g18256));
  NOR2 NOR2_895(.VSS(VSS),.VDD(VDD),.Y(g25311),.A(g24964),.B(g24029));
  NOR2 NOR2_896(.VSS(VSS),.VDD(VDD),.Y(g25343),.A(g24975),.B(g5623));
  NOR2 NOR2_897(.VSS(VSS),.VDD(VDD),.Y(g25357),.A(g24986),.B(g5651));
  NOR2 NOR2_898(.VSS(VSS),.VDD(VDD),.Y(g25372),.A(g24997),.B(g5689));
  NOR2 NOR2_899(.VSS(VSS),.VDD(VDD),.Y(g25389),.A(g25005),.B(g5741));
  NOR2 NOR2_900(.VSS(VSS),.VDD(VDD),.Y(g25418),.A(g24482),.B(g22319));
  NOR2 NOR2_901(.VSS(VSS),.VDD(VDD),.Y(g25426),.A(g24183),.B(g24616));
  NOR2 NOR2_902(.VSS(VSS),.VDD(VDD),.Y(g25429),.A(g24482),.B(g22319));
  NOR2 NOR2_903(.VSS(VSS),.VDD(VDD),.Y(g25450),.A(g16018),.B(g25086));
  NOR2 NOR2_904(.VSS(VSS),.VDD(VDD),.Y(g25451),.A(g16048),.B(g25102));
  NOR2 NOR2_905(.VSS(VSS),.VDD(VDD),.Y(g25452),.A(g16101),.B(g25117));
  NOR2 NOR2_906(.VSS(VSS),.VDD(VDD),.Y(g25523),.A(g20842),.B(g24429));
  NOR2 NOR2_907(.VSS(VSS),.VDD(VDD),.Y(g25539),.A(g25088),.B(g6157));
  NOR2 NOR2_908(.VSS(VSS),.VDD(VDD),.Y(g25569),.A(g24708),.B(g24490));
  NOR2 NOR2_909(.VSS(VSS),.VDD(VDD),.Y(g25589),.A(g20850),.B(g24433));
  NOR2 NOR2_910(.VSS(VSS),.VDD(VDD),.Y(g25605),.A(g25096),.B(g6184));
  NOR2 NOR2_911(.VSS(VSS),.VDD(VDD),.Y(g25631),.A(g24717),.B(g24497));
  NOR2 NOR2_912(.VSS(VSS),.VDD(VDD),.Y(g25648),.A(g24720),.B(g24500));
  NOR2 NOR2_913(.VSS(VSS),.VDD(VDD),.Y(g25668),.A(g20858),.B(g24437));
  NOR2 NOR2_914(.VSS(VSS),.VDD(VDD),.Y(g25684),.A(g25106),.B(g6216));
  NOR2 NOR2_915(.VSS(VSS),.VDD(VDD),.Y(g25699),.A(g24613),.B(g24506));
  NOR2 NOR2_916(.VSS(VSS),.VDD(VDD),.Y(g25708),.A(g24728),.B(g24509));
  NOR2 NOR2_917(.VSS(VSS),.VDD(VDD),.Y(g25725),.A(g24731),.B(g24512));
  NOR2 NOR2_918(.VSS(VSS),.VDD(VDD),.Y(g25745),.A(g20866),.B(g24440));
  NOR2 NOR2_919(.VSS(VSS),.VDD(VDD),.Y(g25761),.A(g25112),.B(g6305));
  NOR2 NOR2_920(.VSS(VSS),.VDD(VDD),.Y(g25764),.A(g25076),.B(g21615));
  NOR2 NOR2_921(.VSS(VSS),.VDD(VDD),.Y(g25772),.A(g24624),.B(g24520));
  NOR2 NOR2_922(.VSS(VSS),.VDD(VDD),.Y(g25781),.A(g24736),.B(g24523));
  NOR2 NOR2_923(.VSS(VSS),.VDD(VDD),.Y(g25798),.A(g24739),.B(g24526));
  NOR2 NOR2_924(.VSS(VSS),.VDD(VDD),.Y(g25818),.A(g25077),.B(g21643));
  NOR2 NOR2_925(.VSS(VSS),.VDD(VDD),.Y(g25826),.A(g24638),.B(g24533));
  NOR2 NOR2_926(.VSS(VSS),.VDD(VDD),.Y(g25835),.A(g24742),.B(g24536));
  NOR3 NOR3_365(.VSS(VSS),.VDD(VDD),.Y(g25852),.A(g4456),.B(g14831),.C(g25078));
  NOR2 NOR2_927(.VSS(VSS),.VDD(VDD),.Y(g25853),.A(g25081),.B(g21674));
  NOR2 NOR2_928(.VSS(VSS),.VDD(VDD),.Y(g25861),.A(g24657),.B(g24546));
  NOR4 NOR4_16(.VSS(VSS),.VDD(VDD),.Y(g25870),.A(g4456),.B(g25078),.C(g18429),.D(g16075));
  NOR3 NOR3_366(.VSS(VSS),.VDD(VDD),.Y(g25873),.A(g4632),.B(g14904),.C(g25082));
  NOR2 NOR2_929(.VSS(VSS),.VDD(VDD),.Y(g25874),.A(g25085),.B(g21703));
  NOR4 NOR4_17(.VSS(VSS),.VDD(VDD),.Y(g25882),.A(g4632),.B(g25082),.C(g18502),.D(g16113));
  NOR3 NOR3_367(.VSS(VSS),.VDD(VDD),.Y(g25885),.A(g4809),.B(g14985),.C(g25091));
  NOR4 NOR4_18(.VSS(VSS),.VDD(VDD),.Y(g25887),.A(g4809),.B(g25091),.C(g18566),.D(g16164));
  NOR3 NOR3_368(.VSS(VSS),.VDD(VDD),.Y(g25890),.A(g4985),.B(g15074),.C(g25099));
  NOR4 NOR4_19(.VSS(VSS),.VDD(VDD),.Y(g25892),.A(g4985),.B(g25099),.C(g18616),.D(g16223));
  NOR2 NOR2_930(.VSS(VSS),.VDD(VDD),.Y(g25932),.A(g25125),.B(g17001));
  NOR2 NOR2_931(.VSS(VSS),.VDD(VDD),.Y(g25935),.A(g25127),.B(g17031));
  NOR2 NOR2_932(.VSS(VSS),.VDD(VDD),.Y(g25938),.A(g25129),.B(g17065));
  NOR2 NOR2_933(.VSS(VSS),.VDD(VDD),.Y(g25940),.A(g24428),.B(g17100));
  NOR2 NOR2_934(.VSS(VSS),.VDD(VDD),.Y(g25941),.A(g24529),.B(g24540));
  NOR2 NOR2_935(.VSS(VSS),.VDD(VDD),.Y(g25943),.A(g24541),.B(g24550));
  NOR2 NOR2_936(.VSS(VSS),.VDD(VDD),.Y(g25944),.A(g24542),.B(g24552));
  NOR2 NOR2_937(.VSS(VSS),.VDD(VDD),.Y(g25946),.A(g24553),.B(g24561));
  NOR2 NOR2_938(.VSS(VSS),.VDD(VDD),.Y(g25947),.A(g24554),.B(g24563));
  NOR2 NOR2_939(.VSS(VSS),.VDD(VDD),.Y(g25948),.A(g24564),.B(g24571));
  NOR2 NOR2_940(.VSS(VSS),.VDD(VDD),.Y(g25949),.A(g24565),.B(g24573));
  NOR2 NOR2_941(.VSS(VSS),.VDD(VDD),.Y(g25950),.A(g24574),.B(g24580));
  NOR2 NOR2_942(.VSS(VSS),.VDD(VDD),.Y(g25962),.A(g24591),.B(g23496));
  NOR2 NOR2_943(.VSS(VSS),.VDD(VDD),.Y(g25967),.A(g24596),.B(g23512));
  NOR2 NOR2_944(.VSS(VSS),.VDD(VDD),.Y(g25974),.A(g24604),.B(g23527));
  NOR2 NOR2_945(.VSS(VSS),.VDD(VDD),.Y(g25979),.A(g24611),.B(g23538));
  NOR2 NOR2_946(.VSS(VSS),.VDD(VDD),.Y(g26025),.A(g25392),.B(g17193));
  NOR2 NOR2_947(.VSS(VSS),.VDD(VDD),.Y(g26031),.A(g25273),.B(g22777));
  NOR2 NOR2_948(.VSS(VSS),.VDD(VDD),.Y(g26037),.A(g25311),.B(g18407));
  NOR2 NOR2_949(.VSS(VSS),.VDD(VDD),.Y(g26041),.A(g25475),.B(g24855));
  NOR2 NOR2_950(.VSS(VSS),.VDD(VDD),.Y(g26042),.A(g25505),.B(g24867));
  NOR2 NOR2_951(.VSS(VSS),.VDD(VDD),.Y(g26043),.A(g25506),.B(g24870));
  NOR2 NOR2_952(.VSS(VSS),.VDD(VDD),.Y(g26044),.A(g25552),.B(g24882));
  NOR2 NOR2_953(.VSS(VSS),.VDD(VDD),.Y(g26045),.A(g25553),.B(g24885));
  NOR2 NOR2_954(.VSS(VSS),.VDD(VDD),.Y(g26046),.A(g25618),.B(g24899));
  NOR2 NOR2_955(.VSS(VSS),.VDD(VDD),.Y(g26047),.A(g25619),.B(g24902));
  NOR2 NOR2_956(.VSS(VSS),.VDD(VDD),.Y(g26048),.A(g25628),.B(g24906));
  NOR2 NOR2_957(.VSS(VSS),.VDD(VDD),.Y(g26049),.A(g25629),.B(g24908));
  NOR2 NOR2_958(.VSS(VSS),.VDD(VDD),.Y(g26050),.A(g25697),.B(g24922));
  NOR2 NOR2_959(.VSS(VSS),.VDD(VDD),.Y(g26055),.A(g25881),.B(g24974));
  NOR2 NOR2_960(.VSS(VSS),.VDD(VDD),.Y(g26081),.A(g25470),.B(g25482));
  NOR2 NOR2_961(.VSS(VSS),.VDD(VDD),.Y(g26083),.A(g25426),.B(g22319));
  NOR2 NOR2_962(.VSS(VSS),.VDD(VDD),.Y(g26084),.A(g25487),.B(g25513));
  NOR3 NOR3_369(.VSS(VSS),.VDD(VDD),.Y(g26087),.A(g6068),.B(g24183),.C(g25319));
  NOR2 NOR2_963(.VSS(VSS),.VDD(VDD),.Y(g26090),.A(g25518),.B(g25560));
  NOR3 NOR3_370(.VSS(VSS),.VDD(VDD),.Y(g26096),.A(g6068),.B(g24183),.C(g25394));
  NOR3 NOR3_371(.VSS(VSS),.VDD(VDD),.Y(g26099),.A(g6068),.B(g24183),.C(g25313));
  NOR2 NOR2_964(.VSS(VSS),.VDD(VDD),.Y(g26103),.A(g25565),.B(g25626));
  NOR3 NOR3_372(.VSS(VSS),.VDD(VDD),.Y(g26107),.A(g6068),.B(g24183),.C(g25383));
  NOR3 NOR3_373(.VSS(VSS),.VDD(VDD),.Y(g26110),.A(g6068),.B(g24183),.C(g25305));
  NOR2 NOR2_965(.VSS(VSS),.VDD(VDD),.Y(g26113),.A(g25426),.B(g22319));
  NOR3 NOR3_374(.VSS(VSS),.VDD(VDD),.Y(g26126),.A(g6068),.B(g24183),.C(g25368));
  NOR3 NOR3_375(.VSS(VSS),.VDD(VDD),.Y(g26137),.A(g6068),.B(g24183),.C(g25355));
  NOR2 NOR2_966(.VSS(VSS),.VDD(VDD),.Y(g26140),.A(g24183),.B(g25430));
  NOR3 NOR3_376(.VSS(VSS),.VDD(VDD),.Y(g26145),.A(g6068),.B(g24183),.C(g25347));
  NOR3 NOR3_377(.VSS(VSS),.VDD(VDD),.Y(g26151),.A(g6068),.B(g24183),.C(g25335));
  NOR3 NOR3_378(.VSS(VSS),.VDD(VDD),.Y(g26154),.A(g6068),.B(g24183),.C(g25329));
  NOR2 NOR2_967(.VSS(VSS),.VDD(VDD),.Y(g26160),.A(g25951),.B(g16162));
  NOR2 NOR2_968(.VSS(VSS),.VDD(VDD),.Y(g26168),.A(g25953),.B(g16212));
  NOR2 NOR2_969(.VSS(VSS),.VDD(VDD),.Y(g26183),.A(g25957),.B(g13270));
  NOR2 NOR2_970(.VSS(VSS),.VDD(VDD),.Y(g26199),.A(g25961),.B(g13291));
  NOR2 NOR2_971(.VSS(VSS),.VDD(VDD),.Y(g26217),.A(g25963),.B(g13320));
  NOR2 NOR2_972(.VSS(VSS),.VDD(VDD),.Y(g26240),.A(g25968),.B(g13340));
  NOR2 NOR2_973(.VSS(VSS),.VDD(VDD),.Y(g26265),.A(g25972),.B(g13360));
  NOR2 NOR2_974(.VSS(VSS),.VDD(VDD),.Y(g26272),.A(g25973),.B(g16423));
  NOR2 NOR2_975(.VSS(VSS),.VDD(VDD),.Y(g26283),.A(g25954),.B(g24486));
  NOR2 NOR2_976(.VSS(VSS),.VDD(VDD),.Y(g26295),.A(g25977),.B(g13385));
  NOR2 NOR2_977(.VSS(VSS),.VDD(VDD),.Y(g26304),.A(g25978),.B(g16451));
  NOR2 NOR2_978(.VSS(VSS),.VDD(VDD),.Y(g26327),.A(g25958),.B(g24493));
  NOR2 NOR2_979(.VSS(VSS),.VDD(VDD),.Y(g26336),.A(g25981),.B(g13481));
  NOR2 NOR2_980(.VSS(VSS),.VDD(VDD),.Y(g26374),.A(g25964),.B(g24503));
  NOR2 NOR2_981(.VSS(VSS),.VDD(VDD),.Y(g26417),.A(g25969),.B(g24515));
  NOR2 NOR2_982(.VSS(VSS),.VDD(VDD),.Y(g26529),.A(g25962),.B(g17001));
  NOR2 NOR2_983(.VSS(VSS),.VDD(VDD),.Y(g26530),.A(g25967),.B(g17031));
  NOR2 NOR2_984(.VSS(VSS),.VDD(VDD),.Y(g26531),.A(g25974),.B(g17065));
  NOR2 NOR2_985(.VSS(VSS),.VDD(VDD),.Y(g26532),.A(g25979),.B(g17100));
  NOR2 NOR2_986(.VSS(VSS),.VDD(VDD),.Y(g26534),.A(g25321),.B(g8869));
  NOR2 NOR2_987(.VSS(VSS),.VDD(VDD),.Y(g26541),.A(g13755),.B(g25269));
  NOR2 NOR2_988(.VSS(VSS),.VDD(VDD),.Y(g26545),.A(g13790),.B(g25277));
  NOR2 NOR2_989(.VSS(VSS),.VDD(VDD),.Y(g26547),.A(g13796),.B(g25278));
  NOR2 NOR2_990(.VSS(VSS),.VDD(VDD),.Y(g26553),.A(g13816),.B(g25282));
  NOR2 NOR2_991(.VSS(VSS),.VDD(VDD),.Y(g26557),.A(g13818),.B(g25286));
  NOR2 NOR2_992(.VSS(VSS),.VDD(VDD),.Y(g26559),.A(g13824),.B(g25287));
  NOR2 NOR2_993(.VSS(VSS),.VDD(VDD),.Y(g26560),.A(g25281),.B(g24559));
  NOR2 NOR2_994(.VSS(VSS),.VDD(VDD),.Y(g26569),.A(g13837),.B(g25290));
  NOR2 NOR2_995(.VSS(VSS),.VDD(VDD),.Y(g26573),.A(g13839),.B(g25294));
  NOR2 NOR2_996(.VSS(VSS),.VDD(VDD),.Y(g26575),.A(g13845),.B(g25295));
  NOR2 NOR2_997(.VSS(VSS),.VDD(VDD),.Y(g26583),.A(g25289),.B(g24569));
  NOR2 NOR2_998(.VSS(VSS),.VDD(VDD),.Y(g26592),.A(g13851),.B(g25300));
  NOR2 NOR2_999(.VSS(VSS),.VDD(VDD),.Y(g26596),.A(g13853),.B(g25304));
  NOR2 NOR2_1000(.VSS(VSS),.VDD(VDD),.Y(g26607),.A(g25299),.B(g24578));
  NOR2 NOR2_1001(.VSS(VSS),.VDD(VDD),.Y(g26616),.A(g13860),.B(g25310));
  NOR2 NOR2_1002(.VSS(VSS),.VDD(VDD),.Y(g26630),.A(g25309),.B(g24585));
  NOR2 NOR2_1003(.VSS(VSS),.VDD(VDD),.Y(g26655),.A(g25328),.B(g17084));
  NOR2 NOR2_1004(.VSS(VSS),.VDD(VDD),.Y(g26659),.A(g25334),.B(g17116));
  NOR2 NOR2_1005(.VSS(VSS),.VDD(VDD),.Y(g26660),.A(g25208),.B(g10024));
  NOR2 NOR2_1006(.VSS(VSS),.VDD(VDD),.Y(g26661),.A(g25337),.B(g17122));
  NOR2 NOR2_1007(.VSS(VSS),.VDD(VDD),.Y(g26664),.A(g25346),.B(g17138));
  NOR2 NOR2_1008(.VSS(VSS),.VDD(VDD),.Y(g26665),.A(g25348),.B(g17143));
  NOR2 NOR2_1009(.VSS(VSS),.VDD(VDD),.Y(g26666),.A(g25216),.B(g10133));
  NOR2 NOR2_1010(.VSS(VSS),.VDD(VDD),.Y(g26667),.A(g25351),.B(g17149));
  NOR2 NOR2_1011(.VSS(VSS),.VDD(VDD),.Y(g26669),.A(g25360),.B(g17161));
  NOR2 NOR2_1012(.VSS(VSS),.VDD(VDD),.Y(g26670),.A(g25362),.B(g17166));
  NOR2 NOR2_1013(.VSS(VSS),.VDD(VDD),.Y(g26671),.A(g25226),.B(g10238));
  NOR2 NOR2_1014(.VSS(VSS),.VDD(VDD),.Y(g26672),.A(g25365),.B(g17172));
  NOR2 NOR2_1015(.VSS(VSS),.VDD(VDD),.Y(g26675),.A(g25375),.B(g17176));
  NOR2 NOR2_1016(.VSS(VSS),.VDD(VDD),.Y(g26676),.A(g25377),.B(g17181));
  NOR2 NOR2_1017(.VSS(VSS),.VDD(VDD),.Y(g26677),.A(g25238),.B(g10340));
  NOR2 NOR2_1018(.VSS(VSS),.VDD(VDD),.Y(g26776),.A(g26042),.B(g10024));
  NOR2 NOR2_1019(.VSS(VSS),.VDD(VDD),.Y(g26781),.A(g26044),.B(g10133));
  NOR2 NOR2_1020(.VSS(VSS),.VDD(VDD),.Y(g26786),.A(g26049),.B(g22777));
  NOR2 NOR2_1021(.VSS(VSS),.VDD(VDD),.Y(g26789),.A(g26046),.B(g10238));
  NOR2 NOR2_1022(.VSS(VSS),.VDD(VDD),.Y(g26795),.A(g26050),.B(g10340));
  NOR2 NOR2_1023(.VSS(VSS),.VDD(VDD),.Y(g26798),.A(g26055),.B(g18407));
  NOR2 NOR2_1024(.VSS(VSS),.VDD(VDD),.Y(g26799),.A(g26158),.B(g25453));
  NOR2 NOR2_1025(.VSS(VSS),.VDD(VDD),.Y(g26800),.A(g26163),.B(g25457));
  NOR2 NOR2_1026(.VSS(VSS),.VDD(VDD),.Y(g26801),.A(g26171),.B(g25461));
  NOR2 NOR2_1027(.VSS(VSS),.VDD(VDD),.Y(g26802),.A(g26188),.B(g25466));
  NOR2 NOR2_1028(.VSS(VSS),.VDD(VDD),.Y(g26803),.A(g15105),.B(g26213));
  NOR2 NOR2_1029(.VSS(VSS),.VDD(VDD),.Y(g26804),.A(g15172),.B(g26235));
  NOR2 NOR2_1030(.VSS(VSS),.VDD(VDD),.Y(g26805),.A(g15173),.B(g26236));
  NOR2 NOR2_1031(.VSS(VSS),.VDD(VDD),.Y(g26806),.A(g15197),.B(g26244));
  NOR2 NOR2_1032(.VSS(VSS),.VDD(VDD),.Y(g26807),.A(g15245),.B(g26261));
  NOR2 NOR2_1033(.VSS(VSS),.VDD(VDD),.Y(g26808),.A(g15246),.B(g26262));
  NOR2 NOR2_1034(.VSS(VSS),.VDD(VDD),.Y(g26809),.A(g15258),.B(g26270));
  NOR2 NOR2_1035(.VSS(VSS),.VDD(VDD),.Y(g26810),.A(g15259),.B(g26271));
  NOR2 NOR2_1036(.VSS(VSS),.VDD(VDD),.Y(g26811),.A(g15283),.B(g26279));
  NOR2 NOR2_1037(.VSS(VSS),.VDD(VDD),.Y(g26812),.A(g15321),.B(g26291));
  NOR2 NOR2_1038(.VSS(VSS),.VDD(VDD),.Y(g26813),.A(g15337),.B(g26302));
  NOR2 NOR2_1039(.VSS(VSS),.VDD(VDD),.Y(g26814),.A(g15338),.B(g26303));
  NOR2 NOR2_1040(.VSS(VSS),.VDD(VDD),.Y(g26815),.A(g15350),.B(g26311));
  NOR2 NOR2_1041(.VSS(VSS),.VDD(VDD),.Y(g26816),.A(g15351),.B(g26312));
  NOR2 NOR2_1042(.VSS(VSS),.VDD(VDD),.Y(g26817),.A(g15375),.B(g26317));
  NOR2 NOR2_1043(.VSS(VSS),.VDD(VDD),.Y(g26818),.A(g15407),.B(g26335));
  NOR2 NOR2_1044(.VSS(VSS),.VDD(VDD),.Y(g26820),.A(g15423),.B(g26346));
  NOR2 NOR2_1045(.VSS(VSS),.VDD(VDD),.Y(g26821),.A(g15424),.B(g26347));
  NOR2 NOR2_1046(.VSS(VSS),.VDD(VDD),.Y(g26822),.A(g15436),.B(g26352));
  NOR2 NOR2_1047(.VSS(VSS),.VDD(VDD),.Y(g26823),.A(g15437),.B(g26353));
  NOR2 NOR2_1048(.VSS(VSS),.VDD(VDD),.Y(g26824),.A(g15491),.B(g26382));
  NOR2 NOR2_1049(.VSS(VSS),.VDD(VDD),.Y(g26825),.A(g15507),.B(g26390));
  NOR2 NOR2_1050(.VSS(VSS),.VDD(VDD),.Y(g26826),.A(g15508),.B(g26391));
  NOR2 NOR2_1051(.VSS(VSS),.VDD(VDD),.Y(g26827),.A(g15577),.B(g26425));
  NOR2 NOR2_1052(.VSS(VSS),.VDD(VDD),.Y(g26869),.A(g26458),.B(g5642));
  NOR2 NOR2_1053(.VSS(VSS),.VDD(VDD),.Y(g26873),.A(g25483),.B(g26260));
  NOR2 NOR2_1054(.VSS(VSS),.VDD(VDD),.Y(g26877),.A(g26140),.B(g22319));
  NOR2 NOR2_1055(.VSS(VSS),.VDD(VDD),.Y(g26878),.A(g26482),.B(g5680));
  NOR2 NOR2_1056(.VSS(VSS),.VDD(VDD),.Y(g26882),.A(g25514),.B(g26301));
  NOR2 NOR2_1057(.VSS(VSS),.VDD(VDD),.Y(g26885),.A(g26140),.B(g22319));
  NOR2 NOR2_1058(.VSS(VSS),.VDD(VDD),.Y(g26887),.A(g26498),.B(g5732));
  NOR2 NOR2_1059(.VSS(VSS),.VDD(VDD),.Y(g26891),.A(g25561),.B(g26345));
  NOR2 NOR2_1060(.VSS(VSS),.VDD(VDD),.Y(g26897),.A(g26513),.B(g5790));
  NOR2 NOR2_1061(.VSS(VSS),.VDD(VDD),.Y(g26901),.A(g25627),.B(g26389));
  NOR2 NOR2_1062(.VSS(VSS),.VDD(VDD),.Y(g26905),.A(g26096),.B(g22319));
  NOR2 NOR2_1063(.VSS(VSS),.VDD(VDD),.Y(g26914),.A(g26107),.B(g22319));
  NOR2 NOR2_1064(.VSS(VSS),.VDD(VDD),.Y(g26988),.A(g24893),.B(g26023));
  NOR2 NOR2_1065(.VSS(VSS),.VDD(VDD),.Y(g26989),.A(g26663),.B(g21913));
  NOR2 NOR2_1066(.VSS(VSS),.VDD(VDD),.Y(g27011),.A(g24916),.B(g26026));
  NOR2 NOR2_1067(.VSS(VSS),.VDD(VDD),.Y(g27012),.A(g26668),.B(g21931));
  NOR2 NOR2_1068(.VSS(VSS),.VDD(VDD),.Y(g27037),.A(g24933),.B(g26028));
  NOR2 NOR2_1069(.VSS(VSS),.VDD(VDD),.Y(g27038),.A(g26674),.B(g20640));
  NOR2 NOR2_1070(.VSS(VSS),.VDD(VDD),.Y(g27051),.A(g4456),.B(g26081));
  NOR2 NOR2_1071(.VSS(VSS),.VDD(VDD),.Y(g27065),.A(g24945),.B(g26029));
  NOR2 NOR2_1072(.VSS(VSS),.VDD(VDD),.Y(g27066),.A(g26024),.B(g20665));
  NOR2 NOR2_1073(.VSS(VSS),.VDD(VDD),.Y(g27078),.A(g4632),.B(g26084));
  NOR2 NOR2_1074(.VSS(VSS),.VDD(VDD),.Y(g27094),.A(g4809),.B(g26090));
  NOR2 NOR2_1075(.VSS(VSS),.VDD(VDD),.Y(g27106),.A(g4985),.B(g26103));
  NOR2 NOR2_1076(.VSS(VSS),.VDD(VDD),.Y(g27120),.A(g26560),.B(g17001));
  NOR2 NOR2_1077(.VSS(VSS),.VDD(VDD),.Y(g27123),.A(g26583),.B(g17031));
  NOR2 NOR2_1078(.VSS(VSS),.VDD(VDD),.Y(g27129),.A(g26607),.B(g17065));
  NOR2 NOR2_1079(.VSS(VSS),.VDD(VDD),.Y(g27131),.A(g26630),.B(g17100));
  NOR2 NOR2_1080(.VSS(VSS),.VDD(VDD),.Y(g27144),.A(g23451),.B(g26052));
  NOR2 NOR2_1081(.VSS(VSS),.VDD(VDD),.Y(g27147),.A(g23458),.B(g26054));
  NOR2 NOR2_1082(.VSS(VSS),.VDD(VDD),.Y(g27149),.A(g23462),.B(g26060));
  NOR2 NOR2_1083(.VSS(VSS),.VDD(VDD),.Y(g27152),.A(g23467),.B(g26062));
  NOR2 NOR2_1084(.VSS(VSS),.VDD(VDD),.Y(g27157),.A(g23471),.B(g26067));
  NOR2 NOR2_1085(.VSS(VSS),.VDD(VDD),.Y(g27160),.A(g23476),.B(g26069));
  NOR2 NOR2_1086(.VSS(VSS),.VDD(VDD),.Y(g27165),.A(g23484),.B(g26074));
  NOR2 NOR2_1087(.VSS(VSS),.VDD(VDD),.Y(g27174),.A(g23494),.B(g26080));
  NOR2 NOR2_1088(.VSS(VSS),.VDD(VDD),.Y(g27175),.A(g26075),.B(g25342));
  NOR2 NOR2_1089(.VSS(VSS),.VDD(VDD),.Y(g27179),.A(g26082),.B(g25356));
  NOR2 NOR2_1090(.VSS(VSS),.VDD(VDD),.Y(g27184),.A(g26085),.B(g25371));
  NOR2 NOR2_1091(.VSS(VSS),.VDD(VDD),.Y(g27188),.A(g26091),.B(g25388));
  NOR2 NOR2_1092(.VSS(VSS),.VDD(VDD),.Y(g27243),.A(g26802),.B(g10340));
  NOR2 NOR2_1093(.VSS(VSS),.VDD(VDD),.Y(g27250),.A(g26955),.B(g26166));
  NOR2 NOR2_1094(.VSS(VSS),.VDD(VDD),.Y(g27251),.A(g26958),.B(g26186));
  NOR2 NOR2_1095(.VSS(VSS),.VDD(VDD),.Y(g27252),.A(g26963),.B(g26207));
  NOR2 NOR2_1096(.VSS(VSS),.VDD(VDD),.Y(g27253),.A(g26965),.B(g26212));
  NOR2 NOR2_1097(.VSS(VSS),.VDD(VDD),.Y(g27254),.A(g26968),.B(g26231));
  NOR2 NOR2_1098(.VSS(VSS),.VDD(VDD),.Y(g27255),.A(g26969),.B(g26233));
  NOR2 NOR2_1099(.VSS(VSS),.VDD(VDD),.Y(g27256),.A(g26970),.B(g26234));
  NOR2 NOR2_1100(.VSS(VSS),.VDD(VDD),.Y(g27257),.A(g26971),.B(g26243));
  NOR2 NOR2_1101(.VSS(VSS),.VDD(VDD),.Y(g27258),.A(g26977),.B(g26257));
  NOR2 NOR2_1102(.VSS(VSS),.VDD(VDD),.Y(g27259),.A(g26978),.B(g26258));
  NOR2 NOR2_1103(.VSS(VSS),.VDD(VDD),.Y(g27260),.A(g26979),.B(g26259));
  NOR2 NOR2_1104(.VSS(VSS),.VDD(VDD),.Y(g27261),.A(g26980),.B(g26263));
  NOR2 NOR2_1105(.VSS(VSS),.VDD(VDD),.Y(g27262),.A(g26981),.B(g26268));
  NOR2 NOR2_1106(.VSS(VSS),.VDD(VDD),.Y(g27263),.A(g26982),.B(g26269));
  NOR2 NOR2_1107(.VSS(VSS),.VDD(VDD),.Y(g27264),.A(g26984),.B(g26278));
  NOR2 NOR2_1108(.VSS(VSS),.VDD(VDD),.Y(g27265),.A(g26993),.B(g26288));
  NOR2 NOR2_1109(.VSS(VSS),.VDD(VDD),.Y(g27266),.A(g26994),.B(g26289));
  NOR2 NOR2_1110(.VSS(VSS),.VDD(VDD),.Y(g27267),.A(g26995),.B(g26290));
  NOR2 NOR2_1111(.VSS(VSS),.VDD(VDD),.Y(g27268),.A(g26996),.B(g26292));
  NOR2 NOR2_1112(.VSS(VSS),.VDD(VDD),.Y(g27269),.A(g26997),.B(g26293));
  NOR2 NOR2_1113(.VSS(VSS),.VDD(VDD),.Y(g27270),.A(g26998),.B(g26298));
  NOR2 NOR2_1114(.VSS(VSS),.VDD(VDD),.Y(g27271),.A(g26999),.B(g26299));
  NOR2 NOR2_1115(.VSS(VSS),.VDD(VDD),.Y(g27272),.A(g27000),.B(g26300));
  NOR2 NOR2_1116(.VSS(VSS),.VDD(VDD),.Y(g27273),.A(g27001),.B(g26307));
  NOR2 NOR2_1117(.VSS(VSS),.VDD(VDD),.Y(g27274),.A(g27002),.B(g26309));
  NOR2 NOR2_1118(.VSS(VSS),.VDD(VDD),.Y(g27275),.A(g27003),.B(g26310));
  NOR2 NOR2_1119(.VSS(VSS),.VDD(VDD),.Y(g27276),.A(g27004),.B(g26316));
  NOR2 NOR2_1120(.VSS(VSS),.VDD(VDD),.Y(g27277),.A(g27005),.B(g26318));
  NOR2 NOR2_1121(.VSS(VSS),.VDD(VDD),.Y(g27278),.A(g27006),.B(g26319));
  NOR2 NOR2_1122(.VSS(VSS),.VDD(VDD),.Y(g27279),.A(g27007),.B(g26324));
  NOR2 NOR2_1123(.VSS(VSS),.VDD(VDD),.Y(g27280),.A(g27008),.B(g26325));
  NOR2 NOR2_1124(.VSS(VSS),.VDD(VDD),.Y(g27281),.A(g27009),.B(g26326));
  NOR2 NOR2_1125(.VSS(VSS),.VDD(VDD),.Y(g27282),.A(g27016),.B(g26332));
  NOR2 NOR2_1126(.VSS(VSS),.VDD(VDD),.Y(g27283),.A(g27017),.B(g26333));
  NOR2 NOR2_1127(.VSS(VSS),.VDD(VDD),.Y(g27284),.A(g27018),.B(g26334));
  NOR2 NOR2_1128(.VSS(VSS),.VDD(VDD),.Y(g27285),.A(g27019),.B(g26339));
  NOR2 NOR2_1129(.VSS(VSS),.VDD(VDD),.Y(g27286),.A(g27020),.B(g26340));
  NOR2 NOR2_1130(.VSS(VSS),.VDD(VDD),.Y(g27287),.A(g27021),.B(g26342));
  NOR2 NOR2_1131(.VSS(VSS),.VDD(VDD),.Y(g27288),.A(g27022),.B(g26343));
  NOR2 NOR2_1132(.VSS(VSS),.VDD(VDD),.Y(g27289),.A(g27023),.B(g26344));
  NOR2 NOR2_1133(.VSS(VSS),.VDD(VDD),.Y(g27290),.A(g27024),.B(g26348));
  NOR2 NOR2_1134(.VSS(VSS),.VDD(VDD),.Y(g27291),.A(g27025),.B(g26350));
  NOR2 NOR2_1135(.VSS(VSS),.VDD(VDD),.Y(g27292),.A(g27026),.B(g26351));
  NOR2 NOR2_1136(.VSS(VSS),.VDD(VDD),.Y(g27293),.A(g27027),.B(g26357));
  NOR2 NOR2_1137(.VSS(VSS),.VDD(VDD),.Y(g27294),.A(g27028),.B(g26361));
  NOR2 NOR2_1138(.VSS(VSS),.VDD(VDD),.Y(g27295),.A(g27029),.B(g26362));
  NOR2 NOR2_1139(.VSS(VSS),.VDD(VDD),.Y(g27296),.A(g27030),.B(g26363));
  NOR2 NOR2_1140(.VSS(VSS),.VDD(VDD),.Y(g27297),.A(g27031),.B(g26365));
  NOR2 NOR2_1141(.VSS(VSS),.VDD(VDD),.Y(g27298),.A(g27032),.B(g26366));
  NOR2 NOR2_1142(.VSS(VSS),.VDD(VDD),.Y(g27299),.A(g27033),.B(g26371));
  NOR2 NOR2_1143(.VSS(VSS),.VDD(VDD),.Y(g27300),.A(g27034),.B(g26372));
  NOR2 NOR2_1144(.VSS(VSS),.VDD(VDD),.Y(g27301),.A(g27035),.B(g26373));
  NOR2 NOR2_1145(.VSS(VSS),.VDD(VDD),.Y(g27302),.A(g27042),.B(g26379));
  NOR2 NOR2_1146(.VSS(VSS),.VDD(VDD),.Y(g27303),.A(g27043),.B(g26380));
  NOR2 NOR2_1147(.VSS(VSS),.VDD(VDD),.Y(g27304),.A(g27044),.B(g26381));
  NOR2 NOR2_1148(.VSS(VSS),.VDD(VDD),.Y(g27305),.A(g27045),.B(g26383));
  NOR2 NOR2_1149(.VSS(VSS),.VDD(VDD),.Y(g27306),.A(g27046),.B(g26384));
  NOR2 NOR2_1150(.VSS(VSS),.VDD(VDD),.Y(g27307),.A(g27047),.B(g26386));
  NOR2 NOR2_1151(.VSS(VSS),.VDD(VDD),.Y(g27308),.A(g27048),.B(g26387));
  NOR2 NOR2_1152(.VSS(VSS),.VDD(VDD),.Y(g27309),.A(g27049),.B(g26388));
  NOR2 NOR2_1153(.VSS(VSS),.VDD(VDD),.Y(g27310),.A(g27050),.B(g26392));
  NOR2 NOR2_1154(.VSS(VSS),.VDD(VDD),.Y(g27311),.A(g27053),.B(g26396));
  NOR2 NOR2_1155(.VSS(VSS),.VDD(VDD),.Y(g27312),.A(g27054),.B(g26397));
  NOR2 NOR2_1156(.VSS(VSS),.VDD(VDD),.Y(g27313),.A(g27055),.B(g26400));
  NOR2 NOR2_1157(.VSS(VSS),.VDD(VDD),.Y(g27314),.A(g27056),.B(g26404));
  NOR2 NOR2_1158(.VSS(VSS),.VDD(VDD),.Y(g27315),.A(g27057),.B(g26405));
  NOR2 NOR2_1159(.VSS(VSS),.VDD(VDD),.Y(g27316),.A(g27058),.B(g26406));
  NOR2 NOR2_1160(.VSS(VSS),.VDD(VDD),.Y(g27317),.A(g27059),.B(g26408));
  NOR2 NOR2_1161(.VSS(VSS),.VDD(VDD),.Y(g27318),.A(g27060),.B(g26409));
  NOR2 NOR2_1162(.VSS(VSS),.VDD(VDD),.Y(g27319),.A(g27061),.B(g26414));
  NOR2 NOR2_1163(.VSS(VSS),.VDD(VDD),.Y(g27320),.A(g27062),.B(g26415));
  NOR2 NOR2_1164(.VSS(VSS),.VDD(VDD),.Y(g27321),.A(g27063),.B(g26416));
  NOR2 NOR2_1165(.VSS(VSS),.VDD(VDD),.Y(g27322),.A(g27070),.B(g26422));
  NOR2 NOR2_1166(.VSS(VSS),.VDD(VDD),.Y(g27323),.A(g27071),.B(g26423));
  NOR2 NOR2_1167(.VSS(VSS),.VDD(VDD),.Y(g27324),.A(g27072),.B(g26424));
  NOR2 NOR2_1168(.VSS(VSS),.VDD(VDD),.Y(g27325),.A(g27073),.B(g26426));
  NOR2 NOR2_1169(.VSS(VSS),.VDD(VDD),.Y(g27326),.A(g27074),.B(g26427));
  NOR2 NOR2_1170(.VSS(VSS),.VDD(VDD),.Y(g27327),.A(g27077),.B(g26432));
  NOR2 NOR2_1171(.VSS(VSS),.VDD(VDD),.Y(g27328),.A(g27080),.B(g26437));
  NOR2 NOR2_1172(.VSS(VSS),.VDD(VDD),.Y(g27329),.A(g27081),.B(g26438));
  NOR2 NOR2_1173(.VSS(VSS),.VDD(VDD),.Y(g27330),.A(g27082),.B(g26441));
  NOR2 NOR2_1174(.VSS(VSS),.VDD(VDD),.Y(g27331),.A(g27083),.B(g26445));
  NOR2 NOR2_1175(.VSS(VSS),.VDD(VDD),.Y(g27332),.A(g27084),.B(g26446));
  NOR2 NOR2_1176(.VSS(VSS),.VDD(VDD),.Y(g27333),.A(g27085),.B(g26447));
  NOR2 NOR2_1177(.VSS(VSS),.VDD(VDD),.Y(g27334),.A(g27086),.B(g26449));
  NOR2 NOR2_1178(.VSS(VSS),.VDD(VDD),.Y(g27335),.A(g27087),.B(g26450));
  NOR2 NOR2_1179(.VSS(VSS),.VDD(VDD),.Y(g27336),.A(g27088),.B(g26455));
  NOR2 NOR2_1180(.VSS(VSS),.VDD(VDD),.Y(g27337),.A(g27089),.B(g26456));
  NOR2 NOR2_1181(.VSS(VSS),.VDD(VDD),.Y(g27338),.A(g27090),.B(g26457));
  NOR2 NOR2_1182(.VSS(VSS),.VDD(VDD),.Y(g27339),.A(g27093),.B(g26464));
  NOR2 NOR2_1183(.VSS(VSS),.VDD(VDD),.Y(g27340),.A(g27096),.B(g26469));
  NOR2 NOR2_1184(.VSS(VSS),.VDD(VDD),.Y(g27341),.A(g27097),.B(g26470));
  NOR2 NOR2_1185(.VSS(VSS),.VDD(VDD),.Y(g27342),.A(g27098),.B(g26473));
  NOR2 NOR2_1186(.VSS(VSS),.VDD(VDD),.Y(g27343),.A(g27099),.B(g26477));
  NOR2 NOR2_1187(.VSS(VSS),.VDD(VDD),.Y(g27344),.A(g27100),.B(g26478));
  NOR2 NOR2_1188(.VSS(VSS),.VDD(VDD),.Y(g27345),.A(g27101),.B(g26479));
  NOR2 NOR2_1189(.VSS(VSS),.VDD(VDD),.Y(g27346),.A(g27105),.B(g26488));
  NOR2 NOR2_1190(.VSS(VSS),.VDD(VDD),.Y(g27347),.A(g27108),.B(g26493));
  NOR2 NOR2_1191(.VSS(VSS),.VDD(VDD),.Y(g27348),.A(g27109),.B(g26494));
  NOR2 NOR2_1192(.VSS(VSS),.VDD(VDD),.Y(g27354),.A(g27112),.B(g26504));
  NOR2 NOR2_1193(.VSS(VSS),.VDD(VDD),.Y(g27414),.A(g26770),.B(g25187));
  NOR3 NOR3_379(.VSS(VSS),.VDD(VDD),.Y(g27415),.A(g23104),.B(g27181),.C(g25128));
  NOR2 NOR2_1194(.VSS(VSS),.VDD(VDD),.Y(g27435),.A(g26777),.B(g25193));
  NOR3 NOR3_380(.VSS(VSS),.VDD(VDD),.Y(g27436),.A(g23118),.B(g27187),.C(g24427));
  NOR2 NOR2_1195(.VSS(VSS),.VDD(VDD),.Y(g27450),.A(g26902),.B(g24613));
  NOR2 NOR2_1196(.VSS(VSS),.VDD(VDD),.Y(g27454),.A(g26783),.B(g25196));
  NOR3 NOR3_381(.VSS(VSS),.VDD(VDD),.Y(g27455),.A(g23127),.B(g26758),.C(g24431));
  NOR2 NOR2_1197(.VSS(VSS),.VDD(VDD),.Y(g27462),.A(g26892),.B(g24622));
  NOR2 NOR2_1198(.VSS(VSS),.VDD(VDD),.Y(g27464),.A(g27178),.B(g25975));
  NOR2 NOR2_1199(.VSS(VSS),.VDD(VDD),.Y(g27466),.A(g26915),.B(g24624));
  NOR2 NOR2_1200(.VSS(VSS),.VDD(VDD),.Y(g27470),.A(g26790),.B(g25198));
  NOR3 NOR3_382(.VSS(VSS),.VDD(VDD),.Y(g27471),.A(g23138),.B(g26764),.C(g24435));
  NOR2 NOR2_1201(.VSS(VSS),.VDD(VDD),.Y(g27478),.A(g26754),.B(g24432));
  NOR2 NOR2_1202(.VSS(VSS),.VDD(VDD),.Y(g27481),.A(g27182),.B(g25980));
  NOR2 NOR2_1203(.VSS(VSS),.VDD(VDD),.Y(g27482),.A(g26906),.B(g24637));
  NOR2 NOR2_1204(.VSS(VSS),.VDD(VDD),.Y(g27485),.A(g26928),.B(g24638));
  NOR3 NOR3_383(.VSS(VSS),.VDD(VDD),.Y(g27492),.A(g24958),.B(g24633),.C(g26771));
  NOR2 NOR2_1205(.VSS(VSS),.VDD(VDD),.Y(g27496),.A(g27185),.B(g25178));
  NOR2 NOR2_1206(.VSS(VSS),.VDD(VDD),.Y(g27501),.A(g26763),.B(g24436));
  NOR2 NOR2_1207(.VSS(VSS),.VDD(VDD),.Y(g27504),.A(g26918),.B(g24656));
  NOR2 NOR2_1208(.VSS(VSS),.VDD(VDD),.Y(g27507),.A(g26941),.B(g24657));
  NOR3 NOR3_384(.VSS(VSS),.VDD(VDD),.Y(g27513),.A(g24969),.B(g24653),.C(g26778));
  NOR2 NOR2_1209(.VSS(VSS),.VDD(VDD),.Y(g27521),.A(g26766),.B(g24439));
  NOR2 NOR2_1210(.VSS(VSS),.VDD(VDD),.Y(g27524),.A(g26931),.B(g24675));
  NOR2 NOR2_1211(.VSS(VSS),.VDD(VDD),.Y(g27527),.A(g26759),.B(g19087));
  NOR2 NOR2_1212(.VSS(VSS),.VDD(VDD),.Y(g27529),.A(g4456),.B(g26873));
  NOR2 NOR2_1213(.VSS(VSS),.VDD(VDD),.Y(g27531),.A(g26760),.B(g25181));
  NOR2 NOR2_1214(.VSS(VSS),.VDD(VDD),.Y(g27532),.A(g26761),.B(g25182));
  NOR3 NOR3_385(.VSS(VSS),.VDD(VDD),.Y(g27538),.A(g24982),.B(g24672),.C(g26784));
  NOR2 NOR2_1215(.VSS(VSS),.VDD(VDD),.Y(g27546),.A(g26769),.B(g24441));
  NOR2 NOR2_1216(.VSS(VSS),.VDD(VDD),.Y(g27549),.A(g26765),.B(g19093));
  NOR2 NOR2_1217(.VSS(VSS),.VDD(VDD),.Y(g27551),.A(g4632),.B(g26882));
  NOR3 NOR3_386(.VSS(VSS),.VDD(VDD),.Y(g27558),.A(g24993),.B(g24691),.C(g26791));
  NOR2 NOR2_1218(.VSS(VSS),.VDD(VDD),.Y(g27563),.A(g26922),.B(g24708));
  NOR2 NOR2_1219(.VSS(VSS),.VDD(VDD),.Y(g27564),.A(g26767),.B(g25184));
  NOR2 NOR2_1220(.VSS(VSS),.VDD(VDD),.Y(g27565),.A(g26768),.B(g19100));
  NOR2 NOR2_1221(.VSS(VSS),.VDD(VDD),.Y(g27567),.A(g4809),.B(g26891));
  NOR2 NOR2_1222(.VSS(VSS),.VDD(VDD),.Y(g27572),.A(g26911),.B(g24717));
  NOR2 NOR2_1223(.VSS(VSS),.VDD(VDD),.Y(g27573),.A(g26773),.B(g25188));
  NOR2 NOR2_1224(.VSS(VSS),.VDD(VDD),.Y(g27574),.A(g26935),.B(g24720));
  NOR2 NOR2_1225(.VSS(VSS),.VDD(VDD),.Y(g27575),.A(g26774),.B(g19107));
  NOR2 NOR2_1226(.VSS(VSS),.VDD(VDD),.Y(g27577),.A(g4985),.B(g26901));
  NOR2 NOR2_1227(.VSS(VSS),.VDD(VDD),.Y(g27579),.A(g26775),.B(g25192));
  NOR2 NOR2_1228(.VSS(VSS),.VDD(VDD),.Y(g27581),.A(g26925),.B(g24728));
  NOR2 NOR2_1229(.VSS(VSS),.VDD(VDD),.Y(g27582),.A(g26944),.B(g24731));
  NOR2 NOR2_1230(.VSS(VSS),.VDD(VDD),.Y(g27584),.A(g26938),.B(g24736));
  NOR2 NOR2_1231(.VSS(VSS),.VDD(VDD),.Y(g27585),.A(g26950),.B(g24739));
  NOR2 NOR2_1232(.VSS(VSS),.VDD(VDD),.Y(g27588),.A(g26947),.B(g24742));
  NOR2 NOR2_1233(.VSS(VSS),.VDD(VDD),.Y(g27594),.A(g27175),.B(g17001));
  NOR2 NOR2_1234(.VSS(VSS),.VDD(VDD),.Y(g27603),.A(g27179),.B(g17031));
  NOR2 NOR2_1235(.VSS(VSS),.VDD(VDD),.Y(g27612),.A(g27184),.B(g17065));
  NOR2 NOR2_1236(.VSS(VSS),.VDD(VDD),.Y(g27621),.A(g27188),.B(g17100));
  NOR2 NOR2_1237(.VSS(VSS),.VDD(VDD),.Y(g27629),.A(g26829),.B(g26051));
  NOR2 NOR2_1238(.VSS(VSS),.VDD(VDD),.Y(g27631),.A(g26833),.B(g26053));
  NOR2 NOR2_1239(.VSS(VSS),.VDD(VDD),.Y(g27655),.A(g26842),.B(g26061));
  NOR2 NOR2_1240(.VSS(VSS),.VDD(VDD),.Y(g27658),.A(g26851),.B(g26068));
  NOR2 NOR2_1241(.VSS(VSS),.VDD(VDD),.Y(g27672),.A(g26799),.B(g10024));
  NOR2 NOR2_1242(.VSS(VSS),.VDD(VDD),.Y(g27678),.A(g26800),.B(g10133));
  NOR2 NOR2_1243(.VSS(VSS),.VDD(VDD),.Y(g27682),.A(g26801),.B(g10238));
  NOR2 NOR2_1244(.VSS(VSS),.VDD(VDD),.Y(g27718),.A(g27251),.B(g10133));
  NOR2 NOR2_1245(.VSS(VSS),.VDD(VDD),.Y(g27722),.A(g27252),.B(g10238));
  NOR2 NOR2_1246(.VSS(VSS),.VDD(VDD),.Y(g27724),.A(g27254),.B(g10340));
  NOR2 NOR2_1247(.VSS(VSS),.VDD(VDD),.Y(g27735),.A(g27394),.B(g26961));
  NOR2 NOR2_1248(.VSS(VSS),.VDD(VDD),.Y(g27736),.A(g27396),.B(g26962));
  NOR2 NOR2_1249(.VSS(VSS),.VDD(VDD),.Y(g27741),.A(g27407),.B(g26966));
  NOR2 NOR2_1250(.VSS(VSS),.VDD(VDD),.Y(g27742),.A(g27409),.B(g26967));
  NOR2 NOR2_1251(.VSS(VSS),.VDD(VDD),.Y(g27746),.A(g27425),.B(g26972));
  NOR2 NOR2_1252(.VSS(VSS),.VDD(VDD),.Y(g27747),.A(g27427),.B(g26973));
  NOR2 NOR2_1253(.VSS(VSS),.VDD(VDD),.Y(g27754),.A(g27446),.B(g26985));
  NOR2 NOR2_1254(.VSS(VSS),.VDD(VDD),.Y(g27755),.A(g27448),.B(g26986));
  NOR2 NOR2_1255(.VSS(VSS),.VDD(VDD),.Y(g27759),.A(g27495),.B(g27052));
  NOR2 NOR2_1256(.VSS(VSS),.VDD(VDD),.Y(g27760),.A(g27509),.B(g27076));
  NOR2 NOR2_1257(.VSS(VSS),.VDD(VDD),.Y(g27761),.A(g27516),.B(g27079));
  NOR2 NOR2_1258(.VSS(VSS),.VDD(VDD),.Y(g27762),.A(g27530),.B(g27091));
  NOR2 NOR2_1259(.VSS(VSS),.VDD(VDD),.Y(g27763),.A(g27534),.B(g27092));
  NOR2 NOR2_1260(.VSS(VSS),.VDD(VDD),.Y(g27764),.A(g27541),.B(g27095));
  NOR2 NOR2_1261(.VSS(VSS),.VDD(VDD),.Y(g27765),.A(g27552),.B(g27103));
  NOR2 NOR2_1262(.VSS(VSS),.VDD(VDD),.Y(g27766),.A(g27554),.B(g27104));
  NOR2 NOR2_1263(.VSS(VSS),.VDD(VDD),.Y(g27767),.A(g27561),.B(g27107));
  NOR2 NOR2_1264(.VSS(VSS),.VDD(VDD),.Y(g27768),.A(g27568),.B(g27110));
  NOR2 NOR2_1265(.VSS(VSS),.VDD(VDD),.Y(g27769),.A(g27570),.B(g27111));
  NOR2 NOR2_1266(.VSS(VSS),.VDD(VDD),.Y(g27771),.A(g27578),.B(g27115));
  NOR2 NOR2_1267(.VSS(VSS),.VDD(VDD),.Y(g27798),.A(g27632),.B(g1223));
  NOR3 NOR3_387(.VSS(VSS),.VDD(VDD),.Y(g27802),.A(g6087),.B(g27632),.C(g25330));
  NOR2 NOR2_1268(.VSS(VSS),.VDD(VDD),.Y(g27810),.A(g27632),.B(g1215));
  NOR3 NOR3_388(.VSS(VSS),.VDD(VDD),.Y(g27811),.A(g6087),.B(g27632),.C(g25404));
  NOR3 NOR3_389(.VSS(VSS),.VDD(VDD),.Y(g27814),.A(g6087),.B(g27632),.C(g25322));
  NOR2 NOR2_1269(.VSS(VSS),.VDD(VDD),.Y(g27823),.A(g27632),.B(g1216));
  NOR3 NOR3_390(.VSS(VSS),.VDD(VDD),.Y(g27824),.A(g6087),.B(g27632),.C(g25399));
  NOR3 NOR3_391(.VSS(VSS),.VDD(VDD),.Y(g27827),.A(g6087),.B(g27632),.C(g25314));
  NOR2 NOR2_1270(.VSS(VSS),.VDD(VDD),.Y(g27834),.A(g27478),.B(g14630));
  NOR2 NOR2_1271(.VSS(VSS),.VDD(VDD),.Y(g27842),.A(g27632),.B(g1217));
  NOR2 NOR2_1272(.VSS(VSS),.VDD(VDD),.Y(g27850),.A(g27501),.B(g14650));
  NOR2 NOR2_1273(.VSS(VSS),.VDD(VDD),.Y(g27854),.A(g27632),.B(g1218));
  NOR3 NOR3_392(.VSS(VSS),.VDD(VDD),.Y(g27855),.A(g6087),.B(g27632),.C(g25385));
  NOR2 NOR2_1274(.VSS(VSS),.VDD(VDD),.Y(g27864),.A(g27632),.B(g1219));
  NOR3 NOR3_393(.VSS(VSS),.VDD(VDD),.Y(g27865),.A(g6087),.B(g27632),.C(g25370));
  NOR2 NOR2_1275(.VSS(VSS),.VDD(VDD),.Y(g27868),.A(g23742),.B(g27632));
  NOR2 NOR2_1276(.VSS(VSS),.VDD(VDD),.Y(g27869),.A(g27632),.B(g25437));
  NOR2 NOR2_1277(.VSS(VSS),.VDD(VDD),.Y(g27875),.A(g27521),.B(g14677));
  NOR2 NOR2_1278(.VSS(VSS),.VDD(VDD),.Y(g27882),.A(g27632),.B(g1220));
  NOR3 NOR3_394(.VSS(VSS),.VDD(VDD),.Y(g27883),.A(g6087),.B(g27632),.C(g25361));
  NOR2 NOR2_1279(.VSS(VSS),.VDD(VDD),.Y(g27886),.A(g27632),.B(g24627));
  NOR2 NOR2_1280(.VSS(VSS),.VDD(VDD),.Y(g27892),.A(g27546),.B(g14711));
  NOR2 NOR2_1281(.VSS(VSS),.VDD(VDD),.Y(g27896),.A(g27632),.B(g1222));
  NOR3 NOR3_395(.VSS(VSS),.VDD(VDD),.Y(g27897),.A(g6087),.B(g27632),.C(g25349));
  NOR3 NOR3_396(.VSS(VSS),.VDD(VDD),.Y(g27900),.A(g6087),.B(g27632),.C(g25338));
  NOR2 NOR2_1282(.VSS(VSS),.VDD(VDD),.Y(g27906),.A(g16127),.B(g27656));
  NOR2 NOR2_1283(.VSS(VSS),.VDD(VDD),.Y(g27911),.A(g16170),.B(g27657));
  NOR2 NOR2_1284(.VSS(VSS),.VDD(VDD),.Y(g27916),.A(g16219),.B(g27659));
  NOR2 NOR2_1285(.VSS(VSS),.VDD(VDD),.Y(g27917),.A(g16220),.B(g27660));
  NOR2 NOR2_1286(.VSS(VSS),.VDD(VDD),.Y(g27925),.A(g16276),.B(g27661));
  NOR2 NOR2_1287(.VSS(VSS),.VDD(VDD),.Y(g27937),.A(g16321),.B(g27666));
  NOR2 NOR2_1288(.VSS(VSS),.VDD(VDD),.Y(g27950),.A(g16367),.B(g27673));
  NOR2 NOR2_1289(.VSS(VSS),.VDD(VDD),.Y(g27962),.A(g16394),.B(g27679));
  NOR2 NOR2_1290(.VSS(VSS),.VDD(VDD),.Y(g27964),.A(g16400),.B(g27680));
  NOR2 NOR2_1291(.VSS(VSS),.VDD(VDD),.Y(g27980),.A(g16428),.B(g27681));
  NOR2 NOR2_1292(.VSS(VSS),.VDD(VDD),.Y(g27997),.A(g16456),.B(g27242));
  NOR2 NOR2_1293(.VSS(VSS),.VDD(VDD),.Y(g28002),.A(g26032),.B(g27246));
  NOR2 NOR2_1294(.VSS(VSS),.VDD(VDD),.Y(g28029),.A(g26033),.B(g27247));
  NOR2 NOR2_1295(.VSS(VSS),.VDD(VDD),.Y(g28059),.A(g26034),.B(g27248));
  NOR2 NOR2_1296(.VSS(VSS),.VDD(VDD),.Y(g28088),.A(g26036),.B(g27249));
  NOR2 NOR2_1297(.VSS(VSS),.VDD(VDD),.Y(g28145),.A(g27629),.B(g17001));
  NOR2 NOR2_1298(.VSS(VSS),.VDD(VDD),.Y(g28146),.A(g27631),.B(g17031));
  NOR2 NOR2_1299(.VSS(VSS),.VDD(VDD),.Y(g28147),.A(g27655),.B(g17065));
  NOR2 NOR2_1300(.VSS(VSS),.VDD(VDD),.Y(g28148),.A(g27658),.B(g17100));
  NOR2 NOR2_1301(.VSS(VSS),.VDD(VDD),.Y(g28157),.A(g13902),.B(g27370));
  NOR2 NOR2_1302(.VSS(VSS),.VDD(VDD),.Y(g28185),.A(g27356),.B(g26845));
  NOR2 NOR2_1303(.VSS(VSS),.VDD(VDD),.Y(g28189),.A(g27359),.B(g26853));
  NOR2 NOR2_1304(.VSS(VSS),.VDD(VDD),.Y(g28191),.A(g27365),.B(g26860));
  NOR2 NOR2_1305(.VSS(VSS),.VDD(VDD),.Y(g28192),.A(g27372),.B(g26866));
  NOR2 NOR2_1306(.VSS(VSS),.VDD(VDD),.Y(g28199),.A(g27250),.B(g10024));
  NOR2 NOR2_1307(.VSS(VSS),.VDD(VDD),.Y(g28321),.A(g27742),.B(g10133));
  NOR2 NOR2_1308(.VSS(VSS),.VDD(VDD),.Y(g28325),.A(g27747),.B(g10238));
  NOR2 NOR2_1309(.VSS(VSS),.VDD(VDD),.Y(g28328),.A(g27755),.B(g10340));
  NOR2 NOR2_1310(.VSS(VSS),.VDD(VDD),.Y(g28342),.A(g15460),.B(g28008));
  NOR2 NOR2_1311(.VSS(VSS),.VDD(VDD),.Y(g28344),.A(g15526),.B(g28027));
  NOR2 NOR2_1312(.VSS(VSS),.VDD(VDD),.Y(g28345),.A(g15527),.B(g28028));
  NOR2 NOR2_1313(.VSS(VSS),.VDD(VDD),.Y(g28346),.A(g15546),.B(g28035));
  NOR2 NOR2_1314(.VSS(VSS),.VDD(VDD),.Y(g28348),.A(g15594),.B(g28050));
  NOR2 NOR2_1315(.VSS(VSS),.VDD(VDD),.Y(g28349),.A(g15595),.B(g28051));
  NOR2 NOR2_1316(.VSS(VSS),.VDD(VDD),.Y(g28350),.A(g15604),.B(g28057));
  NOR2 NOR2_1317(.VSS(VSS),.VDD(VDD),.Y(g28351),.A(g15605),.B(g28058));
  NOR2 NOR2_1318(.VSS(VSS),.VDD(VDD),.Y(g28352),.A(g15624),.B(g28065));
  NOR2 NOR2_1319(.VSS(VSS),.VDD(VDD),.Y(g28353),.A(g15666),.B(g28073));
  NOR2 NOR2_1320(.VSS(VSS),.VDD(VDD),.Y(g28354),.A(g15670),.B(g28079));
  NOR2 NOR2_1321(.VSS(VSS),.VDD(VDD),.Y(g28355),.A(g15671),.B(g28080));
  NOR2 NOR2_1322(.VSS(VSS),.VDD(VDD),.Y(g28356),.A(g15680),.B(g28086));
  NOR2 NOR2_1323(.VSS(VSS),.VDD(VDD),.Y(g28357),.A(g15681),.B(g28087));
  NOR2 NOR2_1324(.VSS(VSS),.VDD(VDD),.Y(g28358),.A(g15700),.B(g28094));
  NOR2 NOR2_1325(.VSS(VSS),.VDD(VDD),.Y(g28360),.A(g15725),.B(g28098));
  NOR2 NOR2_1326(.VSS(VSS),.VDD(VDD),.Y(g28361),.A(g15729),.B(g28104));
  NOR2 NOR2_1327(.VSS(VSS),.VDD(VDD),.Y(g28362),.A(g15730),.B(g28105));
  NOR2 NOR2_1328(.VSS(VSS),.VDD(VDD),.Y(g28363),.A(g15739),.B(g28111));
  NOR2 NOR2_1329(.VSS(VSS),.VDD(VDD),.Y(g28364),.A(g15740),.B(g28112));
  NOR2 NOR2_1330(.VSS(VSS),.VDD(VDD),.Y(g28366),.A(g15765),.B(g28116));
  NOR2 NOR2_1331(.VSS(VSS),.VDD(VDD),.Y(g28367),.A(g15769),.B(g28122));
  NOR2 NOR2_1332(.VSS(VSS),.VDD(VDD),.Y(g28368),.A(g15770),.B(g28123));
  NOR2 NOR2_1333(.VSS(VSS),.VDD(VDD),.Y(g28371),.A(g15793),.B(g28127));
  NOR2 NOR2_1334(.VSS(VSS),.VDD(VDD),.Y(g28392),.A(g27886),.B(g22344));
  NOR2 NOR2_1335(.VSS(VSS),.VDD(VDD),.Y(g28394),.A(g27869),.B(g22344));
  NOR2 NOR2_1336(.VSS(VSS),.VDD(VDD),.Y(g28397),.A(g27869),.B(g22344));
  NOR2 NOR2_1337(.VSS(VSS),.VDD(VDD),.Y(g28400),.A(g27886),.B(g22344));
  NOR2 NOR2_1338(.VSS(VSS),.VDD(VDD),.Y(g28403),.A(g27811),.B(g22344));
  NOR2 NOR2_1339(.VSS(VSS),.VDD(VDD),.Y(g28406),.A(g27824),.B(g22344));
  NOR2 NOR2_1340(.VSS(VSS),.VDD(VDD),.Y(g28409),.A(g24676),.B(g27801));
  NOR2 NOR2_1341(.VSS(VSS),.VDD(VDD),.Y(g28410),.A(g27748),.B(g22344));
  NOR2 NOR2_1342(.VSS(VSS),.VDD(VDD),.Y(g28413),.A(g24695),.B(g27809));
  NOR2 NOR2_1343(.VSS(VSS),.VDD(VDD),.Y(g28414),.A(g27748),.B(g22344));
  NOR2 NOR2_1344(.VSS(VSS),.VDD(VDD),.Y(g28417),.A(g24712),.B(g27830));
  NOR2 NOR2_1345(.VSS(VSS),.VDD(VDD),.Y(g28418),.A(g24723),.B(g27846));
  NOR2 NOR2_1346(.VSS(VSS),.VDD(VDD),.Y(g28420),.A(g16031),.B(g28171));
  NOR2 NOR2_1347(.VSS(VSS),.VDD(VDD),.Y(g28421),.A(g16068),.B(g28176));
  NOR2 NOR2_1348(.VSS(VSS),.VDD(VDD),.Y(g28425),.A(g16133),.B(g28188));
  NOR2 NOR2_1349(.VSS(VSS),.VDD(VDD),.Y(g28449),.A(g27727),.B(g26780));
  NOR2 NOR2_1350(.VSS(VSS),.VDD(VDD),.Y(g28461),.A(g27729),.B(g26787));
  NOR2 NOR2_1351(.VSS(VSS),.VDD(VDD),.Y(g28470),.A(g27671),.B(g28193));
  NOR2 NOR2_1352(.VSS(VSS),.VDD(VDD),.Y(g28473),.A(g27730),.B(g26794));
  NOR2 NOR2_1353(.VSS(VSS),.VDD(VDD),.Y(g28482),.A(g27731),.B(g26797));
  NOR2 NOR2_1354(.VSS(VSS),.VDD(VDD),.Y(g28488),.A(g26755),.B(g27719));
  NOR2 NOR2_1355(.VSS(VSS),.VDD(VDD),.Y(g28489),.A(g26756),.B(g27720));
  NOR2 NOR2_1356(.VSS(VSS),.VDD(VDD),.Y(g28490),.A(g27240),.B(g27721));
  NOR2 NOR2_1357(.VSS(VSS),.VDD(VDD),.Y(g28495),.A(g27244),.B(g27723));
  NOR2 NOR2_1358(.VSS(VSS),.VDD(VDD),.Y(g28499),.A(g26027),.B(g27725));
  NOR2 NOR2_1359(.VSS(VSS),.VDD(VDD),.Y(g28523),.A(g26035),.B(g27732));
  NOR2 NOR2_1360(.VSS(VSS),.VDD(VDD),.Y(g28525),.A(g27245),.B(g27726));
  NOR2 NOR2_1361(.VSS(VSS),.VDD(VDD),.Y(g28528),.A(g26030),.B(g27728));
  NOR2 NOR2_1362(.VSS(VSS),.VDD(VDD),.Y(g28551),.A(g26038),.B(g27733));
  NOR2 NOR2_1363(.VSS(VSS),.VDD(VDD),.Y(g28578),.A(g26039),.B(g27734));
  NOR2 NOR2_1364(.VSS(VSS),.VDD(VDD),.Y(g28606),.A(g26040),.B(g27737));
  NOR2 NOR2_1365(.VSS(VSS),.VDD(VDD),.Y(g28634),.A(g28185),.B(g17001));
  NOR2 NOR2_1366(.VSS(VSS),.VDD(VDD),.Y(g28635),.A(g28189),.B(g17031));
  NOR2 NOR2_1367(.VSS(VSS),.VDD(VDD),.Y(g28636),.A(g28191),.B(g17065));
  NOR2 NOR2_1368(.VSS(VSS),.VDD(VDD),.Y(g28637),.A(g28192),.B(g17100));
  NOR2 NOR2_1369(.VSS(VSS),.VDD(VDD),.Y(g28654),.A(g27770),.B(g27355));
  NOR2 NOR2_1370(.VSS(VSS),.VDD(VDD),.Y(g28656),.A(g27772),.B(g27358));
  NOR2 NOR2_1371(.VSS(VSS),.VDD(VDD),.Y(g28658),.A(g27773),.B(g27364));
  NOR2 NOR2_1372(.VSS(VSS),.VDD(VDD),.Y(g28661),.A(g27775),.B(g27371));
  NOR2 NOR2_1373(.VSS(VSS),.VDD(VDD),.Y(g28668),.A(g27736),.B(g10024));
  NOR2 NOR2_1374(.VSS(VSS),.VDD(VDD),.Y(g28728),.A(g28422),.B(g27904));
  NOR2 NOR2_1375(.VSS(VSS),.VDD(VDD),.Y(g28731),.A(g28423),.B(g27908));
  NOR2 NOR2_1376(.VSS(VSS),.VDD(VDD),.Y(g28732),.A(g14894),.B(g28426));
  NOR2 NOR2_1377(.VSS(VSS),.VDD(VDD),.Y(g28733),.A(g28424),.B(g27909));
  NOR2 NOR2_1378(.VSS(VSS),.VDD(VDD),.Y(g28735),.A(g14957),.B(g28430));
  NOR2 NOR2_1379(.VSS(VSS),.VDD(VDD),.Y(g28736),.A(g28427),.B(g27913));
  NOR2 NOR2_1380(.VSS(VSS),.VDD(VDD),.Y(g28737),.A(g28428),.B(g27914));
  NOR2 NOR2_1381(.VSS(VSS),.VDD(VDD),.Y(g28738),.A(g14975),.B(g28433));
  NOR2 NOR2_1382(.VSS(VSS),.VDD(VDD),.Y(g28739),.A(g28429),.B(g27915));
  NOR2 NOR2_1383(.VSS(VSS),.VDD(VDD),.Y(g28744),.A(g15030),.B(g28439));
  NOR2 NOR2_1384(.VSS(VSS),.VDD(VDD),.Y(g28745),.A(g28431),.B(g27922));
  NOR2 NOR2_1385(.VSS(VSS),.VDD(VDD),.Y(g28746),.A(g15046),.B(g28441));
  NOR2 NOR2_1386(.VSS(VSS),.VDD(VDD),.Y(g28747),.A(g28434),.B(g27923));
  NOR2 NOR2_1387(.VSS(VSS),.VDD(VDD),.Y(g28748),.A(g28435),.B(g27924));
  NOR2 NOR2_1388(.VSS(VSS),.VDD(VDD),.Y(g28749),.A(g15064),.B(g28444));
  NOR2 NOR2_1389(.VSS(VSS),.VDD(VDD),.Y(g28750),.A(g28436),.B(g27926));
  NOR2 NOR2_1390(.VSS(VSS),.VDD(VDD),.Y(g28754),.A(g28440),.B(g27931));
  NOR2 NOR2_1391(.VSS(VSS),.VDD(VDD),.Y(g28758),.A(g15126),.B(g28451));
  NOR2 NOR2_1392(.VSS(VSS),.VDD(VDD),.Y(g28759),.A(g28442),.B(g27935));
  NOR2 NOR2_1393(.VSS(VSS),.VDD(VDD),.Y(g28760),.A(g15142),.B(g28453));
  NOR2 NOR2_1394(.VSS(VSS),.VDD(VDD),.Y(g28761),.A(g28445),.B(g27936));
  NOR2 NOR2_1395(.VSS(VSS),.VDD(VDD),.Y(g28762),.A(g28446),.B(g27938));
  NOR2 NOR2_1396(.VSS(VSS),.VDD(VDD),.Y(g28763),.A(g15160),.B(g28456));
  NOR2 NOR2_1397(.VSS(VSS),.VDD(VDD),.Y(g28767),.A(g28452),.B(g27945));
  NOR2 NOR2_1398(.VSS(VSS),.VDD(VDD),.Y(g28771),.A(g15218),.B(g28463));
  NOR2 NOR2_1399(.VSS(VSS),.VDD(VDD),.Y(g28772),.A(g28454),.B(g27949));
  NOR2 NOR2_1400(.VSS(VSS),.VDD(VDD),.Y(g28773),.A(g15234),.B(g28465));
  NOR2 NOR2_1401(.VSS(VSS),.VDD(VDD),.Y(g28774),.A(g28457),.B(g27951));
  NOR2 NOR2_1402(.VSS(VSS),.VDD(VDD),.Y(g28778),.A(g28464),.B(g27963));
  NOR2 NOR2_1403(.VSS(VSS),.VDD(VDD),.Y(g28782),.A(g15304),.B(g28475));
  NOR2 NOR2_1404(.VSS(VSS),.VDD(VDD),.Y(g28783),.A(g28466),.B(g27968));
  NOR2 NOR2_1405(.VSS(VSS),.VDD(VDD),.Y(g28784),.A(g28468),.B(g27970));
  NOR2 NOR2_1406(.VSS(VSS),.VDD(VDD),.Y(g28788),.A(g28476),.B(g27984));
  NOR2 NOR2_1407(.VSS(VSS),.VDD(VDD),.Y(g28789),.A(g28477),.B(g27985));
  NOR2 NOR2_1408(.VSS(VSS),.VDD(VDD),.Y(g28790),.A(g28478),.B(g27991));
  NOR2 NOR2_1409(.VSS(VSS),.VDD(VDD),.Y(g28794),.A(g28484),.B(g28009));
  NOR2 NOR2_1410(.VSS(VSS),.VDD(VDD),.Y(g28795),.A(g28485),.B(g28015));
  NOR2 NOR2_1411(.VSS(VSS),.VDD(VDD),.Y(g28802),.A(g28492),.B(g28036));
  NOR2 NOR2_1412(.VSS(VSS),.VDD(VDD),.Y(g28803),.A(g28493),.B(g28042));
  NOR2 NOR2_1413(.VSS(VSS),.VDD(VDD),.Y(g28813),.A(g28497),.B(g28066));
  NOR2 NOR2_1414(.VSS(VSS),.VDD(VDD),.Y(g28874),.A(g28657),.B(g16221));
  NOR2 NOR2_1415(.VSS(VSS),.VDD(VDD),.Y(g28886),.A(g28659),.B(g16277));
  NOR2 NOR2_1416(.VSS(VSS),.VDD(VDD),.Y(g28903),.A(g28660),.B(g13295));
  NOR2 NOR2_1417(.VSS(VSS),.VDD(VDD),.Y(g28920),.A(g28662),.B(g13322));
  NOR2 NOR2_1418(.VSS(VSS),.VDD(VDD),.Y(g28941),.A(g28663),.B(g13343));
  NOR3 NOR3_397(.VSS(VSS),.VDD(VDD),.Y(g28954),.A(g26673),.B(g27241),.C(g28323));
  NOR2 NOR2_1419(.VSS(VSS),.VDD(VDD),.Y(g28963),.A(g28664),.B(g13365));
  NOR2 NOR2_1420(.VSS(VSS),.VDD(VDD),.Y(g28982),.A(g28665),.B(g28670));
  NOR2 NOR2_1421(.VSS(VSS),.VDD(VDD),.Y(g28987),.A(g28666),.B(g13390));
  NOR2 NOR2_1422(.VSS(VSS),.VDD(VDD),.Y(g28990),.A(g28667),.B(g16457));
  NOR2 NOR2_1423(.VSS(VSS),.VDD(VDD),.Y(g29009),.A(g28669),.B(g28320));
  NOR2 NOR2_1424(.VSS(VSS),.VDD(VDD),.Y(g29013),.A(g28671),.B(g11607));
  NOR2 NOR2_1425(.VSS(VSS),.VDD(VDD),.Y(g29016),.A(g28672),.B(g13487));
  NOR2 NOR2_1426(.VSS(VSS),.VDD(VDD),.Y(g29031),.A(g28319),.B(g28324));
  NOR2 NOR2_1427(.VSS(VSS),.VDD(VDD),.Y(g29039),.A(g28322),.B(g13500));
  NOR2 NOR2_1428(.VSS(VSS),.VDD(VDD),.Y(g29063),.A(g28326),.B(g28329));
  NOR2 NOR2_1429(.VSS(VSS),.VDD(VDD),.Y(g29064),.A(g28327),.B(g28330));
  NOR2 NOR2_1430(.VSS(VSS),.VDD(VDD),.Y(g29083),.A(g28331),.B(g28333));
  NOR2 NOR2_1431(.VSS(VSS),.VDD(VDD),.Y(g29090),.A(g28332),.B(g28334));
  NOR2 NOR2_1432(.VSS(VSS),.VDD(VDD),.Y(g29097),.A(g28335),.B(g28336));
  NOR2 NOR2_1433(.VSS(VSS),.VDD(VDD),.Y(g29109),.A(g28654),.B(g17001));
  NOR2 NOR2_1434(.VSS(VSS),.VDD(VDD),.Y(g29110),.A(g28656),.B(g17031));
  NOR2 NOR2_1435(.VSS(VSS),.VDD(VDD),.Y(g29111),.A(g28658),.B(g17065));
  NOR2 NOR2_1436(.VSS(VSS),.VDD(VDD),.Y(g29112),.A(g28661),.B(g17100));
  NOR2 NOR2_1437(.VSS(VSS),.VDD(VDD),.Y(g29113),.A(g28381),.B(g8907));
  NOR2 NOR2_1438(.VSS(VSS),.VDD(VDD),.Y(g29126),.A(g28373),.B(g27774));
  NOR2 NOR2_1439(.VSS(VSS),.VDD(VDD),.Y(g29127),.A(g28376),.B(g27779));
  NOR2 NOR2_1440(.VSS(VSS),.VDD(VDD),.Y(g29128),.A(g28380),.B(g27783));
  NOR2 NOR2_1441(.VSS(VSS),.VDD(VDD),.Y(g29129),.A(g28385),.B(g27790));
  NOR2 NOR2_1442(.VSS(VSS),.VDD(VDD),.Y(g29167),.A(g28841),.B(g28396));
  NOR2 NOR2_1443(.VSS(VSS),.VDD(VDD),.Y(g29169),.A(g28843),.B(g28398));
  NOR2 NOR2_1444(.VSS(VSS),.VDD(VDD),.Y(g29170),.A(g28844),.B(g28399));
  NOR2 NOR2_1445(.VSS(VSS),.VDD(VDD),.Y(g29172),.A(g28846),.B(g28401));
  NOR2 NOR2_1446(.VSS(VSS),.VDD(VDD),.Y(g29173),.A(g28847),.B(g28402));
  NOR2 NOR2_1447(.VSS(VSS),.VDD(VDD),.Y(g29178),.A(g28848),.B(g28404));
  NOR2 NOR2_1448(.VSS(VSS),.VDD(VDD),.Y(g29179),.A(g28849),.B(g28405));
  NOR2 NOR2_1449(.VSS(VSS),.VDD(VDD),.Y(g29181),.A(g28850),.B(g28407));
  NOR2 NOR2_1450(.VSS(VSS),.VDD(VDD),.Y(g29182),.A(g28851),.B(g28408));
  NOR2 NOR2_1451(.VSS(VSS),.VDD(VDD),.Y(g29184),.A(g28852),.B(g28411));
  NOR2 NOR2_1452(.VSS(VSS),.VDD(VDD),.Y(g29185),.A(g28853),.B(g28412));
  NOR2 NOR2_1453(.VSS(VSS),.VDD(VDD),.Y(g29187),.A(g28854),.B(g28416));
  NOR2 NOR2_1454(.VSS(VSS),.VDD(VDD),.Y(g29194),.A(g14958),.B(g28881));
  NOR2 NOR2_1455(.VSS(VSS),.VDD(VDD),.Y(g29195),.A(g28880),.B(g28438));
  NOR2 NOR2_1456(.VSS(VSS),.VDD(VDD),.Y(g29197),.A(g15031),.B(g28893));
  NOR2 NOR2_1457(.VSS(VSS),.VDD(VDD),.Y(g29198),.A(g15047),.B(g28898));
  NOR2 NOR2_1458(.VSS(VSS),.VDD(VDD),.Y(g29199),.A(g28892),.B(g28448));
  NOR2 NOR2_1459(.VSS(VSS),.VDD(VDD),.Y(g29201),.A(g15104),.B(g28910));
  NOR2 NOR2_1460(.VSS(VSS),.VDD(VDD),.Y(g29202),.A(g28897),.B(g28450));
  NOR2 NOR2_1461(.VSS(VSS),.VDD(VDD),.Y(g29204),.A(g15127),.B(g28915));
  NOR2 NOR2_1462(.VSS(VSS),.VDD(VDD),.Y(g29205),.A(g15143),.B(g28923));
  NOR2 NOR2_1463(.VSS(VSS),.VDD(VDD),.Y(g29206),.A(g28909),.B(g28459));
  NOR2 NOR2_1464(.VSS(VSS),.VDD(VDD),.Y(g29207),.A(g28914),.B(g28460));
  NOR2 NOR2_1465(.VSS(VSS),.VDD(VDD),.Y(g29209),.A(g15196),.B(g28936));
  NOR2 NOR2_1466(.VSS(VSS),.VDD(VDD),.Y(g29210),.A(g28919),.B(g28462));
  NOR2 NOR2_1467(.VSS(VSS),.VDD(VDD),.Y(g29212),.A(g15219),.B(g28944));
  NOR2 NOR2_1468(.VSS(VSS),.VDD(VDD),.Y(g29213),.A(g15235),.B(g28949));
  NOR2 NOR2_1469(.VSS(VSS),.VDD(VDD),.Y(g29214),.A(g28931),.B(g28469));
  NOR2 NOR2_1470(.VSS(VSS),.VDD(VDD),.Y(g29215),.A(g28935),.B(g28471));
  NOR2 NOR2_1471(.VSS(VSS),.VDD(VDD),.Y(g29216),.A(g28940),.B(g28472));
  NOR2 NOR2_1472(.VSS(VSS),.VDD(VDD),.Y(g29218),.A(g15282),.B(g28966));
  NOR2 NOR2_1473(.VSS(VSS),.VDD(VDD),.Y(g29219),.A(g28948),.B(g28474));
  NOR2 NOR2_1474(.VSS(VSS),.VDD(VDD),.Y(g29221),.A(g15305),.B(g28971));
  NOR2 NOR2_1475(.VSS(VSS),.VDD(VDD),.Y(g29222),.A(g28958),.B(g28479));
  NOR2 NOR2_1476(.VSS(VSS),.VDD(VDD),.Y(g29223),.A(g28962),.B(g28480));
  NOR2 NOR2_1477(.VSS(VSS),.VDD(VDD),.Y(g29224),.A(g28970),.B(g28481));
  NOR2 NOR2_1478(.VSS(VSS),.VDD(VDD),.Y(g29226),.A(g15374),.B(g28997));
  NOR2 NOR2_1479(.VSS(VSS),.VDD(VDD),.Y(g29227),.A(g28986),.B(g28486));
  NOR2 NOR2_1480(.VSS(VSS),.VDD(VDD),.Y(g29228),.A(g28996),.B(g28487));
  NOR2 NOR2_1481(.VSS(VSS),.VDD(VDD),.Y(g29231),.A(g29022),.B(g28494));
  NOR2 NOR2_1482(.VSS(VSS),.VDD(VDD),.Y(g29303),.A(g28716),.B(g19112));
  NOR2 NOR2_1483(.VSS(VSS),.VDD(VDD),.Y(g29313),.A(g28717),.B(g19117));
  NOR2 NOR2_1484(.VSS(VSS),.VDD(VDD),.Y(g29324),.A(g28718),.B(g19124));
  NOR2 NOR2_1485(.VSS(VSS),.VDD(VDD),.Y(g29333),.A(g28719),.B(g19131));
  NOR2 NOR2_1486(.VSS(VSS),.VDD(VDD),.Y(g29340),.A(g28337),.B(g28722));
  NOR2 NOR2_1487(.VSS(VSS),.VDD(VDD),.Y(g29343),.A(g28338),.B(g28724));
  NOR2 NOR2_1488(.VSS(VSS),.VDD(VDD),.Y(g29345),.A(g28339),.B(g28726));
  NOR2 NOR2_1489(.VSS(VSS),.VDD(VDD),.Y(g29347),.A(g28340),.B(g28729));
  NOR2 NOR2_1490(.VSS(VSS),.VDD(VDD),.Y(g29353),.A(g29126),.B(g17001));
  NOR2 NOR2_1491(.VSS(VSS),.VDD(VDD),.Y(g29354),.A(g29127),.B(g17031));
  NOR2 NOR2_1492(.VSS(VSS),.VDD(VDD),.Y(g29355),.A(g29128),.B(g17065));
  NOR2 NOR2_1493(.VSS(VSS),.VDD(VDD),.Y(g29357),.A(g29129),.B(g17100));
  NOR2 NOR2_1494(.VSS(VSS),.VDD(VDD),.Y(g29399),.A(g28834),.B(g28378));
  NOR2 NOR2_1495(.VSS(VSS),.VDD(VDD),.Y(g29403),.A(g28836),.B(g28383));
  NOR2 NOR2_1496(.VSS(VSS),.VDD(VDD),.Y(g29406),.A(g28838),.B(g28387));
  NOR2 NOR2_1497(.VSS(VSS),.VDD(VDD),.Y(g29409),.A(g28840),.B(g28389));
  NOR2 NOR2_1498(.VSS(VSS),.VDD(VDD),.Y(g29552),.A(g29130),.B(g29411));
  NOR2 NOR2_1499(.VSS(VSS),.VDD(VDD),.Y(g29569),.A(g28708),.B(g29174));
  NOR2 NOR2_1500(.VSS(VSS),.VDD(VDD),.Y(g29570),.A(g28709),.B(g29175));
  NOR2 NOR2_1501(.VSS(VSS),.VDD(VDD),.Y(g29571),.A(g28710),.B(g29176));
  NOR2 NOR2_1502(.VSS(VSS),.VDD(VDD),.Y(g29574),.A(g28712),.B(g29180));
  NOR2 NOR2_1503(.VSS(VSS),.VDD(VDD),.Y(g29576),.A(g28713),.B(g29183));
  NOR2 NOR2_1504(.VSS(VSS),.VDD(VDD),.Y(g29577),.A(g28714),.B(g29186));
  NOR2 NOR2_1505(.VSS(VSS),.VDD(VDD),.Y(g29578),.A(g28715),.B(g29188));
  NOR2 NOR2_1506(.VSS(VSS),.VDD(VDD),.Y(g29579),.A(g29399),.B(g17001));
  NOR2 NOR2_1507(.VSS(VSS),.VDD(VDD),.Y(g29580),.A(g29403),.B(g17031));
  NOR2 NOR2_1508(.VSS(VSS),.VDD(VDD),.Y(g29581),.A(g29406),.B(g17065));
  NOR2 NOR2_1509(.VSS(VSS),.VDD(VDD),.Y(g29582),.A(g29409),.B(g17100));
  NOR2 NOR2_1510(.VSS(VSS),.VDD(VDD),.Y(g29606),.A(g13878),.B(g29248));
  NOR2 NOR2_1511(.VSS(VSS),.VDD(VDD),.Y(g29608),.A(g13892),.B(g29251));
  NOR2 NOR2_1512(.VSS(VSS),.VDD(VDD),.Y(g29609),.A(g13900),.B(g29252));
  NOR2 NOR2_1513(.VSS(VSS),.VDD(VDD),.Y(g29611),.A(g13913),.B(g29255));
  NOR2 NOR2_1514(.VSS(VSS),.VDD(VDD),.Y(g29612),.A(g13933),.B(g29256));
  NOR2 NOR2_1515(.VSS(VSS),.VDD(VDD),.Y(g29613),.A(g13941),.B(g29257));
  NOR2 NOR2_1516(.VSS(VSS),.VDD(VDD),.Y(g29616),.A(g13969),.B(g29259));
  NOR2 NOR2_1517(.VSS(VSS),.VDD(VDD),.Y(g29617),.A(g13989),.B(g29260));
  NOR2 NOR2_1518(.VSS(VSS),.VDD(VDD),.Y(g29618),.A(g13997),.B(g29261));
  NOR2 NOR2_1519(.VSS(VSS),.VDD(VDD),.Y(g29620),.A(g14039),.B(g29262));
  NOR2 NOR2_1520(.VSS(VSS),.VDD(VDD),.Y(g29621),.A(g14059),.B(g29263));
  NOR2 NOR2_1521(.VSS(VSS),.VDD(VDD),.Y(g29623),.A(g14130),.B(g29264));
  NOR2 NOR2_1522(.VSS(VSS),.VDD(VDD),.Y(g29663),.A(g29518),.B(g29284));
  NOR2 NOR2_1523(.VSS(VSS),.VDD(VDD),.Y(g29665),.A(g29521),.B(g29289));
  NOR2 NOR2_1524(.VSS(VSS),.VDD(VDD),.Y(g29667),.A(g29524),.B(g29294));
  NOR2 NOR2_1525(.VSS(VSS),.VDD(VDD),.Y(g29669),.A(g29528),.B(g29300));
  NOR2 NOR2_1526(.VSS(VSS),.VDD(VDD),.Y(g29670),.A(g29529),.B(g29302));
  NOR2 NOR2_1527(.VSS(VSS),.VDD(VDD),.Y(g29671),.A(g29534),.B(g29310));
  NOR2 NOR2_1528(.VSS(VSS),.VDD(VDD),.Y(g29672),.A(g29536),.B(g29312));
  NOR2 NOR2_1529(.VSS(VSS),.VDD(VDD),.Y(g29676),.A(g29540),.B(g29320));
  NOR2 NOR2_1530(.VSS(VSS),.VDD(VDD),.Y(g29677),.A(g29543),.B(g29321));
  NOR2 NOR2_1531(.VSS(VSS),.VDD(VDD),.Y(g29678),.A(g29545),.B(g29323));
  NOR2 NOR2_1532(.VSS(VSS),.VDD(VDD),.Y(g29679),.A(g29549),.B(g29329));
  NOR2 NOR2_1533(.VSS(VSS),.VDD(VDD),.Y(g29680),.A(g29553),.B(g29330));
  NOR2 NOR2_1534(.VSS(VSS),.VDD(VDD),.Y(g29681),.A(g29555),.B(g29332));
  NOR2 NOR2_1535(.VSS(VSS),.VDD(VDD),.Y(g29682),.A(g29557),.B(g29336));
  NOR2 NOR2_1536(.VSS(VSS),.VDD(VDD),.Y(g29683),.A(g29559),.B(g29337));
  NOR2 NOR2_1537(.VSS(VSS),.VDD(VDD),.Y(g29684),.A(g29562),.B(g29338));
  NOR2 NOR2_1538(.VSS(VSS),.VDD(VDD),.Y(g29685),.A(g29564),.B(g29341));
  NOR2 NOR2_1539(.VSS(VSS),.VDD(VDD),.Y(g29686),.A(g29566),.B(g29342));
  NOR2 NOR2_1540(.VSS(VSS),.VDD(VDD),.Y(g29687),.A(g29572),.B(g29344));
  NOR2 NOR2_1541(.VSS(VSS),.VDD(VDD),.Y(g29688),.A(g29575),.B(g29346));
  NOR2 NOR2_1542(.VSS(VSS),.VDD(VDD),.Y(g29703),.A(g29583),.B(g1917));
  NOR3 NOR3_398(.VSS(VSS),.VDD(VDD),.Y(g29705),.A(g6104),.B(g29583),.C(g25339));
  NOR2 NOR2_1543(.VSS(VSS),.VDD(VDD),.Y(g29709),.A(g29583),.B(g1909));
  NOR3 NOR3_399(.VSS(VSS),.VDD(VDD),.Y(g29710),.A(g6104),.B(g29583),.C(g25412));
  NOR3 NOR3_400(.VSS(VSS),.VDD(VDD),.Y(g29713),.A(g6104),.B(g29583),.C(g25332));
  NOR2 NOR2_1544(.VSS(VSS),.VDD(VDD),.Y(g29717),.A(g29583),.B(g1910));
  NOR3 NOR3_401(.VSS(VSS),.VDD(VDD),.Y(g29718),.A(g6104),.B(g29583),.C(g25409));
  NOR3 NOR3_402(.VSS(VSS),.VDD(VDD),.Y(g29721),.A(g6104),.B(g29583),.C(g25323));
  NOR2 NOR2_1545(.VSS(VSS),.VDD(VDD),.Y(g29725),.A(g29583),.B(g1911));
  NOR2 NOR2_1546(.VSS(VSS),.VDD(VDD),.Y(g29727),.A(g29583),.B(g1912));
  NOR3 NOR3_403(.VSS(VSS),.VDD(VDD),.Y(g29728),.A(g6104),.B(g29583),.C(g25401));
  NOR2 NOR2_1547(.VSS(VSS),.VDD(VDD),.Y(g29731),.A(g29583),.B(g1913));
  NOR3 NOR3_404(.VSS(VSS),.VDD(VDD),.Y(g29732),.A(g6104),.B(g29583),.C(g25387));
  NOR2 NOR2_1548(.VSS(VSS),.VDD(VDD),.Y(g29735),.A(g23797),.B(g29583));
  NOR2 NOR2_1549(.VSS(VSS),.VDD(VDD),.Y(g29736),.A(g29583),.B(g25444));
  NOR2 NOR2_1550(.VSS(VSS),.VDD(VDD),.Y(g29740),.A(g29583),.B(g1914));
  NOR3 NOR3_405(.VSS(VSS),.VDD(VDD),.Y(g29741),.A(g6104),.B(g29583),.C(g25376));
  NOR2 NOR2_1551(.VSS(VSS),.VDD(VDD),.Y(g29744),.A(g29583),.B(g24641));
  NOR2 NOR2_1552(.VSS(VSS),.VDD(VDD),.Y(g29747),.A(g29583),.B(g1916));
  NOR3 NOR3_406(.VSS(VSS),.VDD(VDD),.Y(g29748),.A(g6104),.B(g29583),.C(g25363));
  NOR3 NOR3_407(.VSS(VSS),.VDD(VDD),.Y(g29751),.A(g6104),.B(g29583),.C(g25352));
  NOR2 NOR2_1553(.VSS(VSS),.VDD(VDD),.Y(g29754),.A(g16178),.B(g29607));
  NOR2 NOR2_1554(.VSS(VSS),.VDD(VDD),.Y(g29755),.A(g16229),.B(g29610));
  NOR2 NOR2_1555(.VSS(VSS),.VDD(VDD),.Y(g29756),.A(g16284),.B(g29614));
  NOR2 NOR2_1556(.VSS(VSS),.VDD(VDD),.Y(g29757),.A(g16285),.B(g29615));
  NOR2 NOR2_1557(.VSS(VSS),.VDD(VDD),.Y(g29758),.A(g16335),.B(g29619));
  NOR2 NOR2_1558(.VSS(VSS),.VDD(VDD),.Y(g29759),.A(g16379),.B(g29622));
  NOR2 NOR2_1559(.VSS(VSS),.VDD(VDD),.Y(g29760),.A(g16411),.B(g29624));
  NOR3 NOR3_408(.VSS(VSS),.VDD(VDD),.Y(g29761),.A(g28707),.B(g28711),.C(g29466));
  NOR2 NOR2_1560(.VSS(VSS),.VDD(VDD),.Y(g29762),.A(g16432),.B(g29625));
  NOR2 NOR2_1561(.VSS(VSS),.VDD(VDD),.Y(g29763),.A(g16438),.B(g29626));
  NOR2 NOR2_1562(.VSS(VSS),.VDD(VDD),.Y(g29764),.A(g16462),.B(g29464));
  NOR2 NOR2_1563(.VSS(VSS),.VDD(VDD),.Y(g29765),.A(g13492),.B(g29465));
  NOR2 NOR2_1564(.VSS(VSS),.VDD(VDD),.Y(g29766),.A(g29467),.B(g19142));
  NOR2 NOR2_1565(.VSS(VSS),.VDD(VDD),.Y(g29767),.A(g29468),.B(g19143));
  NOR2 NOR2_1566(.VSS(VSS),.VDD(VDD),.Y(g29768),.A(g29469),.B(g19146));
  NOR2 NOR2_1567(.VSS(VSS),.VDD(VDD),.Y(g29769),.A(g29470),.B(g19148));
  NOR2 NOR2_1568(.VSS(VSS),.VDD(VDD),.Y(g29770),.A(g29471),.B(g29196));
  NOR2 NOR2_1569(.VSS(VSS),.VDD(VDD),.Y(g29771),.A(g29472),.B(g29200));
  NOR2 NOR2_1570(.VSS(VSS),.VDD(VDD),.Y(g29772),.A(g29473),.B(g29203));
  NOR2 NOR2_1571(.VSS(VSS),.VDD(VDD),.Y(g29773),.A(g29474),.B(g29208));
  NOR2 NOR2_1572(.VSS(VSS),.VDD(VDD),.Y(g29774),.A(g29475),.B(g29211));
  NOR2 NOR2_1573(.VSS(VSS),.VDD(VDD),.Y(g29775),.A(g29476),.B(g29217));
  NOR2 NOR2_1574(.VSS(VSS),.VDD(VDD),.Y(g29776),.A(g29477),.B(g29220));
  NOR2 NOR2_1575(.VSS(VSS),.VDD(VDD),.Y(g29777),.A(g29478),.B(g29225));
  NOR2 NOR2_1576(.VSS(VSS),.VDD(VDD),.Y(g29778),.A(g29479),.B(g29229));
  NOR2 NOR2_1577(.VSS(VSS),.VDD(VDD),.Y(g29779),.A(g13943),.B(g29502));
  NOR2 NOR2_1578(.VSS(VSS),.VDD(VDD),.Y(g29780),.A(g29480),.B(g29232));
  NOR2 NOR2_1579(.VSS(VSS),.VDD(VDD),.Y(g29781),.A(g29481),.B(g29233));
  NOR2 NOR2_1580(.VSS(VSS),.VDD(VDD),.Y(g29782),.A(g29482),.B(g29234));
  NOR2 NOR2_1581(.VSS(VSS),.VDD(VDD),.Y(g29783),.A(g29483),.B(g29235));
  NOR2 NOR2_1582(.VSS(VSS),.VDD(VDD),.Y(g29784),.A(g29484),.B(g29236));
  NOR2 NOR2_1583(.VSS(VSS),.VDD(VDD),.Y(g29785),.A(g29485),.B(g29238));
  NOR2 NOR2_1584(.VSS(VSS),.VDD(VDD),.Y(g29786),.A(g29486),.B(g29239));
  NOR2 NOR2_1585(.VSS(VSS),.VDD(VDD),.Y(g29787),.A(g29487),.B(g29240));
  NOR2 NOR2_1586(.VSS(VSS),.VDD(VDD),.Y(g29788),.A(g29488),.B(g29241));
  NOR2 NOR2_1587(.VSS(VSS),.VDD(VDD),.Y(g29789),.A(g29489),.B(g29242));
  NOR2 NOR2_1588(.VSS(VSS),.VDD(VDD),.Y(g29791),.A(g29490),.B(g29243));
  NOR2 NOR2_1589(.VSS(VSS),.VDD(VDD),.Y(g29912),.A(g24676),.B(g29716));
  NOR2 NOR2_1590(.VSS(VSS),.VDD(VDD),.Y(g29914),.A(g24695),.B(g29724));
  NOR2 NOR2_1591(.VSS(VSS),.VDD(VDD),.Y(g29916),.A(g24712),.B(g29726));
  NOR2 NOR2_1592(.VSS(VSS),.VDD(VDD),.Y(g29918),.A(g29744),.B(g22367));
  NOR2 NOR2_1593(.VSS(VSS),.VDD(VDD),.Y(g29919),.A(g29736),.B(g22367));
  NOR2 NOR2_1594(.VSS(VSS),.VDD(VDD),.Y(g29920),.A(g24723),.B(g29739));
  NOR2 NOR2_1595(.VSS(VSS),.VDD(VDD),.Y(g29921),.A(g29736),.B(g22367));
  NOR2 NOR2_1596(.VSS(VSS),.VDD(VDD),.Y(g29922),.A(g29744),.B(g22367));
  NOR2 NOR2_1597(.VSS(VSS),.VDD(VDD),.Y(g29924),.A(g29710),.B(g22367));
  NOR2 NOR2_1598(.VSS(VSS),.VDD(VDD),.Y(g29926),.A(g29718),.B(g22367));
  NOR2 NOR2_1599(.VSS(VSS),.VDD(VDD),.Y(g29928),.A(g29673),.B(g22367));
  NOR2 NOR2_1600(.VSS(VSS),.VDD(VDD),.Y(g29929),.A(g29673),.B(g22367));
  NOR2 NOR2_1601(.VSS(VSS),.VDD(VDD),.Y(g29936),.A(g16049),.B(g29790));
  NOR2 NOR2_1602(.VSS(VSS),.VDD(VDD),.Y(g29939),.A(g16102),.B(g29792));
  NOR2 NOR2_1603(.VSS(VSS),.VDD(VDD),.Y(g29941),.A(g16182),.B(g29793));
  NOR2 NOR2_1604(.VSS(VSS),.VDD(VDD),.Y(g30010),.A(g29520),.B(g29942));
  NOR2 NOR2_1605(.VSS(VSS),.VDD(VDD),.Y(g30011),.A(g29522),.B(g29944));
  NOR2 NOR2_1606(.VSS(VSS),.VDD(VDD),.Y(g30012),.A(g29523),.B(g29945));
  NOR2 NOR2_1607(.VSS(VSS),.VDD(VDD),.Y(g30013),.A(g29525),.B(g29946));
  NOR2 NOR2_1608(.VSS(VSS),.VDD(VDD),.Y(g30014),.A(g29526),.B(g29947));
  NOR2 NOR2_1609(.VSS(VSS),.VDD(VDD),.Y(g30015),.A(g29527),.B(g29948));
  NOR2 NOR2_1610(.VSS(VSS),.VDD(VDD),.Y(g30016),.A(g29531),.B(g29949));
  NOR2 NOR2_1611(.VSS(VSS),.VDD(VDD),.Y(g30017),.A(g29532),.B(g29950));
  NOR2 NOR2_1612(.VSS(VSS),.VDD(VDD),.Y(g30018),.A(g29533),.B(g29951));
  NOR2 NOR2_1613(.VSS(VSS),.VDD(VDD),.Y(g30019),.A(g29538),.B(g29952));
  NOR2 NOR2_1614(.VSS(VSS),.VDD(VDD),.Y(g30020),.A(g29539),.B(g29953));
  NOR2 NOR2_1615(.VSS(VSS),.VDD(VDD),.Y(g30021),.A(g29541),.B(g29954));
  NOR2 NOR2_1616(.VSS(VSS),.VDD(VDD),.Y(g30022),.A(g29547),.B(g29955));
  NOR2 NOR2_1617(.VSS(VSS),.VDD(VDD),.Y(g30023),.A(g29548),.B(g29956));
  NOR2 NOR2_1618(.VSS(VSS),.VDD(VDD),.Y(g30024),.A(g29550),.B(g29957));
  NOR2 NOR2_1619(.VSS(VSS),.VDD(VDD),.Y(g30025),.A(g29558),.B(g29958));
  NOR2 NOR2_1620(.VSS(VSS),.VDD(VDD),.Y(g30026),.A(g29560),.B(g29959));
  NOR2 NOR2_1621(.VSS(VSS),.VDD(VDD),.Y(g30027),.A(g29565),.B(g29960));
  NOR2 NOR2_1622(.VSS(VSS),.VDD(VDD),.Y(g30028),.A(g29567),.B(g29961));
  NOR2 NOR2_1623(.VSS(VSS),.VDD(VDD),.Y(g30029),.A(g29573),.B(g29962));
  NOR2 NOR2_1624(.VSS(VSS),.VDD(VDD),.Y(g30030),.A(g24676),.B(g29923));
  NOR2 NOR2_1625(.VSS(VSS),.VDD(VDD),.Y(g30031),.A(g24695),.B(g29925));
  NOR2 NOR2_1626(.VSS(VSS),.VDD(VDD),.Y(g30032),.A(g24712),.B(g29927));
  NOR2 NOR2_1627(.VSS(VSS),.VDD(VDD),.Y(g30033),.A(g24723),.B(g29931));
  NOR2 NOR2_1628(.VSS(VSS),.VDD(VDD),.Y(g30053),.A(g29963),.B(g16286));
  NOR2 NOR2_1629(.VSS(VSS),.VDD(VDD),.Y(g30054),.A(g29964),.B(g16336));
  NOR2 NOR2_1630(.VSS(VSS),.VDD(VDD),.Y(g30055),.A(g29965),.B(g13326));
  NOR2 NOR2_1631(.VSS(VSS),.VDD(VDD),.Y(g30056),.A(g29966),.B(g13345));
  NOR2 NOR2_1632(.VSS(VSS),.VDD(VDD),.Y(g30057),.A(g29967),.B(g13368));
  NOR2 NOR2_1633(.VSS(VSS),.VDD(VDD),.Y(g30058),.A(g29968),.B(g13395));
  NOR2 NOR2_1634(.VSS(VSS),.VDD(VDD),.Y(g30059),.A(g29969),.B(g29811));
  NOR2 NOR2_1635(.VSS(VSS),.VDD(VDD),.Y(g30060),.A(g29970),.B(g11612));
  NOR2 NOR2_1636(.VSS(VSS),.VDD(VDD),.Y(g30061),.A(g29971),.B(g13493));
  NOR2 NOR2_1637(.VSS(VSS),.VDD(VDD),.Y(g30062),.A(g29810),.B(g29815));
  NOR2 NOR2_1638(.VSS(VSS),.VDD(VDD),.Y(g30063),.A(g29812),.B(g11637));
  NOR2 NOR2_1639(.VSS(VSS),.VDD(VDD),.Y(g30064),.A(g29813),.B(g13506));
  NOR2 NOR2_1640(.VSS(VSS),.VDD(VDD),.Y(g30065),.A(g29814),.B(g29817));
  NOR2 NOR2_1641(.VSS(VSS),.VDD(VDD),.Y(g30066),.A(g29816),.B(g13517));
  NOR2 NOR2_1642(.VSS(VSS),.VDD(VDD),.Y(g30067),.A(g29818),.B(g29820));
  NOR2 NOR2_1643(.VSS(VSS),.VDD(VDD),.Y(g30068),.A(g29819),.B(g29821));
  NOR2 NOR2_1644(.VSS(VSS),.VDD(VDD),.Y(g30069),.A(g29822),.B(g29828));
  NOR2 NOR2_1645(.VSS(VSS),.VDD(VDD),.Y(g30070),.A(g29827),.B(g29833));
  NOR2 NOR2_1646(.VSS(VSS),.VDD(VDD),.Y(g30071),.A(g29834),.B(g29839));
  NOR2 NOR2_1647(.VSS(VSS),.VDD(VDD),.Y(g30072),.A(g29910),.B(g8947));
  NOR2 NOR2_1648(.VSS(VSS),.VDD(VDD),.Y(g30245),.A(g16074),.B(g30077));
  NOR2 NOR2_1649(.VSS(VSS),.VDD(VDD),.Y(g30246),.A(g16107),.B(g30079));
  NOR2 NOR2_1650(.VSS(VSS),.VDD(VDD),.Y(g30247),.A(g16112),.B(g30080));
  NOR2 NOR2_1651(.VSS(VSS),.VDD(VDD),.Y(g30248),.A(g16139),.B(g30081));
  NOR2 NOR2_1652(.VSS(VSS),.VDD(VDD),.Y(g30249),.A(g16158),.B(g30082));
  NOR2 NOR2_1653(.VSS(VSS),.VDD(VDD),.Y(g30250),.A(g16163),.B(g30083));
  NOR2 NOR2_1654(.VSS(VSS),.VDD(VDD),.Y(g30251),.A(g16198),.B(g30085));
  NOR2 NOR2_1655(.VSS(VSS),.VDD(VDD),.Y(g30252),.A(g16217),.B(g30086));
  NOR2 NOR2_1656(.VSS(VSS),.VDD(VDD),.Y(g30253),.A(g16222),.B(g30087));
  NOR2 NOR2_1657(.VSS(VSS),.VDD(VDD),.Y(g30254),.A(g16242),.B(g30088));
  NOR2 NOR2_1658(.VSS(VSS),.VDD(VDD),.Y(g30255),.A(g16263),.B(g30089));
  NOR2 NOR2_1659(.VSS(VSS),.VDD(VDD),.Y(g30256),.A(g16282),.B(g30090));
  NOR2 NOR2_1660(.VSS(VSS),.VDD(VDD),.Y(g30257),.A(g16290),.B(g30091));
  NOR2 NOR2_1661(.VSS(VSS),.VDD(VDD),.Y(g30258),.A(g16291),.B(g30092));
  NOR2 NOR2_1662(.VSS(VSS),.VDD(VDD),.Y(g30259),.A(g16301),.B(g30093));
  NOR2 NOR2_1663(.VSS(VSS),.VDD(VDD),.Y(g30260),.A(g16322),.B(g30094));
  NOR2 NOR2_1664(.VSS(VSS),.VDD(VDD),.Y(g30261),.A(g16342),.B(g30095));
  NOR2 NOR2_1665(.VSS(VSS),.VDD(VDD),.Y(g30262),.A(g16343),.B(g30096));
  NOR2 NOR2_1666(.VSS(VSS),.VDD(VDD),.Y(g30263),.A(g16344),.B(g30097));
  NOR2 NOR2_1667(.VSS(VSS),.VDD(VDD),.Y(g30264),.A(g16348),.B(g30098));
  NOR2 NOR2_1668(.VSS(VSS),.VDD(VDD),.Y(g30265),.A(g16349),.B(g30099));
  NOR2 NOR2_1669(.VSS(VSS),.VDD(VDD),.Y(g30266),.A(g16359),.B(g30100));
  NOR2 NOR2_1670(.VSS(VSS),.VDD(VDD),.Y(g30267),.A(g16380),.B(g30101));
  NOR2 NOR2_1671(.VSS(VSS),.VDD(VDD),.Y(g30268),.A(g16382),.B(g30102));
  NOR2 NOR2_1672(.VSS(VSS),.VDD(VDD),.Y(g30269),.A(g16386),.B(g30103));
  NOR2 NOR2_1673(.VSS(VSS),.VDD(VDD),.Y(g30270),.A(g16387),.B(g30104));
  NOR2 NOR2_1674(.VSS(VSS),.VDD(VDD),.Y(g30271),.A(g16388),.B(g30105));
  NOR2 NOR2_1675(.VSS(VSS),.VDD(VDD),.Y(g30272),.A(g16392),.B(g30106));
  NOR2 NOR2_1676(.VSS(VSS),.VDD(VDD),.Y(g30273),.A(g16393),.B(g30107));
  NOR2 NOR2_1677(.VSS(VSS),.VDD(VDD),.Y(g30274),.A(g16403),.B(g30108));
  NOR2 NOR2_1678(.VSS(VSS),.VDD(VDD),.Y(g30275),.A(g16413),.B(g30109));
  NOR2 NOR2_1679(.VSS(VSS),.VDD(VDD),.Y(g30276),.A(g16415),.B(g30110));
  NOR2 NOR2_1680(.VSS(VSS),.VDD(VDD),.Y(g30277),.A(g16418),.B(g30111));
  NOR2 NOR2_1681(.VSS(VSS),.VDD(VDD),.Y(g30278),.A(g16420),.B(g30112));
  NOR2 NOR2_1682(.VSS(VSS),.VDD(VDD),.Y(g30279),.A(g16424),.B(g30113));
  NOR2 NOR2_1683(.VSS(VSS),.VDD(VDD),.Y(g30280),.A(g16425),.B(g30114));
  NOR2 NOR2_1684(.VSS(VSS),.VDD(VDD),.Y(g30281),.A(g16426),.B(g30115));
  NOR2 NOR2_1685(.VSS(VSS),.VDD(VDD),.Y(g30282),.A(g16430),.B(g30117));
  NOR2 NOR2_1686(.VSS(VSS),.VDD(VDD),.Y(g30283),.A(g16431),.B(g30118));
  NOR2 NOR2_1687(.VSS(VSS),.VDD(VDD),.Y(g30284),.A(g16444),.B(g29980));
  NOR2 NOR2_1688(.VSS(VSS),.VDD(VDD),.Y(g30285),.A(g16447),.B(g29981));
  NOR2 NOR2_1689(.VSS(VSS),.VDD(VDD),.Y(g30286),.A(g16449),.B(g29982));
  NOR2 NOR2_1690(.VSS(VSS),.VDD(VDD),.Y(g30287),.A(g16452),.B(g29983));
  NOR2 NOR2_1691(.VSS(VSS),.VDD(VDD),.Y(g30288),.A(g16454),.B(g29984));
  NOR2 NOR2_1692(.VSS(VSS),.VDD(VDD),.Y(g30289),.A(g16458),.B(g29985));
  NOR2 NOR2_1693(.VSS(VSS),.VDD(VDD),.Y(g30290),.A(g16459),.B(g29986));
  NOR2 NOR2_1694(.VSS(VSS),.VDD(VDD),.Y(g30291),.A(g16460),.B(g29987));
  NOR2 NOR2_1695(.VSS(VSS),.VDD(VDD),.Y(g30292),.A(g13477),.B(g29988));
  NOR2 NOR2_1696(.VSS(VSS),.VDD(VDD),.Y(g30293),.A(g13480),.B(g29989));
  NOR2 NOR2_1697(.VSS(VSS),.VDD(VDD),.Y(g30294),.A(g13483),.B(g29990));
  NOR2 NOR2_1698(.VSS(VSS),.VDD(VDD),.Y(g30295),.A(g13485),.B(g29991));
  NOR2 NOR2_1699(.VSS(VSS),.VDD(VDD),.Y(g30296),.A(g13488),.B(g29993));
  NOR2 NOR2_1700(.VSS(VSS),.VDD(VDD),.Y(g30297),.A(g13490),.B(g29994));
  NOR2 NOR2_1701(.VSS(VSS),.VDD(VDD),.Y(g30298),.A(g13496),.B(g29995));
  NOR2 NOR2_1702(.VSS(VSS),.VDD(VDD),.Y(g30299),.A(g13499),.B(g29996));
  NOR2 NOR2_1703(.VSS(VSS),.VDD(VDD),.Y(g30300),.A(g13502),.B(g30001));
  NOR2 NOR2_1704(.VSS(VSS),.VDD(VDD),.Y(g30301),.A(g13504),.B(g30002));
  NOR2 NOR2_1705(.VSS(VSS),.VDD(VDD),.Y(g30302),.A(g13513),.B(g30003));
  NOR2 NOR2_1706(.VSS(VSS),.VDD(VDD),.Y(g30303),.A(g13516),.B(g30005));
  NOR2 NOR2_1707(.VSS(VSS),.VDD(VDD),.Y(g30304),.A(g13527),.B(g30007));
  NOR2 NOR2_1708(.VSS(VSS),.VDD(VDD),.Y(g30338),.A(g14297),.B(g30225));
  NOR2 NOR2_1709(.VSS(VSS),.VDD(VDD),.Y(g30341),.A(g14328),.B(g30226));
  NOR2 NOR2_1710(.VSS(VSS),.VDD(VDD),.Y(g30356),.A(g14419),.B(g30227));
  NOR2 NOR2_1711(.VSS(VSS),.VDD(VDD),.Y(g30399),.A(g30116),.B(g30123));
  NOR2 NOR2_1712(.VSS(VSS),.VDD(VDD),.Y(g30400),.A(g29997),.B(g30127));
  NOR2 NOR2_1713(.VSS(VSS),.VDD(VDD),.Y(g30401),.A(g29998),.B(g30128));
  NOR2 NOR2_1714(.VSS(VSS),.VDD(VDD),.Y(g30402),.A(g29999),.B(g30129));
  NOR2 NOR2_1715(.VSS(VSS),.VDD(VDD),.Y(g30403),.A(g30004),.B(g30131));
  NOR2 NOR2_1716(.VSS(VSS),.VDD(VDD),.Y(g30404),.A(g30006),.B(g30132));
  NOR2 NOR2_1717(.VSS(VSS),.VDD(VDD),.Y(g30405),.A(g30008),.B(g30133));
  NOR2 NOR2_1718(.VSS(VSS),.VDD(VDD),.Y(g30406),.A(g30009),.B(g30138));
  NOR2 NOR2_1719(.VSS(VSS),.VDD(VDD),.Y(g30455),.A(g13953),.B(g30216));
  NOR2 NOR2_1720(.VSS(VSS),.VDD(VDD),.Y(g30468),.A(g14007),.B(g30217));
  NOR2 NOR2_1721(.VSS(VSS),.VDD(VDD),.Y(g30470),.A(g14023),.B(g30218));
  NOR2 NOR2_1722(.VSS(VSS),.VDD(VDD),.Y(g30482),.A(g14067),.B(g30219));
  NOR2 NOR2_1723(.VSS(VSS),.VDD(VDD),.Y(g30485),.A(g14098),.B(g30220));
  NOR2 NOR2_1724(.VSS(VSS),.VDD(VDD),.Y(g30487),.A(g14114),.B(g30221));
  NOR2 NOR2_1725(.VSS(VSS),.VDD(VDD),.Y(g30500),.A(g14182),.B(g30222));
  NOR2 NOR2_1726(.VSS(VSS),.VDD(VDD),.Y(g30503),.A(g14213),.B(g30223));
  NOR2 NOR2_1727(.VSS(VSS),.VDD(VDD),.Y(g30505),.A(g14229),.B(g30224));
  NOR2 NOR2_1728(.VSS(VSS),.VDD(VDD),.Y(g30566),.A(g14327),.B(g30398));
  NOR2 NOR2_1729(.VSS(VSS),.VDD(VDD),.Y(g30584),.A(g30412),.B(g2611));
  NOR3 NOR3_409(.VSS(VSS),.VDD(VDD),.Y(g30588),.A(g6119),.B(g30412),.C(g25353));
  NOR2 NOR2_1730(.VSS(VSS),.VDD(VDD),.Y(g30593),.A(g30412),.B(g2603));
  NOR3 NOR3_410(.VSS(VSS),.VDD(VDD),.Y(g30594),.A(g6119),.B(g30412),.C(g25419));
  NOR3 NOR3_411(.VSS(VSS),.VDD(VDD),.Y(g30597),.A(g6119),.B(g30412),.C(g25341));
  NOR2 NOR2_1731(.VSS(VSS),.VDD(VDD),.Y(g30601),.A(g30412),.B(g2604));
  NOR3 NOR3_412(.VSS(VSS),.VDD(VDD),.Y(g30602),.A(g6119),.B(g30412),.C(g25417));
  NOR3 NOR3_413(.VSS(VSS),.VDD(VDD),.Y(g30605),.A(g6119),.B(g30412),.C(g25333));
  NOR2 NOR2_1732(.VSS(VSS),.VDD(VDD),.Y(g30608),.A(g30412),.B(g2605));
  NOR2 NOR2_1733(.VSS(VSS),.VDD(VDD),.Y(g30609),.A(g30412),.B(g2606));
  NOR3 NOR3_414(.VSS(VSS),.VDD(VDD),.Y(g30610),.A(g6119),.B(g30412),.C(g25411));
  NOR2 NOR2_1734(.VSS(VSS),.VDD(VDD),.Y(g30613),.A(g30412),.B(g2607));
  NOR3 NOR3_415(.VSS(VSS),.VDD(VDD),.Y(g30614),.A(g6119),.B(g30412),.C(g25403));
  NOR2 NOR2_1735(.VSS(VSS),.VDD(VDD),.Y(g30617),.A(g23850),.B(g30412));
  NOR2 NOR2_1736(.VSS(VSS),.VDD(VDD),.Y(g30618),.A(g30412),.B(g25449));
  NOR2 NOR2_1737(.VSS(VSS),.VDD(VDD),.Y(g30621),.A(g30412),.B(g2608));
  NOR3 NOR3_416(.VSS(VSS),.VDD(VDD),.Y(g30622),.A(g6119),.B(g30412),.C(g25393));
  NOR2 NOR2_1738(.VSS(VSS),.VDD(VDD),.Y(g30625),.A(g30412),.B(g24660));
  NOR2 NOR2_1739(.VSS(VSS),.VDD(VDD),.Y(g30628),.A(g30412),.B(g2610));
  NOR3 NOR3_417(.VSS(VSS),.VDD(VDD),.Y(g30629),.A(g6119),.B(g30412),.C(g25378));
  NOR3 NOR3_418(.VSS(VSS),.VDD(VDD),.Y(g30632),.A(g6119),.B(g30412),.C(g25366));
  NOR2 NOR2_1740(.VSS(VSS),.VDD(VDD),.Y(g30635),.A(g16108),.B(g30407));
  NOR2 NOR2_1741(.VSS(VSS),.VDD(VDD),.Y(g30636),.A(g16140),.B(g30409));
  NOR2 NOR2_1742(.VSS(VSS),.VDD(VDD),.Y(g30637),.A(g16141),.B(g30410));
  NOR2 NOR2_1743(.VSS(VSS),.VDD(VDD),.Y(g30638),.A(g16159),.B(g30411));
  NOR2 NOR2_1744(.VSS(VSS),.VDD(VDD),.Y(g30639),.A(g16186),.B(g30436));
  NOR2 NOR2_1745(.VSS(VSS),.VDD(VDD),.Y(g30640),.A(g16187),.B(g30437));
  NOR2 NOR2_1746(.VSS(VSS),.VDD(VDD),.Y(g30641),.A(g16188),.B(g30438));
  NOR2 NOR2_1747(.VSS(VSS),.VDD(VDD),.Y(g30642),.A(g16199),.B(g30440));
  NOR2 NOR2_1748(.VSS(VSS),.VDD(VDD),.Y(g30643),.A(g16200),.B(g30441));
  NOR2 NOR2_1749(.VSS(VSS),.VDD(VDD),.Y(g30644),.A(g16218),.B(g30442));
  NOR2 NOR2_1750(.VSS(VSS),.VDD(VDD),.Y(g30645),.A(g16240),.B(g30444));
  NOR2 NOR2_1751(.VSS(VSS),.VDD(VDD),.Y(g30646),.A(g16241),.B(g30445));
  NOR2 NOR2_1752(.VSS(VSS),.VDD(VDD),.Y(g30647),.A(g16251),.B(g30447));
  NOR2 NOR2_1753(.VSS(VSS),.VDD(VDD),.Y(g30648),.A(g16252),.B(g30448));
  NOR2 NOR2_1754(.VSS(VSS),.VDD(VDD),.Y(g30649),.A(g16253),.B(g30449));
  NOR2 NOR2_1755(.VSS(VSS),.VDD(VDD),.Y(g30650),.A(g16264),.B(g30451));
  NOR2 NOR2_1756(.VSS(VSS),.VDD(VDD),.Y(g30651),.A(g16265),.B(g30452));
  NOR2 NOR2_1757(.VSS(VSS),.VDD(VDD),.Y(g30652),.A(g16283),.B(g30453));
  NOR2 NOR2_1758(.VSS(VSS),.VDD(VDD),.Y(g30653),.A(g16289),.B(g30454));
  NOR2 NOR2_1759(.VSS(VSS),.VDD(VDD),.Y(g30654),.A(g16299),.B(g30457));
  NOR2 NOR2_1760(.VSS(VSS),.VDD(VDD),.Y(g30655),.A(g16300),.B(g30458));
  NOR2 NOR2_1761(.VSS(VSS),.VDD(VDD),.Y(g30656),.A(g16310),.B(g30460));
  NOR2 NOR2_1762(.VSS(VSS),.VDD(VDD),.Y(g30657),.A(g16311),.B(g30461));
  NOR2 NOR2_1763(.VSS(VSS),.VDD(VDD),.Y(g30658),.A(g16312),.B(g30462));
  NOR2 NOR2_1764(.VSS(VSS),.VDD(VDD),.Y(g30659),.A(g16323),.B(g30464));
  NOR2 NOR2_1765(.VSS(VSS),.VDD(VDD),.Y(g30660),.A(g16324),.B(g30465));
  NOR2 NOR2_1766(.VSS(VSS),.VDD(VDD),.Y(g30661),.A(g16345),.B(g30467));
  NOR2 NOR2_1767(.VSS(VSS),.VDD(VDD),.Y(g30662),.A(g16347),.B(g30469));
  NOR2 NOR2_1768(.VSS(VSS),.VDD(VDD),.Y(g30663),.A(g16357),.B(g30472));
  NOR2 NOR2_1769(.VSS(VSS),.VDD(VDD),.Y(g30664),.A(g16358),.B(g30473));
  NOR2 NOR2_1770(.VSS(VSS),.VDD(VDD),.Y(g30665),.A(g16368),.B(g30475));
  NOR2 NOR2_1771(.VSS(VSS),.VDD(VDD),.Y(g30666),.A(g16369),.B(g30476));
  NOR2 NOR2_1772(.VSS(VSS),.VDD(VDD),.Y(g30667),.A(g16370),.B(g30477));
  NOR2 NOR2_1773(.VSS(VSS),.VDD(VDD),.Y(g30668),.A(g16381),.B(g30478));
  NOR2 NOR2_1774(.VSS(VSS),.VDD(VDD),.Y(g30669),.A(g16383),.B(g30481));
  NOR2 NOR2_1775(.VSS(VSS),.VDD(VDD),.Y(g30670),.A(g16389),.B(g30484));
  NOR2 NOR2_1776(.VSS(VSS),.VDD(VDD),.Y(g30671),.A(g16391),.B(g30486));
  NOR2 NOR2_1777(.VSS(VSS),.VDD(VDD),.Y(g30672),.A(g16401),.B(g30489));
  NOR2 NOR2_1778(.VSS(VSS),.VDD(VDD),.Y(g30673),.A(g16402),.B(g30490));
  NOR2 NOR2_1779(.VSS(VSS),.VDD(VDD),.Y(g30674),.A(g16414),.B(g30492));
  NOR2 NOR2_1780(.VSS(VSS),.VDD(VDD),.Y(g30675),.A(g16416),.B(g30495));
  NOR2 NOR2_1781(.VSS(VSS),.VDD(VDD),.Y(g30676),.A(g16419),.B(g30496));
  NOR2 NOR2_1782(.VSS(VSS),.VDD(VDD),.Y(g30677),.A(g16421),.B(g30499));
  NOR2 NOR2_1783(.VSS(VSS),.VDD(VDD),.Y(g30678),.A(g16427),.B(g30502));
  NOR2 NOR2_1784(.VSS(VSS),.VDD(VDD),.Y(g30679),.A(g16429),.B(g30504));
  NOR2 NOR2_1785(.VSS(VSS),.VDD(VDD),.Y(g30680),.A(g16443),.B(g30327));
  NOR2 NOR2_1786(.VSS(VSS),.VDD(VDD),.Y(g30681),.A(g16448),.B(g30330));
  NOR2 NOR2_1787(.VSS(VSS),.VDD(VDD),.Y(g30682),.A(g16450),.B(g30333));
  NOR2 NOR2_1788(.VSS(VSS),.VDD(VDD),.Y(g30683),.A(g16453),.B(g30334));
  NOR2 NOR2_1789(.VSS(VSS),.VDD(VDD),.Y(g30684),.A(g16455),.B(g30337));
  NOR3 NOR3_419(.VSS(VSS),.VDD(VDD),.Y(g30685),.A(g29992),.B(g30000),.C(g30372));
  NOR2 NOR2_1790(.VSS(VSS),.VDD(VDD),.Y(g30686),.A(g16461),.B(g30340));
  NOR2 NOR2_1791(.VSS(VSS),.VDD(VDD),.Y(g30687),.A(g13479),.B(g30345));
  NOR2 NOR2_1792(.VSS(VSS),.VDD(VDD),.Y(g30688),.A(g13484),.B(g30348));
  NOR2 NOR2_1793(.VSS(VSS),.VDD(VDD),.Y(g30689),.A(g13486),.B(g30351));
  NOR2 NOR2_1794(.VSS(VSS),.VDD(VDD),.Y(g30690),.A(g13489),.B(g30352));
  NOR2 NOR2_1795(.VSS(VSS),.VDD(VDD),.Y(g30691),.A(g13491),.B(g30355));
  NOR2 NOR2_1796(.VSS(VSS),.VDD(VDD),.Y(g30692),.A(g13498),.B(g30361));
  NOR2 NOR2_1797(.VSS(VSS),.VDD(VDD),.Y(g30693),.A(g13503),.B(g30364));
  NOR2 NOR2_1798(.VSS(VSS),.VDD(VDD),.Y(g30694),.A(g13505),.B(g30367));
  NOR2 NOR2_1799(.VSS(VSS),.VDD(VDD),.Y(g30695),.A(g13515),.B(g30374));
  NOR2 NOR2_1800(.VSS(VSS),.VDD(VDD),.Y(g30699),.A(g13914),.B(g30387));
  NOR2 NOR2_1801(.VSS(VSS),.VDD(VDD),.Y(g30700),.A(g13952),.B(g30388));
  NOR2 NOR2_1802(.VSS(VSS),.VDD(VDD),.Y(g30701),.A(g13970),.B(g30389));
  NOR2 NOR2_1803(.VSS(VSS),.VDD(VDD),.Y(g30702),.A(g14006),.B(g30390));
  NOR2 NOR2_1804(.VSS(VSS),.VDD(VDD),.Y(g30703),.A(g14022),.B(g30391));
  NOR2 NOR2_1805(.VSS(VSS),.VDD(VDD),.Y(g30704),.A(g14040),.B(g30392));
  NOR2 NOR2_1806(.VSS(VSS),.VDD(VDD),.Y(g30705),.A(g14097),.B(g30393));
  NOR2 NOR2_1807(.VSS(VSS),.VDD(VDD),.Y(g30706),.A(g14113),.B(g30394));
  NOR2 NOR2_1808(.VSS(VSS),.VDD(VDD),.Y(g30707),.A(g14131),.B(g30395));
  NOR2 NOR2_1809(.VSS(VSS),.VDD(VDD),.Y(g30708),.A(g14212),.B(g30396));
  NOR2 NOR2_1810(.VSS(VSS),.VDD(VDD),.Y(g30709),.A(g14228),.B(g30397));
  NOR2 NOR2_1811(.VSS(VSS),.VDD(VDD),.Y(g30780),.A(g30625),.B(g22387));
  NOR2 NOR2_1812(.VSS(VSS),.VDD(VDD),.Y(g30783),.A(g30618),.B(g22387));
  NOR2 NOR2_1813(.VSS(VSS),.VDD(VDD),.Y(g30785),.A(g30618),.B(g22387));
  NOR2 NOR2_1814(.VSS(VSS),.VDD(VDD),.Y(g30786),.A(g30625),.B(g22387));
  NOR2 NOR2_1815(.VSS(VSS),.VDD(VDD),.Y(g30787),.A(g30594),.B(g22387));
  NOR2 NOR2_1816(.VSS(VSS),.VDD(VDD),.Y(g30788),.A(g30602),.B(g22387));
  NOR2 NOR2_1817(.VSS(VSS),.VDD(VDD),.Y(g30789),.A(g30575),.B(g22387));
  NOR2 NOR2_1818(.VSS(VSS),.VDD(VDD),.Y(g30790),.A(g30575),.B(g22387));
  NOR2 NOR2_1819(.VSS(VSS),.VDD(VDD),.Y(g30796),.A(g16069),.B(g30696));
  NOR2 NOR2_1820(.VSS(VSS),.VDD(VDD),.Y(g30798),.A(g16134),.B(g30697));
  NOR2 NOR2_1821(.VSS(VSS),.VDD(VDD),.Y(g30801),.A(g16237),.B(g30698));
  NOR2 NOR2_1822(.VSS(VSS),.VDD(VDD),.Y(g30929),.A(g30728),.B(g30736));
  NOR2 NOR2_1823(.VSS(VSS),.VDD(VDD),.Y(g30930),.A(g30735),.B(g30744));
  NOR2 NOR2_1824(.VSS(VSS),.VDD(VDD),.Y(g30931),.A(g30743),.B(g30750));
  NOR2 NOR2_1825(.VSS(VSS),.VDD(VDD),.Y(g30932),.A(g30754),.B(g30757));
  NOR2 NOR2_1826(.VSS(VSS),.VDD(VDD),.Y(g30933),.A(g30755),.B(g30758));
  NOR2 NOR2_1827(.VSS(VSS),.VDD(VDD),.Y(g30934),.A(g30759),.B(g30761));
  NOR2 NOR2_1828(.VSS(VSS),.VDD(VDD),.Y(g30935),.A(g30760),.B(g30762));
  NOR2 NOR2_1829(.VSS(VSS),.VDD(VDD),.Y(g30936),.A(g30763),.B(g30764));
  NOR2 NOR2_1830(.VSS(VSS),.VDD(VDD),.Y(g30954),.A(g30916),.B(g30944));
  NOR2 NOR2_1831(.VSS(VSS),.VDD(VDD),.Y(g30955),.A(g30918),.B(g30945));
  NOR2 NOR2_1832(.VSS(VSS),.VDD(VDD),.Y(g30956),.A(g30919),.B(g30946));
  NOR2 NOR2_1833(.VSS(VSS),.VDD(VDD),.Y(g30957),.A(g30920),.B(g30947));
  NOR2 NOR2_1834(.VSS(VSS),.VDD(VDD),.Y(g30958),.A(g30922),.B(g30948));
  NOR2 NOR2_1835(.VSS(VSS),.VDD(VDD),.Y(g30959),.A(g30923),.B(g30949));
  NOR2 NOR2_1836(.VSS(VSS),.VDD(VDD),.Y(g30960),.A(g30924),.B(g30950));
  NOR2 NOR2_1837(.VSS(VSS),.VDD(VDD),.Y(g30961),.A(g30925),.B(g30951));
  NOR3 NOR3_420(.VSS(VSS),.VDD(VDD),.Y(g30970),.A(g30917),.B(g30921),.C(g30953));

endmodule