module s1585(g6271,g2612,g46,g4205,g886,g6269,g4888,g6266,g93,g4181,g904,g7744,g6256,g4201,g4209,g88,g907,g4175,g9451,g2610,g6278,g10455,g6942,g6270,g1700,g10461,g104,g10459,g6275,g6253,g1203,g4171,g1696,g4212,g1173,g4198,g6926,g10377,g8979,VDD,g743,g4194,g6259,g6285,g8323,g889,g4210,g6264,g3069,g6284,g6842,g919,g18,g8984,g1185,g29,g92,g6283,g10457,g11163,g6280,g2609,g89,g6258,g8563,g8331,g1194,g103,g10801,g11489,g8565,g95,g2604,g2607,g6254,g8328,g8981,g4179,g2355,g31,g4176,g1712,g1188,g4180,g925,g4887,g881,g8318,g6260,g5659,g8976,g6262,g4208,g4204,g895,g8564,g1176,g4172,g8347,g47,g8352,g8561,g872,g910,g4195,g6263,g6955,g8978,g4211,g3007,g5816,g4196,g6273,g94,g6257,g6274,g4191,g8313,g41,g101,g4200,g4215,g913,g42,g10379,g4193,g8062,g5658,g6268,g6281,g4192,g877,g4216,g750,g10465,g2606,g6261,g1961,g1179,g8335,g1182,g4199,g898,g6932,g96,g3327,g4173,g916,g10628,g100,g4202,g6279,g2605,g901,g27,g99,g741,g43,g742,g5105,g6267,g45,g1200,g2648,g4178,g84,g8349,g1960,g8986,g2986,g10463,g87,g30,g6276,g8566,g8316,g82,g892,g2608,g4174,g44,g6282,g6949,g1191,g90,g23,g744,g1957,g9961,g2611,g86,g8271,g1197,g8061,g4203,g6255,g8983,g83,g6920,g109,g2601,g11206,g102,g4214,g6272,g91,g4197,g8340,g4213,g4207,g85,g2602,g922,g8982,g1170,g8562,g5101,g8980,g48,g873,g6277,VSS,g6265,g8977,g2603,g8985,CLOCK,g4177,g4206,g28);
input g46,g886,g93,g904,g88,g907,g1700,g104,g1203,g1696,g1173,VDD,g743,g889,g919,g18,g1185,g29,g92,g89,g1194,g103,g95,g31,g1712,g1188,g925,g881,g895,g1176,g47,g872,g910,g94,g41,g101,g913,g42,g877,g750,g1961,g1179,g1182,g898,g96,g916,g100,g901,g27,g99,g741,g43,g742,g45,g1200,g84,g1960,g87,g30,g82,g892,g44,g1191,g90,g23,g744,g86,g1197,g83,g109,g102,g91,g85,g922,g1170,g48,g873,VSS,CLOCK,g28;
output g6271,g2612,g4205,g6269,g4888,g6266,g4181,g7744,g6256,g4201,g4209,g4175,g9451,g2610,g6278,g10455,g6942,g6270,g10461,g10459,g6275,g6253,g4171,g4212,g4198,g6926,g10377,g8979,g4194,g6259,g6285,g8323,g4210,g6264,g3069,g6284,g6842,g8984,g6283,g10457,g11163,g6280,g2609,g6258,g8563,g8331,g10801,g11489,g8565,g2604,g2607,g6254,g8328,g8981,g4179,g2355,g4176,g4180,g4887,g8318,g6260,g5659,g8976,g6262,g4208,g4204,g8564,g4172,g8347,g8352,g8561,g4195,g6263,g6955,g8978,g4211,g3007,g5816,g4196,g6273,g6257,g6274,g4191,g8313,g4200,g4215,g10379,g4193,g8062,g5658,g6268,g6281,g4192,g4216,g10465,g2606,g6261,g8335,g4199,g6932,g3327,g4173,g10628,g4202,g6279,g2605,g5105,g6267,g2648,g4178,g8349,g8986,g2986,g10463,g6276,g8566,g8316,g2608,g4174,g6282,g6949,g1957,g9961,g2611,g8271,g8061,g4203,g6255,g8983,g6920,g2601,g11206,g4214,g6272,g4197,g8340,g4213,g4207,g2602,g8982,g8562,g5101,g8980,g6277,g6265,g8977,g2603,g8985,g4177,g4206;

  wire g9968,g10200,g3474,g3333,g7021,I5174,I11638,g2418,g7535,g98,g2896,I10834,I17297,g3462,g10763,g7071,I7478,I15263,g5637,g8002,I9574,I8872,g8464,g4908,g8812,I13945,g8408,g10718,I13376,g6462,g8569,g10243,g4746,g4313,g7593,I11444,I13320,I8480,I10904,g76,g5253,g1864,I7260,g6103,g6114,g3626,g4392,g2652,g5528,g9088,g8139,g11438,g9935,g7809,g10390,g6070,g534,g8001,g10449,I4948,I9359,I15335,g6704,I14645,I5684,I11668,g11581,I15225,g10275,g758,g5121,g11646,I13478,I6356,g7882,g8792,g7632,g6236,g1992,I8652,g7719,I9930,I11833,g11246,g7992,I13794,g7119,g9706,g363,g9888,g8639,g4891,g10542,g7113,I15082,I10678,g9958,I12162,g2905,I12776,I9519,g10324,g4585,g8076,I6985,g2895,I11515,g3880,I9773,I13284,g3793,I16295,I15500,g3995,g3411,g10044,I13354,g2179,g10874,I13744,I17681,I16982,g8776,I12126,g2039,g7142,g2645,g2903,I6778,I11701,g7537,I11115,g9903,I5667,g9895,I14257,I7820,g10142,g1089,I5878,g1586,I9174,g7319,g6055,g7618,g6342,I15763,I13027,I4906,g11323,g6706,g7042,I8259,I17112,I12451,g10300,g6387,g2514,g11389,g7242,I17447,I12631,g7749,g6713,g11175,g5878,g11605,I5136,I15589,I5555,g3383,g456,g9809,g5345,g9361,g11416,I8473,g256,g2651,g10220,g11588,g11373,g8616,g7337,g9609,I16496,g8200,g2916,I15491,g10395,I4942,g3219,g5999,g1515,g4943,g2330,g10545,g4305,g3761,g11461,g10199,g9747,I15287,I12229,I11049,g11183,g560,g10187,g11092,g4424,I13293,g4767,g4098,I8436,g4312,g10550,I12616,I8740,g5521,I17161,g5753,I14678,g7848,g3098,I8178,g6739,g6073,g5236,I7923,g8239,g386,g3061,g4360,I8751,I17666,g4164,g9943,g6708,g5598,I16571,I8780,g8279,I12907,g6182,g2650,g2981,I13036,I6436,g4258,I12062,g10878,g4428,g3432,g3037,I7694,g9317,g10679,g6517,g4966,g4373,I7140,I9525,I11420,g2586,I10759,g10866,I6794,I5830,I11494,I17116,g6890,I17395,g2802,g2814,g5104,I5812,g4801,I15609,g10571,g5511,I7909,I4992,g10879,I16735,g8267,g9848,g11304,I12978,I5740,g7048,I5430,I14585,g6554,g7754,I13388,g5052,I15752,I5891,I8730,I7348,g6837,g9269,g8758,g9431,I6037,g2206,g4414,I14642,g7598,I17704,g8174,g1975,g9576,g2970,I6289,g11224,I5403,g2047,g8889,g1601,I7372,g9892,g9266,g4997,g4114,g932,I10078,g182,g11107,g8276,g9868,I7236,g8400,g2256,I17146,I8324,g11046,g5145,g6709,I10858,g3860,g4363,g4400,g4364,g9612,I6448,g1240,g10261,I11261,g7887,I17243,I16641,I13347,g7963,g6030,g5484,I7931,I8877,g4721,I6815,g8154,g7101,g5493,I15353,g7964,g7548,g10482,I7465,g4401,I10150,I8231,g6135,g5169,g9587,I5449,I16015,g7753,g2547,g10320,I12296,g10401,I15229,I8123,I11155,g8390,g4580,I7964,g4156,I8795,g8886,g8795,g3354,g5037,g7915,I11204,g1056,g4673,I9008,g11194,g2838,g5395,g8515,g11455,g6177,g8301,g4589,g8096,g6224,I11659,g10323,I13627,g6099,g7066,g7409,g7946,g10134,g4399,g4492,g1362,I5007,I5593,g9818,g5148,I12226,I5599,g7779,I6989,I7810,g6653,g4458,g9813,I12577,g10698,I15400,g9947,g3997,g7082,g6647,I13660,g4362,I10024,g9990,g8072,I12061,g2707,I10012,I13595,I7205,g587,g553,g4272,I13122,I15617,g6027,I5343,I6220,g5650,I5641,g6796,g5815,g6327,g7567,I10072,g4631,I14370,g3753,I16647,I10144,g5116,g2081,g5421,g9430,I10563,I7109,g1466,g119,g3399,g10667,g9836,g9847,g5981,I9947,g10366,g4836,g8262,g5900,g7536,g9889,I9168,I7752,g5856,g7985,g2228,g6403,I14376,g2864,g7196,g4719,g3095,g8300,g9025,g4242,I11845,g2854,I13822,g10293,g11290,g4715,g4560,g11180,I9483,g7896,I5549,g9362,I17552,I12523,I17486,g10671,I7639,g7273,I9383,I10484,g7269,g3212,g9611,g9700,g1571,g11214,g2208,g5088,g5642,I11725,I13409,g3500,I4900,I7194,g11328,g8363,I13406,g8028,g1537,I11272,g113,g2075,g4445,g10425,I11286,g10733,g2749,g5004,g5497,I7735,g8306,g1645,g11446,I17672,I17188,I15461,I11140,g8148,g11270,I13583,I5677,g10117,g5697,I8514,g7619,g9967,g10883,g11626,I6962,I8328,g6056,g5284,I15704,g2242,g5683,g2904,I14835,g6572,g2246,g9726,g11332,g999,I15994,g8110,g10269,g7259,I5325,g7190,g10235,I6611,g11247,I10520,I12156,g9603,I7405,g8185,g6418,g5103,I6771,I4930,I16051,g6416,I12021,g2177,g7504,I7633,I12779,g5751,g4346,g5838,g5729,I10566,g4950,g9771,g5662,g3937,I15551,g6923,g4785,g8529,I11097,g5167,g1308,g1868,I7984,I9394,I5704,I16332,I16439,g3750,g3911,I6757,g11014,g5009,g2874,I15814,I16616,g11032,g11184,g10972,g5089,g2792,I9783,g11468,I12843,g6859,g5278,g10655,I17470,I11109,g10262,I9869,g2250,g5291,g9733,I5282,g8510,I12174,g4292,I14681,g8736,g3272,I16407,I12598,I17155,I8640,g8315,I15371,g10929,g10050,I10374,g5996,g10911,g3412,g682,g10318,g11430,g7730,g10394,I8476,I17213,g7939,g435,I16298,I17315,g10794,g2302,g4613,I10201,g8754,g4051,I13266,g7243,g5888,g7573,g6990,g5068,g8025,g10970,g35,g4221,g7751,g7845,I17642,g10591,g3121,g1527,I15741,g9474,g10876,I16546,I8996,g10629,I13020,g7217,g10127,g11221,I8590,I12376,g11051,g3512,g8280,g7741,g9950,I13975,g4241,I12040,g1984,I7176,I10538,g6715,I6733,g5994,g10228,g11459,g3737,g8772,I16950,g8701,g11414,I5579,I10831,I8290,I15476,g7317,I16670,g7007,I6432,I9935,I17549,g11338,I12400,g1393,g10621,I15858,g1918,g5879,I13825,g1508,g11633,g11372,I10087,g9865,g8089,g8217,g9653,I17281,g11097,g10702,g4552,g11419,g11650,I16708,g11006,g3765,I15977,g2890,I17234,I9311,g5902,g10797,g11192,I7043,g6084,g5475,g6424,g11263,g11024,g8552,g9010,g10310,g6500,g7127,g5149,g7344,g4229,g6547,g10336,g1610,I13636,g7712,g4440,g2095,I10901,g7610,g5814,I15317,g5800,I15604,I13273,g3908,g5702,g10205,g9828,g7067,I8865,g814,g4223,g11227,g11234,I12454,g5802,I11433,g9602,g6453,g11055,I12460,g1958,g6362,g5626,g2920,g4515,I9557,I10243,g6593,g5587,g8362,g2821,g11630,g10724,g11230,g5527,g4470,g10126,g6287,g3622,I6676,g11249,g8106,g4676,g7256,g4900,I8403,g5486,g4525,g3369,g8358,g4449,g1936,g4182,I12601,g11634,g4228,g2742,g4220,g2164,I4883,I14944,g5992,g2267,I9352,g4352,I16644,I15583,I6428,g4905,I7779,I12046,I16691,I16331,I10388,I14873,I16484,g11411,g2772,g4739,g6438,g5226,g11497,g4441,g3207,g7466,I9662,g5690,g7706,g5813,g4320,g3351,I6761,I7396,g3491,g7911,g5784,g9572,g9831,I11909,g7340,g7527,g2997,g1318,g4048,I14955,I17053,g7430,g586,I5002,g10768,g8266,g4865,g9560,g11057,I9177,g11360,g3015,g10196,g731,g5401,I9905,g9516,g8253,g8199,I17051,g10206,g7615,g8588,g10094,g4526,I13436,g5025,I17394,g6695,g8759,g2755,g11492,I6150,g302,I7118,g8195,I11058,g7820,g9957,g2191,g10589,g4268,g5771,g9424,g7102,g4227,I6233,I5497,g114,g8240,g8073,g10728,g9386,g8093,g6337,g10732,I12910,I11405,g4884,I12137,g7804,I14217,I8529,I6034,g10858,I13260,I8215,g8574,g6077,g9689,g5644,g5514,g8970,g2261,I11879,g4161,I5348,g1327,g3756,g3328,I17327,g8488,I4943,I11351,I8442,g10799,I12759,g7617,I11135,I13991,g4559,g5350,g1776,g9855,I8589,g11145,g10563,g6069,g11613,g2325,g10069,g7775,g7134,g6892,g6323,g8255,g5069,g9605,g8882,I10204,g10711,I13335,g10240,g8483,g1923,I16161,g3397,g2462,g10272,g11047,g4328,I12712,g11499,I16160,g11471,I13332,g11306,I14442,g3528,g4907,g5758,g3119,I5940,I12832,g7522,g7944,g10873,I16261,I10349,g11327,g9291,g5544,I12421,I5600,g7572,g9258,g10579,g7061,g9849,g7656,I14690,g9852,g2647,I14358,g7777,I9368,I12835,g8146,g2014,g9761,g6196,I8576,g5773,I5383,I11191,g10760,g3380,g6221,g6119,I6664,I12424,I16525,g10309,g11463,g10504,g8545,g7085,g5817,g6128,g6887,I14939,g2200,g7265,I13791,I15542,g9817,g8149,g9452,I11817,g8557,g6673,g8425,g4254,I14549,I13714,I16363,g7092,g4456,I16847,g538,g5576,g8449,g1887,g7583,g10731,I7308,g6215,g11064,g11020,I6779,I13612,g8753,g7717,g2309,g4590,g2329,I5060,g9912,g3748,g3688,g6209,I7375,g444,I5725,I5976,g4001,g8648,I16475,g9512,I13545,I16289,g774,I16193,g8152,g3263,g3378,g6515,g11638,g5627,g7742,g10736,g11482,g9723,g1981,g6918,g8605,g2104,I6904,g9915,g4283,I8109,g4353,g1806,g6743,g4052,g4871,g7309,I12948,g2044,g1145,I11408,I5584,g11074,g2171,I5949,g1993,I5612,g2057,g4469,I9688,g4082,g5653,g4609,g709,g5111,g5210,I16623,g10236,g8576,g4538,g1482,g4870,g6198,g9427,g8734,I17261,g3719,g8010,I16635,I13301,I16802,g10497,g11054,g11050,g6661,g6228,g6412,I11608,g6648,I16528,I6421,g8162,I16682,I13538,I15403,g3329,g6983,g6559,g1470,g8424,g6015,g6074,g7503,g8143,I16283,I13233,I4924,g8355,g6527,g9713,I6449,g10784,I14884,g7923,g5917,I13902,I12683,I14127,g3904,I7865,I10477,g6193,g6652,g9923,g7785,g9597,g6111,g10238,g5190,I17306,I9371,I10105,I7707,g4236,I17761,g10150,g8702,g4603,I11037,g778,g2991,I9813,I6851,g10525,g3967,g8190,I13057,g7202,I10063,g10255,g8995,g7671,g9955,g3798,g5703,g8802,g9413,I12538,g956,g8263,g5864,g6841,g766,g6158,g4324,g10664,I15204,I17456,I8561,g8473,I10971,g7299,g4769,g10889,g5126,g9623,g8667,g8683,I17246,g10136,I7829,g521,g7592,g4276,I15452,g4775,I13717,g7733,g6242,g3810,g6529,g10120,I6938,g6741,I8772,g3209,g4088,g6336,g7188,I17701,g10778,g10345,g7585,I5792,I5751,g1781,I8631,I14242,g7051,g11245,g6639,g1998,g4553,I5044,g7402,g3414,g4712,g4476,g6751,I12466,g1982,g1038,g8045,g4308,I5015,g11272,g4989,g10490,I12268,I13669,g11034,I11034,I15266,g4385,I5893,g11506,g10805,I12004,g6325,g7952,g10488,I11079,I8268,g8290,g8415,g9509,I4979,g8875,g5767,I8462,I10659,g7144,I7233,I16944,g2135,g11333,I8004,I12113,I15209,g4096,g6912,g8931,g9535,g5608,g1415,g7786,g4387,g8858,g9409,g4013,g4915,I17698,g632,g6616,g8307,g5349,g3204,I17675,g6395,g9656,g3142,g5085,g2549,I9147,g8295,g5248,I14528,I16277,I5041,g11103,g5746,g4901,I12074,I6168,g7024,I16879,g3382,g8502,I6601,g7004,I15580,I13439,g10530,g6019,g10270,g348,g6088,g2793,g4992,g10154,g431,g11546,g5265,I14424,g6855,g5221,g9357,g5997,I13969,g5203,I8527,g6714,g8988,I8265,g7201,g8230,g11241,I5646,g11627,I11821,g6113,g11642,I6826,g2041,g10901,g6632,g4524,g2239,g3505,g8575,g4490,g7356,g2753,g10312,I16510,g5422,g496,g3991,I16550,g10891,I10698,g6332,g622,g9814,I12045,g6800,I5525,I16979,I15507,I11590,g4990,g7049,I12514,g10432,I15701,g6947,I4869,g2626,g9052,I11360,g11217,g5028,I16518,g4050,I13978,g2209,g8427,g6067,I5297,I16269,g8755,g1845,g8872,g8121,g10360,I10651,g8608,g9489,g11596,g6117,g8599,g2042,g5178,I15744,g1950,g7675,g7999,g7532,I4911,g7041,I10958,g2989,g5947,g9772,g5777,g11453,g9449,I8929,g7107,g2564,g10118,g11287,g1642,g10132,g9643,I9769,g8628,g8951,g10532,I13128,g4575,g8738,I15616,g10445,I4879,g7659,g8957,I16688,I16897,g10165,I16667,g10793,g1311,g248,I5478,g4724,g7519,g2229,g2475,g3385,I16046,g2480,I10006,g7147,I8903,I10810,I17152,g7745,g6752,I5317,I14295,g5189,g4078,I10165,g4319,g9311,I13206,g6156,g2054,I9424,g4505,g5295,I11929,g8136,g10472,g7209,g10551,g10486,g5882,g11377,g1987,I14364,g7814,g5821,g8186,g10141,g3101,g3291,I13314,g5914,g2037,I15176,g6450,I12499,g8589,g8066,I13096,I7659,g6898,g6640,I9779,g11215,I6055,g5938,I13091,g6426,g2012,I14194,I8739,I13307,g9921,g10893,g9995,g1624,g9657,I11122,g9926,g7058,g953,I17258,g8144,g4962,g3731,g6822,g7079,g5490,I7563,I15672,I5827,I8611,g7791,g11470,I11964,g11598,I12335,I10003,I12380,I11183,g8265,I6488,g7676,I5149,I15075,g2444,g11318,I10852,g4351,g6038,g5704,g10303,g611,I12205,g8003,g7633,g9909,g5515,g6319,g5397,g4330,g578,g1687,g1710,g991,I6861,g5919,I11299,g2984,g1663,g8684,g6589,g9739,g10905,g8773,I4903,I16169,g3255,g2827,g8229,g7040,g757,g2175,g874,I13412,g3759,I16577,I8007,g4999,g148,g3424,g10895,g8820,g2833,g1636,I11981,g8319,I11149,I9762,g10665,I12123,I16366,g5299,g213,I6447,g7436,g1059,g1169,I15717,g11335,g6595,I10099,g8161,g11294,I11773,g8718,g7799,g2067,g10161,g4762,g9930,g10346,g8399,g8413,g6485,g9613,g5840,I12418,I7509,g8465,g5830,I15079,g9608,I5916,g10444,g10936,g6621,g10321,I7202,g6312,g8158,g7203,g6888,I16853,g8268,I9896,I9391,g7972,I10898,g10487,I14277,g4348,I15775,g2090,g6566,g6470,I11572,g1098,g7802,g4339,I5410,g4006,g4806,g4464,g5824,g11444,I10289,g11094,I11232,g8270,g11273,g4060,g11160,g10462,g6299,g7780,g4572,g11151,I12553,g7308,g6087,g9732,I8835,I10840,g4421,g4486,g4550,g4969,g5504,I13858,g10620,g11182,g3389,g1607,g8434,g6818,g5147,g3980,g3693,I8543,I16098,g4287,g4430,I7390,g10186,g6200,g4873,g2118,g8477,I15374,g8787,g11286,g10906,g10251,g3003,I12878,I17350,g7470,I13806,I8315,g3391,I5500,I10075,g11426,g11518,g6583,g6625,g4723,I5363,g8641,g7296,g4261,I11450,g2454,I14506,g2022,g5276,g2994,I10521,I13571,g6334,g4396,I13068,I13308,g3913,g1690,g4816,I10861,g4277,g11157,g9416,I15708,g6180,I10702,g1651,g5204,I13868,g9268,g8138,g4437,g11147,I14519,I14561,I17387,g7607,g8532,g6392,g8209,g11462,g8703,g7783,g11208,g11049,g542,g6295,g6716,I9232,g5108,g8704,g10184,I11858,g10580,g9363,I6406,I9988,g7520,g9615,g339,g8814,g11165,g3415,g1872,I14373,I10639,g2271,I16148,I9213,g2353,I10302,g10821,I6654,g9670,g8170,I17510,g4010,g9620,I13869,g10676,g2957,g9097,I13448,g2105,g11169,g10454,g9725,g11503,g10149,g7937,g2909,g7826,I12186,g9861,I16742,I10042,I13618,g7981,g9111,g4967,g7707,I17393,g9683,I8449,g3710,g8600,g9414,I12790,g3938,g10685,I15510,I6988,I16023,I17540,g4130,g374,g11538,g8417,g5588,g6558,I16142,g4760,I10507,g7335,g1564,I13803,g9730,g9808,g4123,g3820,I16632,I6793,g8296,I10258,g10684,I17713,g8153,g11088,g5944,I5105,I7956,g6195,g8251,I9043,I10671,I13504,I12481,g7950,g9667,g11150,g2825,I6373,g2571,I15205,g6204,g589,g6361,g10051,g8880,g9880,I14271,g8181,I6631,g5443,g5317,g3429,I13265,g3086,g7927,g10328,g1462,I15514,g8751,g9,I12556,g6175,g263,g8443,I15072,g1814,g11044,I7743,I5672,I5960,I5847,g11084,g8585,g1032,g7123,I5057,g3400,I10081,I12607,g6315,g7497,I11531,g841,I11740,g7925,g2156,g2623,g1956,g7702,I12019,I15479,g2579,I16214,g4124,g1737,I8900,I5421,g8722,g5803,I17730,I6388,g4960,I5805,g6737,I16000,g6244,g2169,g9890,I12271,I17546,g11330,I16030,g3307,g8652,g7395,g1289,g8100,g8389,I14252,g10528,g7901,g7926,g9802,I15184,g1744,g5783,I9717,g8046,g5292,g7986,g8807,I6784,g794,I9388,g10700,I9575,g11583,g9697,g677,g4958,g7757,g4432,I6792,g11219,g11456,I5632,g2247,g7823,g10257,g8940,g10387,g2204,g631,g10111,g9750,g6904,I13245,I17271,I16863,g9029,g6524,g7324,g11391,g1750,I13894,g8219,g7997,g7245,I13738,g6442,I12517,g2760,I15494,g1419,g8078,g3306,g3260,I5989,g4495,I7899,g9974,g5474,g10933,g1973,g1212,g7983,g2024,g2515,g833,g2348,g8173,I7255,I13373,I8358,g9939,g3726,g10859,g6995,I7630,g5682,g5492,g2163,g3784,g1592,g3507,g818,g378,g7798,g9902,g9343,g4443,I15232,I9665,g11280,g4608,g4080,g5898,g2420,g11235,I6207,g10185,g10558,g6803,I14055,g8135,g8198,g6624,g5844,I12783,g3104,I7269,g6545,g3944,I16379,I5202,I17569,g8336,g6974,g4097,g9511,g10129,g7037,g4465,I15051,g4499,g5747,g64,g6645,g7625,I14385,I12484,g6577,g1357,g8382,I13341,g3050,g11439,g6240,g10715,I6495,g1580,I7790,g7388,g9364,I5126,g1007,I11731,g6994,I16074,g9699,I7280,g11072,I8943,g10536,g5687,g10107,I5979,g704,I7333,g3698,g4485,I12202,g10176,g5568,g10467,I6982,g4260,I16760,I16534,I12993,g11189,g1853,g5005,g3161,g9026,I16679,I9973,g10307,g6901,g6733,g10121,g7975,g4059,g8518,g3811,g2868,g6646,g5774,I10015,g9356,I15832,g3438,I17401,g8644,g10747,g7063,g3105,I14185,I13267,g2914,I13678,g10173,g6181,I9807,g4488,g10515,g3638,I5952,g5031,g572,g2556,g2298,g2126,I6094,g10311,g10875,I11767,g9835,g2103,I6110,I14531,g2655,g2731,g8441,g4471,g2843,I5237,g6879,g11309,g868,g9735,g10217,I11956,g2322,g9767,g6499,I9132,I10807,g7816,g5688,I17164,g10668,g2799,g9419,I14858,I7840,g5903,g8155,I17142,I11936,g8846,I16723,g635,I5765,g3164,g11589,g476,g6538,g4717,g7509,g2758,I6894,g11021,g2352,g3696,g4895,g9862,g3246,g10365,I15377,g8435,g10042,g4436,g10431,I6145,g1216,g6106,g2855,I15804,g3875,I13809,g8210,g10950,I17237,g2158,g4263,g6109,I9571,g4988,g1231,I9845,g2013,g5001,I14537,g1101,I17684,g6146,g6488,g8444,I11656,I6302,I11235,g2979,I5737,g1428,g2227,g7651,g9527,g8804,g762,g4671,g10625,g7886,I16145,I5565,g4116,I12038,g7687,I13272,g8844,g4541,I5850,I16720,g8179,g11483,g962,g11357,I13030,I6772,I12502,g11655,g4412,g5918,g6306,g8065,g4125,g7638,g10849,g756,g7467,I14876,I5815,g9365,g8629,I17534,I6513,g2779,g9094,I5716,g8097,I14786,g4564,g11349,g4061,g6321,I15395,g1896,I4985,g5592,g7582,I11587,I14499,g9768,g7614,g3829,I12106,I7244,g9876,g6619,I13418,I7417,g11017,g5781,g8757,g7670,I8671,g8801,I10343,g11404,g10057,g8615,g5533,I14967,g9952,g6363,g5300,g1424,g1050,g6343,g1292,g3732,g5179,I8728,g7471,g4359,I7651,I9224,I6469,g6161,g7496,I5922,I13639,g4089,g7320,g6172,g6844,g3094,I6240,g2733,g7515,I12986,g6183,I16793,I11540,g8948,g2082,g5693,I15497,I7713,g3087,g2005,g6698,I12171,g8273,g10762,I10643,I10120,g3791,g8119,g4638,g5596,g7604,g7132,g6687,I17633,g5822,g9150,I11836,g8849,g5763,g2222,g3704,I9111,I14525,g5035,g10503,I8551,g6951,g2987,g4636,g4288,I6264,g4601,g2347,g7629,g7001,I15554,I5995,I5459,g1648,I7276,I5336,g5935,g4265,g5525,g4972,I6747,I9684,I12403,I6106,g7464,g6793,g1113,I14264,g5099,g2098,I12144,g10163,I17104,g11069,I11662,I10910,g7683,g6584,g11178,I7322,I7321,I8080,g10494,I7612,g11043,g10553,I15956,I5880,I10756,g9508,I15448,g7227,g11279,g6218,g3077,g4418,g5804,g3970,g2275,g8547,I14709,g10436,g9641,I16286,I7763,I6156,g3941,g5625,I6805,I15054,I16817,I13197,g8567,I15725,g9962,g9261,g4321,I5245,g582,g7736,I5451,g7945,I7014,I16258,g11478,g10484,I14388,g8643,g1955,I7453,g3009,g11172,I10924,g8291,g11289,g4736,g3226,I8308,I13529,g2812,g4732,g6798,g7627,I12930,I16032,g3752,g7413,g2431,g3428,g8272,g8609,I7556,g162,I10724,I10963,g2510,I8848,g10087,g11226,g2046,I5576,g9583,I15782,g8412,g7697,g1149,I14989,g3373,g940,g2818,g2338,g6308,g6463,I4941,g10612,I4973,I8647,g5110,g6104,g11282,I7642,I13224,I7432,I14948,g10442,I15453,g3906,g3141,g9601,g2891,g1681,I9007,g8656,I9893,g2944,g6915,I6200,I17503,g5623,g3538,I10541,g3348,g10349,g6536,g826,g11284,g10576,I8418,I13574,g11100,I14097,I9981,g5536,g10214,I5077,g11435,I13812,g8769,I15962,g10405,I13489,I15214,I14701,I16060,g4081,g1549,g3108,g7674,I11211,I8831,I15060,g11610,I15464,g10937,I5662,g2902,g3305,g6406,I12592,g5699,g2889,g6179,g6289,g7441,g4463,g8008,g11594,g3768,g2341,I7729,g7750,I6125,I17444,g6297,g3706,I5406,g5664,g11209,g5823,g2074,I11665,g10367,g4340,g4948,g746,I13621,g8784,g8285,I12081,g3685,g5212,I5095,I12805,I7435,g6546,I5231,g1531,I8237,g3352,I16360,g10820,g1791,I15971,g3437,g10754,g4103,g7098,g5499,I13400,g10101,g10577,g11256,g9389,g1630,g10758,g9953,g10289,g8811,g9776,g6035,g4961,g9966,g6672,g55,g7511,g5529,g8777,I9789,g8128,I12363,g876,g6662,g7765,g7587,g5741,g2084,g4335,g4323,g506,I9984,g6905,g3458,I11387,g7772,g5530,I16664,g1765,I5932,I15974,g557,I9096,g9621,g10546,g8677,I13338,I15880,g416,g3321,g2007,g4347,g6916,g5446,I15635,I9594,g2950,g3982,g7636,I16067,g1861,g305,g3996,g6776,g10231,g10155,g3585,I11790,g11077,g8032,g5684,I15965,g2778,g3770,g3068,g10534,g5503,g7516,g1657,g6805,I12838,g10510,I12942,g7367,g2166,I16808,g3394,I11602,g7824,g3423,g2240,g10226,I17176,I11707,I10816,g6856,g9648,g1618,I13907,g7770,g3540,g10544,I10607,I14083,g8631,I12496,I12559,I17419,g11167,I15694,g8442,g6170,I9901,g10305,I17092,g10696,g7987,g11315,g11513,g4252,I12282,g11651,I11737,g4478,g11029,I12550,g8360,g7725,g4411,I5391,g10352,g10295,g8711,g261,I7852,I13589,I10795,I14805,I15308,g9534,g8125,g7226,g6133,g9894,I8787,g5127,g6895,I8116,I15993,I5858,g8341,g5481,g7990,g7445,g9366,I8650,g4425,g2016,I12067,I12919,I5469,I17400,g5091,g6105,g5518,I15302,I11498,g7389,I12265,g6359,I7749,I9883,I13323,g6052,I16586,I9720,I10920,I15523,g4121,g8960,I8234,I13648,I10996,I13773,g2554,I11599,g3363,g5082,g8651,g1377,I13962,g8693,g9875,I7837,g3978,g2389,g10317,g2906,g4170,I12115,g4677,g4378,g8791,g3519,g2800,I11071,g3417,g5314,I14444,g7766,I14570,I14005,g6967,I14831,I11704,g4619,g3738,g6439,g4882,g4543,I15269,I5221,I11159,g11510,I4780,I6273,g8748,g1857,I10221,I16799,g8709,g9553,g11366,g3775,g3330,g272,g4725,g8234,g6833,g2339,g4770,I4917,I6007,I17466,I13720,g4327,g2115,I12933,g1546,g5648,I10421,g4475,g7260,g8922,I10535,g8974,g6778,g3910,g3536,g11601,g5787,g1499,g6724,I12003,g2759,g3463,I11973,g2088,g2268,g9599,g8715,I8154,g580,g4358,g4944,I10739,I5229,g11420,I12463,I7131,I7210,I15224,g6934,g6054,g2334,g10753,I15898,g3862,g8892,I5128,g7897,g11451,g8710,g8250,g5643,g7800,g6145,g2203,g1125,I16458,I10096,g6617,I8797,g4951,g4417,g7574,I11188,I11947,I16781,g4755,g9763,g11632,g7538,I10334,g4483,I9020,g2873,g7145,I8761,g8516,g10887,g7360,I13952,g3633,g7302,I11278,g6305,g4839,I6370,g4484,g8845,g9904,I15443,g1974,g9853,I13010,g8873,g8015,g9676,g2186,g2850,g4376,g4903,g8311,g5006,I5502,g9882,I6338,I14202,g9883,g9944,I11456,g7054,I11255,g8115,I9759,g5633,g8236,g8123,I11921,g8431,g10556,g1304,g4511,g8193,g1965,g1878,g166,g1371,g9312,g1707,g2106,g8364,I13469,g10808,I9243,g9925,g3335,g10722,g8059,g4285,g4563,I8282,g9843,g9900,I16008,I10132,g8921,g6112,g10433,g10871,g1245,I11680,g8538,g6398,I15592,I9006,I12638,g4748,I7683,g1962,g11255,I6350,I15380,g10351,I9567,I15386,g5318,I8429,I11303,I6316,g9109,I8513,g4976,I10804,g6397,g8245,I11641,g4885,g10325,g530,g5214,g7355,g8168,g6944,g10692,g2776,g10894,g6037,g6939,I9625,I17228,I9776,g11423,I6867,g10862,g5228,g9584,I5284,g5013,g5151,g10313,I13990,g7303,I8642,I10613,g8664,g10013,g10353,I10891,I12493,g2945,g11213,g8818,I9550,I13816,g10288,g11081,g6858,g7240,I17519,g3877,g5478,I15733,I10355,I9205,g7588,I15441,I6880,g2070,I16184,g1133,g8339,I16772,g754,I16787,g5176,I16101,I6118,g7376,g8768,g6075,g4869,I14379,g4730,g5789,I10846,g7580,g4266,g8287,g6036,I6898,I6799,g7815,g4939,g5124,g9729,I8934,I6111,g5778,g39,I15320,g6696,I17739,g11479,g8329,I13230,g293,I5427,I13017,g11602,I8247,g2321,I4929,g4190,I5332,g6163,g5759,I16673,g11012,g8484,g10974,I8624,I6549,g4616,g2120,g8972,g10890,I4997,g3390,g5552,g7350,g10496,g2541,g7904,I6046,I13403,g6320,g10848,I14140,g5201,g2214,I9479,I13708,g5402,I11898,g7347,g9710,g6862,g5546,I17613,g7426,g5000,g5259,g9076,g11311,g8640,g8381,g11486,I7104,g3407,I13351,g7378,g10299,g7755,g5081,g2363,I11112,g11629,I16468,g11149,g6471,g9432,I17410,g9738,I12647,g3008,I13013,g3999,g5512,I6121,g10652,g7186,I10391,g6294,I6748,g421,g11624,g617,g9928,g8942,I12026,I14503,I11698,g4345,g9774,g3682,g8067,g7225,I13522,I14540,I12475,I13099,g5098,I4873,I7363,g6925,g6091,g8770,g6154,g11166,g2862,g7935,g11586,I5734,g5032,g8939,g3416,g7819,g10691,I9851,I12415,I16080,g6330,g10752,I5203,g1753,I17657,g8172,g4592,g6787,g6816,g1458,I8061,g3012,g2988,g7205,g2644,g9931,I14010,g6622,g6758,I16038,g2555,I10030,I12409,I12849,g5304,g2034,I8180,g6688,g6686,g6523,g4824,g6121,g8159,g8706,g2775,g8933,g10512,I17052,g6948,g8523,I9915,g4497,g8423,I13394,g2410,g4963,g10339,g8480,g8498,g6318,g4606,I16580,g7740,I5588,I14973,g9760,I13615,g588,I16607,g10148,g4738,g3799,g5012,g1654,g8771,I6022,I6832,g8445,g10720,I9854,g2077,I6565,I11686,g11571,I11942,g11275,g2124,g3304,g10931,g7938,g4069,g8385,g7821,g8799,g10599,g7422,I5611,I5295,g810,I14558,g10853,I7864,I10111,g10167,g7106,g4105,I12574,I17296,g2305,g2744,g6853,I16081,I11312,I15290,I12248,g10125,g10770,g11242,g6873,g6775,I12875,I10771,I17158,g3517,I16626,I7559,g9672,I6686,g8303,I13729,g2235,I11974,g11539,I8577,g5934,g9350,I5164,I11982,I14543,g7996,I10461,g2479,g4275,I5926,g4217,g9829,g6692,g11397,g1047,I16920,g10795,g8023,g11557,g7818,g7662,I13451,g5205,g10370,I6068,I5518,I11889,g11415,I6102,g5752,g4380,g2296,g8632,g8104,I15855,g6794,I9938,g10441,I7782,g581,g10322,I12180,g9610,g11402,I15718,g3274,g4394,g3345,g4567,I12604,I5943,g8778,I8298,g8476,I12613,g6291,g3093,g6521,g11239,g5851,g8049,g5074,g10581,g2349,g2424,g5277,g6399,g10247,g585,I13077,I9377,g11220,g9741,g10860,g6127,g6801,g6812,I7402,I14903,g10663,g6563,I9658,I11228,g2345,g10593,g8124,g10471,g11144,I6726,I15177,g8401,I8752,I5240,g6900,g7705,g10804,g6860,g8790,g8133,g4883,g8160,I10557,g3763,I11423,I5957,g1669,g11556,g10541,g2863,g5875,I15530,I8641,g5539,I15999,I10168,g6580,g11625,g4912,I14675,I7564,g3912,I5315,g8006,g11148,I11907,g9388,I8133,I16717,I11222,g549,I7342,g3533,I5501,g2499,g7586,g11440,g8191,g2456,g11237,I5592,I15299,I17290,g10025,g11085,g6861,g10440,g8293,g2043,g5040,I11932,g10766,g11437,g7589,g3749,I10885,g10276,I5186,I6186,g9598,I15314,g2794,I5652,g2774,I13051,I12232,g10384,g7761,g10822,g7899,g579,g9965,I6856,g5983,g10302,g6760,g4811,I16273,g34,g11495,g5472,g10265,g6443,g2754,I14109,g5320,I9162,I16052,I13765,g5216,I10620,g9690,g8337,g3813,g9647,g1453,g6085,g3247,g6928,g5720,g6560,I7577,I11671,g11158,g3431,I17459,g9313,g4921,I9558,g2943,I5486,I6137,I7166,I11915,g299,I11611,g2224,g7591,I5357,g7693,g4761,g8284,g3539,g11319,g10646,g4094,g2819,g11429,I6560,g2752,I15088,I7462,g4823,I8406,g7394,g8992,g9125,g7971,I10508,g6819,g11607,g7759,g4453,g11225,g4296,I14232,g7637,I8520,g2939,I13302,g7550,g3736,g4232,g5392,g5113,g5396,g5073,I6322,g11413,g7623,g2310,I15085,g6322,g4875,I12562,g11019,g7902,g4186,I7291,g643,g4262,I7185,g6249,I13258,I9016,g5620,g5117,g9423,I15899,g466,g2837,g2757,g10527,I6690,g5023,g5112,I8085,I11166,g11441,g9316,g9240,I12508,g2593,g591,I5085,g6809,g6197,g11146,g2215,g8879,g7064,I9114,I6580,I7411,I9171,I10456,g5391,g11073,I14210,g7872,g7917,g7,g10680,I10274,g6528,g9664,g4454,I9443,I14265,g6164,g10357,g10666,g6251,g8042,g6003,g8767,I12261,g5726,g6745,g7688,g10727,I6881,I6381,g10699,g3506,g11326,g4053,g10498,g8785,g10751,g3261,g11427,g11496,I14279,I6507,g3819,g7235,I11575,g5769,g566,g6956,g4640,g7336,g2212,I8858,I6019,I6323,g4513,I13959,I8820,g4162,I11728,I6091,I15778,g486,g7039,g6040,g8334,g5029,g6789,g10330,g3903,g6813,g10092,g8472,g2162,g713,g1555,g8775,g4554,g6891,I5276,g5649,g700,g6050,g5279,g10116,I8031,I15190,I10117,g11022,g5114,g9645,g3010,g2949,g4913,g5264,I6911,g9914,I9117,g10892,I12165,I16039,g755,g2405,I11143,g5192,g11612,g7116,g7387,g2221,I10560,I7154,I9734,g4674,g2391,g5072,I10946,g4314,g6594,I5371,g4273,g8225,g7301,g10596,I11467,I10706,g1983,I6409,I9647,g10140,g9707,I6715,g8440,I9287,g10485,I11447,g11038,g8559,g8535,g9205,I8256,I16467,g10363,g10122,g6635,I5618,g9204,g5883,I13723,g7921,g2110,g10408,I13645,I10234,g7416,g11590,g6078,g4450,g9694,g2432,I9229,g8638,g4583,g11277,g7385,g6871,g7323,g369,g7601,g9820,g2539,I16613,g10555,I5351,g7956,I9259,g7599,g8971,g2719,g5701,g6927,g8346,g3792,g2351,g4253,I6836,I11692,g2537,g5285,I4783,g8428,I6077,I5710,g8414,g7139,g5845,I15293,g6447,g3663,g9884,g3979,g2880,g11059,g5698,g10439,g7763,I7157,I5171,g11079,g9082,g11317,g11156,g5171,g10882,g5725,g7929,I17687,g11159,I7800,I14449,I14906,g4533,g6575,g4225,g7288,I6944,g7626,g8436,g7936,g7721,I15749,g10396,g802,g6046,I15247,g2548,g11454,I8669,g3138,g8595,I11584,g6293,g6571,g4722,I11997,g10783,g4444,g8069,I11797,g3530,g5507,g2270,g8969,g1713,I8815,g8134,g2194,g5768,g5187,g2654,g2791,g5857,I7648,g5150,I9409,I17662,g9742,g5036,g6062,g11066,I9531,g8131,I12015,g9490,g2550,I13544,I11065,I13788,I16024,I6487,g6238,g6872,g11344,I5517,g2743,I12999,I11330,g11617,I7345,g10382,g7852,g9341,g5668,I9839,I16058,I14534,g2343,g11348,g9339,I7423,g8579,g11384,g10868,g287,I11566,g5007,I6138,g6482,g11560,I16805,g11395,g5736,g10690,I15039,I8985,g2096,g11550,I9863,g8622,I6929,I5120,I10828,g7293,g9586,g7796,g8551,g3751,I7935,g2411,g9704,I14979,g8176,g722,I11242,I5539,g5696,g1810,I12799,g10263,I7719,g10738,g1092,g7345,I12307,g11434,I13837,g11091,g6326,I14209,g10233,g3743,g8592,g10031,I14312,g10529,I6085,g4581,I17460,g11296,g1598,g4503,g1083,I5605,g3381,I17149,g4219,g4317,g7762,g1080,I7360,g11152,g11095,I16280,g8947,g4896,g7315,g8958,I16111,g32,g2100,I5127,g11345,g5222,I12809,g10119,g3200,I6133,g3102,g8837,g11450,I12239,g6060,g9525,I17334,g11216,g11393,g2451,g6731,g5674,I13735,g6884,g11407,I15665,g1153,g10331,g8479,g5041,g8944,g4165,I7182,g5862,I10198,I13766,I11534,g7420,g4772,I17568,g1736,I16072,g5740,g6191,I12245,I12825,I13236,g10043,g11310,g2223,I12857,g5094,g3271,I11674,g10739,g8721,g5547,g3387,g3343,I14179,g11210,I11348,g5689,g10523,I8228,g6432,I17307,g6155,g6086,I9699,g2832,g6755,g7571,g7729,g6834,g950,g3473,I17265,g5252,g10670,I10589,g10777,g3089,g11480,g278,g10253,g875,g6885,I13023,g7213,I10437,g2677,g7410,I9591,g5889,I14112,g9533,I6177,g8403,g3939,I16175,I6802,g6674,g4361,g6452,I6702,g10195,g9515,I12216,I11459,g5708,g5874,g7602,g7879,I10159,g6984,g4535,g11611,g6542,g2097,g8570,g8946,g6081,g11548,g2629,I15172,I17567,I8663,g2008,g10443,g10481,g8705,I4891,g4079,I5713,g1932,g6628,g5220,g6227,I8973,g8437,g2211,g10294,I11914,I12520,I15792,g554,I12012,I9329,I6163,I7760,I7330,I8729,g4338,g4369,g8526,g11421,g258,g2380,g10881,I9123,g4733,g5348,g936,I15305,I12286,g1324,I12627,I16492,g6199,g3110,g10548,g7263,g3988,g9897,g7210,g255,g2248,I13888,g1321,g4716,I6671,g11334,g5232,I17337,I15526,I6598,I8869,I5292,g10973,g8749,I7369,I9265,g9886,g7953,g10292,g6764,g2000,g11274,I12168,g9779,I7216,I5005,I15879,I16059,g11584,g9085,I17377,g7597,I13965,I12357,g8333,g5676,I11528,g5818,I6126,g10827,g4787,g10192,g7390,g10479,g7595,g3529,g5193,g9554,g9644,g8943,g569,I7766,g5980,g58,g11325,I6477,g5737,g7883,I16217,g8187,g2368,g4747,I5020,I9798,g11442,I11722,g1724,g10788,g2317,I9612,I6013,I11759,I12412,I9544,I5986,g491,g11058,I13086,I6260,g8309,I11127,g10264,g4835,g11276,g8555,g4566,g1504,g10735,g11390,g11243,I14522,g7606,g10402,I12490,g7122,g3705,g11388,I11841,I7002,g11369,I4935,g5469,I14822,g6627,g2892,I5031,g2154,g11331,g5482,g7546,I5992,I13586,g11604,g11101,g2253,g2028,g10358,I15759,I6043,g4521,g8760,g9420,I5516,g4904,g6311,g8350,g6552,g10371,g8611,g3205,g4122,g9124,g10669,g10033,g7884,g7663,g11262,g4332,I11824,g8938,g9804,g5287,g10578,g2061,g6444,I10984,I15238,I17482,g7289,g5700,I5053,g7685,I12159,g11399,I16610,g5891,g11543,g11572,I14405,g8930,g4291,g8823,g10250,g1615,g4239,g8949,g11070,I15829,g296,g9785,g3318,g3056,g9777,g1270,I6924,I17368,g3120,g4986,I12085,I7662,g4502,I7843,g5416,g6205,g4919,I5283,I8803,g237,g8163,g10007,I6454,g7221,g10277,g10171,g8617,g11425,g6941,g2449,g2225,g4142,g4545,g7622,g9588,g8448,g269,I9585,g6539,g7011,g4000,g10855,I7450,I13482,g9919,I8011,I12274,g3879,I14397,g7704,g4398,g8029,g658,I12813,I16376,g3326,g10661,g9703,I5073,g11473,g411,g266,g4879,g3460,g6562,I7677,I15983,I14982,g9893,g6840,I11082,I6484,g11418,g7782,g1882,I10937,g5639,g2232,g9331,g5619,g11639,g3413,g6839,g605,g49,g4084,I10753,g10483,g1766,I9099,g7009,g3434,g8383,g4379,I7680,g10284,I13329,g7658,I11926,g7311,g73,I15675,g3055,g6032,I11510,g6681,g7286,g3268,g8486,I11901,I13048,I11106,I6777,g5275,I9188,g3070,g2522,g8779,g4306,g3635,g6581,g6744,g11582,I13445,g8558,I11989,I9240,I7284,g10501,g2689,I9446,g7549,I16178,g11040,g7603,g8380,g2726,I13083,I6385,g5811,g9353,I17365,g7764,g1015,g583,g7342,I12047,I12436,g9964,g11023,g10139,g9951,g321,g5904,g6435,g2344,g8354,g11112,g8330,g4163,g2091,g7912,g3992,I7671,g3396,I6124,g7758,g2771,I10384,g5624,g6699,g2450,g9579,I5311,g7446,g10867,g4315,g4968,I5184,I5510,I11593,g7890,g10478,I10770,I5204,g7979,g4159,g6717,g11603,g11061,I15199,I11653,g8197,g7442,g2919,g7292,I10573,I12916,g8416,I8479,I14866,g5894,g4734,g5107,I8670,I17669,g9757,I14303,g10158,g8774,g9864,g2125,g2337,I5629,g275,g3392,g2167,I6498,I14130,g8989,g10088,g4577,g11616,g10001,I17374,g5887,g40,g7200,I17416,g2911,g2436,g944,I4980,I9108,I14355,I11623,g8297,g5790,g11592,g10423,I10090,g4994,I13828,g8043,I13893,g8305,I10427,g6763,g2202,g6137,g6446,I13360,g5123,I7685,I5378,g6237,g6178,g6203,g7928,g10492,g9845,I9090,g2273,I15968,g2218,g5617,I15565,g3773,g7738,g4343,g7316,g9519,I11995,g9569,g11036,g6186,g11502,g3563,g11308,I6461,I12953,I9062,I11713,g1265,I12069,g8377,I10362,I7323,I12529,g11109,g4998,g2406,I9744,g6667,g7620,I15241,g11577,I15890,g4496,I7225,g4735,g2234,g3943,g5943,g7984,g7805,g4185,g2507,g11376,I15210,g5706,g7539,g9887,g7068,g1738,g9837,I7099,I6838,g10470,g11652,g5613,I16956,g4763,g3733,g6970,I17505,g6472,g10500,g7611,g7110,g10242,g5199,g10172,g7361,g3624,I10663,I9279,g9563,g6126,I16850,I6648,g8660,I15986,g7998,I15215,g10315,g7797,I8677,g10283,g7711,I7272,g3290,g2540,I5824,I9433,g6532,I5265,I8715,I6553,g8806,g3344,g7305,I7691,g6881,g2884,g11394,g11508,g5166,g6115,I6144,g11622,I17461,I6225,I17100,I8711,I11716,I16108,g1595,g3213,g6241,g5661,g11292,g6728,g9932,g8252,g9448,g6300,g8782,g108,I11363,I8465,I4951,g4892,g664,I7996,g2245,I10519,g9340,I7546,g8789,I14443,g5542,g10946,g2255,g9782,g6051,I9282,g9355,g4366,g11060,g4752,I14751,g11541,g8888,I13857,g10056,g2233,g6746,g1368,g11403,I12318,g2015,I5913,g11574,g9856,g7722,g10296,g1280,g9942,g7219,g9349,g7330,g6917,g4189,g6742,g6210,g5096,I10394,g8568,g10826,g3981,g1811,I17305,g1900,g2021,g7631,I15485,g10491,g9866,g8764,g7808,g1990,g2840,I8337,g7270,I4955,g3362,I13840,I15171,g11010,g4678,g3433,I9857,g1019,g11205,I13695,g10559,g9526,g471,I16025,g3769,g1360,g10865,g11244,g7931,g11491,g2252,g5686,g9360,I5218,I11501,I5070,I5248,g11143,g4498,g6618,g4226,I6347,I15311,I9221,g6136,I16938,g4395,I4987,I17692,g7182,g7594,I15716,g5669,g8731,I5540,g6002,g3709,g9507,g4753,g7363,g11519,g11498,I6287,I6770,g8630,I8024,g8260,g8324,g10348,I5866,I8851,g9619,I17321,I17522,I12406,g10582,g11080,g8338,g10380,g8819,g8312,g4129,I7408,I6587,g11504,I5655,I9995,g9600,I9402,g5500,g6048,g5444,g6382,g2883,I9102,g8376,g6838,g2985,g3353,g8321,I13661,g8332,g10362,I5754,g7088,g7732,I12114,g7349,g10524,g2502,g10949,I15992,I12039,g9418,g7790,g2796,g3744,g7187,g5654,I9144,g10434,g1945,I10630,g2809,g7739,g3520,g7307,I14239,g7010,g3817,g4604,I10849,g7510,g7669,g10138,g6469,g11026,I13433,g1141,g6943,g5197,g9736,g9993,g11093,g5510,I16784,g7843,I5690,g7246,g2669,I8563,g8478,g2038,I5264,g4754,g2938,g7547,g201,g6551,g481,I10162,g6889,g8375,g2331,g9354,g1011,g11316,I7833,g4126,I12690,g11623,g11452,g7192,I7315,I6217,g11398,g5024,g2829,g8405,I6097,g5274,I6109,g6537,g10191,g8233,g2056,g6353,I8854,I6065,g3186,I10251,I16811,I17413,I16187,g8,g2172,I12193,g7359,g6799,I13194,g7034,I8164,I14272,I6196,g4297,g4953,I5358,g4355,g7351,I9822,I6504,g4438,I12397,g1756,g4501,g6718,g2701,g5010,g8247,g10564,g8469,I10710,g7406,g6697,g5881,g10047,g9773,g8796,g6893,g10314,g3812,I9608,g1218,g4233,g10969,g10764,I9948,g1980,g5602,I11629,g7596,g9582,g1314,I8535,g2478,g1828,g123,g9833,g8936,g2072,g11608,g7958,I8805,I7447,g5657,I9872,g695,I6812,g2220,I10927,I15536,I17240,g8482,g4370,I17362,g8816,g5727,I9440,g11591,I12215,g8325,g6804,I14087,g5912,I17493,g11443,g7920,g4298,I17610,g5403,I10499,g10506,I6661,I5263,g7756,I17283,g5272,I12457,g11177,g4713,g4728,I7035,g7295,I10322,g4222,I5719,g6150,g1490,I7710,I12862,g3718,g11353,g3062,g630,g8378,g5251,g7334,I16311,I10952,g2080,g2184,I14888,g6509,g3582,g7374,g8934,I9068,g3143,g6792,g8507,I15193,g6810,I14101,g1567,g1383,g4344,g6348,I11800,g5030,g8694,g10411,g8653,g3998,g8053,g9260,g7657,I11241,g7502,I10308,g3790,I5006,I11119,I17616,I5210,I5731,g7053,I12913,I6309,g10400,g7889,I11061,g11011,g5039,g4880,g2877,I13209,g10297,g7031,g6478,I6917,g2861,I16592,I17302,g965,g8987,g798,g5672,g3946,I14672,g2251,g6120,g1086,g563,g7784,I7426,g4188,g2238,g7465,I17513,I17356,I15365,I8651,g9891,g9872,g9391,I7536,g7379,g11312,I12099,I11970,g1217,g8140,I8379,I6310,I7096,I6199,g7978,I14687,I7086,g5491,I6557,g11400,g8147,g4455,g654,g7326,g2662,I16814,I9816,I6247,I15826,g11197,g10742,g861,I12433,I16629,g2867,g10424,g11099,I12442,g3439,g7794,g7329,I5098,g1317,g1963,g6506,g11170,g9506,g11232,g2534,g6938,g7812,g10156,I11338,I8211,I13561,g6847,I15586,g10932,I10108,g7366,g8891,I14933,g1474,g8719,I11810,g11511,g9668,g1762,g4003,I5034,g5895,g7026,g8625,g7581,g10177,g10554,g7947,g1494,g7512,g2264,g8103,g6797,I9156,g3287,g1964,g6910,I13747,g8294,I7163,I12020,g4375,I14315,g8670,I10813,g8726,g9696,g4840,g9024,g9705,g1065,I4965,g1260,g131,g3425,g5638,I14976,I13105,g10635,g10775,g8167,I9296,I12384,g9273,g3662,g8955,I16763,g3066,I5946,g3076,I11342,I7223,I4956,g2860,g11028,g10717,g5122,g2506,I8303,g2079,g6824,g5742,g9110,I9380,g6094,g4482,I17194,I6468,I8892,g2807,I5484,I11794,I14045,I10509,g8713,g6508,g7684,I16209,g7070,g8654,g207,g8645,g2496,I15033,g3365,g6666,I10293,g5309,g4278,g6870,g8361,g6001,g2797,g11086,g5034,g11490,g6565,g7959,g4112,g1300,g1577,I14319,g5880,g6655,g1988,g4507,g9860,g3522,g3252,g1801,I13212,g5480,g8877,g6906,g6815,g11656,g9421,g8314,g2399,g2524,g11300,I9801,g61,g9352,I12138,g8780,g7803,g4064,g11212,g9658,g2509,g3537,g366,g6550,g8887,g8487,I11519,g10093,g9151,g6043,g8624,g8920,g2858,g4487,I10299,g7556,g4056,g1633,I6879,g782,I5887,I15412,g10271,g4756,I16769,g5721,I12867,g5522,I10503,g2531,g8511,g7033,g1110,g7008,g2959,g6116,g8803,g11561,I7973,g5250,g6134,I15219,g7673,g6310,g8815,g2635,g6396,g11098,g5470,I5613,I17288,I11354,I14862,I13568,g5557,g5225,g10884,g8500,g8388,g6108,g4168,g3783,I12580,g8950,I6630,I13285,g4789,g11155,g8040,I8967,g8890,g2434,I12511,g11597,g8421,I13901,g5083,g10429,I9349,g9934,g4231,g6843,g7994,I5445,g9642,I6990,g6344,g7682,g10904,I12035,I7264,g976,g1407,I8575,I4820,g6596,I9749,I14612,g11153,g7059,g5273,I15891,g4255,g7608,g7710,I13732,g115,g5043,g8462,I13415,I11975,g4452,g9662,I16775,g4837,I11472,g8169,g10203,I9421,g10204,I9105,I13819,g11071,g10430,g6786,I13514,g6535,g11620,g4480,g38,g8206,g8011,I13915,g318,g5180,g7136,g7893,I4996,g1972,g8044,I15347,g7919,g2340,g6707,I16088,I7295,I5818,g3427,I13089,g10178,g4372,g6225,I13370,g6877,I10979,I12369,g9719,g9896,g8056,I11937,I13546,I6282,g9028,I15424,g2018,g4783,I10855,g9832,I13711,I9655,g8928,g5231,g11200,g11096,g7038,I11563,g9591,g3976,g8953,I15356,g8075,g4354,g8446,I17179,g2808,I14827,g6445,g11469,g6465,g4256,g10574,g6620,g2824,g8728,I17170,g7437,g2299,g11268,g5593,I6789,g7143,I8385,I8626,g1524,g10514,g5569,I11176,g9758,I14216,g6169,g10227,I7381,g2174,I13908,g6875,I5530,g6479,g6235,g10495,I10837,g4011,I10762,I5879,g3426,g7380,g345,I13887,I5025,g6039,I17255,g4280,I15632,I13577,g11618,I15068,I4961,g9819,g2107,I5316,g11347,I9268,g5062,I8139,I11391,g2207,I8293,g9905,g11576,I11734,I7022,g8429,I6025,g4393,I4964,g5691,I10021,g6298,g10333,g5494,g11240,g8965,g8606,g11307,g6823,g7072,g4682,I11882,g9740,g6125,I16196,I16656,g6971,I10825,I13506,I11046,g2789,I17424,g3714,I13876,g10522,g2852,g11065,g11185,g7906,I5998,g5217,g4166,g8095,g5660,I9706,g4681,g8994,I16220,g7524,g8745,g10157,g1346,g8512,g8881,I14964,g9454,g9585,I8262,g2254,I14914,g7913,g8542,I8036,g8157,g10019,g3040,g5471,g8108,g2990,g11447,g10852,g8941,g6933,g7204,g9770,g4530,g1077,g9945,g5695,g10706,I6417,g11222,I5067,g10110,I17359,g9727,g6339,g6386,I10526,g5707,g3475,I12196,g4729,g3566,g2379,I9536,g6720,I17198,g2728,g11409,g2094,g10508,g4008,I5142,g6341,g5756,g6836,g1023,g3370,g686,I6590,I15157,I16543,g7924,g5601,g9660,g10773,I7048,I10305,g6585,g5757,g5263,g7885,g10947,g5808,g8659,g10538,g5066,g4329,g4586,g9717,g4802,I17277,g10886,g10131,I9737,g11336,I13039,g8868,g8572,I6294,I9452,g5685,I10180,I8250,g3715,g6454,g7073,g2078,g7291,g9709,I6955,g7463,I9886,I10009,g7029,g315,g3722,g4881,I5892,g10863,g5595,I13580,g6433,I10623,g7727,I17318,g7542,g7735,I12366,I11992,g11337,g7045,g3060,g11188,g5718,I5192,g11352,g4224,g2913,g2069,I9290,g5735,g10623,I8989,g8081,g8020,g351,g11293,g10825,g9346,I16500,g1041,g5809,g7792,g5866,g4479,g10913,g7277,g2517,g5796,I6538,I13227,g8099,g786,g158,g8838,g7771,I14582,g7776,g4293,I11581,g3521,g9367,I10057,g5941,I9539,I15418,g9698,g8602,I14136,g4615,g6351,g1850,I14090,g6475,g2117,g4104,g2750,g1909,g1104,I13188,g11196,g186,g5723,g5877,g5594,I14415,g8343,g4838,I10685,I5450,g9680,I8089,g7089,g9328,g10427,g7961,I9248,I8763,g3720,I10514,g7321,g4264,I10237,g7224,g4461,g8876,I8351,g4342,g2971,I13992,I14958,g11505,g2764,g9922,g9711,I8771,g11545,I12143,g1137,g10075,g2947,I12293,g8798,g10480,g11018,I10027,g2004,g11501,I17209,I13767,g8357,g8213,I14326,g2086,g4388,g7521,g3047,g9840,I10769,g10662,I13895,g5286,g3222,g5477,I6528,I8481,g3735,I13250,g7056,g5209,I7366,g10114,g3531,g3262,I9165,g6578,g5254,I9632,g3331,I13630,I12075,g5998,g11428,I6088,g3418,I12448,g7214,g10137,g3112,g7847,g11266,g5655,I6187,I16373,g11037,g4557,g7724,g4639,g8506,g7272,g2765,g10608,I5571,I7716,I7793,I5620,I11543,I17525,g8952,g7384,I16236,g11063,g7236,I6324,I10689,g8964,g3372,I9677,I4786,g10493,g2346,g6389,g11636,g5524,I15338,g6176,I11076,I14776,g9839,g4274,g1703,I6166,g5233,I6546,g2820,g357,I7726,I16514,g10198,g7338,I15244,g7138,I17742,I15568,g4898,g7949,I15729,I17752,I14249,I14203,g7332,g8117,g5656,I12846,g10388,g2839,g9863,g1730,g6807,g67,g4140,g2942,g5090,g7313,g5843,I11306,I15811,I12214,g2085,g5748,g7613,g10201,g5541,g4591,g3697,g8937,g10083,g11433,I6360,g6360,g11405,g2395,I13949,g5219,I5789,g7333,I12183,g6712,g5513,I9617,g11068,g7435,g10745,g9415,I9829,I6968,I8192,g11035,g6185,g7954,g10343,I6049,g6960,g2542,g2435,I14567,g11218,g5913,g7357,g9948,g8080,g9673,I6424,I7017,g9824,g10421,g3727,I11043,g5230,g11102,g5033,g8991,g11168,g11621,g3914,I11677,g7672,I9792,g7813,I9087,I15256,g8805,g4670,g8744,g1341,g6831,g8968,g309,g5354,g4614,I11961,g3109,I17312,g7731,I7029,g6638,g8407,g8800,g7449,g10900,g6303,g5269,I5840,I15368,g2846,g9531,g9596,I9013,g10456,g10174,I5341,g2195,g7557,g7306,I7886,g3459,g7650,I14494,I14607,g11644,I16843,g7268,g6534,g6679,I6080,g8275,I14367,I9040,I15281,g10885,I14555,g3228,g6732,g2501,I11620,g10549,I13933,I8839,g1062,g5640,g2445,g4542,I4954,g4250,g5901,I10531,I15520,g7876,I9150,I15430,g3440,g7810,g6464,I9605,I11614,I13877,g8283,g2940,I14133,g11173,I11710,g8509,I11483,g4584,g2369,I13239,I17555,g8501,g8254,I8716,I5023,g10239,I10228,g2180,I15595,I11318,I11068,I13295,g1997,g8359,g5100,g4991,g3273,g10562,I9138,g4368,g259,g6555,g8612,g4536,g5003,g6929,g7903,I11869,g7044,I11280,g5646,I14349,I7684,I15864,I15181,g4128,I10733,g7789,g2557,g5572,g9927,g8041,g7206,g5174,I17719,g10372,g11481,I9120,g5680,I8098,g7023,I17274,I13430,g6553,I9135,I10598,I14485,g3301,g8281,g4777,I6010,g2003,g5852,g9555,I8204,g6909,g4605,I13513,I17707,g5739,I6443,g36,g3284,g9590,g7768,I10156,g3221,I16387,I14799,g10531,g4610,g668,g8610,I6343,g11295,I12153,I13463,g4420,g3368,g9714,g7773,I5279,I16604,g7579,g9410,g9946,g2646,g4587,I14352,g5095,I9216,g153,I10801,g6588,g6902,g2569,I10716,g2804,I6351,g4995,I5689,I11719,g11554,I9652,g10781,g2885,g9107,g178,g10761,g3584,I17084,g4868,g6629,g10910,g552,g6586,I14421,g1117,I12223,g8054,g8317,I8625,I11085,I11935,I6576,g5195,g9589,g8327,g8430,I9194,g4996,g3983,I14330,g2025,g10383,I14439,g11161,I4850,g6288,g8304,g9528,g10743,g7878,I8664,I9202,I15870,I16766,g3106,g4063,g11340,g8129,g8151,g11487,g5867,I12002,I16044,I10864,g6736,I17381,g9846,g8122,I9860,g8505,I7586,g10926,g8098,g3940,g4467,g5629,I5418,I6474,g8932,g4127,g1163,g10104,g10080,I7562,I11644,I11333,g10389,g7339,g6730,g2089,g4117,g9359,g7541,g10902,I12595,g324,g6911,I6914,g9693,g9764,g10869,g6090,g4576,I6976,g11540,g5590,g5106,g10857,I10282,g3388,g5681,g6561,g1284,g4561,g10600,I12258,g9345,I13956,g9425,I5649,g6059,g7331,I13797,g10634,g10426,g4935,I10138,g3723,I6742,g5526,g8635,I13294,g6657,I11778,g6068,I5258,I15421,I17537,g5425,I6395,g9335,g1989,I6714,g829,I10549,g6845,g1166,g8192,g8246,g8601,g2578,I16017,I8662,I6965,I17070,g3977,g5825,I12571,g4333,g6957,I6694,g2303,g9223,g6049,g7294,g4975,I11508,g8402,I12372,g5404,g11075,I6001,g9850,g5498,I14596,g254,g4781,g11087,g10258,g9916,g7325,g10248,I6666,I12678,g4259,g10557,g4382,g5128,I17678,I7054,I16009,g5519,I5080,g2372,g5846,g2482,I6958,g2963,I17173,g4949,g3107,I16778,g9718,g6649,g10249,g6345,g10649,g5755,g6058,g3876,g7748,g11030,I10412,g5144,g837,g4942,g6656,g8626,g4158,g11314,g10759,I10286,g10643,I6825,I11262,g9100,g4866,g8004,g8647,g7050,I13248,g10707,I9159,g6829,g7743,I5271,I11683,g6365,g3419,g9871,g7648,g4087,I16121,g10260,I16537,g2068,I6535,g6440,g6913,g281,g5191,g4257,g9270,I12796,g10583,g7062,I12445,I5460,g7888,I7606,g9937,g6358,g8351,I11008,g6425,I16066,g5837,g2560,g382,g4234,g6385,g5772,g4481,I11786,g6314,g1394,g10035,g9938,g6693,g7523,g6907,g7075,g10750,g2960,I6403,g8175,g9899,I5342,g11104,I12128,g10856,g7297,g3729,g6719,g4821,g7898,g8156,g5678,g2374,I14382,g5839,g8725,I13290,g8655,g7137,g11653,g11027,g5743,g4049,g11599,g6411,g406,g7500,I5982,I6907,g2493,g8439,g3485,I15235,I15908,g7787,g5415,I12068,g7103,g4731,I9498,I9180,g8517,g11303,g2276,I13076,g4286,g10948,g4620,g7774,g3524,I12093,g7689,I5230,g3716,I8770,I10069,I15539,g7692,g5679,g7443,I16660,g8546,I9514,I6167,I7938,g2433,g2851,g10734,g11269,g7966,g4439,g6507,g5694,g5258,I17231,g5611,g1074,g9815,g8474,I17340,I5675,I16601,I11345,g4311,I7889,g9877,g6525,g790,I10045,g11509,g3479,g9411,g6089,g6729,g3332,g6317,g599,g3878,g9666,I7143,g7230,I16239,g5008,I12339,g2373,g10193,g10182,I11225,I10147,I15503,g6071,I7803,I16427,g1540,g8929,g2130,I12939,g7257,g2121,g8241,g2101,g8085,g6407,g5915,g3942,I10789,g3621,g10539,g7284,I12786,g11039,I5843,I13391,g2116,g1914,g10223,g9594,g9618,g9722,g6582,g5002,g10771,g11547,I6061,g5651,g3206,g5445,g9954,g6516,I16540,g6852,g5200,g7988,g8410,g7960,g6903,I14309,I17773,g7559,I12583,g10301,g10809,g1520,g3766,I11904,I10974,g8116,g9737,g4057,g79,g10864,g2335,g9822,I5722,g10355,g6346,g2111,I9848,g5942,I13554,I7006,g10386,I11326,I9695,g2614,g7028,I9126,g10285,g2745,I12532,g5858,g4426,g7022,g6461,I6716,g8118,I12094,g6141,I5676,I13078,I14176,g5268,g7696,g9505,g7211,g8344,I10370,g8127,g8463,g5724,I6543,I9293,g4784,g4794,I12053,I5494,I6028,I10917,g8183,I5935,I17636,g4773,g1356,g4914,g2354,g3630,g8235,g2642,g2201,g2503,I15892,I15989,g10716,g7318,g10282,g2217,g10469,g5812,I15250,I7357,g10502,g5705,g10888,g1157,g10638,g6501,g3814,g9412,I17450,g4834,I9065,g8519,I5973,g8141,g3088,g4235,I8796,g2198,g5502,g4007,g6846,I6467,I12060,g4109,g5738,g3405,g6252,g2980,I15807,I11746,g8286,I5475,g9616,g8783,g1675,g9941,g10897,I11560,g9342,g3406,I10907,g6590,g10453,I16867,g516,I15045,g5859,g8178,g11350,g4593,g5109,g9091,g5172,g9665,I13800,g3818,g8925,I16796,I11394,g8470,g2315,g4500,I15323,I15442,g10782,g3398,g6735,g11267,g5993,g5115,g4959,I17402,g8967,g10422,I7354,I9308,g10344,g10741,I10819,g6417,g8975,g2937,I9875,I15329,g1071,I8179,I7757,g8874,I6941,g10877,g9422,I12326,g6352,g10725,I16053,g2161,g7635,I13166,g4617,g6502,g6863,g8411,I15768,g10437,I8147,I15482,I13109,g5266,I14188,I14116,I14793,I10084,g10446,g2962,g2060,I14361,g6207,I8762,g1,I9833,g3807,I4972,g126,g5770,g9450,I6136,g7801,I12255,g8730,g9881,g3044,g3379,g2951,g4067,I16016,g2446,g5227,g1528,g7679,g4083,I6996,g5647,g8326,g9348,g9834,g5652,g257,I5089,I8253,I7311,g7806,g7908,I14779,I10189,g8840,g6806,g6000,I11293,g4294,g11052,g7605,g9392,g3052,g4473,g7948,g11254,g10543,g11305,g5899,g7526,I14094,g8259,g2185,I17710,g6368,I16574,g986,I5106,g8220,I9826,g5202,g1786,I5441,g7708,g8101,g7590,g8406,I16469,I11397,g4718,g1336,g4791,g10854,I13466,g4504,g4973,g7630,g3772,g2643,g8177,g4675,g8432,g3909,g8203,g10304,g6144,g3861,I17384,g2396,I13043,I8885,g9309,g7822,g7569,g5605,g7723,g5063,g6526,I17724,I11814,g4558,g11056,g9272,I8591,g6187,g11343,g5281,g9781,g10872,g11448,g9870,I16479,g584,I13382,g9778,I4920,I17108,I15517,g4397,I15639,g10898,g2170,g9702,g8541,g8365,I13300,g10934,g6710,g4419,I14713,g6567,I9458,g1351,g17,I5084,g8150,g9838,g7967,g11648,g10590,g1583,g4523,I12770,g4389,g2356,I16531,g2108,g6041,I7916,g448,I10331,g3011,g9851,I4928,I12303,g9529,g6171,g6194,g8598,I15036,g3532,g6107,I5485,g9918,g6302,g7508,g1478,g7686,I7674,g9290,g6184,g7851,g9691,g7932,g5418,I13659,I15350,I9588,g3393,g7244,g9830,I7033,g11171,g6556,g3974,g5820,g7421,g5849,I7420,I12765,g2159,I11383,I6616,I11100,g6557,g8109,g6404,g9766,g10726,g8132,g10039,g231,g3144,g426,g5732,I14340,g7624,g8739,g6131,g10451,I11524,g5308,I11509,g2381,I15601,g4820,g4897,g10570,g1003,g882,I17584,g11203,I8724,g11258,g8825,g2872,I6489,g3334,g4334,g5257,g7354,g10535,g4070,g8269,g6874,g7993,g4427,g3118,g10560,I15063,g6876,g5479,I9046,g11228,I8911,I13834,g4099,g5360,g2131,g1570,g6564,g1718,g1941,g4737,g4872,g4459,g2538,g4055,g5483,I15817,g11174,g1968,g10870,g9532,g3583,g9692,g6347,g1432,g4322,I11005,I10123,g9765,g8508,I11249,g10347,g10686,I9185,g1854,g6243,g9679,I5395,I13553,g3523,g11341,g7895,g2274,g1389,g6950,g10737,I6337,I10941,g8732,g11005,g8074,g8418,I10177,I12354,I9766,I11029,I9320,I14509,I6531,g525,g10567,g3497,g11600,g8839,g2521,I9712,I11162,I12177,g11381,g3322,I11569,g8475,I7303,g11615,g9592,g10681,I10051,g4435,g5641,I14123,g7965,g7279,g5508,g4565,g1296,g7621,I5135,I8605,g10278,g4047,g6896,g8680,I5092,g7146,g8274,I12439,g11181,I9338,g10342,I5867,g4054,I8676,g4514,g7850,g1121,g4451,g1905,g5538,I12526,g6304,g6220,g1711,I15042,g10594,I10655,I17746,g1380,I11807,g2640,I9427,g5616,g5671,I8528,I10033,g10143,g1027,I15275,g9874,g1068,g7970,I8311,I9953,g4749,g8513,g2269,g5842,g9780,I8136,I6256,g5026,g8264,g11619,I13900,I16650,g2908,g8218,g8604,I13552,g3816,g4757,I10546,I16105,g11111,g10414,I6523,g1660,g9009,g6522,g7989,g10164,g5745,g10489,g6734,I9598,g11449,I9023,g4270,g4106,g4271,g11500,g845,g5184,I15467,I13485,g8282,g11640,g7560,I10610,I4886,g9980,I7213,g4243,I7288,g8485,I14391,g11445,g5143,I12322,I13397,g10391,g6420,g2328,I7009,I17504,g3717,g7534,I7746,g7191,g10701,g9959,g7328,g8700,I4978,g2226,g10392,g9351,I12565,g7678,g4187,g127,g1604,g6931,g2544,I5104,g3422,g5535,g2297,I15861,g7057,g6544,g4920,I16953,I13259,g11186,I14697,g7853,I7441,g883,g7846,g5042,g6290,I11829,g2316,I11743,g2076,I16172,I9731,I8414,g6122,g10521,g5419,g9746,g8302,g11176,I7523,g9338,g2562,g11614,g5826,g3436,g4878,I5513,I15736,I12190,g9920,g1486,g2304,g7505,g2777,I10888,I17249,I12544,I12989,g7934,g9963,g8404,g6825,I12251,g5801,g8793,g10254,g10130,I16001,g7916,g3386,I15907,g9595,g11204,I13421,I11916,I10495,g8884,g7478,g2958,I7456,I11464,g6791,I11605,I7876,g10912,g11233,g7310,g8137,g7473,g7027,I6760,I5707,I9276,g4630,g2071,g1678,I14400,g2197,I16007,g5731,g4607,I6639,g7793,g11067,g7030,I17182,g5485,g6548,g7530,I13242,g5173,g10361,g2045,g5260,g5589,g9731,g2364,g6748,g7962,I11275,g11657,g5645,I12056,g10279,g8550,g968,g6063,g11464,g5987,g8781,g3496,I8606,g11387,g10385,g33,I11477,I7240,I10633,I16685,I6979,g4381,g4336,g9827,g10477,g11231,g2055,g8184,g4300,g12,g2847,g3636,g4309,g4068,I15900,g2249,g7183,g10166,I11180,I16031,g4556,g6549,g2773,I7487,g3461,g6324,I5970,I10171,g3774,I12360,g6919,I14573,g6531,I14224,g4416,g9651,g3742,I15608,g4788,I10153,g3762,g5119,g5531,g5027,g5722,I13785,I17191,g174,I11950,g7069,g4894,I16087,g11016,I15427,I7946,I15451,g8737,I11214,g3945,g9646,g8299,g8451,g10194,g857,g6083,g5305,I9305,I6844,I6288,g10533,g2119,g11248,g8699,g10378,I17487,I8333,g8014,g7767,g7941,I6569,g2421,g5791,g11514,g7232,I7351,I17344,g6239,g5501,g5067,g9192,I14105,g70,g8009,I15820,g1095,I12029,g11229,g546,g7035,I12822,I10873,g4522,g5532,g9751,g3395,I16461,I8275,g6307,I5165,g2881,g10381,I13002,g6772,g2795,g7189,g2955,g10291,g959,g10909,g10626,I15389,I11094,I16292,g8077,g7891,I13280,I10553,I9620,g8735,g8194,g1223,I14579,I16095,g6573,I9727,g8752,g10475,g4899,g3631,g1796,g5591,g8707,I10048,I7593,g9271,I15296,g7825,g11595,g6513,g8649,I7817,I7112,g10074,g6777,I15798,g7460,g7951,g5097,g8935,I11783,g8145,g7558,I13592,g4477,g9453,g7055,g6759,I5865,I5728,I6143,g3404,I8396,g6216,g7769,I9559,I13457,g4365,g8055,g11635,g11587,g8750,I8421,g2882,g1436,I12853,I15437,g1374,I5561,I15278,I14802,g10368,g135,I5036,g10032,g6749,g6868,g5196,g6530,g6093,g7781,I9810,g4141,g8278,g7543,I16356,I9032,g9745,g8847,g10779,I8456,g6817,g4618,I12694,g11431,I12279,I5837,g7844,I16065,g8674,I9923,I7999,g6354,g7807,g6166,g4289,g6633,I6188,g10170,g9734,g3364,g4371,g10935,I17528,I6208,g9655,g9624,g6045,g5361,g2210,g8627,g11573,g5911,g10687,g5509,I7034,g2157,g9910,I15559,g10326,g9358,g110,g5534,g2941,I8717,g8051,I12076,g10537,g4831,g3336,g5353,g11199,g11558,g2083,g4474,g575,g11283,g7894,g8481,I11635,I7920,g354,g452,g7212,I14684,g4295,g11223,g928,g10290,I16181,g3374,g9867,g11009,g7220,g7362,g10211,g8214,g11406,g2965,I7771,g6082,I12817,g6820,g11164,I5529,g3771,g37,I17770,g7454,I6818,g8743,g1333,I6209,g7314,I12108,g5673,g6247,g11041,g1621,g4512,I5833,I14614,I10693,g2845,g9614,I17531,I15257,g3041,g11585,g1543,I14918,g9807,I7387,g8322,I5254,g4,g8039,g2511,g5848,g4827,g7241,I12344,g6790,I11146,g10851,g3051,g5420,g11264,g5663,g4987,g11297,g5241,g3546,g1589,g9267,g11211,I12136,g10169,g5586,g3337,g7141,g9663,g5886,g2516,g1759,I15200,g10746,g6878,g9347,g4602,g6301,I9093,g5125,g2419,g1991,g7910,g11417,I4859,g6355,g4331,g2168,I13776,g11201,I4910,g7907,g7957,g10359,I16203,I7224,I13560,I11596,g2438,g7431,g11401,g11408,I11238,g5603,g8450,g10769,I14204,g1440,g3254,g5424,I10314,I4912,I13005,I16307,I14182,g6857,g3684,I6074,I16370,g5984,I9491,g10796,g7458,I8545,g4267,g11187,g4669,g8973,I10060,g6826,I6159,g5597,g6313,g10133,I8515,I12586,g8387,g1235,g4970,g7126,g333,I5468,g6756,g8556,g11302,g8094,g11202,g10063,g6747,g2518,I10398,g2050,g4508,g6757,I10843,g5223,I7697,g11025,I15258,g3695,g10683,I13090,g4391,g4062,g7501,I17494,I17185,g10642,I13364,g6400,g6286,g11207,g2258,g9622,g9762,g4230,g4534,g6338,I9208,I12793,g8797,g9604,g11320,g10197,g1976,I9199,g3275,g10234,g590,I9141,g6914,I5296,g10899,I16941,I13831,I15562,g1733,g9812,g6869,I6031,g8870,I12568,g11190,I15615,I10601,I7825,g4771,g7414,I17324,g9103,g7218,g11424,g2620,I9362,I5366,I12235,g6634,I8126,g5245,g4941,g2803,g5728,g6031,g6246,g4144,g2123,g5255,g4065,I5470,I9237,I5013,g6431,g8697,g10153,I7300,g6309,g7264,I12541,I7151,g7439,g10616,g2844,I5862,g8614,g1400,I11279,g6248,g8419,g2336,I17268,I6317,g4974,I7378,I6821,g290,g8954,I9673,g2956,g11162,g10507,g3708,g7078,I9302,I12478,g10373,I13539,g7544,g4325,g7231,g5218,I13741,I4777,I14270,g4066,g5473,I10248,g5863,I6193,g8961,g5177,g6886,I16149,I14077,g11045,g10772,g650,g10350,I6016,I4938,I10445,g1403,g7726,g1999,I8778,g7358,I10141,I14473,g9530,I7336,g7076,g1129,I15607,g4807,g6684,g8060,g5910,g10513,g822,I9053,g6576,g9949,g5555,g995,g4727,g11313,g6044,g8560,g6641,g6924,I13523,g6514,g8712,g9825,I6888,g5948,g3863,I5111,g8826,g1444,g8447,g10058,g4491,g9936,g97,g7570,g10630,g6935,I5591,g10850,I11804,g197,I8604,g6468,g7562,I15980,g6448,g2023,g7131,I16124,I11289,I5798,g11154,g5754,g6165,g4889,g7918,I5324,g8927,I5929,g9859,I8161,g6080,I17485,g3683,I15470,g5344,g3632,g9310,g4377,g3874,g7933,I6224,g6795,I11367,g4472,I11243,g2530,g10458,I11953,I15220,g10168,g7453,I12652,g11645,I14236,g6705,g6118,I13666,g9721,I7061,g1044,g461,I11505,g6245,I15253,g10374,I17438,g6702,I11296,g6202,g5937,g10327,g11015,I14306,g8353,g8308,g9754,I12289,g869,g11083,g2727,g4562,g4160,g6828,g10448,g6064,g1215,g8810,g9728,g3625,g5520,I6398,I14278,I6480,I8490,g5118,g4095,g8571,g3113,I16856,I17347,g7348,I9786,g6540,g8966,g7760,g6481,I13326,g6449,g1397,g8261,I11315,I13515,I12505,g10259,I5308,g9390,I15795,g8813,g7525,g1411,g8292,I14694,g10923,I11617,g8742,g9769,g4238,g6430,g5423,g4506,g7880,I13909,I13125,g4282,g1255,g6980,I12904,g8048,I13867,I8340,I16859,I12871,g2099,g2508,g9994,g8130,g3092,g5256,g4582,g1771,I6201,g5390,g8924,g4237,g8613,g2763,g9898,g8642,g7609,g3071,g8289,I10296,g3907,g8298,I12829,g105,I7863,I6870,g7661,g5810,g7074,g7425,I10174,g6014,g4940,g10682,I12936,g7531,g10329,I9273,I8320,g7036,g1840,g3435,I7906,g8817,I15458,g4468,I8487,I11752,g5543,g6427,g11299,I7444,g7540,g8724,I16739,g8727,g5734,g4720,g4279,g10604,g9823,I16086,I15415,g8603,g9265,g5892,g2190,g4804,g7298,I9795,I13606,g11609,g6388,I13531,g4367,g5319,g3664,g10244,I7459,I13859,g9908,g7995,g3067,g5744,g8553,g6882,g4637,g6092,I7191,g8962,g9447,I7732,I9642,g2834,I10317,g4374,g4774,I9415,g8788,g2695,I17543,g9826,g4954,I14668,I9486,I8779,g192,g6671,g2155,I12472,g2213,g1250,I8982,g7677,g11106,g10595,g10159,g5762,g2002,g336,g8963,I13642,g5050,I7064,g8990,I8506,g11301,I13878,g225,I5014,g3220,g3323,g2638,I12901,g3371,I14477,g4143,I5435,g10509,g7849,g10316,g7660,g10908,I5821,g8623,g2798,I5909,g5168,g636,g4549,g6296,g9857,g1741,I13385,I12103,g6854,g7922,g7415,I5638,g1035,I11967,g2918,g11288,g10658,g1834,g2912,I12242,g9428,g2350,I11173,g10674,g2160,I4986,g6213,g10232,g11484,I10931,g8822,g52,g3767,I9836,g2649,g9671,I9956,g4460,g9344,g4759,g8885,I7468,g7197,g6711,I11103,g2243,I11357,g10802,I14080,I17500,g4588,g3734,g10729,g170,g7285,g1386,g11553,g8070,g10040,I14602,I13427,g7943,I11908,I17216,I10584,g11488,g8733,I17716,g11033,g5296,g6835,g5545,I11873,g8196,g7681,I14409,g11579,g6543,g8695,I5424,I15359,g6821,g6226,g7450,g10806,g8842,I6952,g1727,I10736,g7459,g10971,g8007,g5198,g5051,I15688,I15548,g10622,g10505,g3281,I5619,g139,I10930,g5604,I13203,g5548,g11108,g7479,I11412,g627,g5540,g2390,g9869,g5890,g501,g10499,I6921,I11647,g4952,I10822,g10473,g9873,g11654,I6971,g10034,g4977,g4442,g11637,I16589,g10765,g8786,g2528,I14613,I11252,g391,g11062,g7977,g4299,g5185,g8923,g4113,g2525,g6694,g2871,g8650,I11011,g10175,g6100,g8956,I5064,g6079,I15432,g9257,I16206,g10460,I17736,g4680,I10949,g4009,g11329,g7290,g3384,I14961,g11552,g8573,I11537,I11055,I4966,I10186,g5011,g4413,g10468,g5615,g9030,I13624,I7875,g7616,g9842,I10018,g7032,g6689,I9084,g4819,I10195,I17558,g6830,g5183,g7140,g4115,I15431,I6762,I8880,g4004,g2001,g11191,g1891,g7287,I11021,I10966,g5797,I12981,g3292,g7555,g6680,I17206,g6700,g6880,g10098,g3627,g10697,g2563,g2259,g4290,g6541,I14299,g11324,g511,g2382,I9576,g4073,g10675,g6814,I5323,I15272,g6206,g7304,I9505,g6214,I9680,I15771,g10375,I10102,g10190,g6750,g4457,I9461,g4077,g8716,g718,g11110,g9715,g5733,g5188,g8036,g5417,g6703,I10114,g9256,g7718,g6192,I11489,g8729,I5373,g6292,g9654,g10450,I9946,I9510,g9593,g6740,I13367,I11980,g736,g8926,g7457,g1160,g312,g5670,g10308,I17225,g10435,g4184,g11643,I7429,I5438,I5570,g8708,g7533,I17331,g5893,g11007,I11201,g8342,g9607,g2437,g10354,g11466,g8582,g9901,g9759,g8409,g2961,g2617,g7444,I5185,g5573,I10054,I14855,I11440,g330,I15362,g7612,g3516,g2237,g5665,g6350,I5050,g7093,I8199,I17219,g9650,I10932,g2917,I9399,I9077,g10135,I14552,I15162,g2178,g6591,g8878,I16871,g865,g5398,g9308,I11217,I5809,g4768,g2998,g3703,g6231,g5897,g2187,I13633,g4902,I16947,g4893,g8765,g9879,I17282,g4520,g6930,I9842,g7148,g11647,g2132,I5024,g6217,g10128,I17492,I8495,g11410,g5182,g6123,I10378,I17407,I5116,I12430,g7817,g7060,I15872,g6157,I15326,g10798,g4076,g10065,g3776,I6414,I8499,g2241,g11593,g6788,g11555,g4058,I17755,g6827,g7322,g4529,I9001,I15823,g9917,g8883,I6947,g327,g8717,g9429,g10189,I5886,g6026,g4886,g11412,I15048,g7930,g9652,g8221,g4933,I5035,g6140,I12634,g5556,g7680,g3266,g6623,I13559,I8811,g4876,g4971,g9669,g2006,g8824,I10666,g8426,g10803,I6391,g8843,g8050,g4093,g1666,g1561,g10780,g4877,g4307,g8438,g10428,I8738,g3208,g2230,g6434,g7133,g6574,g4766,I16553,I9332,g6413,g9027,g9940,g2199,I9669,g10268,I13357,g3629,g7124,I7513,g2236,g7795,I15196,I6331,I10682,I6643,g2641,g10776,g5405,g7703,I15871,I12762,g3800,g10712,I8750,I10240,g6660,g10252,g8024,g11465,I12009,g7900,g1672,I13505,g8348,I11269,g9573,g401,g1627,g7472,g2653,g5853,g3764,g7386,g2790,g2725,g7300,I7701,I12087,g6333,g11346,g11457,g1534,g7940,g5795,g6738,g10598,g11578,g7976,g8384,I11578,I15341,g11253,g7737,g11339,g6410,g9510,g1994,g10188,I12199,g6162,I6439,g8841,I12644,g5181,I16598,g3038,g4890,I8278,g8688,g10179,g143,g11472,g6441,g10907,g8019,I7636,g7584,g10619,I11169,I13454,g11342,g10744,g7353,I6932,g5489,I17586,g11432,I14119,I7414,g7734,g5632,g10896,g5692,g2306,g6587,g10807,g10511,g10624,I16676,I5352,g7905,g9885,g6451,g5175,g11396,I9191,g8320,g10376,g8379,g3721,g10792,g9913,g10719,g4828,g2031,g4779,g7327,g5884,g2173,I9074,g9708,I12487,I7399,g853,g9263,g10818,I13475,I6510,g3111,g4316,g1558,g5766,I7339,g11082,g6644,g9841,g5782,I11207,g11474,g10787,g10393,g10280,g9695,g6883,g8720,I12150,I13309,g9417,g7369,g11351,I13674,g5788,g11053,I5795,I11322,I17767,g2216,I14323,g6329,g8102,I15787,g7909,g6110,g3815,I17289,g11458,g3097,g11649,I15344,g11631,I9317,g219,g9557,g11008,g4726,g2087,g7025,g691,g10183,I6738,I5224,g1361,I11632,g5936,I13344,g5270,I5966,g4934,g4169,g7271,g5537,g10267,g3518,g8827,g10241,g11291,g8461,I9804,g6132,g7440,I11650,I13609,g9108,I5658,I9346,g2632,I5399,g10420,I6754,g6723,I6999,I9880,g8310,g5523,g9878,g5819,g6961,g9385,g2756,g7052,I17758,g5084,g8687,g3905,g26,g6016,g11559,I6891,g639,g11467,g4012,g4758,I10592,I7877,g5213,g3375,I12145,g11392,g6316,I10340,I12547,I15127,I8919,I11309,g10369,g6098,I7668,I5388,g4786,g9956,g4005,I6173,g7403,g11575,g9775,g10266,I12655,I11626,g10800,g10091,I7654,I8842,g4548,g7788,g5876,g10287,I17563,g2109,g4489,I12427,I7173,I5372,I6178,g878,g11460,g5995,g5280,g8018,g2853,g5170,I12208,g6701,g7709,g10306,g6503,g4466,g10160,I5198,g11322,g4429,g262,g10298,g2826,g11628,g11198,g7438,g6832,g1552,g8356,g8763,I8804,g8063,g7811,g4803,g9079,g3545,g2481,I10991,I13918,g9384,g10880,g5780,g7942,g5666,g7237,I17733,g4240,g6663,I8678,I9866,g11236,I6052,g10447,I7625,g10417,g11260,g8120,g3747,g11278,g5224,g360,I11417,I6183,I14418,I16432,g8433,g10062,I16638,g5102,g10561,g11031,g11363,I11198,I4876,g9984,I7070,g9522,g11281,I8503,I10183,I4894,g4310,I14412,g3628,g10466,g8607,g5885,g4874,I17252,g3989,I13117,g6331,I15332,g971,g10552,g8420,g7377,g7545,g4537,I7393,I10325,g2543,g8548,g8869,I16037,I16790,I6520,g7047,g2748,g3634,g10928,g7368,g8226,I10648,I12610,g11048,g10256,g7364,g5827,g4251,g8047,g5850,g4932,g8248,g1574,g4714,g3039,g6364,g4765,g1330,g2529,g8105,I11152,g10730,g8554,g10474,g9536,I13779,g3623,g10145,I8562,g8345,g7125,g2219,g3681,I5304,g9720,g6072,I7665,g8696,g1512,I6517,g10064,g10319,g8821,g4780,g2342,I4866,g8671,g6405,I14211,I16200,I8240,I10352,g8499,g9387,I10036,g5575,g2102,g6208,I14191,I7858,g2257,g6569,g7258,g4167,g7346,I13131,I4995,g8068,I13114,g3707,g3757,g1849,I14228,g6097,g5215,g6124,I11756,I16507,g2040,I15409,g4822,g2439,g11507,g2260,I6876,g6897,g8079,I13521,g1927,g4390,g11436,I6277,g10584,g7352,I8039,g2915,g11641,g6201,g1684,I9029,g8171,g8288,g6811,g7065,I13460,g6102,g8766,I6806,I17516,g1053,g9929,g9566,I11770,g10705,I5695,g5262,I13249,I12086,g6727,I15756,I14970,I16190,I11194,g11179,I8889,I13317,I11689,g9556,g10597,g5836,I6746,g9844,I9153,g9724,g9661,g6023,g2613,g11271,g10334,g7477,g9907,I5528,g7343,g3430,g10208,g9274,g2011,g6101,g4906,g5271,I16583,g5044,I5804,g1721,I11024,g11321,I10367,g4672,g6670,g10476,g6802,g6993,g7600,I6624,g2828,g6234,g5120,I12133,g10162,g3544,g8828,g22,g10785,g3096,I16413,I9326,I13191,g9960,I11996,I17121,g6894,g10518,g7020,I5854,g3408,g7561,g10592,g947,g7664,I12092,g6808,I4971,I9129,I16079,g11515,g9911,g5047,g8180,g11485,g6771,I15959,g6349,g8871,g9617,g8663,g3971,g6076,I17202,g5794,g8514,g4510,I15801,I17585,g2455,g2817,g260,g6922,g9473,g10673,I9581,g9686,I15057,I8786,g11380,g5612,g6053,g3214,I5047,g2244,I15284,g6335,I12032,g10356,g2231,g5075,g9659,g4431,g9292,g3103,g7982,g2500,g2713,I9365,g9712,g7746,g5841,g2751,g6626,I11695,g1448,g7427,g5730,g849,g6190,g2561,I16255,I15545,g3694,I15473,g5618,I6767,I11132,I10278,I5919,I17124,g1206,g10927,g11544,g2683,I9080,g11512,I12971,I10914,I15187,I5606,g6940,g7747,g10281,g4386,g3661,I6071,g11252,g7077,I17441,g2196,g1639,g4544,g9854,g5865,g8366,g4551,g7043,g6340,I13941,g3359,g3730,g10207,g6047,g7476,I6040,g4805,g4867,g7375,I17695,I12107,g2570,g3586,I8788,g10547,g11193,g8848,g1959,g11354,g6042,g3543,g8033,g9821,g9858,g8959,g11042,I8544,I16416,I13274,I8285,g7649,I13886,g7752,g8277,I5801,I7076,g10672,g1822,g6654,I15406,g2907,g2946,I15598,I7600,g2181,g1227,I10135,I13537,g10041,g6423,g5426,g5249,g6568,g6328,g10202,g6964,g4318,I6665,g11257,g7046,g8182,g673,I13782,I13726,g4596,I17096,g11195,g5628,g3782,g5211,g11298,I10093,g11238,g4790,g5982,g5630,I6679,I6176,g4679,g2801,g727,I5626,g1209,g7955,g8945,I13283,g8723,I13442,g253,g1848,g5847,g9803,g9987,g4555,g10721,g6419,g11076,g4284,g4337,g11422,g8471,g2112,g4509,g5779,g11259,g11013,g2859,I17435,I10381,I15488,g8107,g5267,g8747,g4415,g2320,g5719,g4218,I5461,g440,g4183,I16487,I14910,I17295,g5229,g6480,g11551,I16330,g2910,g4993,I12535,I9639,g9173,I5963,g10452,I13379,g7720,I17453,I9341,I14263,I9602,g7991,g7135,g7432,g5186,g4384,g3760,I9253,g3513,g9933,I7952,g9701,g11475,I12641,g4776,g2888,I14218,g5916,I7384,g9649,I16252,g6061,I6501,g4764,g7365,I11436,g3758,g1107,g2205,g9716,I15392,I5604,I5251,g11078,I15383,g7184,g9606,g9259,I12388,I10713,g3637,g16,g3804,I13424,g9816,g5476,g8993,I12300,g6685,I13530,g4281,g7185,g2813,g7312,g7728,I13200,g5896,g7341,g10723,g6921,g11285,g284,g8224,g2176,g7568,g4782,g6250,g3728,I16264,g10332,I9754,I5414,g3227,I14564,g5677,g9262,g7096,g5194,g8794,I12751,g11542,g2272,g9906,g342,I10719,g7628,I9965,g7195,I10729,I5289,g9106,g11606,g646,g2017,g3975,g8756,g10540,I7249,g1747,I5101,I8614,g2523,I10039,g2407,g10767,g4778,I8388,I5166,g4326,g3215,g10364,I7438,I10129,g4518,g6095,g8000,I10434,g5146,g11265,I15669,g10740,I17749,g11105,I17764,I16114,g10627,g6908,g2639,I7776,g5675,g10229,g9426,g806,g4269,I11427,I10192,g9924,g8549,I9992,g11549,g3828,g6057,I15691,I13185,g5949,g6533,g6219,g4002,I14040,g7980,g6096,g5078,g10695,g10230,g5567,g1365,g7778,I11088,I6901,g6570,I16045,g5574,g3253,g6149,g8698,g4383,g2952,g6151,g8164,g5614,g2948,g10633,I12773,I17591,g10903,g4102,g3257,g10526,I6226,g2073,g8071,g2964,I9056,g10930,g8746,g8520,I16595,g7914,g2732,I12120,I6572,g7892,I17371,g981,g10791,g11261,I5137,I6363,g243,I12589,I9323,g10335,g8052,g4711,I13255,g10115,I8410,g2165,I5538,I7220,I10231,g4519,I12127,g10575,g10464,I9256,g1969,g2459,I9564,g3267,I12469,g3987,I10126,g6592,g10786,I6827,g4341,g7877,g3256,g10286,g6899,I15698,I14546,g4462,g7634,g10708,g7130,I17353,g7278,I8050,I6299,I14452,I8827,I13682,g396,I13102,g10774,I14490,g6579,I15878,g10438,I17390,g7419,I16073,g1275,I6330,g745,I11263,g9324,g5805,g5667,g10861,I10066,g7881,g4157,g8126,g8064,g5301,g8005,I6837,g10237,I9475,g5288,g10819,g9264,g7097,I14394,g8422,I6367,g2122,g10639,I7847,g770,g8714,I7318,g5038,g3990,g8244,g8646,g10079,g10144,g6954,g3501,g5261,I6807,g8142,g5631,g8249,g11580,I15114,I11091,g8386,I15906;
//# 77 inputs
//# 150 outputs
//# 534 D-type flipflops
//# 6324 inverters
//# 3448 gates (1619 ANDs + 968 NANDs + 710 ORs + 151 NORs)
//
//
//
  MSFF DFF_0(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1289),.DATA(g5660));
  MSFF DFF_1(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1882),.DATA(g9349));
  MSFF DFF_2(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g312),.DATA(g5644));
  MSFF DFF_3(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g452),.DATA(g11257));
  MSFF DFF_4(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g123),.DATA(g8272));
  MSFF DFF_5(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g207),.DATA(g7315));
  MSFF DFF_6(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g713),.DATA(g9345));
  MSFF DFF_7(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1153),.DATA(g6304));
  MSFF DFF_8(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1209),.DATA(g10873));
  MSFF DFF_9(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1744),.DATA(g5663));
  MSFF DFF_10(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1558),.DATA(g7349));
  MSFF DFF_11(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g695),.DATA(g9343));
  MSFF DFF_12(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g461),.DATA(g11467));
  MSFF DFF_13(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g940),.DATA(g8572));
  MSFF DFF_14(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g976),.DATA(g11471));
  MSFF DFF_15(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g709),.DATA(g8432));
  MSFF DFF_16(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1092),.DATA(g6810));
  MSFF DFF_17(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1574),.DATA(g7354));
  MSFF DFF_18(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1864),.DATA(g7816));
  MSFF DFF_19(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g369),.DATA(g11439));
  MSFF DFF_20(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1580),.DATA(g7356));
  MSFF DFF_21(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1736),.DATA(g6846));
  MSFF DFF_22(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g39),.DATA(g10774));
  MSFF DFF_23(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1651),.DATA(g11182));
  MSFF DFF_24(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1424),.DATA(g7330));
  MSFF DFF_25(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1737),.DATA(g1736));
  MSFF DFF_26(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1672),.DATA(g11037));
  MSFF DFF_27(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1077),.DATA(g6805));
  MSFF DFF_28(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1231),.DATA(g8279));
  MSFF DFF_29(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g4),.DATA(g8079));
  MSFF DFF_30(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g774),.DATA(g7785));
  MSFF DFF_31(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1104),.DATA(g6815));
  MSFF DFF_32(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1304),.DATA(g7290));
  MSFF DFF_33(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g243),.DATA(g7325));
  MSFF DFF_34(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1499),.DATA(g8447));
  MSFF DFF_35(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1044),.DATA(g7789));
  MSFF DFF_36(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1444),.DATA(g8987));
  MSFF DFF_37(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g757),.DATA(g11179));
  MSFF DFF_38(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g786),.DATA(g8436));
  MSFF DFF_39(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1543),.DATA(g7344));
  MSFF DFF_40(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g552),.DATA(g11045));
  MSFF DFF_41(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g315),.DATA(g5645));
  MSFF DFF_42(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1534),.DATA(g7341));
  MSFF DFF_43(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g622),.DATA(g9338));
  MSFF DFF_44(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1927),.DATA(g9354));
  MSFF DFF_45(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1660),.DATA(g11033));
  MSFF DFF_46(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g278),.DATA(g7765));
  MSFF DFF_47(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1436),.DATA(g8989));
  MSFF DFF_48(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g718),.DATA(g8433));
  MSFF DFF_49(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g76),.DATA(g7775));
  MSFF DFF_50(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g554),.DATA(g11047));
  MSFF DFF_51(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g496),.DATA(g11333));
  MSFF DFF_52(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g981),.DATA(g11472));
  MSFF DFF_53(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g878),.DATA(g4896));
  MSFF DFF_54(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g590),.DATA(g5653));
  MSFF DFF_55(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g829),.DATA(g4182));
  MSFF DFF_56(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1095),.DATA(g6811));
  MSFF DFF_57(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g704),.DATA(g9344));
  MSFF DFF_58(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1265),.DATA(g7302));
  MSFF DFF_59(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1786),.DATA(g7814));
  MSFF DFF_60(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g682),.DATA(g8429));
  MSFF DFF_61(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1296),.DATA(g7292));
  MSFF DFF_62(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g587),.DATA(g6295));
  MSFF DFF_63(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g52),.DATA(g7777));
  MSFF DFF_64(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g646),.DATA(g8065));
  MSFF DFF_65(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g327),.DATA(g5649));
  MSFF DFF_66(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1389),.DATA(g6836));
  MSFF DFF_67(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1371),.DATA(g7311));
  MSFF DFF_68(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1956),.DATA(g1955));
  MSFF DFF_69(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1675),.DATA(g11038));
  MSFF DFF_70(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g354),.DATA(g11508));
  MSFF DFF_71(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g113),.DATA(g7285));
  MSFF DFF_72(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g639),.DATA(g8063));
  MSFF DFF_73(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1684),.DATA(g11041));
  MSFF DFF_74(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1639),.DATA(g8448));
  MSFF DFF_75(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1791),.DATA(g8080));
  MSFF DFF_76(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g248),.DATA(g7323));
  MSFF DFF_77(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1707),.DATA(g4907));
  MSFF DFF_78(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1759),.DATA(g5668));
  MSFF DFF_79(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g351),.DATA(g11507));
  MSFF DFF_80(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1957),.DATA(g1956));
  MSFF DFF_81(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1604),.DATA(g7364));
  MSFF DFF_82(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1098),.DATA(g6812));
  MSFF DFF_83(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g932),.DATA(g8570));
  MSFF DFF_84(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g126),.DATA(g5642));
  MSFF DFF_85(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1896),.DATA(g8282));
  MSFF DFF_86(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g736),.DATA(g8435));
  MSFF DFF_87(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1019),.DATA(g7807));
  MSFF DFF_88(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1362),.DATA(g7305));
  MSFF DFF_89(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g745),.DATA(g2639));
  MSFF DFF_90(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1419),.DATA(g7332));
  MSFF DFF_91(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g58),.DATA(g7779));
  MSFF DFF_92(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g32),.DATA(g11397));
  MSFF DFF_93(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g876),.DATA(g878));
  MSFF DFF_94(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1086),.DATA(g6808));
  MSFF DFF_95(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1486),.DATA(g8444));
  MSFF DFF_96(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1730),.DATA(g10881));
  MSFF DFF_97(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1504),.DATA(g7328));
  MSFF DFF_98(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1470),.DATA(g8440));
  MSFF DFF_99(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g822),.DATA(g8437));
  MSFF DFF_100(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g583),.DATA(g6291));
  MSFF DFF_101(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1678),.DATA(g11039));
  MSFF DFF_102(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g174),.DATA(g8423));
  MSFF DFF_103(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1766),.DATA(g7810));
  MSFF DFF_104(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1801),.DATA(g8450));
  MSFF DFF_105(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g186),.DATA(g7317));
  MSFF DFF_106(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g959),.DATA(g11403));
  MSFF DFF_107(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1169),.DATA(g6314));
  MSFF DFF_108(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1007),.DATA(g7806));
  MSFF DFF_109(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1407),.DATA(g8993));
  MSFF DFF_110(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1059),.DATA(g7794));
  MSFF DFF_111(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1868),.DATA(g7817));
  MSFF DFF_112(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g758),.DATA(g6797));
  MSFF DFF_113(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1718),.DATA(g6337));
  MSFF DFF_114(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g396),.DATA(g11265));
  MSFF DFF_115(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1015),.DATA(g7808));
  MSFF DFF_116(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g38),.DATA(g10872));
  MSFF DFF_117(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g632),.DATA(g5655));
  MSFF DFF_118(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1415),.DATA(g7335));
  MSFF DFF_119(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1227),.DATA(g8278));
  MSFF DFF_120(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1721),.DATA(g10878));
  MSFF DFF_121(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g882),.DATA(g883));
  MSFF DFF_122(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g16),.DATA(g4906));
  MSFF DFF_123(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g284),.DATA(g7767));
  MSFF DFF_124(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g426),.DATA(g11256));
  MSFF DFF_125(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g219),.DATA(g7310));
  MSFF DFF_126(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1216),.DATA(g1360));
  MSFF DFF_127(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g806),.DATA(g7289));
  MSFF DFF_128(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1428),.DATA(g8992));
  MSFF DFF_129(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g579),.DATA(g6287));
  MSFF DFF_130(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1564),.DATA(g7351));
  MSFF DFF_131(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1741),.DATA(g5662));
  MSFF DFF_132(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g225),.DATA(g7309));
  MSFF DFF_133(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g281),.DATA(g7766));
  MSFF DFF_134(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1308),.DATA(g11627));
  MSFF DFF_135(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g611),.DATA(g9930));
  MSFF DFF_136(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g631),.DATA(g5654));
  MSFF DFF_137(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1217),.DATA(g9823));
  MSFF DFF_138(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1589),.DATA(g7359));
  MSFF DFF_139(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1466),.DATA(g8439));
  MSFF DFF_140(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1571),.DATA(g7353));
  MSFF DFF_141(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1861),.DATA(g7815));
  MSFF DFF_142(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1365),.DATA(g7307));
  MSFF DFF_143(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1448),.DATA(g11594));
  MSFF DFF_144(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1711),.DATA(g6335));
  MSFF DFF_145(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1133),.DATA(g6309));
  MSFF DFF_146(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1333),.DATA(g11635));
  MSFF DFF_147(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g153),.DATA(g8426));
  MSFF DFF_148(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g962),.DATA(g11404));
  MSFF DFF_149(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g766),.DATA(g6799));
  MSFF DFF_150(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g588),.DATA(g6296));
  MSFF DFF_151(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g486),.DATA(g11331));
  MSFF DFF_152(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g471),.DATA(g11469));
  MSFF DFF_153(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1397),.DATA(g7322));
  MSFF DFF_154(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g580),.DATA(g6288));
  MSFF DFF_155(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1950),.DATA(g8288));
  MSFF DFF_156(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g756),.DATA(g755));
  MSFF DFF_157(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g635),.DATA(g5656));
  MSFF DFF_158(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1101),.DATA(g6814));
  MSFF DFF_159(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g549),.DATA(g11044));
  MSFF DFF_160(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1041),.DATA(g7788));
  MSFF DFF_161(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g105),.DATA(g11180));
  MSFF DFF_162(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1669),.DATA(g11036));
  MSFF DFF_163(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1368),.DATA(g7308));
  MSFF DFF_164(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1531),.DATA(g7340));
  MSFF DFF_165(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1458),.DATA(g7327));
  MSFF DFF_166(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g572),.DATA(g10877));
  MSFF DFF_167(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1011),.DATA(g7805));
  MSFF DFF_168(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g33),.DATA(g10867));
  MSFF DFF_169(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1411),.DATA(g7331));
  MSFF DFF_170(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1074),.DATA(g6813));
  MSFF DFF_171(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g444),.DATA(g11259));
  MSFF DFF_172(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1474),.DATA(g8441));
  MSFF DFF_173(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1080),.DATA(g6806));
  MSFF DFF_174(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1713),.DATA(g6336));
  MSFF DFF_175(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g333),.DATA(g5651));
  MSFF DFF_176(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g269),.DATA(g7762));
  MSFF DFF_177(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g401),.DATA(g11266));
  MSFF DFF_178(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1857),.DATA(g11409));
  MSFF DFF_179(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g9),.DATA(g7336));
  MSFF DFF_180(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g664),.DATA(g8782));
  MSFF DFF_181(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g965),.DATA(g11405));
  MSFF DFF_182(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1400),.DATA(g7324));
  MSFF DFF_183(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g309),.DATA(g5652));
  MSFF DFF_184(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g814),.DATA(g8077));
  MSFF DFF_185(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g231),.DATA(g7319));
  MSFF DFF_186(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g557),.DATA(g11048));
  MSFF DFF_187(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g586),.DATA(g6294));
  MSFF DFF_188(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g869),.DATA(g875));
  MSFF DFF_189(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1383),.DATA(g7316));
  MSFF DFF_190(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g158),.DATA(g8425));
  MSFF DFF_191(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g627),.DATA(g5657));
  MSFF DFF_192(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1023),.DATA(g7799));
  MSFF DFF_193(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g259),.DATA(g7755));
  MSFF DFF_194(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1361),.DATA(g1206));
  MSFF DFF_195(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1327),.DATA(g11633));
  MSFF DFF_196(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g654),.DATA(g8067));
  MSFF DFF_197(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g293),.DATA(g7770));
  MSFF DFF_198(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1346),.DATA(g11656));
  MSFF DFF_199(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1633),.DATA(g8873));
  MSFF DFF_200(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1753),.DATA(g5666));
  MSFF DFF_201(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1508),.DATA(g7329));
  MSFF DFF_202(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1240),.DATA(g7297));
  MSFF DFF_203(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g538),.DATA(g11326));
  MSFF DFF_204(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g416),.DATA(g11269));
  MSFF DFF_205(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g542),.DATA(g11325));
  MSFF DFF_206(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1681),.DATA(g11040));
  MSFF DFF_207(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g374),.DATA(g11440));
  MSFF DFF_208(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g563),.DATA(g11050));
  MSFF DFF_209(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1914),.DATA(g8284));
  MSFF DFF_210(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g530),.DATA(g11328));
  MSFF DFF_211(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g575),.DATA(g11052));
  MSFF DFF_212(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1936),.DATA(g9355));
  MSFF DFF_213(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g55),.DATA(g7778));
  MSFF DFF_214(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1117),.DATA(g6299));
  MSFF DFF_215(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1317),.DATA(g1356));
  MSFF DFF_216(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g357),.DATA(g11509));
  MSFF DFF_217(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g386),.DATA(g11263));
  MSFF DFF_218(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1601),.DATA(g7363));
  MSFF DFF_219(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g553),.DATA(g11046));
  MSFF DFF_220(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g166),.DATA(g7747));
  MSFF DFF_221(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g501),.DATA(g11334));
  MSFF DFF_222(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g262),.DATA(g7758));
  MSFF DFF_223(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1840),.DATA(g8694));
  MSFF DFF_224(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g70),.DATA(g7783));
  MSFF DFF_225(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g318),.DATA(g5646));
  MSFF DFF_226(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1356),.DATA(g6818));
  MSFF DFF_227(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g794),.DATA(g6800));
  MSFF DFF_228(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g36),.DATA(g10870));
  MSFF DFF_229(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g302),.DATA(g7773));
  MSFF DFF_230(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g342),.DATA(g11513));
  MSFF DFF_231(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1250),.DATA(g7299));
  MSFF DFF_232(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1163),.DATA(g6301));
  MSFF DFF_233(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1810),.DATA(g2044));
  MSFF DFF_234(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1032),.DATA(g7800));
  MSFF DFF_235(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1432),.DATA(g8990));
  MSFF DFF_236(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1053),.DATA(g7792));
  MSFF DFF_237(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1453),.DATA(g7326));
  MSFF DFF_238(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g363),.DATA(g11511));
  MSFF DFF_239(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g330),.DATA(g5650));
  MSFF DFF_240(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1157),.DATA(g6303));
  MSFF DFF_241(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1357),.DATA(g6330));
  MSFF DFF_242(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g35),.DATA(g10869));
  MSFF DFF_243(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g928),.DATA(g8569));
  MSFF DFF_244(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g261),.DATA(g7757));
  MSFF DFF_245(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g516),.DATA(g11337));
  MSFF DFF_246(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g254),.DATA(g7759));
  MSFF DFF_247(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g778),.DATA(g8076));
  MSFF DFF_248(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g861),.DATA(g4190));
  MSFF DFF_249(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1627),.DATA(g8871));
  MSFF DFF_250(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1292),.DATA(g7293));
  MSFF DFF_251(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g290),.DATA(g7769));
  MSFF DFF_252(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1850),.DATA(g5671));
  MSFF DFF_253(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g770),.DATA(g7288));
  MSFF DFF_254(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1583),.DATA(g7357));
  MSFF DFF_255(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g466),.DATA(g11468));
  MSFF DFF_256(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1561),.DATA(g7350));
  MSFF DFF_257(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1527),.DATA(g4899));
  MSFF DFF_258(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1546),.DATA(g7345));
  MSFF DFF_259(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g287),.DATA(g7768));
  MSFF DFF_260(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g560),.DATA(g11049));
  MSFF DFF_261(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g617),.DATA(g8780));
  MSFF DFF_262(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g17),.DATA(g4894));
  MSFF DFF_263(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g336),.DATA(g11653));
  MSFF DFF_264(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g456),.DATA(g11466));
  MSFF DFF_265(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g305),.DATA(g5643));
  MSFF DFF_266(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g345),.DATA(g11642));
  MSFF DFF_267(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g8),.DATA(g2613));
  MSFF DFF_268(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1771),.DATA(g7811));
  MSFF DFF_269(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g865),.DATA(g8275));
  MSFF DFF_270(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g255),.DATA(g7751));
  MSFF DFF_271(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1945),.DATA(g9356));
  MSFF DFF_272(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1738),.DATA(g5661));
  MSFF DFF_273(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1478),.DATA(g8442));
  MSFF DFF_274(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1035),.DATA(g7787));
  MSFF DFF_275(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1959),.DATA(g4217));
  MSFF DFF_276(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1690),.DATA(g6844));
  MSFF DFF_277(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1482),.DATA(g8443));
  MSFF DFF_278(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1110),.DATA(g6817));
  MSFF DFF_279(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g296),.DATA(g7771));
  MSFF DFF_280(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1663),.DATA(g11034));
  MSFF DFF_281(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g700),.DATA(g8431));
  MSFF DFF_282(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1762),.DATA(g5669));
  MSFF DFF_283(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g360),.DATA(g11510));
  MSFF DFF_284(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g192),.DATA(g6837));
  MSFF DFF_285(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1657),.DATA(g10875));
  MSFF DFF_286(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g722),.DATA(g9346));
  MSFF DFF_287(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g61),.DATA(g7780));
  MSFF DFF_288(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g566),.DATA(g11051));
  MSFF DFF_289(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1394),.DATA(g7809));
  MSFF DFF_290(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1089),.DATA(g6809));
  MSFF DFF_291(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g883),.DATA(g4897));
  MSFF DFF_292(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1071),.DATA(g6804));
  MSFF DFF_293(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g986),.DATA(g11473));
  MSFF DFF_294(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g971),.DATA(g11470));
  MSFF DFF_295(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1955),.DATA(g6338));
  MSFF DFF_296(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g143),.DATA(g7746));
  MSFF DFF_297(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1814),.DATA(g9825));
  MSFF DFF_298(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1038),.DATA(g7797));
  MSFF DFF_299(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1212),.DATA(g1217));
  MSFF DFF_300(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1918),.DATA(g9353));
  MSFF DFF_301(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g782),.DATA(g8273));
  MSFF DFF_302(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1822),.DATA(g9826));
  MSFF DFF_303(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g237),.DATA(g7306));
  MSFF DFF_304(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g746),.DATA(g2638));
  MSFF DFF_305(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1062),.DATA(g7795));
  MSFF DFF_306(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1462),.DATA(g8438));
  MSFF DFF_307(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g178),.DATA(g7748));
  MSFF DFF_308(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g366),.DATA(g11512));
  MSFF DFF_309(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g837),.DATA(g4184));
  MSFF DFF_310(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g599),.DATA(g9819));
  MSFF DFF_311(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1854),.DATA(g11408));
  MSFF DFF_312(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g944),.DATA(g11398));
  MSFF DFF_313(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1941),.DATA(g8287));
  MSFF DFF_314(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g170),.DATA(g8422));
  MSFF DFF_315(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1520),.DATA(g7334));
  MSFF DFF_316(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g686),.DATA(g9342));
  MSFF DFF_317(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g953),.DATA(g11401));
  MSFF DFF_318(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1958),.DATA(g6339));
  MSFF DFF_319(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g40),.DATA(g10775));
  MSFF DFF_320(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1765),.DATA(g3329));
  MSFF DFF_321(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1733),.DATA(g10882));
  MSFF DFF_322(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1270),.DATA(g7303));
  MSFF DFF_323(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1610),.DATA(g6845));
  MSFF DFF_324(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1796),.DATA(g8280));
  MSFF DFF_325(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1324),.DATA(g11632));
  MSFF DFF_326(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1540),.DATA(g7343));
  MSFF DFF_327(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1377),.DATA(g7312));
  MSFF DFF_328(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1206),.DATA(g4898));
  MSFF DFF_329(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g491),.DATA(g11332));
  MSFF DFF_330(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1849),.DATA(g5670));
  MSFF DFF_331(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g213),.DATA(g7313));
  MSFF DFF_332(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1781),.DATA(g7813));
  MSFF DFF_333(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1900),.DATA(g9351));
  MSFF DFF_334(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1245),.DATA(g7298));
  MSFF DFF_335(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g108),.DATA(g11593));
  MSFF DFF_336(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g630),.DATA(g7287));
  MSFF DFF_337(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g148),.DATA(g8427));
  MSFF DFF_338(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g833),.DATA(g4183));
  MSFF DFF_339(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1923),.DATA(g8285));
  MSFF DFF_340(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g936),.DATA(g8571));
  MSFF DFF_341(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1215),.DATA(g6315));
  MSFF DFF_342(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1314),.DATA(g11629));
  MSFF DFF_343(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g849),.DATA(g4187));
  MSFF DFF_344(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1336),.DATA(g11654));
  MSFF DFF_345(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g272),.DATA(g7763));
  MSFF DFF_346(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1806),.DATA(g8573));
  MSFF DFF_347(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g826),.DATA(g8568));
  MSFF DFF_348(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1065),.DATA(g7796));
  MSFF DFF_349(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1887),.DATA(g8281));
  MSFF DFF_350(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g37),.DATA(g10871));
  MSFF DFF_351(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g968),.DATA(g11406));
  MSFF DFF_352(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1845),.DATA(g5673));
  MSFF DFF_353(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1137),.DATA(g6310));
  MSFF DFF_354(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1891),.DATA(g9350));
  MSFF DFF_355(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1255),.DATA(g7300));
  MSFF DFF_356(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g257),.DATA(g7753));
  MSFF DFF_357(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g874),.DATA(g9821));
  MSFF DFF_358(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g591),.DATA(g9818));
  MSFF DFF_359(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g731),.DATA(g9347));
  MSFF DFF_360(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g636),.DATA(g8781));
  MSFF DFF_361(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1218),.DATA(g8276));
  MSFF DFF_362(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g605),.DATA(g9820));
  MSFF DFF_363(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g79),.DATA(g7776));
  MSFF DFF_364(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g182),.DATA(g7749));
  MSFF DFF_365(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g950),.DATA(g11400));
  MSFF DFF_366(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1129),.DATA(g6308));
  MSFF DFF_367(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g857),.DATA(g4189));
  MSFF DFF_368(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g448),.DATA(g11258));
  MSFF DFF_369(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1828),.DATA(g9827));
  MSFF DFF_370(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1727),.DATA(g10880));
  MSFF DFF_371(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1592),.DATA(g7360));
  MSFF DFF_372(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1703),.DATA(g6843));
  MSFF DFF_373(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1932),.DATA(g8286));
  MSFF DFF_374(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1624),.DATA(g8870));
  MSFF DFF_375(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g26),.DATA(g4885));
  MSFF DFF_376(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1068),.DATA(g6803));
  MSFF DFF_377(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g578),.DATA(g6286));
  MSFF DFF_378(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g440),.DATA(g11260));
  MSFF DFF_379(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g476),.DATA(g11338));
  MSFF DFF_380(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g119),.DATA(g7745));
  MSFF DFF_381(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g668),.DATA(g9340));
  MSFF DFF_382(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g139),.DATA(g8418));
  MSFF DFF_383(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1149),.DATA(g6305));
  MSFF DFF_384(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g34),.DATA(g10868));
  MSFF DFF_385(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1848),.DATA(g7366));
  MSFF DFF_386(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g263),.DATA(g7760));
  MSFF DFF_387(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g818),.DATA(g8274));
  MSFF DFF_388(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1747),.DATA(g5664));
  MSFF DFF_389(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g802),.DATA(g6802));
  MSFF DFF_390(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g275),.DATA(g7764));
  MSFF DFF_391(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1524),.DATA(g7338));
  MSFF DFF_392(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1577),.DATA(g7355));
  MSFF DFF_393(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g810),.DATA(g7786));
  MSFF DFF_394(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g391),.DATA(g11264));
  MSFF DFF_395(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g658),.DATA(g9339));
  MSFF DFF_396(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1386),.DATA(g7318));
  MSFF DFF_397(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g253),.DATA(g7750));
  MSFF DFF_398(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g875),.DATA(g9822));
  MSFF DFF_399(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1125),.DATA(g6307));
  MSFF DFF_400(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g201),.DATA(g7304));
  MSFF DFF_401(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1280),.DATA(g7295));
  MSFF DFF_402(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1083),.DATA(g6807));
  MSFF DFF_403(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g650),.DATA(g8066));
  MSFF DFF_404(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1636),.DATA(g8874));
  MSFF DFF_405(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g853),.DATA(g4188));
  MSFF DFF_406(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g421),.DATA(g11270));
  MSFF DFF_407(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g762),.DATA(g6798));
  MSFF DFF_408(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g956),.DATA(g11402));
  MSFF DFF_409(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g378),.DATA(g11441));
  MSFF DFF_410(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1756),.DATA(g5667));
  MSFF DFF_411(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g589),.DATA(g6297));
  MSFF DFF_412(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g841),.DATA(g4185));
  MSFF DFF_413(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1027),.DATA(g7798));
  MSFF DFF_414(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1003),.DATA(g7803));
  MSFF DFF_415(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1403),.DATA(g8991));
  MSFF DFF_416(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1145),.DATA(g6312));
  MSFF DFF_417(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1107),.DATA(g6816));
  MSFF DFF_418(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1223),.DATA(g8277));
  MSFF DFF_419(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g406),.DATA(g11267));
  MSFF DFF_420(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1811),.DATA(g11185));
  MSFF DFF_421(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1642),.DATA(g11183));
  MSFF DFF_422(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1047),.DATA(g7790));
  MSFF DFF_423(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1654),.DATA(g10874));
  MSFF DFF_424(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g197),.DATA(g6835));
  MSFF DFF_425(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1595),.DATA(g7361));
  MSFF DFF_426(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1537),.DATA(g7342));
  MSFF DFF_427(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g727),.DATA(g8434));
  MSFF DFF_428(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g999),.DATA(g7804));
  MSFF DFF_429(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g798),.DATA(g6801));
  MSFF DFF_430(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g481),.DATA(g11324));
  MSFF DFF_431(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g754),.DATA(g4895));
  MSFF DFF_432(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1330),.DATA(g11634));
  MSFF DFF_433(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g845),.DATA(g4186));
  MSFF DFF_434(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g790),.DATA(g8567));
  MSFF DFF_435(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1512),.DATA(g8449));
  MSFF DFF_436(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g114),.DATA(g113));
  MSFF DFF_437(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1490),.DATA(g8445));
  MSFF DFF_438(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1166),.DATA(g6300));
  MSFF DFF_439(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1056),.DATA(g7793));
  MSFF DFF_440(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g348),.DATA(g11506));
  MSFF DFF_441(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g868),.DATA(g874));
  MSFF DFF_442(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1260),.DATA(g7301));
  MSFF DFF_443(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g260),.DATA(g7756));
  MSFF DFF_444(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g131),.DATA(g8420));
  MSFF DFF_445(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g7),.DATA(g2731));
  MSFF DFF_446(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g258),.DATA(g7754));
  MSFF DFF_447(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g521),.DATA(g11330));
  MSFF DFF_448(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1318),.DATA(g11630));
  MSFF DFF_449(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1872),.DATA(g9348));
  MSFF DFF_450(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g677),.DATA(g9341));
  MSFF DFF_451(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g582),.DATA(g6290));
  MSFF DFF_452(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1393),.DATA(g7320));
  MSFF DFF_453(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1549),.DATA(g7346));
  MSFF DFF_454(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g947),.DATA(g11399));
  MSFF DFF_455(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1834),.DATA(g9895));
  MSFF DFF_456(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1598),.DATA(g7362));
  MSFF DFF_457(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1121),.DATA(g6306));
  MSFF DFF_458(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1321),.DATA(g11631));
  MSFF DFF_459(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g506),.DATA(g11335));
  MSFF DFF_460(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g546),.DATA(g11043));
  MSFF DFF_461(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1909),.DATA(g9352));
  MSFF DFF_462(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g755),.DATA(g6298));
  MSFF DFF_463(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1552),.DATA(g7347));
  MSFF DFF_464(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g584),.DATA(g6292));
  MSFF DFF_465(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1687),.DATA(g11042));
  MSFF DFF_466(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1586),.DATA(g7358));
  MSFF DFF_467(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g324),.DATA(g5648));
  MSFF DFF_468(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1141),.DATA(g6311));
  MSFF DFF_469(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1570),.DATA(g4900));
  MSFF DFF_470(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1341),.DATA(g11655));
  MSFF DFF_471(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1710),.DATA(g4901));
  MSFF DFF_472(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1645),.DATA(g11184));
  MSFF DFF_473(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g115),.DATA(g7321));
  MSFF DFF_474(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g135),.DATA(g8419));
  MSFF DFF_475(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g525),.DATA(g11329));
  MSFF DFF_476(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g581),.DATA(g6289));
  MSFF DFF_477(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1607),.DATA(g7365));
  MSFF DFF_478(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g321),.DATA(g5647));
  MSFF DFF_479(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g67),.DATA(g7782));
  MSFF DFF_480(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1275),.DATA(g11443));
  MSFF DFF_481(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1311),.DATA(g11628));
  MSFF DFF_482(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1615),.DATA(g8868));
  MSFF DFF_483(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g382),.DATA(g11442));
  MSFF DFF_484(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1374),.DATA(g6825));
  MSFF DFF_485(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g266),.DATA(g7761));
  MSFF DFF_486(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1284),.DATA(g7294));
  MSFF DFF_487(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1380),.DATA(g7314));
  MSFF DFF_488(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g673),.DATA(g8428));
  MSFF DFF_489(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1853),.DATA(g5672));
  MSFF DFF_490(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g162),.DATA(g8424));
  MSFF DFF_491(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g411),.DATA(g11268));
  MSFF DFF_492(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g431),.DATA(g11262));
  MSFF DFF_493(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1905),.DATA(g8283));
  MSFF DFF_494(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1515),.DATA(g7333));
  MSFF DFF_495(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1630),.DATA(g8872));
  MSFF DFF_496(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g49),.DATA(g7774));
  MSFF DFF_497(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g991),.DATA(g7802));
  MSFF DFF_498(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1300),.DATA(g7291));
  MSFF DFF_499(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g339),.DATA(g11505));
  MSFF DFF_500(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g256),.DATA(g7752));
  MSFF DFF_501(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1750),.DATA(g5665));
  MSFF DFF_502(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g585),.DATA(g6293));
  MSFF DFF_503(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1440),.DATA(g8988));
  MSFF DFF_504(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1666),.DATA(g11035));
  MSFF DFF_505(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1528),.DATA(g7339));
  MSFF DFF_506(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1351),.DATA(g11657));
  MSFF DFF_507(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1648),.DATA(g11181));
  MSFF DFF_508(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g127),.DATA(g8421));
  MSFF DFF_509(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1618),.DATA(g11611));
  MSFF DFF_510(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1235),.DATA(g7296));
  MSFF DFF_511(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g299),.DATA(g7772));
  MSFF DFF_512(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g435),.DATA(g11261));
  MSFF DFF_513(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g64),.DATA(g7781));
  MSFF DFF_514(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1555),.DATA(g7348));
  MSFF DFF_515(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g995),.DATA(g7801));
  MSFF DFF_516(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1621),.DATA(g8869));
  MSFF DFF_517(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1113),.DATA(g6313));
  MSFF DFF_518(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g643),.DATA(g8064));
  MSFF DFF_519(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1494),.DATA(g8446));
  MSFF DFF_520(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1567),.DATA(g7352));
  MSFF DFF_521(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g691),.DATA(g8430));
  MSFF DFF_522(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g534),.DATA(g11327));
  MSFF DFF_523(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1776),.DATA(g7812));
  MSFF DFF_524(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g569),.DATA(g10876));
  MSFF DFF_525(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1160),.DATA(g6302));
  MSFF DFF_526(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1360),.DATA(g9824));
  MSFF DFF_527(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1050),.DATA(g7791));
  MSFF DFF_528(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1),.DATA(g8078));
  MSFF DFF_529(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g511),.DATA(g11336));
  MSFF DFF_530(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1724),.DATA(g10879));
  MSFF DFF_531(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g12),.DATA(g7337));
  MSFF DFF_532(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g1878),.DATA(g8695));
  MSFF DFF_533(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(g73),.DATA(g7784));
//
  NOT NOT1_0(.VSS(VSS),.VDD(VDD),.Y(I8854),.A(g4500));
  NOT NOT1_1(.VSS(VSS),.VDD(VDD),.Y(g5652),.A(I9117));
  NOT NOT1_2(.VSS(VSS),.VDD(VDD),.Y(I12913),.A(g7845));
  NOT NOT1_3(.VSS(VSS),.VDD(VDD),.Y(g11354),.A(I17179));
  NOT NOT1_4(.VSS(VSS),.VDD(VDD),.Y(g6837),.A(I10891));
  NOT NOT1_5(.VSS(VSS),.VDD(VDD),.Y(I10941),.A(g6555));
  NOT NOT1_6(.VSS(VSS),.VDD(VDD),.Y(I6979),.A(g2888));
  NOT NOT1_7(.VSS(VSS),.VDD(VDD),.Y(g5843),.A(I9458));
  NOT NOT1_8(.VSS(VSS),.VDD(VDD),.Y(g2771),.A(I5854));
  NOT NOT1_9(.VSS(VSS),.VDD(VDD),.Y(g3537),.A(g3164));
  NOT NOT1_10(.VSS(VSS),.VDD(VDD),.Y(g6062),.A(I9699));
  NOT NOT1_11(.VSS(VSS),.VDD(VDD),.Y(I9984),.A(g5529));
  NOT NOT1_12(.VSS(VSS),.VDD(VDD),.Y(I14382),.A(g8886));
  NOT NOT1_13(.VSS(VSS),.VDD(VDD),.Y(g7706),.A(I12335));
  NOT NOT1_14(.VSS(VSS),.VDD(VDD),.Y(I13618),.A(g8345));
  NOT NOT1_15(.VSS(VSS),.VDD(VDD),.Y(I15181),.A(g9968));
  NOT NOT1_16(.VSS(VSS),.VDD(VDD),.Y(g6620),.A(I10573));
  NOT NOT1_17(.VSS(VSS),.VDD(VDD),.Y(I12436),.A(g7659));
  NOT NOT1_18(.VSS(VSS),.VDD(VDD),.Y(g5193),.A(g4682));
  NOT NOT1_19(.VSS(VSS),.VDD(VDD),.Y(g6462),.A(I10394));
  NOT NOT1_20(.VSS(VSS),.VDD(VDD),.Y(g8925),.A(I14252));
  NOT NOT1_21(.VSS(VSS),.VDD(VDD),.Y(I14519),.A(g9106));
  NOT NOT1_22(.VSS(VSS),.VDD(VDD),.Y(g10289),.A(I15691));
  NOT NOT1_23(.VSS(VSS),.VDD(VDD),.Y(I14176),.A(g8784));
  NOT NOT1_24(.VSS(VSS),.VDD(VDD),.Y(I14185),.A(g8790));
  NOT NOT1_25(.VSS(VSS),.VDD(VDD),.Y(g11181),.A(I16944));
  NOT NOT1_26(.VSS(VSS),.VDD(VDD),.Y(I14675),.A(g9263));
  NOT NOT1_27(.VSS(VSS),.VDD(VDD),.Y(g2299),.A(g1707));
  NOT NOT1_28(.VSS(VSS),.VDD(VDD),.Y(I12607),.A(g7633));
  NOT NOT1_29(.VSS(VSS),.VDD(VDD),.Y(g3272),.A(g2450));
  NOT NOT1_30(.VSS(VSS),.VDD(VDD),.Y(g2547),.A(g23));
  NOT NOT1_31(.VSS(VSS),.VDD(VDD),.Y(g9291),.A(g8892));
  NOT NOT1_32(.VSS(VSS),.VDD(VDD),.Y(I6001),.A(g2548));
  NOT NOT1_33(.VSS(VSS),.VDD(VDD),.Y(I7048),.A(g2807));
  NOT NOT1_34(.VSS(VSS),.VDD(VDD),.Y(g10309),.A(I15733));
  NOT NOT1_35(.VSS(VSS),.VDD(VDD),.Y(g7029),.A(I11180));
  NOT NOT1_36(.VSS(VSS),.VDD(VDD),.Y(g4440),.A(g4130));
  NOT NOT1_37(.VSS(VSS),.VDD(VDD),.Y(I9544),.A(g5024));
  NOT NOT1_38(.VSS(VSS),.VDD(VDD),.Y(g10288),.A(I15688));
  NOT NOT1_39(.VSS(VSS),.VDD(VDD),.Y(I12274),.A(g7110));
  NOT NOT1_40(.VSS(VSS),.VDD(VDD),.Y(I9483),.A(g5050));
  NOT NOT1_41(.VSS(VSS),.VDD(VDD),.Y(g7787),.A(I12526));
  NOT NOT1_42(.VSS(VSS),.VDD(VDD),.Y(I6676),.A(g2759));
  NOT NOT1_43(.VSS(VSS),.VDD(VDD),.Y(I8520),.A(g4338));
  NOT NOT1_44(.VSS(VSS),.VDD(VDD),.Y(g10571),.A(I16236));
  NOT NOT1_45(.VSS(VSS),.VDD(VDD),.Y(I17692),.A(g11596));
  NOT NOT1_46(.VSS(VSS),.VDD(VDD),.Y(I17761),.A(g11652));
  NOT NOT1_47(.VSS(VSS),.VDD(VDD),.Y(I13469),.A(g8147));
  NOT NOT1_48(.VSS(VSS),.VDD(VDD),.Y(g9344),.A(I14537));
  NOT NOT1_49(.VSS(VSS),.VDD(VDD),.Y(g7956),.A(g7432));
  NOT NOT1_50(.VSS(VSS),.VDD(VDD),.Y(g3417),.A(I6624));
  NOT NOT1_51(.VSS(VSS),.VDD(VDD),.Y(g4323),.A(g4130));
  NOT NOT1_52(.VSS(VSS),.VDD(VDD),.Y(I11286),.A(g6551));
  NOT NOT1_53(.VSS(VSS),.VDD(VDD),.Y(I8031),.A(g3540));
  NOT NOT1_54(.VSS(VSS),.VDD(VDD),.Y(g7675),.A(I12300));
  NOT NOT1_55(.VSS(VSS),.VDD(VDD),.Y(g8320),.A(I13344));
  NOT NOT1_56(.VSS(VSS),.VDD(VDD),.Y(I12565),.A(g7388));
  NOT NOT1_57(.VSS(VSS),.VDD(VDD),.Y(I16644),.A(g10865));
  NOT NOT1_58(.VSS(VSS),.VDD(VDD),.Y(I11306),.A(g6731));
  NOT NOT1_59(.VSS(VSS),.VDD(VDD),.Y(g1981),.A(g650));
  NOT NOT1_60(.VSS(VSS),.VDD(VDD),.Y(I7333),.A(g3729));
  NOT NOT1_61(.VSS(VSS),.VDD(VDD),.Y(I13039),.A(g8054));
  NOT NOT1_62(.VSS(VSS),.VDD(VDD),.Y(g3982),.A(g3052));
  NOT NOT1_63(.VSS(VSS),.VDD(VDD),.Y(g6249),.A(I10006));
  NOT NOT1_64(.VSS(VSS),.VDD(VDD),.Y(g9259),.A(g8892));
  NOT NOT1_65(.VSS(VSS),.VDD(VDD),.Y(I15190),.A(g9974));
  NOT NOT1_66(.VSS(VSS),.VDD(VDD),.Y(g11426),.A(I17331));
  NOT NOT1_67(.VSS(VSS),.VDD(VDD),.Y(g9819),.A(I14958));
  NOT NOT1_68(.VSS(VSS),.VDD(VDD),.Y(g8277),.A(I13203));
  NOT NOT1_69(.VSS(VSS),.VDD(VDD),.Y(I5050),.A(g1216));
  NOT NOT1_70(.VSS(VSS),.VDD(VDD),.Y(I5641),.A(g546));
  NOT NOT1_71(.VSS(VSS),.VDD(VDD),.Y(g5121),.A(g4682));
  NOT NOT1_72(.VSS(VSS),.VDD(VDD),.Y(g1997),.A(g798));
  NOT NOT1_73(.VSS(VSS),.VDD(VDD),.Y(g3629),.A(g3228));
  NOT NOT1_74(.VSS(VSS),.VDD(VDD),.Y(g3328),.A(I6501));
  NOT NOT1_75(.VSS(VSS),.VDD(VDD),.Y(I12641),.A(g7709));
  NOT NOT1_76(.VSS(VSS),.VDD(VDD),.Y(g5670),.A(I9171));
  NOT NOT1_77(.VSS(VSS),.VDD(VDD),.Y(g6842),.A(I10898));
  NOT NOT1_78(.VSS(VSS),.VDD(VDD),.Y(g8617),.A(g8465));
  NOT NOT1_79(.VSS(VSS),.VDD(VDD),.Y(I15520),.A(g10035));
  NOT NOT1_80(.VSS(VSS),.VDD(VDD),.Y(I7396),.A(g4102));
  NOT NOT1_81(.VSS(VSS),.VDD(VDD),.Y(I7803),.A(g3820));
  NOT NOT1_82(.VSS(VSS),.VDD(VDD),.Y(g3330),.A(I6507));
  NOT NOT1_83(.VSS(VSS),.VDD(VDD),.Y(g2991),.A(I6233));
  NOT NOT1_84(.VSS(VSS),.VDD(VDD),.Y(I9461),.A(g4940));
  NOT NOT1_85(.VSS(VSS),.VDD(VDD),.Y(g2244),.A(I5251));
  NOT NOT1_86(.VSS(VSS),.VDD(VDD),.Y(g6192),.A(I9923));
  NOT NOT1_87(.VSS(VSS),.VDD(VDD),.Y(g6298),.A(I10153));
  NOT NOT1_88(.VSS(VSS),.VDD(VDD),.Y(g6085),.A(I9734));
  NOT NOT1_89(.VSS(VSS),.VDD(VDD),.Y(I12153),.A(g6874));
  NOT NOT1_90(.VSS(VSS),.VDD(VDD),.Y(g4351),.A(I7630));
  NOT NOT1_91(.VSS(VSS),.VDD(VDD),.Y(I11677),.A(g7056));
  NOT NOT1_92(.VSS(VSS),.VDD(VDD),.Y(g10687),.A(I16356));
  NOT NOT1_93(.VSS(VSS),.VDD(VDD),.Y(g4530),.A(I7935));
  NOT NOT1_94(.VSS(VSS),.VDD(VDD),.Y(g8516),.A(I13717));
  NOT NOT1_95(.VSS(VSS),.VDD(VDD),.Y(g5232),.A(g4640));
  NOT NOT1_96(.VSS(VSS),.VDD(VDD),.Y(I13975),.A(g8588));
  NOT NOT1_97(.VSS(VSS),.VDD(VDD),.Y(g2078),.A(g135));
  NOT NOT1_98(.VSS(VSS),.VDD(VDD),.Y(I8911),.A(g4565));
  NOT NOT1_99(.VSS(VSS),.VDD(VDD),.Y(g2340),.A(g1918));
  NOT NOT1_100(.VSS(VSS),.VDD(VDD),.Y(g7684),.A(g7148));
  NOT NOT1_101(.VSS(VSS),.VDD(VDD),.Y(I12409),.A(g7501));
  NOT NOT1_102(.VSS(VSS),.VDD(VDD),.Y(g7745),.A(I12400));
  NOT NOT1_103(.VSS(VSS),.VDD(VDD),.Y(g8987),.A(I14382));
  NOT NOT1_104(.VSS(VSS),.VDD(VDD),.Y(g11546),.A(g11519));
  NOT NOT1_105(.VSS(VSS),.VDD(VDD),.Y(I10729),.A(g5935));
  NOT NOT1_106(.VSS(VSS),.VDD(VDD),.Y(g5253),.A(g4346));
  NOT NOT1_107(.VSS(VSS),.VDD(VDD),.Y(g7338),.A(I11662));
  NOT NOT1_108(.VSS(VSS),.VDD(VDD),.Y(I7509),.A(g3566));
  NOT NOT1_109(.VSS(VSS),.VDD(VDD),.Y(I9427),.A(g4963));
  NOT NOT1_110(.VSS(VSS),.VDD(VDD),.Y(g3800),.A(g3292));
  NOT NOT1_111(.VSS(VSS),.VDD(VDD),.Y(I15088),.A(g9832));
  NOT NOT1_112(.VSS(VSS),.VDD(VDD),.Y(g2907),.A(I6074));
  NOT NOT1_113(.VSS(VSS),.VDD(VDD),.Y(g7791),.A(I12538));
  NOT NOT1_114(.VSS(VSS),.VDD(VDD),.Y(I11143),.A(g6446));
  NOT NOT1_115(.VSS(VSS),.VDD(VDD),.Y(g6854),.A(I10920));
  NOT NOT1_116(.VSS(VSS),.VDD(VDD),.Y(g11088),.A(I16871));
  NOT NOT1_117(.VSS(VSS),.VDD(VDD),.Y(g7309),.A(I11575));
  NOT NOT1_118(.VSS(VSS),.VDD(VDD),.Y(g8299),.A(I13255));
  NOT NOT1_119(.VSS(VSS),.VDD(VDD),.Y(I9046),.A(g4736));
  NOT NOT1_120(.VSS(VSS),.VDD(VDD),.Y(g6941),.A(g6503));
  NOT NOT1_121(.VSS(VSS),.VDD(VDD),.Y(g2435),.A(g201));
  NOT NOT1_122(.VSS(VSS),.VDD(VDD),.Y(I14439),.A(g8969));
  NOT NOT1_123(.VSS(VSS),.VDD(VDD),.Y(g4010),.A(g3144));
  NOT NOT1_124(.VSS(VSS),.VDD(VDD),.Y(g2082),.A(g1371));
  NOT NOT1_125(.VSS(VSS),.VDD(VDD),.Y(I6932),.A(g2850));
  NOT NOT1_126(.VSS(VSS),.VDD(VDD),.Y(I7662),.A(g3336));
  NOT NOT1_127(.VSS(VSS),.VDD(VDD),.Y(I9446),.A(g5052));
  NOT NOT1_128(.VSS(VSS),.VDD(VDD),.Y(g5519),.A(g4811));
  NOT NOT1_129(.VSS(VSS),.VDD(VDD),.Y(g5740),.A(I9302));
  NOT NOT1_130(.VSS(VSS),.VDD(VDD),.Y(I5289),.A(g49));
  NOT NOT1_131(.VSS(VSS),.VDD(VDD),.Y(I9514),.A(g5094));
  NOT NOT1_132(.VSS(VSS),.VDD(VDD),.Y(g7808),.A(I12589));
  NOT NOT1_133(.VSS(VSS),.VDD(VDD),.Y(g2482),.A(I5565));
  NOT NOT1_134(.VSS(VSS),.VDD(VDD),.Y(I5658),.A(g560));
  NOT NOT1_135(.VSS(VSS),.VDD(VDD),.Y(I15497),.A(g10119));
  NOT NOT1_136(.VSS(VSS),.VDD(VDD),.Y(I6624),.A(g2629));
  NOT NOT1_137(.VSS(VSS),.VDD(VDD),.Y(g8892),.A(I14242));
  NOT NOT1_138(.VSS(VSS),.VDD(VDD),.Y(I11169),.A(g6481));
  NOT NOT1_139(.VSS(VSS),.VDD(VDD),.Y(g3213),.A(I6388));
  NOT NOT1_140(.VSS(VSS),.VDD(VDD),.Y(I6068),.A(g2227));
  NOT NOT1_141(.VSS(VSS),.VDD(VDD),.Y(g11497),.A(I17510));
  NOT NOT1_142(.VSS(VSS),.VDD(VDD),.Y(I13791),.A(g8518));
  NOT NOT1_143(.VSS(VSS),.VDD(VDD),.Y(I16867),.A(g10913));
  NOT NOT1_144(.VSS(VSS),.VDD(VDD),.Y(I10349),.A(g6215));
  NOT NOT1_145(.VSS(VSS),.VDD(VDD),.Y(g10260),.A(g10125));
  NOT NOT1_146(.VSS(VSS),.VDD(VDD),.Y(g7759),.A(I12442));
  NOT NOT1_147(.VSS(VSS),.VDD(VDD),.Y(I8473),.A(g4577));
  NOT NOT1_148(.VSS(VSS),.VDD(VDD),.Y(I14349),.A(g8958));
  NOT NOT1_149(.VSS(VSS),.VDD(VDD),.Y(g6708),.A(I10689));
  NOT NOT1_150(.VSS(VSS),.VDD(VDD),.Y(g10668),.A(g10563));
  NOT NOT1_151(.VSS(VSS),.VDD(VDD),.Y(I5271),.A(g70));
  NOT NOT1_152(.VSS(VSS),.VDD(VDD),.Y(I9191),.A(g5546));
  NOT NOT1_153(.VSS(VSS),.VDD(VDD),.Y(I9391),.A(g5013));
  NOT NOT1_154(.VSS(VSS),.VDD(VDD),.Y(g6219),.A(g5426));
  NOT NOT1_155(.VSS(VSS),.VDD(VDD),.Y(I15250),.A(g9980));
  NOT NOT1_156(.VSS(VSS),.VDD(VDD),.Y(I17100),.A(g11221));
  NOT NOT1_157(.VSS(VSS),.VDD(VDD),.Y(I14906),.A(g9508));
  NOT NOT1_158(.VSS(VSS),.VDD(VDD),.Y(g9825),.A(I14976));
  NOT NOT1_159(.VSS(VSS),.VDD(VDD),.Y(g7201),.A(I11427));
  NOT NOT1_160(.VSS(VSS),.VDD(VDD),.Y(I14083),.A(g8747));
  NOT NOT1_161(.VSS(VSS),.VDD(VDD),.Y(g10195),.A(I15559));
  NOT NOT1_162(.VSS(VSS),.VDD(VDD),.Y(I8324),.A(g4794));
  NOT NOT1_163(.VSS(VSS),.VDD(VDD),.Y(g6031),.A(I9642));
  NOT NOT1_164(.VSS(VSS),.VDD(VDD),.Y(g2915),.A(I6094));
  NOT NOT1_165(.VSS(VSS),.VDD(VDD),.Y(I13666),.A(g8292));
  NOT NOT1_166(.VSS(VSS),.VDD(VDD),.Y(I9695),.A(g5212));
  NOT NOT1_167(.VSS(VSS),.VDD(VDD),.Y(I11363),.A(g6595));
  NOT NOT1_168(.VSS(VSS),.VDD(VDD),.Y(I11217),.A(g6529));
  NOT NOT1_169(.VSS(VSS),.VDD(VDD),.Y(g6431),.A(g6145));
  NOT NOT1_170(.VSS(VSS),.VDD(VDD),.Y(g6252),.A(I10015));
  NOT NOT1_171(.VSS(VSS),.VDD(VDD),.Y(g4172),.A(I7333));
  NOT NOT1_172(.VSS(VSS),.VDD(VDD),.Y(g6812),.A(I10846));
  NOT NOT1_173(.VSS(VSS),.VDD(VDD),.Y(g8991),.A(I14394));
  NOT NOT1_174(.VSS(VSS),.VDD(VDD),.Y(g4372),.A(I7677));
  NOT NOT1_175(.VSS(VSS),.VDD(VDD),.Y(g7049),.A(I11228));
  NOT NOT1_176(.VSS(VSS),.VDD(VDD),.Y(I6576),.A(g2617));
  NOT NOT1_177(.VSS(VSS),.VDD(VDD),.Y(g10525),.A(g10499));
  NOT NOT1_178(.VSS(VSS),.VDD(VDD),.Y(g10488),.A(I16101));
  NOT NOT1_179(.VSS(VSS),.VDD(VDD),.Y(I10566),.A(g5904));
  NOT NOT1_180(.VSS(VSS),.VDD(VDD),.Y(I13478),.A(g8191));
  NOT NOT1_181(.VSS(VSS),.VDD(VDD),.Y(g5586),.A(I8996));
  NOT NOT1_182(.VSS(VSS),.VDD(VDD),.Y(g8709),.A(g8674));
  NOT NOT1_183(.VSS(VSS),.VDD(VDD),.Y(g2214),.A(g115));
  NOT NOT1_184(.VSS(VSS),.VDD(VDD),.Y(I9536),.A(g5008));
  NOT NOT1_185(.VSS(VSS),.VDD(VDD),.Y(g6176),.A(I9905));
  NOT NOT1_186(.VSS(VSS),.VDD(VDD),.Y(g4618),.A(g3829));
  NOT NOT1_187(.VSS(VSS),.VDD(VDD),.Y(I15296),.A(g9995));
  NOT NOT1_188(.VSS(VSS),.VDD(VDD),.Y(g4143),.A(I7291));
  NOT NOT1_189(.VSS(VSS),.VDD(VDD),.Y(I7381),.A(g4078));
  NOT NOT1_190(.VSS(VSS),.VDD(VDD),.Y(I9159),.A(g5033));
  NOT NOT1_191(.VSS(VSS),.VDD(VDD),.Y(g11339),.A(I17142));
  NOT NOT1_192(.VSS(VSS),.VDD(VDD),.Y(g8140),.A(I13017));
  NOT NOT1_193(.VSS(VSS),.VDD(VDD),.Y(I16979),.A(g11088));
  NOT NOT1_194(.VSS(VSS),.VDD(VDD),.Y(I16496),.A(g10707));
  NOT NOT1_195(.VSS(VSS),.VDD(VDD),.Y(g8078),.A(I12936));
  NOT NOT1_196(.VSS(VSS),.VDD(VDD),.Y(I7847),.A(g3435));
  NOT NOT1_197(.VSS(VSS),.VDD(VDD),.Y(I9359),.A(g5576));
  NOT NOT1_198(.VSS(VSS),.VDD(VDD),.Y(g8340),.A(I13400));
  NOT NOT1_199(.VSS(VSS),.VDD(VDD),.Y(g2110),.A(I5002));
  NOT NOT1_200(.VSS(VSS),.VDD(VDD),.Y(I15338),.A(g10013));
  NOT NOT1_201(.VSS(VSS),.VDD(VDD),.Y(g6405),.A(g6133));
  NOT NOT1_202(.VSS(VSS),.VDD(VDD),.Y(g8478),.A(I13678));
  NOT NOT1_203(.VSS(VSS),.VDD(VDD),.Y(I16111),.A(g10385));
  NOT NOT1_204(.VSS(VSS),.VDD(VDD),.Y(g4282),.A(g4013));
  NOT NOT1_205(.VSS(VSS),.VDD(VDD),.Y(g11644),.A(I17736));
  NOT NOT1_206(.VSS(VSS),.VDD(VDD),.Y(g7604),.A(I12162));
  NOT NOT1_207(.VSS(VSS),.VDD(VDD),.Y(g9768),.A(g9432));
  NOT NOT1_208(.VSS(VSS),.VDD(VDD),.Y(g4566),.A(g3753));
  NOT NOT1_209(.VSS(VSS),.VDD(VDD),.Y(g7098),.A(I11333));
  NOT NOT1_210(.VSS(VSS),.VDD(VDD),.Y(g10893),.A(I16641));
  NOT NOT1_211(.VSS(VSS),.VDD(VDD),.Y(I4961),.A(g254));
  NOT NOT1_212(.VSS(VSS),.VDD(VDD),.Y(g4988),.A(I8358));
  NOT NOT1_213(.VSS(VSS),.VDD(VDD),.Y(g6286),.A(I10117));
  NOT NOT1_214(.VSS(VSS),.VDD(VDD),.Y(g8959),.A(I14326));
  NOT NOT1_215(.VSS(VSS),.VDD(VDD),.Y(I13580),.A(g8338));
  NOT NOT1_216(.VSS(VSS),.VDD(VDD),.Y(I9016),.A(g4722));
  NOT NOT1_217(.VSS(VSS),.VDD(VDD),.Y(I6398),.A(g2335));
  NOT NOT1_218(.VSS(VSS),.VDD(VDD),.Y(g8517),.A(I13720));
  NOT NOT1_219(.VSS(VSS),.VDD(VDD),.Y(g3348),.A(g2733));
  NOT NOT1_220(.VSS(VSS),.VDD(VDD),.Y(I15060),.A(g9696));
  NOT NOT1_221(.VSS(VSS),.VDD(VDD),.Y(I15968),.A(g10408));
  NOT NOT1_222(.VSS(VSS),.VDD(VDD),.Y(I5332),.A(g756));
  NOT NOT1_223(.VSS(VSS),.VDD(VDD),.Y(g8482),.A(g8329));
  NOT NOT1_224(.VSS(VSS),.VDD(VDD),.Y(g2002),.A(g818));
  NOT NOT1_225(.VSS(VSS),.VDD(VDD),.Y(I10138),.A(g5677));
  NOT NOT1_226(.VSS(VSS),.VDD(VDD),.Y(g11060),.A(g10937));
  NOT NOT1_227(.VSS(VSS),.VDD(VDD),.Y(I17407),.A(g11417));
  NOT NOT1_228(.VSS(VSS),.VDD(VDD),.Y(I12303),.A(g7242));
  NOT NOT1_229(.VSS(VSS),.VDD(VDD),.Y(g5645),.A(I9096));
  NOT NOT1_230(.VSS(VSS),.VDD(VDD),.Y(I15855),.A(g10336));
  NOT NOT1_231(.VSS(VSS),.VDD(VDD),.Y(g2824),.A(I5932));
  NOT NOT1_232(.VSS(VSS),.VDD(VDD),.Y(g11197),.A(g11112));
  NOT NOT1_233(.VSS(VSS),.VDD(VDD),.Y(g4555),.A(I7964));
  NOT NOT1_234(.VSS(VSS),.VDD(VDD),.Y(g5691),.A(g5236));
  NOT NOT1_235(.VSS(VSS),.VDD(VDD),.Y(I9642),.A(g5229));
  NOT NOT1_236(.VSS(VSS),.VDD(VDD),.Y(g7539),.A(I11953));
  NOT NOT1_237(.VSS(VSS),.VDD(VDD),.Y(g7896),.A(I12678));
  NOT NOT1_238(.VSS(VSS),.VDD(VDD),.Y(g8656),.A(I13941));
  NOT NOT1_239(.VSS(VSS),.VDD(VDD),.Y(g9887),.A(I15068));
  NOT NOT1_240(.VSS(VSS),.VDD(VDD),.Y(I8199),.A(g4013));
  NOT NOT1_241(.VSS(VSS),.VDD(VDD),.Y(g6974),.A(g6365));
  NOT NOT1_242(.VSS(VSS),.VDD(VDD),.Y(g6270),.A(I10069));
  NOT NOT1_243(.VSS(VSS),.VDD(VDD),.Y(I14415),.A(g8940));
  NOT NOT1_244(.VSS(VSS),.VDD(VDD),.Y(g3260),.A(I6428));
  NOT NOT1_245(.VSS(VSS),.VDD(VDD),.Y(g11411),.A(I17274));
  NOT NOT1_246(.VSS(VSS),.VDD(VDD),.Y(I10852),.A(g6751));
  NOT NOT1_247(.VSS(VSS),.VDD(VDD),.Y(g10042),.A(I15253));
  NOT NOT1_248(.VSS(VSS),.VDD(VDD),.Y(g10255),.A(g10139));
  NOT NOT1_249(.VSS(VSS),.VDD(VDD),.Y(g6073),.A(I9712));
  NOT NOT1_250(.VSS(VSS),.VDD(VDD),.Y(g10189),.A(I15545));
  NOT NOT1_251(.VSS(VSS),.VDD(VDD),.Y(I4903),.A(g259));
  NOT NOT1_252(.VSS(VSS),.VDD(VDD),.Y(g2877),.A(I6025));
  NOT NOT1_253(.VSS(VSS),.VDD(VDD),.Y(I11531),.A(g7126));
  NOT NOT1_254(.VSS(VSS),.VDD(VDD),.Y(g10679),.A(g10584));
  NOT NOT1_255(.VSS(VSS),.VDD(VDD),.Y(g6796),.A(g6252));
  NOT NOT1_256(.VSS(VSS),.VDD(VDD),.Y(I8900),.A(g4560));
  NOT NOT1_257(.VSS(VSS),.VDD(VDD),.Y(I16735),.A(g10855));
  NOT NOT1_258(.VSS(VSS),.VDD(VDD),.Y(g1968),.A(g369));
  NOT NOT1_259(.VSS(VSS),.VDD(VDD),.Y(g5879),.A(I9498));
  NOT NOT1_260(.VSS(VSS),.VDD(VDD),.Y(I10963),.A(g6793));
  NOT NOT1_261(.VSS(VSS),.VDD(VDD),.Y(g10270),.A(g10156));
  NOT NOT1_262(.VSS(VSS),.VDD(VDD),.Y(g3463),.A(g3256));
  NOT NOT1_263(.VSS(VSS),.VDD(VDD),.Y(g7268),.A(I11505));
  NOT NOT1_264(.VSS(VSS),.VDD(VDD),.Y(g7362),.A(I11734));
  NOT NOT1_265(.VSS(VSS),.VDD(VDD),.Y(I11740),.A(g7030));
  NOT NOT1_266(.VSS(VSS),.VDD(VDD),.Y(g10188),.A(I15542));
  NOT NOT1_267(.VSS(VSS),.VDD(VDD),.Y(I12174),.A(g6939));
  NOT NOT1_268(.VSS(VSS),.VDD(VDD),.Y(I12796),.A(g7543));
  NOT NOT1_269(.VSS(VSS),.VDD(VDD),.Y(g5659),.A(I9138));
  NOT NOT1_270(.VSS(VSS),.VDD(VDD),.Y(g7419),.A(g7206));
  NOT NOT1_271(.VSS(VSS),.VDD(VDD),.Y(I15503),.A(g10044));
  NOT NOT1_272(.VSS(VSS),.VDD(VDD),.Y(I17441),.A(g11445));
  NOT NOT1_273(.VSS(VSS),.VDD(VDD),.Y(g6980),.A(I11127));
  NOT NOT1_274(.VSS(VSS),.VDD(VDD),.Y(I17206),.A(g11323));
  NOT NOT1_275(.VSS(VSS),.VDD(VDD),.Y(g4113),.A(I7255));
  NOT NOT1_276(.VSS(VSS),.VDD(VDD),.Y(g6069),.A(I9706));
  NOT NOT1_277(.VSS(VSS),.VDD(VDD),.Y(g11503),.A(I17528));
  NOT NOT1_278(.VSS(VSS),.VDD(VDD),.Y(g7052),.A(I11235));
  NOT NOT1_279(.VSS(VSS),.VDD(VDD),.Y(g8110),.A(g7996));
  NOT NOT1_280(.VSS(VSS),.VDD(VDD),.Y(g2556),.A(g186));
  NOT NOT1_281(.VSS(VSS),.VDD(VDD),.Y(g4313),.A(g3586));
  NOT NOT1_282(.VSS(VSS),.VDD(VDD),.Y(I16196),.A(g10496));
  NOT NOT1_283(.VSS(VSS),.VDD(VDD),.Y(I7817),.A(g3399));
  NOT NOT1_284(.VSS(VSS),.VDD(VDD),.Y(g8310),.A(I13314));
  NOT NOT1_285(.VSS(VSS),.VDD(VDD),.Y(g10460),.A(I15971));
  NOT NOT1_286(.VSS(VSS),.VDD(VDD),.Y(g2222),.A(g158));
  NOT NOT1_287(.VSS(VSS),.VDD(VDD),.Y(I11953),.A(g6907));
  NOT NOT1_288(.VSS(VSS),.VDD(VDD),.Y(I13373),.A(g8226));
  NOT NOT1_289(.VSS(VSS),.VDD(VDD),.Y(I6818),.A(g2758));
  NOT NOT1_290(.VSS(VSS),.VDD(VDD),.Y(g4202),.A(I7423));
  NOT NOT1_291(.VSS(VSS),.VDD(VDD),.Y(I6867),.A(g2949));
  NOT NOT1_292(.VSS(VSS),.VDD(VDD),.Y(I9880),.A(g5405));
  NOT NOT1_293(.VSS(VSS),.VDD(VDD),.Y(g10093),.A(I15326));
  NOT NOT1_294(.VSS(VSS),.VDD(VDD),.Y(I10484),.A(g6155));
  NOT NOT1_295(.VSS(VSS),.VDD(VDD),.Y(g9845),.A(g9679));
  NOT NOT1_296(.VSS(VSS),.VDD(VDD),.Y(g3720),.A(I6888));
  NOT NOT1_297(.VSS(VSS),.VDD(VDD),.Y(g10267),.A(g10130));
  NOT NOT1_298(.VSS(VSS),.VDD(VDD),.Y(g10294),.A(I15704));
  NOT NOT1_299(.VSS(VSS),.VDD(VDD),.Y(I11800),.A(g7246));
  NOT NOT1_300(.VSS(VSS),.VDD(VDD),.Y(g4908),.A(g4396));
  NOT NOT1_301(.VSS(VSS),.VDD(VDD),.Y(g5111),.A(I8499));
  NOT NOT1_302(.VSS(VSS),.VDD(VDD),.Y(g11450),.A(I17407));
  NOT NOT1_303(.VSS(VSS),.VDD(VDD),.Y(I13800),.A(g8500));
  NOT NOT1_304(.VSS(VSS),.VDD(VDD),.Y(g5275),.A(g4371));
  NOT NOT1_305(.VSS(VSS),.VDD(VDD),.Y(I11417),.A(g6638));
  NOT NOT1_306(.VSS(VSS),.VDD(VDD),.Y(I17758),.A(g11647));
  NOT NOT1_307(.VSS(VSS),.VDD(VDD),.Y(g3318),.A(g2245));
  NOT NOT1_308(.VSS(VSS),.VDD(VDD),.Y(g11315),.A(I17108));
  NOT NOT1_309(.VSS(VSS),.VDD(VDD),.Y(g4094),.A(g2744));
  NOT NOT1_310(.VSS(VSS),.VDD(VDD),.Y(I17435),.A(g11454));
  NOT NOT1_311(.VSS(VSS),.VDD(VDD),.Y(g10065),.A(I15293));
  NOT NOT1_312(.VSS(VSS),.VDD(VDD),.Y(I5092),.A(g32));
  NOT NOT1_313(.VSS(VSS),.VDD(VDD),.Y(g8002),.A(I12832));
  NOT NOT1_314(.VSS(VSS),.VDD(VDD),.Y(g5615),.A(I9043));
  NOT NOT1_315(.VSS(VSS),.VDD(VDD),.Y(g4567),.A(g3374));
  NOT NOT1_316(.VSS(VSS),.VDD(VDD),.Y(I8259),.A(g4590));
  NOT NOT1_317(.VSS(VSS),.VDD(VDD),.Y(g11202),.A(g11112));
  NOT NOT1_318(.VSS(VSS),.VDD(VDD),.Y(g7728),.A(I12369));
  NOT NOT1_319(.VSS(VSS),.VDD(VDD),.Y(g6287),.A(I10120));
  NOT NOT1_320(.VSS(VSS),.VDD(VDD),.Y(I14312),.A(g8814));
  NOT NOT1_321(.VSS(VSS),.VDD(VDD),.Y(I9612),.A(g5149));
  NOT NOT1_322(.VSS(VSS),.VDD(VDD),.Y(g10875),.A(I16595));
  NOT NOT1_323(.VSS(VSS),.VDD(VDD),.Y(I9243),.A(g5245));
  NOT NOT1_324(.VSS(VSS),.VDD(VDD),.Y(g11055),.A(g10950));
  NOT NOT1_325(.VSS(VSS),.VDD(VDD),.Y(g3393),.A(g3144));
  NOT NOT1_326(.VSS(VSS),.VDD(VDD),.Y(g9807),.A(g9490));
  NOT NOT1_327(.VSS(VSS),.VDD(VDD),.Y(g11111),.A(g10974));
  NOT NOT1_328(.VSS(VSS),.VDD(VDD),.Y(g4776),.A(g3586));
  NOT NOT1_329(.VSS(VSS),.VDD(VDD),.Y(I9935),.A(g5477));
  NOT NOT1_330(.VSS(VSS),.VDD(VDD),.Y(g4593),.A(I8004));
  NOT NOT1_331(.VSS(VSS),.VDD(VDD),.Y(I11964),.A(g6910));
  NOT NOT1_332(.VSS(VSS),.VDD(VDD),.Y(I7441),.A(g3473));
  NOT NOT1_333(.VSS(VSS),.VDD(VDD),.Y(I15986),.A(g10417));
  NOT NOT1_334(.VSS(VSS),.VDD(VDD),.Y(g3971),.A(I7104));
  NOT NOT1_335(.VSS(VSS),.VDD(VDD),.Y(g7070),.A(I11289));
  NOT NOT1_336(.VSS(VSS),.VDD(VDD),.Y(g2237),.A(g713));
  NOT NOT1_337(.VSS(VSS),.VDD(VDD),.Y(g6399),.A(I10305));
  NOT NOT1_338(.VSS(VSS),.VDD(VDD),.Y(g5284),.A(g4376));
  NOT NOT1_339(.VSS(VSS),.VDD(VDD),.Y(I11423),.A(g6488));
  NOT NOT1_340(.VSS(VSS),.VDD(VDD),.Y(g7470),.A(g6927));
  NOT NOT1_341(.VSS(VSS),.VDD(VDD),.Y(I15741),.A(g10260));
  NOT NOT1_342(.VSS(VSS),.VDD(VDD),.Y(g7897),.A(g7712));
  NOT NOT1_343(.VSS(VSS),.VDD(VDD),.Y(g7025),.A(g6400));
  NOT NOT1_344(.VSS(VSS),.VDD(VDD),.Y(I6370),.A(g2356));
  NOT NOT1_345(.VSS(VSS),.VDD(VDD),.Y(g7425),.A(g7214));
  NOT NOT1_346(.VSS(VSS),.VDD(VDD),.Y(I11587),.A(g6828));
  NOT NOT1_347(.VSS(VSS),.VDD(VDD),.Y(g2844),.A(I5966));
  NOT NOT1_348(.VSS(VSS),.VDD(VDD),.Y(I12553),.A(g7676));
  NOT NOT1_349(.VSS(VSS),.VDD(VDD),.Y(I12862),.A(g7638));
  NOT NOT1_350(.VSS(VSS),.VDD(VDD),.Y(I8215),.A(g3981));
  NOT NOT1_351(.VSS(VSS),.VDD(VDD),.Y(I10813),.A(g6397));
  NOT NOT1_352(.VSS(VSS),.VDD(VDD),.Y(g11384),.A(I17209));
  NOT NOT1_353(.VSS(VSS),.VDD(VDD),.Y(I14799),.A(g9661));
  NOT NOT1_354(.VSS(VSS),.VDD(VDD),.Y(I6821),.A(g3015));
  NOT NOT1_355(.VSS(VSS),.VDD(VDD),.Y(g2194),.A(g47));
  NOT NOT1_356(.VSS(VSS),.VDD(VDD),.Y(g10160),.A(I15476));
  NOT NOT1_357(.VSS(VSS),.VDD(VDD),.Y(g6797),.A(I10801));
  NOT NOT1_358(.VSS(VSS),.VDD(VDD),.Y(g11067),.A(g10974));
  NOT NOT1_359(.VSS(VSS),.VDD(VDD),.Y(g9342),.A(I14531));
  NOT NOT1_360(.VSS(VSS),.VDD(VDD),.Y(I12326),.A(g7246));
  NOT NOT1_361(.VSS(VSS),.VDD(VDD),.Y(g8928),.A(I14257));
  NOT NOT1_362(.VSS(VSS),.VDD(VDD),.Y(g3121),.A(g2462));
  NOT NOT1_363(.VSS(VSS),.VDD(VDD),.Y(I16280),.A(g10537));
  NOT NOT1_364(.VSS(VSS),.VDD(VDD),.Y(g4160),.A(I7303));
  NOT NOT1_365(.VSS(VSS),.VDD(VDD),.Y(g3321),.A(I6484));
  NOT NOT1_366(.VSS(VSS),.VDD(VDD),.Y(g2089),.A(I4917));
  NOT NOT1_367(.VSS(VSS),.VDD(VDD),.Y(g4933),.A(I8298));
  NOT NOT1_368(.VSS(VSS),.VDD(VDD),.Y(I14973),.A(g9733));
  NOT NOT1_369(.VSS(VSS),.VDD(VDD),.Y(g2731),.A(I5789));
  NOT NOT1_370(.VSS(VSS),.VDD(VDD),.Y(I16688),.A(g10800));
  NOT NOT1_371(.VSS(VSS),.VDD(VDD),.Y(I11543),.A(g6881));
  NOT NOT1_372(.VSS(VSS),.VDD(VDD),.Y(g5420),.A(g4300));
  NOT NOT1_373(.VSS(VSS),.VDD(VDD),.Y(I15801),.A(g10282));
  NOT NOT1_374(.VSS(VSS),.VDD(VDD),.Y(I12948),.A(g8019));
  NOT NOT1_375(.VSS(VSS),.VDD(VDD),.Y(g10455),.A(I15956));
  NOT NOT1_376(.VSS(VSS),.VDD(VDD),.Y(g8064),.A(I12910));
  NOT NOT1_377(.VSS(VSS),.VDD(VDD),.Y(g4521),.A(g3586));
  NOT NOT1_378(.VSS(VSS),.VDD(VDD),.Y(I14805),.A(g9360));
  NOT NOT1_379(.VSS(VSS),.VDD(VDD),.Y(g6291),.A(I10132));
  NOT NOT1_380(.VSS(VSS),.VDD(VDD),.Y(g2557),.A(g1840));
  NOT NOT1_381(.VSS(VSS),.VDD(VDD),.Y(g4050),.A(I7163));
  NOT NOT1_382(.VSS(VSS),.VDD(VDD),.Y(I13117),.A(g7904));
  NOT NOT1_383(.VSS(VSS),.VDD(VDD),.Y(I12904),.A(g7985));
  NOT NOT1_384(.VSS(VSS),.VDD(VDD),.Y(I4873),.A(g105));
  NOT NOT1_385(.VSS(VSS),.VDD(VDD),.Y(g8785),.A(I14090));
  NOT NOT1_386(.VSS(VSS),.VDD(VDD),.Y(g4450),.A(g3914));
  NOT NOT1_387(.VSS(VSS),.VDD(VDD),.Y(g5794),.A(I9394));
  NOT NOT1_388(.VSS(VSS),.VDD(VDD),.Y(g9097),.A(g8892));
  NOT NOT1_389(.VSS(VSS),.VDD(VDD),.Y(g2071),.A(I4873));
  NOT NOT1_390(.VSS(VSS),.VDD(VDD),.Y(g7678),.A(I12307));
  NOT NOT1_391(.VSS(VSS),.VDD(VDD),.Y(g6144),.A(I9857));
  NOT NOT1_392(.VSS(VSS),.VDD(VDD),.Y(I11569),.A(g6821));
  NOT NOT1_393(.VSS(VSS),.VDD(VDD),.Y(g3253),.A(I6417));
  NOT NOT1_394(.VSS(VSS),.VDD(VDD),.Y(I7743),.A(g3762));
  NOT NOT1_395(.VSS(VSS),.VDD(VDD),.Y(g6344),.A(I10251));
  NOT NOT1_396(.VSS(VSS),.VDD(VDD),.Y(g3938),.A(g2991));
  NOT NOT1_397(.VSS(VSS),.VDD(VDD),.Y(g7331),.A(I11641));
  NOT NOT1_398(.VSS(VSS),.VDD(VDD),.Y(I15196),.A(g9974));
  NOT NOT1_399(.VSS(VSS),.VDD(VDD),.Y(g9354),.A(I14567));
  NOT NOT1_400(.VSS(VSS),.VDD(VDD),.Y(g10201),.A(g10175));
  NOT NOT1_401(.VSS(VSS),.VDD(VDD),.Y(g7406),.A(I11786));
  NOT NOT1_402(.VSS(VSS),.VDD(VDD),.Y(g10277),.A(I15675));
  NOT NOT1_403(.VSS(VSS),.VDD(VDD),.Y(g2242),.A(I5245));
  NOT NOT1_404(.VSS(VSS),.VDD(VDD),.Y(I9213),.A(g4944));
  NOT NOT1_405(.VSS(VSS),.VDD(VDD),.Y(g3909),.A(g2920));
  NOT NOT1_406(.VSS(VSS),.VDD(VDD),.Y(I6106),.A(g2116));
  NOT NOT1_407(.VSS(VSS),.VDD(VDD),.Y(g7635),.A(I12245));
  NOT NOT1_408(.VSS(VSS),.VDD(VDD),.Y(I4869),.A(g253));
  NOT NOT1_409(.VSS(VSS),.VDD(VDD),.Y(I13568),.A(g8343));
  NOT NOT1_410(.VSS(VSS),.VDD(VDD),.Y(I13747),.A(g8299));
  NOT NOT1_411(.VSS(VSS),.VDD(VDD),.Y(I15526),.A(g10051));
  NOT NOT1_412(.VSS(VSS),.VDD(VDD),.Y(g8563),.A(I13782));
  NOT NOT1_413(.VSS(VSS),.VDD(VDD),.Y(g10075),.A(I15302));
  NOT NOT1_414(.VSS(VSS),.VDD(VDD),.Y(g4724),.A(g3586));
  NOT NOT1_415(.VSS(VSS),.VDD(VDD),.Y(g6259),.A(I10036));
  NOT NOT1_416(.VSS(VSS),.VDD(VDD),.Y(g4179),.A(I7354));
  NOT NOT1_417(.VSS(VSS),.VDD(VDD),.Y(g7766),.A(I12463));
  NOT NOT1_418(.VSS(VSS),.VDD(VDD),.Y(I5722),.A(g2075));
  NOT NOT1_419(.VSS(VSS),.VDD(VDD),.Y(g7682),.A(g7148));
  NOT NOT1_420(.VSS(VSS),.VDD(VDD),.Y(I13242),.A(g8267));
  NOT NOT1_421(.VSS(VSS),.VDD(VDD),.Y(I17500),.A(g11478));
  NOT NOT1_422(.VSS(VSS),.VDD(VDD),.Y(g6694),.A(I10663));
  NOT NOT1_423(.VSS(VSS),.VDD(VDD),.Y(g4379),.A(g3698));
  NOT NOT1_424(.VSS(VSS),.VDD(VDD),.Y(g3519),.A(g3164));
  NOT NOT1_425(.VSS(VSS),.VDD(VDD),.Y(g7801),.A(I12568));
  NOT NOT1_426(.VSS(VSS),.VDD(VDD),.Y(g7305),.A(I11563));
  NOT NOT1_427(.VSS(VSS),.VDD(VDD),.Y(I7411),.A(g4140));
  NOT NOT1_428(.VSS(VSS),.VDD(VDD),.Y(g8295),.A(I13239));
  NOT NOT1_429(.VSS(VSS),.VDD(VDD),.Y(g2955),.A(I6156));
  NOT NOT1_430(.VSS(VSS),.VDD(VDD),.Y(I8136),.A(g4144));
  NOT NOT1_431(.VSS(VSS),.VDD(VDD),.Y(g5628),.A(I9062));
  NOT NOT1_432(.VSS(VSS),.VDD(VDD),.Y(I6061),.A(g2246));
  NOT NOT1_433(.VSS(VSS),.VDD(VDD),.Y(I12183),.A(g7007));
  NOT NOT1_434(.VSS(VSS),.VDD(VDD),.Y(g6852),.A(I10914));
  NOT NOT1_435(.VSS(VSS),.VDD(VDD),.Y(I11814),.A(g7196));
  NOT NOT1_436(.VSS(VSS),.VDD(VDD),.Y(g5515),.A(g4429));
  NOT NOT1_437(.VSS(VSS),.VDD(VDD),.Y(I6461),.A(g2261));
  NOT NOT1_438(.VSS(VSS),.VDD(VDD),.Y(g5630),.A(I9068));
  NOT NOT1_439(.VSS(VSS),.VDD(VDD),.Y(I12397),.A(g7284));
  NOT NOT1_440(.VSS(VSS),.VDD(VDD),.Y(I4917),.A(g584));
  NOT NOT1_441(.VSS(VSS),.VDD(VDD),.Y(g2254),.A(g131));
  NOT NOT1_442(.VSS(VSS),.VDD(VDD),.Y(g2814),.A(I5916));
  NOT NOT1_443(.VSS(VSS),.VDD(VDD),.Y(g11402),.A(I17249));
  NOT NOT1_444(.VSS(VSS),.VDD(VDD),.Y(g4289),.A(g4013));
  NOT NOT1_445(.VSS(VSS),.VDD(VDD),.Y(g7748),.A(I12409));
  NOT NOT1_446(.VSS(VSS),.VDD(VDD),.Y(g4777),.A(g3992));
  NOT NOT1_447(.VSS(VSS),.VDD(VDD),.Y(I11807),.A(g6854));
  NOT NOT1_448(.VSS(VSS),.VDD(VDD),.Y(g11457),.A(I17424));
  NOT NOT1_449(.VSS(VSS),.VDD(VDD),.Y(I9090),.A(g5567));
  NOT NOT1_450(.VSS(VSS),.VDD(VDD),.Y(g4835),.A(I8192));
  NOT NOT1_451(.VSS(VSS),.VDD(VDD),.Y(I14400),.A(g8891));
  NOT NOT1_452(.VSS(VSS),.VDD(VDD),.Y(g2350),.A(I5424));
  NOT NOT1_453(.VSS(VSS),.VDD(VDD),.Y(g7755),.A(I12430));
  NOT NOT1_454(.VSS(VSS),.VDD(VDD),.Y(g9267),.A(g8892));
  NOT NOT1_455(.VSS(VSS),.VDD(VDD),.Y(g9312),.A(I14509));
  NOT NOT1_456(.VSS(VSS),.VDD(VDD),.Y(I13639),.A(g8321));
  NOT NOT1_457(.VSS(VSS),.VDD(VDD),.Y(g2038),.A(g1776));
  NOT NOT1_458(.VSS(VSS),.VDD(VDD),.Y(I8943),.A(g4585));
  NOT NOT1_459(.VSS(VSS),.VDD(VDD),.Y(I16763),.A(g10890));
  NOT NOT1_460(.VSS(VSS),.VDD(VDD),.Y(I12933),.A(g7899));
  NOT NOT1_461(.VSS(VSS),.VDD(VDD),.Y(g7226),.A(I11464));
  NOT NOT1_462(.VSS(VSS),.VDD(VDD),.Y(g8089),.A(g7934));
  NOT NOT1_463(.VSS(VSS),.VDD(VDD),.Y(g10352),.A(I15820));
  NOT NOT1_464(.VSS(VSS),.VDD(VDD),.Y(g2438),.A(g243));
  NOT NOT1_465(.VSS(VSS),.VDD(VDD),.Y(I11293),.A(g6516));
  NOT NOT1_466(.VSS(VSS),.VDD(VDD),.Y(I13230),.A(g8244));
  NOT NOT1_467(.VSS(VSS),.VDD(VDD),.Y(g2773),.A(I5858));
  NOT NOT1_468(.VSS(VSS),.VDD(VDD),.Y(g4271),.A(g3971));
  NOT NOT1_469(.VSS(VSS),.VDD(VDD),.Y(I6904),.A(g2820));
  NOT NOT1_470(.VSS(VSS),.VDD(VDD),.Y(I12508),.A(g7731));
  NOT NOT1_471(.VSS(VSS),.VDD(VDD),.Y(I11638),.A(g6948));
  NOT NOT1_472(.VSS(VSS),.VDD(VDD),.Y(I12634),.A(g7727));
  NOT NOT1_473(.VSS(VSS),.VDD(VDD),.Y(g10155),.A(I15461));
  NOT NOT1_474(.VSS(VSS),.VDD(VDD),.Y(I17613),.A(g11550));
  NOT NOT1_475(.VSS(VSS),.VDD(VDD),.Y(g10822),.A(I16534));
  NOT NOT1_476(.VSS(VSS),.VDD(VDD),.Y(I4786),.A(g109));
  NOT NOT1_477(.VSS(VSS),.VDD(VDD),.Y(I6046),.A(g2218));
  NOT NOT1_478(.VSS(VSS),.VDD(VDD),.Y(I9056),.A(g4753));
  NOT NOT1_479(.VSS(VSS),.VDD(VDD),.Y(g6951),.A(I11097));
  NOT NOT1_480(.VSS(VSS),.VDD(VDD),.Y(g10266),.A(g10129));
  NOT NOT1_481(.VSS(VSS),.VDD(VDD),.Y(I8228),.A(g4468));
  NOT NOT1_482(.VSS(VSS),.VDD(VDD),.Y(I14005),.A(g8631));
  NOT NOT1_483(.VSS(VSS),.VDD(VDD),.Y(g10170),.A(g10118));
  NOT NOT1_484(.VSS(VSS),.VDD(VDD),.Y(I8465),.A(g4807));
  NOT NOT1_485(.VSS(VSS),.VDD(VDD),.Y(I16660),.A(g10793));
  NOT NOT1_486(.VSS(VSS),.VDD(VDD),.Y(g7045),.A(g6435));
  NOT NOT1_487(.VSS(VSS),.VDD(VDD),.Y(I10538),.A(g5910));
  NOT NOT1_488(.VSS(VSS),.VDD(VDD),.Y(I8934),.A(g4271));
  NOT NOT1_489(.VSS(VSS),.VDD(VDD),.Y(I5424),.A(g910));
  NOT NOT1_490(.VSS(VSS),.VDD(VDD),.Y(I5795),.A(g2462));
  NOT NOT1_491(.VSS(VSS),.VDD(VDD),.Y(g7445),.A(I11845));
  NOT NOT1_492(.VSS(VSS),.VDD(VDD),.Y(g6114),.A(I9795));
  NOT NOT1_493(.VSS(VSS),.VDD(VDD),.Y(I5737),.A(g2100));
  NOT NOT1_494(.VSS(VSS),.VDD(VDD),.Y(I6403),.A(g2337));
  NOT NOT1_495(.VSS(VSS),.VDD(VDD),.Y(I5809),.A(g2356));
  NOT NOT1_496(.VSS(VSS),.VDD(VDD),.Y(g6314),.A(I10201));
  NOT NOT1_497(.VSS(VSS),.VDD(VDD),.Y(I7713),.A(g3750));
  NOT NOT1_498(.VSS(VSS),.VDD(VDD),.Y(g9761),.A(g9454));
  NOT NOT1_499(.VSS(VSS),.VDD(VDD),.Y(I11841),.A(g7226));
  NOT NOT1_500(.VSS(VSS),.VDD(VDD),.Y(I11992),.A(g7058));
  NOT NOT1_501(.VSS(VSS),.VDD(VDD),.Y(I11391),.A(g6387));
  NOT NOT1_502(.VSS(VSS),.VDD(VDD),.Y(I9851),.A(g5405));
  NOT NOT1_503(.VSS(VSS),.VDD(VDD),.Y(g2212),.A(g686));
  NOT NOT1_504(.VSS(VSS),.VDD(VDD),.Y(I13391),.A(g8178));
  NOT NOT1_505(.VSS(VSS),.VDD(VDD),.Y(g6870),.A(I10952));
  NOT NOT1_506(.VSS(VSS),.VDD(VDD),.Y(g4674),.A(I8050));
  NOT NOT1_507(.VSS(VSS),.VDD(VDD),.Y(g8948),.A(I14299));
  NOT NOT1_508(.VSS(VSS),.VDD(VDD),.Y(g3141),.A(g2563));
  NOT NOT1_509(.VSS(VSS),.VDD(VDD),.Y(I6391),.A(g2478));
  NOT NOT1_510(.VSS(VSS),.VDD(VDD),.Y(I5672),.A(g569));
  NOT NOT1_511(.VSS(VSS),.VDD(VDD),.Y(I15688),.A(g10207));
  NOT NOT1_512(.VSS(VSS),.VDD(VDD),.Y(g5040),.A(I8421));
  NOT NOT1_513(.VSS(VSS),.VDD(VDD),.Y(I5077),.A(g35));
  NOT NOT1_514(.VSS(VSS),.VDD(VDD),.Y(g1983),.A(g750));
  NOT NOT1_515(.VSS(VSS),.VDD(VDD),.Y(g6825),.A(I10873));
  NOT NOT1_516(.VSS(VSS),.VDD(VDD),.Y(g3710),.A(g3215));
  NOT NOT1_517(.VSS(VSS),.VDD(VDD),.Y(g7369),.A(g7273));
  NOT NOT1_518(.VSS(VSS),.VDD(VDD),.Y(g7602),.A(I12156));
  NOT NOT1_519(.VSS(VSS),.VDD(VDD),.Y(g10167),.A(I15497));
  NOT NOT1_520(.VSS(VSS),.VDD(VDD),.Y(g10194),.A(g10062));
  NOT NOT1_521(.VSS(VSS),.VDD(VDD),.Y(g10589),.A(I16252));
  NOT NOT1_522(.VSS(VSS),.VDD(VDD),.Y(I16550),.A(g10726));
  NOT NOT1_523(.VSS(VSS),.VDD(VDD),.Y(g4541),.A(I7946));
  NOT NOT1_524(.VSS(VSS),.VDD(VDD),.Y(g7007),.A(I11146));
  NOT NOT1_525(.VSS(VSS),.VDD(VDD),.Y(I17371),.A(g11410));
  NOT NOT1_526(.VSS(VSS),.VDD(VDD),.Y(I17234),.A(g11353));
  NOT NOT1_527(.VSS(VSS),.VDD(VDD),.Y(g7920),.A(g7516));
  NOT NOT1_528(.VSS(VSS),.VDD(VDD),.Y(I11578),.A(g6824));
  NOT NOT1_529(.VSS(VSS),.VDD(VDD),.Y(I12574),.A(g7522));
  NOT NOT1_530(.VSS(VSS),.VDD(VDD),.Y(g10524),.A(g10458));
  NOT NOT1_531(.VSS(VSS),.VDD(VDD),.Y(g2229),.A(g162));
  NOT NOT1_532(.VSS(VSS),.VDD(VDD),.Y(I15157),.A(g9931));
  NOT NOT1_533(.VSS(VSS),.VDD(VDD),.Y(I16307),.A(g10589));
  NOT NOT1_534(.VSS(VSS),.VDD(VDD),.Y(g4332),.A(g4130));
  NOT NOT1_535(.VSS(VSS),.VDD(VDD),.Y(I12205),.A(g6993));
  NOT NOT1_536(.VSS(VSS),.VDD(VDD),.Y(g7767),.A(I12466));
  NOT NOT1_537(.VSS(VSS),.VDD(VDD),.Y(I6159),.A(g2123));
  NOT NOT1_538(.VSS(VSS),.VDD(VDD),.Y(g11157),.A(g10950));
  NOT NOT1_539(.VSS(VSS),.VDD(VDD),.Y(g4680),.A(g3829));
  NOT NOT1_540(.VSS(VSS),.VDD(VDD),.Y(g6136),.A(I9845));
  NOT NOT1_541(.VSS(VSS),.VDD(VDD),.Y(g8150),.A(I13039));
  NOT NOT1_542(.VSS(VSS),.VDD(VDD),.Y(g4209),.A(I7444));
  NOT NOT1_543(.VSS(VSS),.VDD(VDD),.Y(g4353),.A(I7636));
  NOT NOT1_544(.VSS(VSS),.VDD(VDD),.Y(g5666),.A(I9159));
  NOT NOT1_545(.VSS(VSS),.VDD(VDD),.Y(g6336),.A(I10231));
  NOT NOT1_546(.VSS(VSS),.VDD(VDD),.Y(g8350),.A(I13430));
  NOT NOT1_547(.VSS(VSS),.VDD(VDD),.Y(I13586),.A(g8356));
  NOT NOT1_548(.VSS(VSS),.VDD(VDD),.Y(g10119),.A(I15365));
  NOT NOT1_549(.VSS(VSS),.VDD(VDD),.Y(I8337),.A(g4352));
  NOT NOT1_550(.VSS(VSS),.VDD(VDD),.Y(g8438),.A(I13612));
  NOT NOT1_551(.VSS(VSS),.VDD(VDD),.Y(g6594),.A(I10560));
  NOT NOT1_552(.VSS(VSS),.VDD(VDD),.Y(g11066),.A(g10974));
  NOT NOT1_553(.VSS(VSS),.VDD(VDD),.Y(g4802),.A(g3337));
  NOT NOT1_554(.VSS(VSS),.VDD(VDD),.Y(I13442),.A(g8182));
  NOT NOT1_555(.VSS(VSS),.VDD(VDD),.Y(g8009),.A(I12849));
  NOT NOT1_556(.VSS(VSS),.VDD(VDD),.Y(I5304),.A(g79));
  NOT NOT1_557(.VSS(VSS),.VDD(VDD),.Y(g10118),.A(I15362));
  NOT NOT1_558(.VSS(VSS),.VDD(VDD),.Y(I6016),.A(g2201));
  NOT NOT1_559(.VSS(VSS),.VDD(VDD),.Y(I6757),.A(g2732));
  NOT NOT1_560(.VSS(VSS),.VDD(VDD),.Y(g7793),.A(I12544));
  NOT NOT1_561(.VSS(VSS),.VDD(VDD),.Y(I9279),.A(g5314));
  NOT NOT1_562(.VSS(VSS),.VDD(VDD),.Y(g5648),.A(I9105));
  NOT NOT1_563(.VSS(VSS),.VDD(VDD),.Y(g6806),.A(I10828));
  NOT NOT1_564(.VSS(VSS),.VDD(VDD),.Y(g5875),.A(g5361));
  NOT NOT1_565(.VSS(VSS),.VDD(VDD),.Y(g6943),.A(I11079));
  NOT NOT1_566(.VSS(VSS),.VDD(VDD),.Y(I16269),.A(g10558));
  NOT NOT1_567(.VSS(VSS),.VDD(VDD),.Y(I9720),.A(g5248));
  NOT NOT1_568(.VSS(VSS),.VDD(VDD),.Y(I12592),.A(g7445));
  NOT NOT1_569(.VSS(VSS),.VDD(VDD),.Y(g10616),.A(I16289));
  NOT NOT1_570(.VSS(VSS),.VDD(VDD),.Y(g4558),.A(g3880));
  NOT NOT1_571(.VSS(VSS),.VDD(VDD),.Y(g5655),.A(I9126));
  NOT NOT1_572(.VSS(VSS),.VDD(VDD),.Y(I13615),.A(g8333));
  NOT NOT1_573(.VSS(VSS),.VDD(VDD),.Y(g7415),.A(I11797));
  NOT NOT1_574(.VSS(VSS),.VDD(VDD),.Y(g7227),.A(I11467));
  NOT NOT1_575(.VSS(VSS),.VDD(VDD),.Y(I9872),.A(g5557));
  NOT NOT1_576(.VSS(VSS),.VDD(VDD),.Y(g10313),.A(I15741));
  NOT NOT1_577(.VSS(VSS),.VDD(VDD),.Y(I5926),.A(g2172));
  NOT NOT1_578(.VSS(VSS),.VDD(VDD),.Y(I13720),.A(g8358));
  NOT NOT1_579(.VSS(VSS),.VDD(VDD),.Y(I9652),.A(g5426));
  NOT NOT1_580(.VSS(VSS),.VDD(VDD),.Y(I5754),.A(g2304));
  NOT NOT1_581(.VSS(VSS),.VDD(VDD),.Y(I10991),.A(g6759));
  NOT NOT1_582(.VSS(VSS),.VDD(VDD),.Y(I15763),.A(g10244));
  NOT NOT1_583(.VSS(VSS),.VDD(VDD),.Y(I11275),.A(g6502));
  NOT NOT1_584(.VSS(VSS),.VDD(VDD),.Y(g10276),.A(I15672));
  NOT NOT1_585(.VSS(VSS),.VDD(VDD),.Y(g11511),.A(I17552));
  NOT NOT1_586(.VSS(VSS),.VDD(VDD),.Y(g4901),.A(I8268));
  NOT NOT1_587(.VSS(VSS),.VDD(VDD),.Y(I7760),.A(g3768));
  NOT NOT1_588(.VSS(VSS),.VDD(VDD),.Y(I16670),.A(g10797));
  NOT NOT1_589(.VSS(VSS),.VDD(VDD),.Y(I11746),.A(g6857));
  NOT NOT1_590(.VSS(VSS),.VDD(VDD),.Y(I13430),.A(g8241));
  NOT NOT1_591(.VSS(VSS),.VDD(VDD),.Y(g10305),.A(I15725));
  NOT NOT1_592(.VSS(VSS),.VDD(VDD),.Y(g10254),.A(g10196));
  NOT NOT1_593(.VSS(VSS),.VDD(VDD),.Y(g4511),.A(g3586));
  NOT NOT1_594(.VSS(VSS),.VDD(VDD),.Y(g10900),.A(I16656));
  NOT NOT1_595(.VSS(VSS),.VDD(VDD),.Y(g9576),.A(I14713));
  NOT NOT1_596(.VSS(VSS),.VDD(VDD),.Y(g2837),.A(g2130));
  NOT NOT1_597(.VSS(VSS),.VDD(VDD),.Y(g10466),.A(I15989));
  NOT NOT1_598(.VSS(VSS),.VDD(VDD),.Y(g5884),.A(I9505));
  NOT NOT1_599(.VSS(VSS),.VDD(VDD),.Y(I5044),.A(g1182));
  NOT NOT1_600(.VSS(VSS),.VDD(VDD),.Y(g6433),.A(I10349));
  NOT NOT1_601(.VSS(VSS),.VDD(VDD),.Y(g5839),.A(I9452));
  NOT NOT1_602(.VSS(VSS),.VDD(VDD),.Y(g8229),.A(g7826));
  NOT NOT1_603(.VSS(VSS),.VDD(VDD),.Y(I6654),.A(g2952));
  NOT NOT1_604(.VSS(VSS),.VDD(VDD),.Y(g8993),.A(I14400));
  NOT NOT1_605(.VSS(VSS),.VDD(VDD),.Y(g2620),.A(g1998));
  NOT NOT1_606(.VSS(VSS),.VDD(VDD),.Y(I12846),.A(g7685));
  NOT NOT1_607(.VSS(VSS),.VDD(VDD),.Y(g2462),.A(I5555));
  NOT NOT1_608(.VSS(VSS),.VDD(VDD),.Y(g9349),.A(I14552));
  NOT NOT1_609(.VSS(VSS),.VDD(VDD),.Y(I8815),.A(g4471));
  NOT NOT1_610(.VSS(VSS),.VDD(VDD),.Y(g10101),.A(I15335));
  NOT NOT1_611(.VSS(VSS),.VDD(VDD),.Y(g10177),.A(I15523));
  NOT NOT1_612(.VSS(VSS),.VDD(VDD),.Y(I16667),.A(g10780));
  NOT NOT1_613(.VSS(VSS),.VDD(VDD),.Y(I13806),.A(g8478));
  NOT NOT1_614(.VSS(VSS),.VDD(VDD),.Y(I7220),.A(g3213));
  NOT NOT1_615(.VSS(VSS),.VDD(VDD),.Y(I5862),.A(g2537));
  NOT NOT1_616(.VSS(VSS),.VDD(VDD),.Y(I9598),.A(g5120));
  NOT NOT1_617(.VSS(VSS),.VDD(VDD),.Y(I7779),.A(g3774));
  NOT NOT1_618(.VSS(VSS),.VDD(VDD),.Y(I17724),.A(g11625));
  NOT NOT1_619(.VSS(VSS),.VDD(VDD),.Y(g6845),.A(I10907));
  NOT NOT1_620(.VSS(VSS),.VDD(VDD),.Y(g7502),.A(I11882));
  NOT NOT1_621(.VSS(VSS),.VDD(VDD),.Y(I8154),.A(g3636));
  NOT NOT1_622(.VSS(VSS),.VDD(VDD),.Y(I10584),.A(g5864));
  NOT NOT1_623(.VSS(VSS),.VDD(VDD),.Y(I17359),.A(g11372));
  NOT NOT1_624(.VSS(VSS),.VDD(VDD),.Y(g3545),.A(I6733));
  NOT NOT1_625(.VSS(VSS),.VDD(VDD),.Y(I15314),.A(g10007));
  NOT NOT1_626(.VSS(VSS),.VDD(VDD),.Y(g11550),.A(I17591));
  NOT NOT1_627(.VSS(VSS),.VDD(VDD),.Y(I15287),.A(g9980));
  NOT NOT1_628(.VSS(VSS),.VDD(VDD),.Y(g6195),.A(g5426));
  NOT NOT1_629(.VSS(VSS),.VDD(VDD),.Y(I7423),.A(g3331));
  NOT NOT1_630(.VSS(VSS),.VDD(VDD),.Y(g6137),.A(I9848));
  NOT NOT1_631(.VSS(VSS),.VDD(VDD),.Y(g5667),.A(I9162));
  NOT NOT1_632(.VSS(VSS),.VDD(VDD),.Y(g6395),.A(I10293));
  NOT NOT1_633(.VSS(VSS),.VDD(VDD),.Y(g3380),.A(I6576));
  NOT NOT1_634(.VSS(VSS),.VDD(VDD),.Y(g5143),.A(g4682));
  NOT NOT1_635(.VSS(VSS),.VDD(VDD),.Y(g6337),.A(I10234));
  NOT NOT1_636(.VSS(VSS),.VDD(VDD),.Y(I16487),.A(g10771));
  NOT NOT1_637(.VSS(VSS),.VDD(VDD),.Y(g6913),.A(I11021));
  NOT NOT1_638(.VSS(VSS),.VDD(VDD),.Y(g10064),.A(I15290));
  NOT NOT1_639(.VSS(VSS),.VDD(VDD),.Y(g11287),.A(g11207));
  NOT NOT1_640(.VSS(VSS),.VDD(VDD),.Y(I15085),.A(g9720));
  NOT NOT1_641(.VSS(VSS),.VDD(VDD),.Y(g2249),.A(g127));
  NOT NOT1_642(.VSS(VSS),.VDD(VDD),.Y(I9625),.A(g5405));
  NOT NOT1_643(.VSS(VSS),.VDD(VDD),.Y(g4580),.A(g3880));
  NOT NOT1_644(.VSS(VSS),.VDD(VDD),.Y(I10759),.A(g5803));
  NOT NOT1_645(.VSS(VSS),.VDD(VDD),.Y(g11307),.A(I17092));
  NOT NOT1_646(.VSS(VSS),.VDD(VDD),.Y(g11076),.A(I16843));
  NOT NOT1_647(.VSS(VSS),.VDD(VDD),.Y(I9232),.A(g4944));
  NOT NOT1_648(.VSS(VSS),.VDD(VDD),.Y(g7188),.A(I11408));
  NOT NOT1_649(.VSS(VSS),.VDD(VDD),.Y(g7689),.A(I12322));
  NOT NOT1_650(.VSS(VSS),.VDD(VDD),.Y(I17121),.A(g11231));
  NOT NOT1_651(.VSS(VSS),.VDD(VDD),.Y(g11596),.A(g11580));
  NOT NOT1_652(.VSS(VSS),.VDD(VDD),.Y(g7388),.A(I11773));
  NOT NOT1_653(.VSS(VSS),.VDD(VDD),.Y(I10114),.A(g5768));
  NOT NOT1_654(.VSS(VSS),.VDD(VDD),.Y(I9253),.A(g5052));
  NOT NOT1_655(.VSS(VSS),.VDD(VDD),.Y(I9938),.A(g5478));
  NOT NOT1_656(.VSS(VSS),.VDD(VDD),.Y(g10874),.A(I16592));
  NOT NOT1_657(.VSS(VSS),.VDD(VDD),.Y(g11054),.A(g10950));
  NOT NOT1_658(.VSS(VSS),.VDD(VDD),.Y(g6807),.A(I10831));
  NOT NOT1_659(.VSS(VSS),.VDD(VDD),.Y(I9813),.A(g5241));
  NOT NOT1_660(.VSS(VSS),.VDD(VDD),.Y(I6417),.A(g2344));
  NOT NOT1_661(.VSS(VSS),.VDD(VDD),.Y(g5693),.A(I9224));
  NOT NOT1_662(.VSS(VSS),.VDD(VDD),.Y(g11243),.A(g11112));
  NOT NOT1_663(.VSS(VSS),.VDD(VDD),.Y(I17344),.A(g11369));
  NOT NOT1_664(.VSS(VSS),.VDD(VDD),.Y(g3507),.A(g3307));
  NOT NOT1_665(.VSS(VSS),.VDD(VDD),.Y(g4262),.A(g4013));
  NOT NOT1_666(.VSS(VSS),.VDD(VDD),.Y(g2298),.A(I5336));
  NOT NOT1_667(.VSS(VSS),.VDD(VDD),.Y(g2085),.A(I4903));
  NOT NOT1_668(.VSS(VSS),.VDD(VDD),.Y(I7665),.A(g3732));
  NOT NOT1_669(.VSS(VSS),.VDD(VDD),.Y(g10630),.A(I16311));
  NOT NOT1_670(.VSS(VSS),.VDD(VDD),.Y(g11431),.A(I17344));
  NOT NOT1_671(.VSS(VSS),.VDD(VDD),.Y(g6859),.A(I10937));
  NOT NOT1_672(.VSS(VSS),.VDD(VDD),.Y(g7028),.A(g6407));
  NOT NOT1_673(.VSS(VSS),.VDD(VDD),.Y(I6982),.A(g2889));
  NOT NOT1_674(.VSS(VSS),.VDD(VDD),.Y(g6266),.A(I10057));
  NOT NOT1_675(.VSS(VSS),.VDD(VDD),.Y(I15269),.A(g9993));
  NOT NOT1_676(.VSS(VSS),.VDD(VDD),.Y(g10166),.A(I15494));
  NOT NOT1_677(.VSS(VSS),.VDD(VDD),.Y(g7030),.A(I11183));
  NOT NOT1_678(.VSS(VSS),.VDD(VDD),.Y(I12583),.A(g7546));
  NOT NOT1_679(.VSS(VSS),.VDD(VDD),.Y(I9519),.A(g4998));
  NOT NOT1_680(.VSS(VSS),.VDD(VDD),.Y(g8062),.A(I12904));
  NOT NOT1_681(.VSS(VSS),.VDD(VDD),.Y(g7430),.A(g7221));
  NOT NOT1_682(.VSS(VSS),.VDD(VDD),.Y(I15341),.A(g10019));
  NOT NOT1_683(.VSS(VSS),.VDD(VDD),.Y(I5414),.A(g904));
  NOT NOT1_684(.VSS(VSS),.VDD(VDD),.Y(I16286),.A(g10540));
  NOT NOT1_685(.VSS(VSS),.VDD(VDD),.Y(I7999),.A(g4114));
  NOT NOT1_686(.VSS(VSS),.VDD(VDD),.Y(g2854),.A(I5986));
  NOT NOT1_687(.VSS(VSS),.VDD(VDD),.Y(I17173),.A(g11293));
  NOT NOT1_688(.VSS(VSS),.VDD(VDD),.Y(I5946),.A(g2176));
  NOT NOT1_689(.VSS(VSS),.VDD(VDD),.Y(I10849),.A(g6734));
  NOT NOT1_690(.VSS(VSS),.VDD(VDD),.Y(g11341),.A(I17146));
  NOT NOT1_691(.VSS(VSS),.VDD(VDD),.Y(I7633),.A(g3474));
  NOT NOT1_692(.VSS(VSS),.VDD(VDD),.Y(g4889),.A(I8240));
  NOT NOT1_693(.VSS(VSS),.VDD(VDD),.Y(g2941),.A(I6118));
  NOT NOT1_694(.VSS(VSS),.VDD(VDD),.Y(g6248),.A(I10003));
  NOT NOT1_695(.VSS(VSS),.VDD(VDD),.Y(g11655),.A(I17767));
  NOT NOT1_696(.VSS(VSS),.VDD(VDD),.Y(g9258),.A(g8892));
  NOT NOT1_697(.VSS(VSS),.VDD(VDD),.Y(g3905),.A(g2920));
  NOT NOT1_698(.VSS(VSS),.VDD(VDD),.Y(g10892),.A(I16638));
  NOT NOT1_699(.VSS(VSS),.VDD(VDD),.Y(g9818),.A(I14955));
  NOT NOT1_700(.VSS(VSS),.VDD(VDD),.Y(g9352),.A(I14561));
  NOT NOT1_701(.VSS(VSS),.VDD(VDD),.Y(I7303),.A(g3262));
  NOT NOT1_702(.VSS(VSS),.VDD(VDD),.Y(I8293),.A(g4779));
  NOT NOT1_703(.VSS(VSS),.VDD(VDD),.Y(I10398),.A(g5820));
  NOT NOT1_704(.VSS(VSS),.VDD(VDD),.Y(I13475),.A(g8173));
  NOT NOT1_705(.VSS(VSS),.VDD(VDD),.Y(g11180),.A(I16941));
  NOT NOT1_706(.VSS(VSS),.VDD(VDD),.Y(g7826),.A(I12627));
  NOT NOT1_707(.VSS(VSS),.VDD(VDD),.Y(g3628),.A(g3111));
  NOT NOT1_708(.VSS(VSS),.VDD(VDD),.Y(g6255),.A(I10024));
  NOT NOT1_709(.VSS(VSS),.VDD(VDD),.Y(g4175),.A(I7342));
  NOT NOT1_710(.VSS(VSS),.VDD(VDD),.Y(g6081),.A(g4977));
  NOT NOT1_711(.VSS(VSS),.VDD(VDD),.Y(g6815),.A(I10855));
  NOT NOT1_712(.VSS(VSS),.VDD(VDD),.Y(I10141),.A(g5683));
  NOT NOT1_713(.VSS(VSS),.VDD(VDD),.Y(g4375),.A(g3638));
  NOT NOT1_714(.VSS(VSS),.VDD(VDD),.Y(I10804),.A(g6388));
  NOT NOT1_715(.VSS(VSS),.VDD(VDD),.Y(I5513),.A(g255));
  NOT NOT1_716(.VSS(VSS),.VDD(VDD),.Y(g3630),.A(I6789));
  NOT NOT1_717(.VSS(VSS),.VDD(VDD),.Y(g8788),.A(I14097));
  NOT NOT1_718(.VSS(VSS),.VDD(VDD),.Y(I11222),.A(g6533));
  NOT NOT1_719(.VSS(VSS),.VDD(VDD),.Y(I12282),.A(g7113));
  NOT NOT1_720(.VSS(VSS),.VDD(VDD),.Y(I15335),.A(g10007));
  NOT NOT1_721(.VSS(VSS),.VDD(VDD),.Y(I16601),.A(g10806));
  NOT NOT1_722(.VSS(VSS),.VDD(VDD),.Y(g5113),.A(I8503));
  NOT NOT1_723(.VSS(VSS),.VDD(VDD),.Y(g6692),.A(I10659));
  NOT NOT1_724(.VSS(VSS),.VDD(VDD),.Y(I16187),.A(g10492));
  NOT NOT1_725(.VSS(VSS),.VDD(VDD),.Y(g6097),.A(I9754));
  NOT NOT1_726(.VSS(VSS),.VDD(VDD),.Y(I7732),.A(g3758));
  NOT NOT1_727(.VSS(VSS),.VDD(VDD),.Y(g7910),.A(g7460));
  NOT NOT1_728(.VSS(VSS),.VDD(VDD),.Y(I12357),.A(g7147));
  NOT NOT1_729(.VSS(VSS),.VDD(VDD),.Y(g2219),.A(g94));
  NOT NOT1_730(.VSS(VSS),.VDD(VDD),.Y(g9893),.A(I15082));
  NOT NOT1_731(.VSS(VSS),.VDD(VDD),.Y(g2640),.A(g1984));
  NOT NOT1_732(.VSS(VSS),.VDD(VDD),.Y(g6154),.A(I9875));
  NOT NOT1_733(.VSS(VSS),.VDD(VDD),.Y(g4285),.A(g3688));
  NOT NOT1_734(.VSS(VSS),.VDD(VDD),.Y(g6354),.A(g5867));
  NOT NOT1_735(.VSS(VSS),.VDD(VDD),.Y(g2031),.A(g1690));
  NOT NOT1_736(.VSS(VSS),.VDD(VDD),.Y(g10907),.A(I16673));
  NOT NOT1_737(.VSS(VSS),.VDD(VDD),.Y(g5202),.A(g4640));
  NOT NOT1_738(.VSS(VSS),.VDD(VDD),.Y(g6960),.A(I11112));
  NOT NOT1_739(.VSS(VSS),.VDD(VDD),.Y(I15694),.A(g10234));
  NOT NOT1_740(.VSS(VSS),.VDD(VDD),.Y(I5378),.A(g1857));
  NOT NOT1_741(.VSS(VSS),.VDD(VDD),.Y(g2431),.A(I5510));
  NOT NOT1_742(.VSS(VSS),.VDD(VDD),.Y(I15965),.A(g10405));
  NOT NOT1_743(.VSS(VSS),.VDD(VDD),.Y(g2252),.A(I5271));
  NOT NOT1_744(.VSS(VSS),.VDD(VDD),.Y(g2812),.A(g2158));
  NOT NOT1_745(.VSS(VSS),.VDD(VDD),.Y(I7240),.A(g2824));
  NOT NOT1_746(.VSS(VSS),.VDD(VDD),.Y(g7609),.A(I12177));
  NOT NOT1_747(.VSS(VSS),.VDD(VDD),.Y(I10135),.A(g6249));
  NOT NOT1_748(.VSS(VSS),.VDD(VDD),.Y(g7308),.A(I11572));
  NOT NOT1_749(.VSS(VSS),.VDD(VDD),.Y(g8192),.A(I13117));
  NOT NOT1_750(.VSS(VSS),.VDD(VDD),.Y(g2958),.A(I6163));
  NOT NOT1_751(.VSS(VSS),.VDD(VDD),.Y(g8085),.A(g7932));
  NOT NOT1_752(.VSS(VSS),.VDD(VDD),.Y(g10074),.A(I15299));
  NOT NOT1_753(.VSS(VSS),.VDD(VDD),.Y(g5094),.A(I8462));
  NOT NOT1_754(.VSS(VSS),.VDD(VDD),.Y(I13347),.A(g8122));
  NOT NOT1_755(.VSS(VSS),.VDD(VDD),.Y(g2176),.A(g82));
  NOT NOT1_756(.VSS(VSS),.VDD(VDD),.Y(g9026),.A(I14415));
  NOT NOT1_757(.VSS(VSS),.VDD(VDD),.Y(g8485),.A(g8341));
  NOT NOT1_758(.VSS(VSS),.VDD(VDD),.Y(g4184),.A(I7369));
  NOT NOT1_759(.VSS(VSS),.VDD(VDD),.Y(g5494),.A(g4412));
  NOT NOT1_760(.VSS(VSS),.VDD(VDD),.Y(g3750),.A(I6941));
  NOT NOT1_761(.VSS(VSS),.VDD(VDD),.Y(g2005),.A(g928));
  NOT NOT1_762(.VSS(VSS),.VDD(VDD),.Y(g7883),.A(g7689));
  NOT NOT1_763(.VSS(VSS),.VDD(VDD),.Y(I7043),.A(g2908));
  NOT NOT1_764(.VSS(VSS),.VDD(VDD),.Y(g4384),.A(I7707));
  NOT NOT1_765(.VSS(VSS),.VDD(VDD),.Y(I9141),.A(g5402));
  NOT NOT1_766(.VSS(VSS),.VDD(VDD),.Y(I9860),.A(g5405));
  NOT NOT1_767(.VSS(VSS),.VDD(VDD),.Y(g5567),.A(I8982));
  NOT NOT1_768(.VSS(VSS),.VDD(VDD),.Y(g4339),.A(g4144));
  NOT NOT1_769(.VSS(VSS),.VDD(VDD),.Y(I9341),.A(g5013));
  NOT NOT1_770(.VSS(VSS),.VDD(VDD),.Y(g10238),.A(g10191));
  NOT NOT1_771(.VSS(VSS),.VDD(VDD),.Y(I16169),.A(g10448));
  NOT NOT1_772(.VSS(VSS),.VDD(VDD),.Y(I9525),.A(g5001));
  NOT NOT1_773(.VSS(VSS),.VDD(VDD),.Y(I14361),.A(g8951));
  NOT NOT1_774(.VSS(VSS),.VDD(VDD),.Y(g2829),.A(I5943));
  NOT NOT1_775(.VSS(VSS),.VDD(VDD),.Y(g11619),.A(I17675));
  NOT NOT1_776(.VSS(VSS),.VDD(VDD),.Y(g2765),.A(g2184));
  NOT NOT1_777(.VSS(VSS),.VDD(VDD),.Y(g9821),.A(I14964));
  NOT NOT1_778(.VSS(VSS),.VDD(VDD),.Y(g11502),.A(I17525));
  NOT NOT1_779(.VSS(VSS),.VDD(VDD),.Y(g7758),.A(I12439));
  NOT NOT1_780(.VSS(VSS),.VDD(VDD),.Y(I5916),.A(g2217));
  NOT NOT1_781(.VSS(VSS),.VDD(VDD),.Y(I13236),.A(g8245));
  NOT NOT1_782(.VSS(VSS),.VDD(VDD),.Y(g7066),.A(I11275));
  NOT NOT1_783(.VSS(VSS),.VDD(VDD),.Y(g7589),.A(I12099));
  NOT NOT1_784(.VSS(VSS),.VDD(VDD),.Y(g4424),.A(g3688));
  NOT NOT1_785(.VSS(VSS),.VDD(VDD),.Y(g3040),.A(g2135));
  NOT NOT1_786(.VSS(VSS),.VDD(VDD),.Y(g4737),.A(g3440));
  NOT NOT1_787(.VSS(VSS),.VDD(VDD),.Y(I11351),.A(g6698));
  NOT NOT1_788(.VSS(VSS),.VDD(VDD),.Y(I13952),.A(g8451));
  NOT NOT1_789(.VSS(VSS),.VDD(VDD),.Y(g5593),.A(I9013));
  NOT NOT1_790(.VSS(VSS),.VDD(VDD),.Y(g6112),.A(I9789));
  NOT NOT1_791(.VSS(VSS),.VDD(VDD),.Y(I13351),.A(g8214));
  NOT NOT1_792(.VSS(VSS),.VDD(VDD),.Y(g6218),.A(I9965));
  NOT NOT1_793(.VSS(VSS),.VDD(VDD),.Y(g6267),.A(I10060));
  NOT NOT1_794(.VSS(VSS),.VDD(VDD),.Y(g3440),.A(g3041));
  NOT NOT1_795(.VSS(VSS),.VDD(VDD),.Y(g6312),.A(I10195));
  NOT NOT1_796(.VSS(VSS),.VDD(VDD),.Y(g11618),.A(I17672));
  NOT NOT1_797(.VSS(VSS),.VDD(VDD),.Y(g9984),.A(I15184));
  NOT NOT1_798(.VSS(VSS),.VDD(VDD),.Y(I11821),.A(g7205));
  NOT NOT1_799(.VSS(VSS),.VDD(VDD),.Y(g10176),.A(I15520));
  NOT NOT1_800(.VSS(VSS),.VDD(VDD),.Y(g10185),.A(g10040));
  NOT NOT1_801(.VSS(VSS),.VDD(VDD),.Y(g10675),.A(g10574));
  NOT NOT1_802(.VSS(VSS),.VDD(VDD),.Y(I16479),.A(g10767));
  NOT NOT1_803(.VSS(VSS),.VDD(VDD),.Y(g10092),.A(I15323));
  NOT NOT1_804(.VSS(VSS),.VDD(VDD),.Y(I10048),.A(g5734));
  NOT NOT1_805(.VSS(VSS),.VDD(VDD),.Y(I16363),.A(g10599));
  NOT NOT1_806(.VSS(VSS),.VDD(VDD),.Y(I16217),.A(g10501));
  NOT NOT1_807(.VSS(VSS),.VDD(VDD),.Y(g3323),.A(g2157));
  NOT NOT1_808(.VSS(VSS),.VDD(VDD),.Y(I15278),.A(g10033));
  NOT NOT1_809(.VSS(VSS),.VDD(VDD),.Y(g7571),.A(I12035));
  NOT NOT1_810(.VSS(VSS),.VDD(VDD),.Y(g7365),.A(I11743));
  NOT NOT1_811(.VSS(VSS),.VDD(VDD),.Y(g2733),.A(I5795));
  NOT NOT1_812(.VSS(VSS),.VDD(VDD),.Y(g4077),.A(I7202));
  NOT NOT1_813(.VSS(VSS),.VDD(VDD),.Y(g6001),.A(I9625));
  NOT NOT1_814(.VSS(VSS),.VDD(VDD),.Y(g7048),.A(I11225));
  NOT NOT1_815(.VSS(VSS),.VDD(VDD),.Y(g10154),.A(I15458));
  NOT NOT1_816(.VSS(VSS),.VDD(VDD),.Y(g2270),.A(I5311));
  NOT NOT1_817(.VSS(VSS),.VDD(VDD),.Y(I5798),.A(g2085));
  NOT NOT1_818(.VSS(VSS),.VDD(VDD),.Y(I17240),.A(g11395));
  NOT NOT1_819(.VSS(VSS),.VDD(VDD),.Y(g7711),.A(I12344));
  NOT NOT1_820(.VSS(VSS),.VDD(VDD),.Y(g4523),.A(g3546));
  NOT NOT1_821(.VSS(VSS),.VDD(VDD),.Y(I10221),.A(g6117));
  NOT NOT1_822(.VSS(VSS),.VDD(VDD),.Y(I11790),.A(g7246));
  NOT NOT1_823(.VSS(VSS),.VDD(VDD),.Y(g8520),.A(I13729));
  NOT NOT1_824(.VSS(VSS),.VDD(VDD),.Y(g6293),.A(I10138));
  NOT NOT1_825(.VSS(VSS),.VDD(VDD),.Y(g11469),.A(I17444));
  NOT NOT1_826(.VSS(VSS),.VDD(VDD),.Y(g8219),.A(g7826));
  NOT NOT1_827(.VSS(VSS),.VDD(VDD),.Y(g2225),.A(I5210));
  NOT NOT1_828(.VSS(VSS),.VDD(VDD),.Y(g8640),.A(g8512));
  NOT NOT1_829(.VSS(VSS),.VDD(VDD),.Y(g10935),.A(g10827));
  NOT NOT1_830(.VSS(VSS),.VDD(VDD),.Y(g2610),.A(I5731));
  NOT NOT1_831(.VSS(VSS),.VDD(VDD),.Y(g2073),.A(I4879));
  NOT NOT1_832(.VSS(VSS),.VDD(VDD),.Y(g2796),.A(g2276));
  NOT NOT1_833(.VSS(VSS),.VDD(VDD),.Y(g11468),.A(I17441));
  NOT NOT1_834(.VSS(VSS),.VDD(VDD),.Y(g11039),.A(I16778));
  NOT NOT1_835(.VSS(VSS),.VDD(VDD),.Y(I6851),.A(g2937));
  NOT NOT1_836(.VSS(VSS),.VDD(VDD),.Y(g4205),.A(I7432));
  NOT NOT1_837(.VSS(VSS),.VDD(VDD),.Y(I7697),.A(g3743));
  NOT NOT1_838(.VSS(VSS),.VDD(VDD),.Y(I10613),.A(g6000));
  NOT NOT1_839(.VSS(VSS),.VDD(VDD),.Y(I11873),.A(g6863));
  NOT NOT1_840(.VSS(VSS),.VDD(VDD),.Y(g10883),.A(g10809));
  NOT NOT1_841(.VSS(VSS),.VDD(VDD),.Y(I17755),.A(g11646));
  NOT NOT1_842(.VSS(VSS),.VDD(VDD),.Y(g7333),.A(I11647));
  NOT NOT1_843(.VSS(VSS),.VDD(VDD),.Y(g9106),.A(I14439));
  NOT NOT1_844(.VSS(VSS),.VDD(VDD),.Y(I7210),.A(g2798));
  NOT NOT1_845(.VSS(VSS),.VDD(VDD),.Y(g7774),.A(I12487));
  NOT NOT1_846(.VSS(VSS),.VDD(VDD),.Y(g5521),.A(g4530));
  NOT NOT1_847(.VSS(VSS),.VDD(VDD),.Y(g3528),.A(g3164));
  NOT NOT1_848(.VSS(VSS),.VDD(VDD),.Y(g8958),.A(I14323));
  NOT NOT1_849(.VSS(VSS),.VDD(VDD),.Y(I16580),.A(g10826));
  NOT NOT1_850(.VSS(VSS),.VDD(VDD),.Y(I17770),.A(g11649));
  NOT NOT1_851(.VSS(VSS),.VDD(VDD),.Y(g11038),.A(I16775));
  NOT NOT1_852(.VSS(VSS),.VDD(VDD),.Y(g5050),.A(I8429));
  NOT NOT1_853(.VSS(VSS),.VDD(VDD),.Y(g2124),.A(I5050));
  NOT NOT1_854(.VSS(VSS),.VDD(VDD),.Y(g3351),.A(I6535));
  NOT NOT1_855(.VSS(VSS),.VDD(VDD),.Y(g5641),.A(I9084));
  NOT NOT1_856(.VSS(VSS),.VDD(VDD),.Y(I17563),.A(g11492));
  NOT NOT1_857(.VSS(VSS),.VDD(VDD),.Y(g2980),.A(g1983));
  NOT NOT1_858(.VSS(VSS),.VDD(VDD),.Y(g6727),.A(g5997));
  NOT NOT1_859(.VSS(VSS),.VDD(VDD),.Y(g8376),.A(I13478));
  NOT NOT1_860(.VSS(VSS),.VDD(VDD),.Y(I5632),.A(g932));
  NOT NOT1_861(.VSS(VSS),.VDD(VDD),.Y(I5095),.A(g37));
  NOT NOT1_862(.VSS(VSS),.VDD(VDD),.Y(I6260),.A(g2025));
  NOT NOT1_863(.VSS(VSS),.VDD(VDD),.Y(g2069),.A(I4869));
  NOT NOT1_864(.VSS(VSS),.VDD(VDD),.Y(I9111),.A(g5596));
  NOT NOT1_865(.VSS(VSS),.VDD(VDD),.Y(g7196),.A(I11420));
  NOT NOT1_866(.VSS(VSS),.VDD(VDD),.Y(g4551),.A(g3946));
  NOT NOT1_867(.VSS(VSS),.VDD(VDD),.Y(I15601),.A(g10173));
  NOT NOT1_868(.VSS(VSS),.VDD(VDD),.Y(I9311),.A(g4915));
  NOT NOT1_869(.VSS(VSS),.VDD(VDD),.Y(I15187),.A(g9968));
  NOT NOT1_870(.VSS(VSS),.VDD(VDD),.Y(g7803),.A(I12574));
  NOT NOT1_871(.VSS(VSS),.VDD(VDD),.Y(I12248),.A(g7098));
  NOT NOT1_872(.VSS(VSS),.VDD(VDD),.Y(I13209),.A(g8198));
  NOT NOT1_873(.VSS(VSS),.VDD(VDD),.Y(g4499),.A(g3546));
  NOT NOT1_874(.VSS(VSS),.VDD(VDD),.Y(I8848),.A(g4490));
  NOT NOT1_875(.VSS(VSS),.VDD(VDD),.Y(g2540),.A(I5655));
  NOT NOT1_876(.VSS(VSS),.VDD(VDD),.Y(g7538),.A(I11950));
  NOT NOT1_877(.VSS(VSS),.VDD(VDD),.Y(I13834),.A(g8488));
  NOT NOT1_878(.VSS(VSS),.VDD(VDD),.Y(I5579),.A(g1197));
  NOT NOT1_879(.VSS(VSS),.VDD(VDD),.Y(g7780),.A(I12505));
  NOT NOT1_880(.VSS(VSS),.VDD(VDD),.Y(g5724),.A(I9268));
  NOT NOT1_881(.VSS(VSS),.VDD(VDD),.Y(g9027),.A(I14418));
  NOT NOT1_882(.VSS(VSS),.VDD(VDD),.Y(g2206),.A(I5171));
  NOT NOT1_883(.VSS(VSS),.VDD(VDD),.Y(I12779),.A(g7608));
  NOT NOT1_884(.VSS(VSS),.VDD(VDD),.Y(g10729),.A(g10630));
  NOT NOT1_885(.VSS(VSS),.VDD(VDD),.Y(g6703),.A(I10678));
  NOT NOT1_886(.VSS(VSS),.VDD(VDD),.Y(I9174),.A(g4903));
  NOT NOT1_887(.VSS(VSS),.VDD(VDD),.Y(I5719),.A(g2072));
  NOT NOT1_888(.VSS(VSS),.VDD(VDD),.Y(g10577),.A(g10526));
  NOT NOT1_889(.VSS(VSS),.VDD(VDD),.Y(I17767),.A(g11648));
  NOT NOT1_890(.VSS(VSS),.VDD(VDD),.Y(g7509),.A(I11889));
  NOT NOT1_891(.VSS(VSS),.VDD(VDD),.Y(g9427),.A(g9079));
  NOT NOT1_892(.VSS(VSS),.VDD(VDD),.Y(I10033),.A(g5693));
  NOT NOT1_893(.VSS(VSS),.VDD(VDD),.Y(I7820),.A(g3811));
  NOT NOT1_894(.VSS(VSS),.VDD(VDD),.Y(I10234),.A(g6114));
  NOT NOT1_895(.VSS(VSS),.VDD(VDD),.Y(g4754),.A(g3440));
  NOT NOT1_896(.VSS(VSS),.VDD(VDD),.Y(I16531),.A(g10720));
  NOT NOT1_897(.VSS(VSS),.VDD(VDD),.Y(g10439),.A(g10334));
  NOT NOT1_898(.VSS(VSS),.VDD(VDD),.Y(I11021),.A(g6398));
  NOT NOT1_899(.VSS(VSS),.VDD(VDD),.Y(I12081),.A(g6934));
  NOT NOT1_900(.VSS(VSS),.VDD(VDD),.Y(g5878),.A(g5309));
  NOT NOT1_901(.VSS(VSS),.VDD(VDD),.Y(g6932),.A(I11058));
  NOT NOT1_902(.VSS(VSS),.VDD(VDD),.Y(g7662),.A(I12279));
  NOT NOT1_903(.VSS(VSS),.VDD(VDD),.Y(g4273),.A(g4013));
  NOT NOT1_904(.VSS(VSS),.VDD(VDD),.Y(I16178),.A(g10490));
  NOT NOT1_905(.VSS(VSS),.VDD(VDD),.Y(I12786),.A(g7622));
  NOT NOT1_906(.VSS(VSS),.VDD(VDD),.Y(I17633),.A(g11578));
  NOT NOT1_907(.VSS(VSS),.VDD(VDD),.Y(g5658),.A(I9135));
  NOT NOT1_908(.VSS(VSS),.VDD(VDD),.Y(g5777),.A(I9365));
  NOT NOT1_909(.VSS(VSS),.VDD(VDD),.Y(I10795),.A(g6123));
  NOT NOT1_910(.VSS(VSS),.VDD(VDD),.Y(I13726),.A(g8375));
  NOT NOT1_911(.VSS(VSS),.VDD(VDD),.Y(g7467),.A(g7148));
  NOT NOT1_912(.VSS(VSS),.VDD(VDD),.Y(g1990),.A(g774));
  NOT NOT1_913(.VSS(VSS),.VDD(VDD),.Y(I6118),.A(g2248));
  NOT NOT1_914(.VSS(VSS),.VDD(VDD),.Y(g8225),.A(g7826));
  NOT NOT1_915(.VSS(VSS),.VDD(VDD),.Y(I17191),.A(g11315));
  NOT NOT1_916(.VSS(VSS),.VDD(VDD),.Y(I17719),.A(g11623));
  NOT NOT1_917(.VSS(VSS),.VDD(VDD),.Y(I11614),.A(g6838));
  NOT NOT1_918(.VSS(VSS),.VDD(VDD),.Y(g8610),.A(g8483));
  NOT NOT1_919(.VSS(VSS),.VDD(VDD),.Y(I6367),.A(g2045));
  NOT NOT1_920(.VSS(VSS),.VDD(VDD),.Y(I9180),.A(g4905));
  NOT NOT1_921(.VSS(VSS),.VDD(VDD),.Y(I12647),.A(g7711));
  NOT NOT1_922(.VSS(VSS),.VDD(VDD),.Y(I16676),.A(g10798));
  NOT NOT1_923(.VSS(VSS),.VDD(VDD),.Y(I16685),.A(g10785));
  NOT NOT1_924(.VSS(VSS),.VDD(VDD),.Y(I11436),.A(g6488));
  NOT NOT1_925(.VSS(VSS),.VDD(VDD),.Y(I9380),.A(g5013));
  NOT NOT1_926(.VSS(VSS),.VDD(VDD),.Y(g10349),.A(I15811));
  NOT NOT1_927(.VSS(VSS),.VDD(VDD),.Y(g9345),.A(I14540));
  NOT NOT1_928(.VSS(VSS),.VDD(VDD),.Y(I16953),.A(g11082));
  NOT NOT1_929(.VSS(VSS),.VDD(VDD),.Y(I13436),.A(g8187));
  NOT NOT1_930(.VSS(VSS),.VDD(VDD),.Y(I9591),.A(g5095));
  NOT NOT1_931(.VSS(VSS),.VDD(VDD),.Y(I16373),.A(g10593));
  NOT NOT1_932(.VSS(VSS),.VDD(VDD),.Y(g4444),.A(I7800));
  NOT NOT1_933(.VSS(VSS),.VDD(VDD),.Y(g8473),.A(I13669));
  NOT NOT1_934(.VSS(VSS),.VDD(VDD),.Y(g2199),.A(g48));
  NOT NOT1_935(.VSS(VSS),.VDD(VDD),.Y(g11410),.A(I17271));
  NOT NOT1_936(.VSS(VSS),.VDD(VDD),.Y(g2399),.A(g605));
  NOT NOT1_937(.VSS(VSS),.VDD(VDD),.Y(g9763),.A(I14906));
  NOT NOT1_938(.VSS(VSS),.VDD(VDD),.Y(g7093),.A(I11326));
  NOT NOT1_939(.VSS(VSS),.VDD(VDD),.Y(I12999),.A(g7844));
  NOT NOT1_940(.VSS(VSS),.VDD(VDD),.Y(g3372),.A(g3121));
  NOT NOT1_941(.VSS(VSS),.VDD(VDD),.Y(I10514),.A(g6154));
  NOT NOT1_942(.VSS(VSS),.VDD(VDD),.Y(I12380),.A(g7204));
  NOT NOT1_943(.VSS(VSS),.VDD(VDD),.Y(g10906),.A(I16670));
  NOT NOT1_944(.VSS(VSS),.VDD(VDD),.Y(I15479),.A(g10091));
  NOT NOT1_945(.VSS(VSS),.VDD(VDD),.Y(I13320),.A(g8096));
  NOT NOT1_946(.VSS(VSS),.VDD(VDD),.Y(g10083),.A(I15311));
  NOT NOT1_947(.VSS(VSS),.VDD(VDD),.Y(I9020),.A(g4773));
  NOT NOT1_948(.VSS(VSS),.VDD(VDD),.Y(g8124),.A(g8011));
  NOT NOT1_949(.VSS(VSS),.VDD(VDD),.Y(g10284),.A(g10167));
  NOT NOT1_950(.VSS(VSS),.VDD(VDD),.Y(g7256),.A(I11489));
  NOT NOT1_951(.VSS(VSS),.VDD(VDD),.Y(g8980),.A(I14361));
  NOT NOT1_952(.VSS(VSS),.VDD(VDD),.Y(g7816),.A(I12613));
  NOT NOT1_953(.VSS(VSS),.VDD(VDD),.Y(g8324),.A(I13354));
  NOT NOT1_954(.VSS(VSS),.VDD(VDD),.Y(g11479),.A(I17470));
  NOT NOT1_955(.VSS(VSS),.VDD(VDD),.Y(I6193),.A(g2155));
  NOT NOT1_956(.VSS(VSS),.VDD(VDD),.Y(I11593),.A(g6830));
  NOT NOT1_957(.VSS(VSS),.VDD(VDD),.Y(g3143),.A(I6363));
  NOT NOT1_958(.VSS(VSS),.VDD(VDD),.Y(g11363),.A(I17188));
  NOT NOT1_959(.VSS(VSS),.VDD(VDD),.Y(g3343),.A(g2779));
  NOT NOT1_960(.VSS(VSS),.VDD(VDD),.Y(I11122),.A(g6450));
  NOT NOT1_961(.VSS(VSS),.VDD(VDD),.Y(g2797),.A(g2524));
  NOT NOT1_962(.VSS(VSS),.VDD(VDD),.Y(I13122),.A(g7966));
  NOT NOT1_963(.VSS(VSS),.VDD(VDD),.Y(I6549),.A(g2838));
  NOT NOT1_964(.VSS(VSS),.VDD(VDD),.Y(g4543),.A(g3946));
  NOT NOT1_965(.VSS(VSS),.VDD(VDD),.Y(I10421),.A(g5826));
  NOT NOT1_966(.VSS(VSS),.VDD(VDD),.Y(I11464),.A(g6443));
  NOT NOT1_967(.VSS(VSS),.VDD(VDD),.Y(g3566),.A(I6738));
  NOT NOT1_968(.VSS(VSS),.VDD(VDD),.Y(I6971),.A(g2882));
  NOT NOT1_969(.VSS(VSS),.VDD(VDD),.Y(g6716),.A(g5949));
  NOT NOT1_970(.VSS(VSS),.VDD(VDD),.Y(I14421),.A(g8944));
  NOT NOT1_971(.VSS(VSS),.VDD(VDD),.Y(g2245),.A(I5254));
  NOT NOT1_972(.VSS(VSS),.VDD(VDD),.Y(g6149),.A(I9866));
  NOT NOT1_973(.VSS(VSS),.VDD(VDD),.Y(g3988),.A(g3121));
  NOT NOT1_974(.VSS(VSS),.VDD(VDD),.Y(I6686),.A(g3015));
  NOT NOT1_975(.VSS(VSS),.VDD(VDD),.Y(g6349),.A(I10258));
  NOT NOT1_976(.VSS(VSS),.VDD(VDD),.Y(g7847),.A(I12638));
  NOT NOT1_977(.VSS(VSS),.VDD(VDD),.Y(g3693),.A(g2920));
  NOT NOT1_978(.VSS(VSS),.VDD(VDD),.Y(I11034),.A(g6629));
  NOT NOT1_979(.VSS(VSS),.VDD(VDD),.Y(I10012),.A(g5543));
  NOT NOT1_980(.VSS(VSS),.VDD(VDD),.Y(g3334),.A(I6517));
  NOT NOT1_981(.VSS(VSS),.VDD(VDD),.Y(I5725),.A(g2079));
  NOT NOT1_982(.VSS(VSS),.VDD(VDD),.Y(g7685),.A(g7148));
  NOT NOT1_983(.VSS(VSS),.VDD(VDD),.Y(g7197),.A(I11423));
  NOT NOT1_984(.VSS(VSS),.VDD(VDD),.Y(I11641),.A(g6960));
  NOT NOT1_985(.VSS(VSS),.VDD(VDD),.Y(I11797),.A(g6852));
  NOT NOT1_986(.VSS(VSS),.VDD(VDD),.Y(g5997),.A(I9617));
  NOT NOT1_987(.VSS(VSS),.VDD(VDD),.Y(I15580),.A(g10155));
  NOT NOT1_988(.VSS(VSS),.VDD(VDD),.Y(I13797),.A(g8473));
  NOT NOT1_989(.VSS(VSS),.VDD(VDD),.Y(I6598),.A(g2623));
  NOT NOT1_990(.VSS(VSS),.VDD(VDD),.Y(g7021),.A(I11162));
  NOT NOT1_991(.VSS(VSS),.VDD(VDD),.Y(g4729),.A(g3586));
  NOT NOT1_992(.VSS(VSS),.VDD(VDD),.Y(g4961),.A(I8333));
  NOT NOT1_993(.VSS(VSS),.VDD(VDD),.Y(g7421),.A(I11807));
  NOT NOT1_994(.VSS(VSS),.VDD(VDD),.Y(g10139),.A(I15415));
  NOT NOT1_995(.VSS(VSS),.VDD(VDD),.Y(g2344),.A(I5410));
  NOT NOT1_996(.VSS(VSS),.VDD(VDD),.Y(I8211),.A(g3566));
  NOT NOT1_997(.VSS(VSS),.VDD(VDD),.Y(I9905),.A(g5300));
  NOT NOT1_998(.VSS(VSS),.VDD(VDD),.Y(g6398),.A(I10302));
  NOT NOT1_999(.VSS(VSS),.VDD(VDD),.Y(I10541),.A(g6176));
  NOT NOT1_1000(.VSS(VSS),.VDD(VDD),.Y(I6121),.A(g2121));
  NOT NOT1_1001(.VSS(VSS),.VDD(VDD),.Y(g1963),.A(g110));
  NOT NOT1_1002(.VSS(VSS),.VDD(VDD),.Y(I17324),.A(g11347));
  NOT NOT1_1003(.VSS(VSS),.VDD(VDD),.Y(g7263),.A(I11498));
  NOT NOT1_1004(.VSS(VSS),.VDD(VDD),.Y(I14473),.A(g8921));
  NOT NOT1_1005(.VSS(VSS),.VDD(VDD),.Y(g2207),.A(I5174));
  NOT NOT1_1006(.VSS(VSS),.VDD(VDD),.Y(g10138),.A(I15412));
  NOT NOT1_1007(.VSS(VSS),.VDD(VDD),.Y(I17701),.A(g11617));
  NOT NOT1_1008(.VSS(VSS),.VDD(VDD),.Y(I10789),.A(g5867));
  NOT NOT1_1009(.VSS(VSS),.VDD(VDD),.Y(I12448),.A(g7530));
  NOT NOT1_1010(.VSS(VSS),.VDD(VDD),.Y(I13409),.A(g8141));
  NOT NOT1_1011(.VSS(VSS),.VDD(VDD),.Y(I17534),.A(g11495));
  NOT NOT1_1012(.VSS(VSS),.VDD(VDD),.Y(g3792),.A(I7017));
  NOT NOT1_1013(.VSS(VSS),.VDD(VDD),.Y(g5353),.A(I8820));
  NOT NOT1_1014(.VSS(VSS),.VDD(VDD),.Y(g8849),.A(g8745));
  NOT NOT1_1015(.VSS(VSS),.VDD(VDD),.Y(g2259),.A(I5292));
  NOT NOT1_1016(.VSS(VSS),.VDD(VDD),.Y(g6241),.A(I9992));
  NOT NOT1_1017(.VSS(VSS),.VDD(VDD),.Y(g2819),.A(g2159));
  NOT NOT1_1018(.VSS(VSS),.VDD(VDD),.Y(I11408),.A(g6405));
  NOT NOT1_1019(.VSS(VSS),.VDD(VDD),.Y(I12505),.A(g7728));
  NOT NOT1_1020(.VSS(VSS),.VDD(VDD),.Y(I11635),.A(g6947));
  NOT NOT1_1021(.VSS(VSS),.VDD(VDD),.Y(I10724),.A(g6096));
  NOT NOT1_1022(.VSS(VSS),.VDD(VDD),.Y(g11084),.A(I16863));
  NOT NOT1_1023(.VSS(VSS),.VDD(VDD),.Y(g4885),.A(I8228));
  NOT NOT1_1024(.VSS(VSS),.VDD(VDD),.Y(g4414),.A(I7752));
  NOT NOT1_1025(.VSS(VSS),.VDD(VDD),.Y(I10325),.A(g6003));
  NOT NOT1_1026(.VSS(VSS),.VDD(VDD),.Y(g11110),.A(g10974));
  NOT NOT1_1027(.VSS(VSS),.VDD(VDD),.Y(g3621),.A(I6754));
  NOT NOT1_1028(.VSS(VSS),.VDD(VDD),.Y(I6938),.A(g2854));
  NOT NOT1_1029(.VSS(VSS),.VDD(VDD),.Y(I7668),.A(g3733));
  NOT NOT1_1030(.VSS(VSS),.VDD(VDD),.Y(g2852),.A(I5982));
  NOT NOT1_1031(.VSS(VSS),.VDD(VDD),.Y(I7840),.A(g3431));
  NOT NOT1_1032(.VSS(VSS),.VDD(VDD),.Y(I16543),.A(g10747));
  NOT NOT1_1033(.VSS(VSS),.VDD(VDD),.Y(g10852),.A(g10740));
  NOT NOT1_1034(.VSS(VSS),.VDD(VDD),.Y(g8781),.A(I14080));
  NOT NOT1_1035(.VSS(VSS),.VDD(VDD),.Y(I8614),.A(g4414));
  NOT NOT1_1036(.VSS(VSS),.VDD(VDD),.Y(I10920),.A(g6733));
  NOT NOT1_1037(.VSS(VSS),.VDD(VDD),.Y(I10535),.A(g5867));
  NOT NOT1_1038(.VSS(VSS),.VDD(VDD),.Y(I12026),.A(g7119));
  NOT NOT1_1039(.VSS(VSS),.VDD(VDD),.Y(I10434),.A(g5843));
  NOT NOT1_1040(.VSS(VSS),.VDD(VDD),.Y(g11179),.A(I16938));
  NOT NOT1_1041(.VSS(VSS),.VDD(VDD),.Y(g2701),.A(g2040));
  NOT NOT1_1042(.VSS(VSS),.VDD(VDD),.Y(g3113),.A(I6343));
  NOT NOT1_1043(.VSS(VSS),.VDD(VDD),.Y(g7562),.A(g6984));
  NOT NOT1_1044(.VSS(VSS),.VDD(VDD),.Y(I14358),.A(g8950));
  NOT NOT1_1045(.VSS(VSS),.VDD(VDD),.Y(I7390),.A(g4087));
  NOT NOT1_1046(.VSS(VSS),.VDD(VDD),.Y(I10828),.A(g6708));
  NOT NOT1_1047(.VSS(VSS),.VDD(VDD),.Y(I10946),.A(g6548));
  NOT NOT1_1048(.VSS(VSS),.VDD(VDD),.Y(g8797),.A(I14116));
  NOT NOT1_1049(.VSS(VSS),.VDD(VDD),.Y(g6644),.A(I10601));
  NOT NOT1_1050(.VSS(VSS),.VDD(VDD),.Y(g4513),.A(g3546));
  NOT NOT1_1051(.VSS(VSS),.VDD(VDD),.Y(g7631),.A(I12235));
  NOT NOT1_1052(.VSS(VSS),.VDD(VDD),.Y(I5171),.A(g1419));
  NOT NOT1_1053(.VSS(VSS),.VDD(VDD),.Y(g7723),.A(I12354));
  NOT NOT1_1054(.VSS(VSS),.VDD(VDD),.Y(g6119),.A(I9810));
  NOT NOT1_1055(.VSS(VSS),.VDD(VDD),.Y(I9973),.A(g5502));
  NOT NOT1_1056(.VSS(VSS),.VDD(VDD),.Y(g7817),.A(I12616));
  NOT NOT1_1057(.VSS(VSS),.VDD(VDD),.Y(g5901),.A(g5361));
  NOT NOT1_1058(.VSS(VSS),.VDD(VDD),.Y(I4920),.A(g260));
  NOT NOT1_1059(.VSS(VSS),.VDD(VDD),.Y(g8291),.A(I13227));
  NOT NOT1_1060(.VSS(VSS),.VDD(VDD),.Y(g11373),.A(I17198));
  NOT NOT1_1061(.VSS(VSS),.VDD(VDD),.Y(g3094),.A(I6302));
  NOT NOT1_1062(.VSS(VSS),.VDD(VDD),.Y(g6258),.A(I10033));
  NOT NOT1_1063(.VSS(VSS),.VDD(VDD),.Y(g4178),.A(I7351));
  NOT NOT1_1064(.VSS(VSS),.VDD(VDD),.Y(g4436),.A(g3638));
  NOT NOT1_1065(.VSS(VSS),.VDD(VDD),.Y(g6818),.A(I10864));
  NOT NOT1_1066(.VSS(VSS),.VDD(VDD),.Y(g4679),.A(g4013));
  NOT NOT1_1067(.VSS(VSS),.VDD(VDD),.Y(g11654),.A(I17764));
  NOT NOT1_1068(.VSS(VSS),.VDD(VDD),.Y(g4378),.A(I7697));
  NOT NOT1_1069(.VSS(VSS),.VDD(VDD),.Y(g7605),.A(I12165));
  NOT NOT1_1070(.VSS(VSS),.VDD(VDD),.Y(g5511),.A(I8934));
  NOT NOT1_1071(.VSS(VSS),.VDD(VDD),.Y(I11575),.A(g6823));
  NOT NOT1_1072(.VSS(VSS),.VDD(VDD),.Y(g3518),.A(g3164));
  NOT NOT1_1073(.VSS(VSS),.VDD(VDD),.Y(I10682),.A(g6051));
  NOT NOT1_1074(.VSS(VSS),.VDD(VDD),.Y(g10576),.A(g10524));
  NOT NOT1_1075(.VSS(VSS),.VDD(VDD),.Y(I9040),.A(g4794));
  NOT NOT1_1076(.VSS(VSS),.VDD(VDD),.Y(g8144),.A(I13027));
  NOT NOT1_1077(.VSS(VSS),.VDD(VDD),.Y(g8344),.A(I13412));
  NOT NOT1_1078(.VSS(VSS),.VDD(VDD),.Y(g6717),.A(I10706));
  NOT NOT1_1079(.VSS(VSS),.VDD(VDD),.Y(I9440),.A(g5078));
  NOT NOT1_1080(.VSS(VSS),.VDD(VDD),.Y(g11417),.A(I17302));
  NOT NOT1_1081(.VSS(VSS),.VDD(VDD),.Y(I13711),.A(g8342));
  NOT NOT1_1082(.VSS(VSS),.VDD(VDD),.Y(I16814),.A(g10910));
  NOT NOT1_1083(.VSS(VSS),.VDD(VDD),.Y(I12433),.A(g7657));
  NOT NOT1_1084(.VSS(VSS),.VDD(VDD),.Y(g4335),.A(I7612));
  NOT NOT1_1085(.VSS(VSS),.VDD(VDD),.Y(I9123),.A(g4890));
  NOT NOT1_1086(.VSS(VSS),.VDD(VDD),.Y(I11109),.A(g6464));
  NOT NOT1_1087(.VSS(VSS),.VDD(VDD),.Y(g7751),.A(I12418));
  NOT NOT1_1088(.VSS(VSS),.VDD(VDD),.Y(g4182),.A(I7363));
  NOT NOT1_1089(.VSS(VSS),.VDD(VDD),.Y(I9323),.A(g5620));
  NOT NOT1_1090(.VSS(VSS),.VDD(VDD),.Y(I13109),.A(g7981));
  NOT NOT1_1091(.VSS(VSS),.VDD(VDD),.Y(g4288),.A(g4130));
  NOT NOT1_1092(.VSS(VSS),.VDD(VDD),.Y(I11537),.A(g7144));
  NOT NOT1_1093(.VSS(VSS),.VDD(VDD),.Y(g4382),.A(g3638));
  NOT NOT1_1094(.VSS(VSS),.VDD(VDD),.Y(I16772),.A(g10887));
  NOT NOT1_1095(.VSS(VSS),.VDD(VDD),.Y(g3776),.A(g2579));
  NOT NOT1_1096(.VSS(VSS),.VDD(VDD),.Y(g6893),.A(I10991));
  NOT NOT1_1097(.VSS(VSS),.VDD(VDD),.Y(g5574),.A(g4300));
  NOT NOT1_1098(.VSS(VSS),.VDD(VDD),.Y(g5864),.A(I9483));
  NOT NOT1_1099(.VSS(VSS),.VDD(VDD),.Y(g10200),.A(g10169));
  NOT NOT1_1100(.VSS(VSS),.VDD(VDD),.Y(g8694),.A(I13975));
  NOT NOT1_1101(.VSS(VSS),.VDD(VDD),.Y(g2825),.A(I5935));
  NOT NOT1_1102(.VSS(VSS),.VDD(VDD),.Y(g2650),.A(g2006));
  NOT NOT1_1103(.VSS(VSS),.VDD(VDD),.Y(g10608),.A(I16283));
  NOT NOT1_1104(.VSS(VSS),.VDD(VDD),.Y(g10115),.A(I15353));
  NOT NOT1_1105(.VSS(VSS),.VDD(VDD),.Y(g6386),.A(I10282));
  NOT NOT1_1106(.VSS(VSS),.VDD(VDD),.Y(g7585),.A(I12081));
  NOT NOT1_1107(.VSS(VSS),.VDD(VDD),.Y(I17447),.A(g11457));
  NOT NOT1_1108(.VSS(VSS),.VDD(VDD),.Y(I5684),.A(g572));
  NOT NOT1_1109(.VSS(VSS),.VDD(VDD),.Y(I8061),.A(g3381));
  NOT NOT1_1110(.VSS(VSS),.VDD(VDD),.Y(g4805),.A(g3337));
  NOT NOT1_1111(.VSS(VSS),.VDD(VDD),.Y(I7163),.A(g2643));
  NOT NOT1_1112(.VSS(VSS),.VDD(VDD),.Y(I5963),.A(g2179));
  NOT NOT1_1113(.VSS(VSS),.VDD(VDD),.Y(I7810),.A(g3799));
  NOT NOT1_1114(.VSS(VSS),.VDD(VDD),.Y(g7041),.A(g6427));
  NOT NOT1_1115(.VSS(VSS),.VDD(VDD),.Y(I7363),.A(g4005));
  NOT NOT1_1116(.VSS(VSS),.VDD(VDD),.Y(I16638),.A(g10863));
  NOT NOT1_1117(.VSS(VSS),.VDD(VDD),.Y(g2008),.A(g971));
  NOT NOT1_1118(.VSS(VSS),.VDD(VDD),.Y(I13606),.A(g8311));
  NOT NOT1_1119(.VSS(VSS),.VDD(VDD),.Y(I12971),.A(g8039));
  NOT NOT1_1120(.VSS(VSS),.VDD(VDD),.Y(I11303),.A(g6526));
  NOT NOT1_1121(.VSS(VSS),.VDD(VDD),.Y(g6274),.A(I10081));
  NOT NOT1_1122(.VSS(VSS),.VDD(VDD),.Y(I7432),.A(g3663));
  NOT NOT1_1123(.VSS(VSS),.VDD(VDD),.Y(g6426),.A(I10340));
  NOT NOT1_1124(.VSS(VSS),.VDD(VDD),.Y(g11423),.A(I17324));
  NOT NOT1_1125(.VSS(VSS),.VDD(VDD),.Y(g2336),.A(g1900));
  NOT NOT1_1126(.VSS(VSS),.VDD(VDD),.Y(I16416),.A(g10664));
  NOT NOT1_1127(.VSS(VSS),.VDD(VDD),.Y(I12369),.A(g7189));
  NOT NOT1_1128(.VSS(VSS),.VDD(VDD),.Y(I9875),.A(g5278));
  NOT NOT1_1129(.VSS(VSS),.VDD(VDD),.Y(I7453),.A(g3708));
  NOT NOT1_1130(.VSS(VSS),.VDD(VDD),.Y(g6170),.A(g5426));
  NOT NOT1_1131(.VSS(VSS),.VDD(VDD),.Y(I14506),.A(g8923));
  NOT NOT1_1132(.VSS(VSS),.VDD(VDD),.Y(g7673),.A(I12296));
  NOT NOT1_1133(.VSS(VSS),.VDD(VDD),.Y(I9655),.A(g5173));
  NOT NOT1_1134(.VSS(VSS),.VDD(VDD),.Y(g6125),.A(I9822));
  NOT NOT1_1135(.VSS(VSS),.VDD(VDD),.Y(I5707),.A(g2418));
  NOT NOT1_1136(.VSS(VSS),.VDD(VDD),.Y(g8886),.A(I14228));
  NOT NOT1_1137(.VSS(VSS),.VDD(VDD),.Y(g3521),.A(g3164));
  NOT NOT1_1138(.VSS(VSS),.VDD(VDD),.Y(g8951),.A(I14306));
  NOT NOT1_1139(.VSS(VSS),.VDD(VDD),.Y(I16510),.A(g10712));
  NOT NOT1_1140(.VSS(VSS),.VDD(VDD),.Y(g5262),.A(g4353));
  NOT NOT1_1141(.VSS(VSS),.VDD(VDD),.Y(g3050),.A(I6260));
  NOT NOT1_1142(.VSS(VSS),.VDD(VDD),.Y(I11091),.A(g6657));
  NOT NOT1_1143(.VSS(VSS),.VDD(VDD),.Y(g10973),.A(I16720));
  NOT NOT1_1144(.VSS(VSS),.VDD(VDD),.Y(g5736),.A(I9296));
  NOT NOT1_1145(.VSS(VSS),.VDD(VDD),.Y(g6984),.A(g6382));
  NOT NOT1_1146(.VSS(VSS),.VDD(VDD),.Y(g6280),.A(I10099));
  NOT NOT1_1147(.VSS(VSS),.VDD(VDD),.Y(g6939),.A(I11071));
  NOT NOT1_1148(.VSS(VSS),.VDD(VDD),.Y(g7669),.A(I12286));
  NOT NOT1_1149(.VSS(VSS),.VDD(VDD),.Y(I17246),.A(g11341));
  NOT NOT1_1150(.VSS(VSS),.VDD(VDD),.Y(g11543),.A(g11519));
  NOT NOT1_1151(.VSS(VSS),.VDD(VDD),.Y(g3996),.A(g3144));
  NOT NOT1_1152(.VSS(VSS),.VDD(VDD),.Y(g10184),.A(g10039));
  NOT NOT1_1153(.VSS(VSS),.VDD(VDD),.Y(I12412),.A(g7520));
  NOT NOT1_1154(.VSS(VSS),.VDD(VDD),.Y(I8403),.A(g4264));
  NOT NOT1_1155(.VSS(VSS),.VDD(VDD),.Y(g10674),.A(g10584));
  NOT NOT1_1156(.VSS(VSS),.VDD(VDD),.Y(g8314),.A(I13326));
  NOT NOT1_1157(.VSS(VSS),.VDD(VDD),.Y(g5623),.A(I9053));
  NOT NOT1_1158(.VSS(VSS),.VDD(VDD),.Y(g7772),.A(I12481));
  NOT NOT1_1159(.VSS(VSS),.VDD(VDD),.Y(I7157),.A(g3015));
  NOT NOT1_1160(.VSS(VSS),.VDD(VDD),.Y(g7058),.A(I11255));
  NOT NOT1_1161(.VSS(VSS),.VDD(VDD),.Y(I12133),.A(g6870));
  NOT NOT1_1162(.VSS(VSS),.VDD(VDD),.Y(I5957),.A(g2178));
  NOT NOT1_1163(.VSS(VSS),.VDD(VDD),.Y(I7357),.A(g4077));
  NOT NOT1_1164(.VSS(VSS),.VDD(VDD),.Y(g2122),.A(I5044));
  NOT NOT1_1165(.VSS(VSS),.VDD(VDD),.Y(g2228),.A(g28));
  NOT NOT1_1166(.VSS(VSS),.VDD(VDD),.Y(g7531),.A(I11929));
  NOT NOT1_1167(.VSS(VSS),.VDD(VDD),.Y(g4095),.A(I7233));
  NOT NOT1_1168(.VSS(VSS),.VDD(VDD),.Y(g9554),.A(I14697));
  NOT NOT1_1169(.VSS(VSS),.VDD(VDD),.Y(g8870),.A(I14182));
  NOT NOT1_1170(.VSS(VSS),.VDD(VDD),.Y(g2322),.A(I5378));
  NOT NOT1_1171(.VSS(VSS),.VDD(VDD),.Y(I10927),.A(g6755));
  NOT NOT1_1172(.VSS(VSS),.VDD(VDD),.Y(g7458),.A(g7123));
  NOT NOT1_1173(.VSS(VSS),.VDD(VDD),.Y(g5889),.A(I9514));
  NOT NOT1_1174(.VSS(VSS),.VDD(VDD),.Y(I12229),.A(g7070));
  NOT NOT1_1175(.VSS(VSS),.VDD(VDD),.Y(I6962),.A(g2791));
  NOT NOT1_1176(.VSS(VSS),.VDD(VDD),.Y(g4495),.A(I7886));
  NOT NOT1_1177(.VSS(VSS),.VDD(VDD),.Y(I9839),.A(g5226));
  NOT NOT1_1178(.VSS(VSS),.VDD(VDD),.Y(g2230),.A(g704));
  NOT NOT1_1179(.VSS(VSS),.VDD(VDD),.Y(g4437),.A(g3345));
  NOT NOT1_1180(.VSS(VSS),.VDD(VDD),.Y(g4102),.A(I7244));
  NOT NOT1_1181(.VSS(VSS),.VDD(VDD),.Y(I17591),.A(g11514));
  NOT NOT1_1182(.VSS(VSS),.VDD(VDD),.Y(g4208),.A(I7441));
  NOT NOT1_1183(.VSS(VSS),.VDD(VDD),.Y(g7890),.A(g7479));
  NOT NOT1_1184(.VSS(VSS),.VDD(VDD),.Y(g8650),.A(I13933));
  NOT NOT1_1185(.VSS(VSS),.VDD(VDD),.Y(I13840),.A(g8488));
  NOT NOT1_1186(.VSS(VSS),.VDD(VDD),.Y(I16586),.A(g10850));
  NOT NOT1_1187(.VSS(VSS),.VDD(VDD),.Y(g3379),.A(g3121));
  NOT NOT1_1188(.VSS(VSS),.VDD(VDD),.Y(I15568),.A(g10094));
  NOT NOT1_1189(.VSS(VSS),.VDD(VDD),.Y(g10934),.A(g10827));
  NOT NOT1_1190(.VSS(VSS),.VDD(VDD),.Y(g6106),.A(I9773));
  NOT NOT1_1191(.VSS(VSS),.VDD(VDD),.Y(g5175),.A(g4682));
  NOT NOT1_1192(.VSS(VSS),.VDD(VDD),.Y(g6306),.A(I10177));
  NOT NOT1_1193(.VSS(VSS),.VDD(VDD),.Y(g7505),.A(g7148));
  NOT NOT1_1194(.VSS(VSS),.VDD(VDD),.Y(g3878),.A(g2920));
  NOT NOT1_1195(.VSS(VSS),.VDD(VDD),.Y(g11242),.A(g11112));
  NOT NOT1_1196(.VSS(VSS),.VDD(VDD),.Y(I5098),.A(g38));
  NOT NOT1_1197(.VSS(VSS),.VDD(VDD),.Y(g8008),.A(I12846));
  NOT NOT1_1198(.VSS(VSS),.VDD(VDD),.Y(I10240),.A(g5937));
  NOT NOT1_1199(.VSS(VSS),.VDD(VDD),.Y(g7011),.A(g6503));
  NOT NOT1_1200(.VSS(VSS),.VDD(VDD),.Y(g4719),.A(g3586));
  NOT NOT1_1201(.VSS(VSS),.VDD(VDD),.Y(g10692),.A(I16363));
  NOT NOT1_1202(.VSS(VSS),.VDD(VDD),.Y(g5651),.A(I9114));
  NOT NOT1_1203(.VSS(VSS),.VDD(VDD),.Y(I6587),.A(g2620));
  NOT NOT1_1204(.VSS(VSS),.VDD(VDD),.Y(I10648),.A(g6030));
  NOT NOT1_1205(.VSS(VSS),.VDD(VDD),.Y(I15814),.A(g10202));
  NOT NOT1_1206(.VSS(VSS),.VDD(VDD),.Y(g8336),.A(I13388));
  NOT NOT1_1207(.VSS(VSS),.VDD(VDD),.Y(I14903),.A(g9507));
  NOT NOT1_1208(.VSS(VSS),.VDD(VDD),.Y(I5833),.A(g2103));
  NOT NOT1_1209(.VSS(VSS),.VDD(VDD),.Y(g6387),.A(g6121));
  NOT NOT1_1210(.VSS(VSS),.VDD(VDD),.Y(g5285),.A(g4355));
  NOT NOT1_1211(.VSS(VSS),.VDD(VDD),.Y(g6461),.A(I10391));
  NOT NOT1_1212(.VSS(VSS),.VDD(VDD),.Y(I15807),.A(g10284));
  NOT NOT1_1213(.VSS(VSS),.VDD(VDD),.Y(I15974),.A(g10411));
  NOT NOT1_1214(.VSS(VSS),.VDD(VDD),.Y(I8858),.A(g4506));
  NOT NOT1_1215(.VSS(VSS),.VDD(VDD),.Y(g2550),.A(g1834));
  NOT NOT1_1216(.VSS(VSS),.VDD(VDD),.Y(g7074),.A(I11299));
  NOT NOT1_1217(.VSS(VSS),.VDD(VDD),.Y(I16720),.A(g10854));
  NOT NOT1_1218(.VSS(VSS),.VDD(VDD),.Y(g3271),.A(I6443));
  NOT NOT1_1219(.VSS(VSS),.VDD(VDD),.Y(g10400),.A(g10348));
  NOT NOT1_1220(.VSS(VSS),.VDD(VDD),.Y(g2845),.A(g2168));
  NOT NOT1_1221(.VSS(VSS),.VDD(VDD),.Y(I9282),.A(g5633));
  NOT NOT1_1222(.VSS(VSS),.VDD(VDD),.Y(I15639),.A(g10179));
  NOT NOT1_1223(.VSS(VSS),.VDD(VDD),.Y(I10563),.A(g6043));
  NOT NOT1_1224(.VSS(VSS),.VDD(VDD),.Y(I5584),.A(g1200));
  NOT NOT1_1225(.VSS(VSS),.VDD(VDD),.Y(g10214),.A(I15586));
  NOT NOT1_1226(.VSS(VSS),.VDD(VDD),.Y(g9490),.A(g9324));
  NOT NOT1_1227(.VSS(VSS),.VDD(VDD),.Y(g9823),.A(I14970));
  NOT NOT1_1228(.VSS(VSS),.VDD(VDD),.Y(g2195),.A(g83));
  NOT NOT1_1229(.VSS(VSS),.VDD(VDD),.Y(g4265),.A(g3664));
  NOT NOT1_1230(.VSS(VSS),.VDD(VDD),.Y(I15293),.A(g10001));
  NOT NOT1_1231(.VSS(VSS),.VDD(VDD),.Y(I9988),.A(g5526));
  NOT NOT1_1232(.VSS(VSS),.VDD(VDD),.Y(g6427),.A(I10343));
  NOT NOT1_1233(.VSS(VSS),.VDD(VDD),.Y(I12627),.A(g7697));
  NOT NOT1_1234(.VSS(VSS),.VDD(VDD),.Y(g2395),.A(g231));
  NOT NOT1_1235(.VSS(VSS),.VDD(VDD),.Y(g2891),.A(I6055));
  NOT NOT1_1236(.VSS(VSS),.VDD(VDD),.Y(g5184),.A(g4682));
  NOT NOT1_1237(.VSS(VSS),.VDD(VDD),.Y(g2337),.A(I5395));
  NOT NOT1_1238(.VSS(VSS),.VDD(VDD),.Y(I11483),.A(g6567));
  NOT NOT1_1239(.VSS(VSS),.VDD(VDD),.Y(g2913),.A(I6088));
  NOT NOT1_1240(.VSS(VSS),.VDD(VDD),.Y(g10329),.A(I15775));
  NOT NOT1_1241(.VSS(VSS),.VDD(VDD),.Y(g10207),.A(g10186));
  NOT NOT1_1242(.VSS(VSS),.VDD(VDD),.Y(g4442),.A(g3638));
  NOT NOT1_1243(.VSS(VSS),.VDD(VDD),.Y(I6985),.A(g2890));
  NOT NOT1_1244(.VSS(VSS),.VDD(VDD),.Y(g6904),.A(I11008));
  NOT NOT1_1245(.VSS(VSS),.VDD(VDD),.Y(g6200),.A(I9935));
  NOT NOT1_1246(.VSS(VSS),.VDD(VDD),.Y(g11638),.A(I17724));
  NOT NOT1_1247(.VSS(VSS),.VDD(VDD),.Y(g10539),.A(I16184));
  NOT NOT1_1248(.VSS(VSS),.VDD(VDD),.Y(g4786),.A(I8154));
  NOT NOT1_1249(.VSS(VSS),.VDD(VDD),.Y(g6046),.A(I9669));
  NOT NOT1_1250(.VSS(VSS),.VDD(VDD),.Y(g8065),.A(I12913));
  NOT NOT1_1251(.VSS(VSS),.VDD(VDD),.Y(g3799),.A(I7022));
  NOT NOT1_1252(.VSS(VSS),.VDD(VDD),.Y(I8315),.A(g4788));
  NOT NOT1_1253(.VSS(VSS),.VDD(VDD),.Y(I8811),.A(g4465));
  NOT NOT1_1254(.VSS(VSS),.VDD(VDD),.Y(g6446),.A(I10370));
  NOT NOT1_1255(.VSS(VSS),.VDD(VDD),.Y(g8122),.A(I12981));
  NOT NOT1_1256(.VSS(VSS),.VDD(VDD),.Y(g3981),.A(I7118));
  NOT NOT1_1257(.VSS(VSS),.VDD(VDD),.Y(g8465),.A(g8289));
  NOT NOT1_1258(.VSS(VSS),.VDD(VDD),.Y(g9529),.A(I14672));
  NOT NOT1_1259(.VSS(VSS),.VDD(VDD),.Y(g4164),.A(I7311));
  NOT NOT1_1260(.VSS(VSS),.VDD(VDD),.Y(g10538),.A(I16181));
  NOT NOT1_1261(.VSS(VSS),.VDD(VDD),.Y(g4233),.A(g3698));
  NOT NOT1_1262(.VSS(VSS),.VDD(VDD),.Y(g5424),.A(I8865));
  NOT NOT1_1263(.VSS(VSS),.VDD(VDD),.Y(g9348),.A(I14549));
  NOT NOT1_1264(.VSS(VSS),.VDD(VDD),.Y(I11326),.A(g6660));
  NOT NOT1_1265(.VSS(VSS),.VDD(VDD),.Y(I13949),.A(g8451));
  NOT NOT1_1266(.VSS(VSS),.VDD(VDD),.Y(g6403),.A(g6128));
  NOT NOT1_1267(.VSS(VSS),.VDD(VDD),.Y(I13326),.A(g8203));
  NOT NOT1_1268(.VSS(VSS),.VDD(VDD),.Y(I9804),.A(g5417));
  NOT NOT1_1269(.VSS(VSS),.VDD(VDD),.Y(g6145),.A(I9860));
  NOT NOT1_1270(.VSS(VSS),.VDD(VDD),.Y(g2859),.A(I5995));
  NOT NOT1_1271(.VSS(VSS),.VDD(VDD),.Y(g3997),.A(I7131));
  NOT NOT1_1272(.VSS(VSS),.VDD(VDD),.Y(I15510),.A(g10035));
  NOT NOT1_1273(.VSS(VSS),.VDD(VDD),.Y(g9355),.A(I14570));
  NOT NOT1_1274(.VSS(VSS),.VDD(VDD),.Y(I9792),.A(g5403));
  NOT NOT1_1275(.VSS(VSS),.VDD(VDD),.Y(I6832),.A(g2909));
  NOT NOT1_1276(.VSS(VSS),.VDD(VDD),.Y(g4454),.A(g3914));
  NOT NOT1_1277(.VSS(VSS),.VDD(VDD),.Y(g8033),.A(I12875));
  NOT NOT1_1278(.VSS(VSS),.VDD(VDD),.Y(g11510),.A(I17549));
  NOT NOT1_1279(.VSS(VSS),.VDD(VDD),.Y(g6191),.A(g5446));
  NOT NOT1_1280(.VSS(VSS),.VDD(VDD),.Y(g7569),.A(I12029));
  NOT NOT1_1281(.VSS(VSS),.VDD(VDD),.Y(g5672),.A(I9177));
  NOT NOT1_1282(.VSS(VSS),.VDD(VDD),.Y(g4296),.A(I7559));
  NOT NOT1_1283(.VSS(VSS),.VDD(VDD),.Y(I11904),.A(g6902));
  NOT NOT1_1284(.VSS(VSS),.VDD(VDD),.Y(I10633),.A(g6015));
  NOT NOT1_1285(.VSS(VSS),.VDD(VDD),.Y(I10898),.A(g6735));
  NOT NOT1_1286(.VSS(VSS),.VDD(VDD),.Y(g5231),.A(g4640));
  NOT NOT1_1287(.VSS(VSS),.VDD(VDD),.Y(I17318),.A(g11340));
  NOT NOT1_1288(.VSS(VSS),.VDD(VDD),.Y(g3332),.A(I6513));
  NOT NOT1_1289(.VSS(VSS),.VDD(VDD),.Y(I11252),.A(g6542));
  NOT NOT1_1290(.VSS(VSS),.VDD(VDD),.Y(g10241),.A(g10192));
  NOT NOT1_1291(.VSS(VSS),.VDD(VDD),.Y(g9260),.A(g8892));
  NOT NOT1_1292(.VSS(VSS),.VDD(VDD),.Y(g6695),.A(I10666));
  NOT NOT1_1293(.VSS(VSS),.VDD(VDD),.Y(I10719),.A(g6003));
  NOT NOT1_1294(.VSS(VSS),.VDD(VDD),.Y(I13621),.A(g8315));
  NOT NOT1_1295(.VSS(VSS),.VDD(VDD),.Y(g5643),.A(I9090));
  NOT NOT1_1296(.VSS(VSS),.VDD(VDD),.Y(g3353),.A(g3121));
  NOT NOT1_1297(.VSS(VSS),.VDD(VDD),.Y(I7735),.A(g3759));
  NOT NOT1_1298(.VSS(VSS),.VDD(VDD),.Y(I6507),.A(g2808));
  NOT NOT1_1299(.VSS(VSS),.VDD(VDD),.Y(I14191),.A(g8795));
  NOT NOT1_1300(.VSS(VSS),.VDD(VDD),.Y(g8096),.A(I12953));
  NOT NOT1_1301(.VSS(VSS),.VDD(VDD),.Y(g2248),.A(g99));
  NOT NOT1_1302(.VSS(VSS),.VDD(VDD),.Y(g11578),.A(I17616));
  NOT NOT1_1303(.VSS(VSS),.VDD(VDD),.Y(g2342),.A(I5406));
  NOT NOT1_1304(.VSS(VSS),.VDD(VDD),.Y(I7782),.A(g3775));
  NOT NOT1_1305(.VSS(VSS),.VDD(VDD),.Y(g6107),.A(I9776));
  NOT NOT1_1306(.VSS(VSS),.VDD(VDD),.Y(I17540),.A(g11498));
  NOT NOT1_1307(.VSS(VSS),.VDD(VDD),.Y(I12857),.A(g7638));
  NOT NOT1_1308(.VSS(VSS),.VDD(VDD),.Y(g11014),.A(I16735));
  NOT NOT1_1309(.VSS(VSS),.VDD(VDD),.Y(g6307),.A(I10180));
  NOT NOT1_1310(.VSS(VSS),.VDD(VDD),.Y(g3744),.A(g3307));
  NOT NOT1_1311(.VSS(VSS),.VDD(VDD),.Y(g6536),.A(I10456));
  NOT NOT1_1312(.VSS(VSS),.VDD(VDD),.Y(I4883),.A(g581));
  NOT NOT1_1313(.VSS(VSS),.VDD(VDD),.Y(g5205),.A(g4366));
  NOT NOT1_1314(.VSS(VSS),.VDD(VDD),.Y(I15586),.A(g10159));
  NOT NOT1_1315(.VSS(VSS),.VDD(VDD),.Y(I8880),.A(g4537));
  NOT NOT1_1316(.VSS(VSS),.VDD(VDD),.Y(g2255),.A(I5276));
  NOT NOT1_1317(.VSS(VSS),.VDD(VDD),.Y(I5728),.A(g2084));
  NOT NOT1_1318(.VSS(VSS),.VDD(VDD),.Y(g7688),.A(g7148));
  NOT NOT1_1319(.VSS(VSS),.VDD(VDD),.Y(I12793),.A(g7619));
  NOT NOT1_1320(.VSS(VSS),.VDD(VDD),.Y(g2481),.A(g882));
  NOT NOT1_1321(.VSS(VSS),.VDD(VDD),.Y(I9202),.A(g4915));
  NOT NOT1_1322(.VSS(VSS),.VDD(VDD),.Y(g8195),.A(I13122));
  NOT NOT1_1323(.VSS(VSS),.VDD(VDD),.Y(g7976),.A(I12776));
  NOT NOT1_1324(.VSS(VSS),.VDD(VDD),.Y(g8137),.A(I13010));
  NOT NOT1_1325(.VSS(VSS),.VDD(VDD),.Y(g8891),.A(I14239));
  NOT NOT1_1326(.VSS(VSS),.VDD(VDD),.Y(g8337),.A(I13391));
  NOT NOT1_1327(.VSS(VSS),.VDD(VDD),.Y(g10235),.A(g10189));
  NOT NOT1_1328(.VSS(VSS),.VDD(VDD),.Y(g4012),.A(I7154));
  NOT NOT1_1329(.VSS(VSS),.VDD(VDD),.Y(I11183),.A(g6507));
  NOT NOT1_1330(.VSS(VSS),.VDD(VDD),.Y(I16193),.A(g10485));
  NOT NOT1_1331(.VSS(VSS),.VDD(VDD),.Y(g11442),.A(I17377));
  NOT NOT1_1332(.VSS(VSS),.VDD(VDD),.Y(g2097),.A(I4935));
  NOT NOT1_1333(.VSS(VSS),.VDD(VDD),.Y(I12765),.A(g7638));
  NOT NOT1_1334(.VSS(VSS),.VDD(VDD),.Y(g10683),.A(g10612));
  NOT NOT1_1335(.VSS(VSS),.VDD(VDD),.Y(g5742),.A(I9308));
  NOT NOT1_1336(.VSS(VSS),.VDD(VDD),.Y(g2726),.A(g2021));
  NOT NOT1_1337(.VSS(VSS),.VDD(VDD),.Y(g4412),.A(I7746));
  NOT NOT1_1338(.VSS(VSS),.VDD(VDD),.Y(I11397),.A(g6713));
  NOT NOT1_1339(.VSS(VSS),.VDD(VDD),.Y(I13397),.A(g8138));
  NOT NOT1_1340(.VSS(VSS),.VDD(VDD),.Y(g2154),.A(I5067));
  NOT NOT1_1341(.VSS(VSS),.VDD(VDD),.Y(g6016),.A(I9632));
  NOT NOT1_1342(.VSS(VSS),.VDD(VDD),.Y(I12690),.A(g7555));
  NOT NOT1_1343(.VSS(VSS),.VDD(VDD),.Y(g4189),.A(I7384));
  NOT NOT1_1344(.VSS(VSS),.VDD(VDD),.Y(I5070),.A(g1194));
  NOT NOT1_1345(.VSS(VSS),.VDD(VDD),.Y(g2960),.A(I6173));
  NOT NOT1_1346(.VSS(VSS),.VDD(VDD),.Y(I10861),.A(g6694));
  NOT NOT1_1347(.VSS(VSS),.VDD(VDD),.Y(I10573),.A(g5980));
  NOT NOT1_1348(.VSS(VSS),.VDD(VDD),.Y(I9567),.A(g5556));
  NOT NOT1_1349(.VSS(VSS),.VDD(VDD),.Y(g8807),.A(I14140));
  NOT NOT1_1350(.VSS(VSS),.VDD(VDD),.Y(I14573),.A(g9029));
  NOT NOT1_1351(.VSS(VSS),.VDD(VDD),.Y(g4888),.A(I8237));
  NOT NOT1_1352(.VSS(VSS),.VDD(VDD),.Y(g7126),.A(I11367));
  NOT NOT1_1353(.VSS(VSS),.VDD(VDD),.Y(I13933),.A(g8505));
  NOT NOT1_1354(.VSS(VSS),.VDD(VDD),.Y(I17377),.A(g11412));
  NOT NOT1_1355(.VSS(VSS),.VDD(VDD),.Y(g7326),.A(I11626));
  NOT NOT1_1356(.VSS(VSS),.VDD(VDD),.Y(I10045),.A(g5727));
  NOT NOT1_1357(.VSS(VSS),.VDD(VDD),.Y(g6115),.A(I9798));
  NOT NOT1_1358(.VSS(VSS),.VDD(VDD),.Y(g6251),.A(I10012));
  NOT NOT1_1359(.VSS(VSS),.VDD(VDD),.Y(g4171),.A(I7330));
  NOT NOT1_1360(.VSS(VSS),.VDD(VDD),.Y(g6315),.A(I10204));
  NOT NOT1_1361(.VSS(VSS),.VDD(VDD),.Y(g6811),.A(I10843));
  NOT NOT1_1362(.VSS(VSS),.VDD(VDD),.Y(I15275),.A(g9994));
  NOT NOT1_1363(.VSS(VSS),.VDD(VDD),.Y(g4371),.A(I7674));
  NOT NOT1_1364(.VSS(VSS),.VDD(VDD),.Y(I14045),.A(g8603));
  NOT NOT1_1365(.VSS(VSS),.VDD(VDD),.Y(I17739),.A(g11641));
  NOT NOT1_1366(.VSS(VSS),.VDD(VDD),.Y(g4429),.A(I7779));
  NOT NOT1_1367(.VSS(VSS),.VDD(VDD),.Y(g4787),.A(g3423));
  NOT NOT1_1368(.VSS(VSS),.VDD(VDD),.Y(I8982),.A(g4728));
  NOT NOT1_1369(.VSS(VSS),.VDD(VDD),.Y(g11041),.A(I16784));
  NOT NOT1_1370(.VSS(VSS),.VDD(VDD),.Y(g10882),.A(I16616));
  NOT NOT1_1371(.VSS(VSS),.VDD(VDD),.Y(g5754),.A(I9332));
  NOT NOT1_1372(.VSS(VSS),.VDD(VDD),.Y(I9776),.A(g5353));
  NOT NOT1_1373(.VSS(VSS),.VDD(VDD),.Y(I10099),.A(g5800));
  NOT NOT1_1374(.VSS(VSS),.VDD(VDD),.Y(I16475),.A(g10765));
  NOT NOT1_1375(.VSS(VSS),.VDD(VDD),.Y(g6447),.A(g6166));
  NOT NOT1_1376(.VSS(VSS),.VDD(VDD),.Y(I10388),.A(g5830));
  NOT NOT1_1377(.VSS(VSS),.VDD(VDD),.Y(I8234),.A(g4232));
  NOT NOT1_1378(.VSS(VSS),.VDD(VDD),.Y(g7760),.A(I12445));
  NOT NOT1_1379(.VSS(VSS),.VDD(VDD),.Y(I14388),.A(g8924));
  NOT NOT1_1380(.VSS(VSS),.VDD(VDD),.Y(I8328),.A(g4801));
  NOT NOT1_1381(.VSS(VSS),.VDD(VDD),.Y(I17146),.A(g11305));
  NOT NOT1_1382(.VSS(VSS),.VDD(VDD),.Y(I16863),.A(g10972));
  NOT NOT1_1383(.VSS(VSS),.VDD(VDD),.Y(g3092),.A(g2181));
  NOT NOT1_1384(.VSS(VSS),.VDD(VDD),.Y(I14701),.A(g9291));
  NOT NOT1_1385(.VSS(VSS),.VDD(VDD),.Y(I10251),.A(g6126));
  NOT NOT1_1386(.VSS(VSS),.VDD(VDD),.Y(I14534),.A(g9290));
  NOT NOT1_1387(.VSS(VSS),.VDD(VDD),.Y(g4281),.A(g3586));
  NOT NOT1_1388(.VSS(VSS),.VDD(VDD),.Y(I9965),.A(g5493));
  NOT NOT1_1389(.VSS(VSS),.VDD(VDD),.Y(g5613),.A(g4840));
  NOT NOT1_1390(.VSS(VSS),.VDD(VDD),.Y(g6874),.A(I10958));
  NOT NOT1_1391(.VSS(VSS),.VDD(VDD),.Y(g8142),.A(I13023));
  NOT NOT1_1392(.VSS(VSS),.VDD(VDD),.Y(g2112),.A(g639));
  NOT NOT1_1393(.VSS(VSS),.VDD(VDD),.Y(g8342),.A(I13406));
  NOT NOT1_1394(.VSS(VSS),.VDD(VDD),.Y(g2218),.A(g85));
  NOT NOT1_1395(.VSS(VSS),.VDD(VDD),.Y(I15983),.A(g10414));
  NOT NOT1_1396(.VSS(VSS),.VDD(VDD),.Y(g2267),.A(I5304));
  NOT NOT1_1397(.VSS(VSS),.VDD(VDD),.Y(I17698),.A(g11616));
  NOT NOT1_1398(.VSS(VSS),.VDD(VDD),.Y(g11035),.A(I16766));
  NOT NOT1_1399(.VSS(VSS),.VDD(VDD),.Y(g8255),.A(g7986));
  NOT NOT1_1400(.VSS(VSS),.VDD(VDD),.Y(g8081),.A(g8000));
  NOT NOT1_1401(.VSS(VSS),.VDD(VDD),.Y(g8481),.A(g8324));
  NOT NOT1_1402(.VSS(VSS),.VDD(VDD),.Y(g2001),.A(g814));
  NOT NOT1_1403(.VSS(VSS),.VDD(VDD),.Y(g7608),.A(I12174));
  NOT NOT1_1404(.VSS(VSS),.VDD(VDD),.Y(g7924),.A(g7470));
  NOT NOT1_1405(.VSS(VSS),.VDD(VDD),.Y(I5406),.A(g898));
  NOT NOT1_1406(.VSS(VSS),.VDD(VDD),.Y(g7220),.A(I11456));
  NOT NOT1_1407(.VSS(VSS),.VDD(VDD),.Y(g5572),.A(I8989));
  NOT NOT1_1408(.VSS(VSS),.VDD(VDD),.Y(g5862),.A(I9479));
  NOT NOT1_1409(.VSS(VSS),.VDD(VDD),.Y(I12245),.A(g7093));
  NOT NOT1_1410(.VSS(VSS),.VDD(VDD),.Y(g7779),.A(I12502));
  NOT NOT1_1411(.VSS(VSS),.VDD(VDD),.Y(I4780),.A(g872));
  NOT NOT1_1412(.VSS(VSS),.VDD(VDD),.Y(I6040),.A(g2216));
  NOT NOT1_1413(.VSS(VSS),.VDD(VDD),.Y(g6595),.A(I10563));
  NOT NOT1_1414(.VSS(VSS),.VDD(VDD),.Y(g10584),.A(g10522));
  NOT NOT1_1415(.VSS(VSS),.VDD(VDD),.Y(I15517),.A(g10051));
  NOT NOT1_1416(.VSS(VSS),.VDD(VDD),.Y(I13574),.A(g8360));
  NOT NOT1_1417(.VSS(VSS),.VDD(VDD),.Y(g2329),.A(I5383));
  NOT NOT1_1418(.VSS(VSS),.VDD(VDD),.Y(g8354),.A(I13442));
  NOT NOT1_1419(.VSS(VSS),.VDD(VDD),.Y(I14140),.A(g8717));
  NOT NOT1_1420(.VSS(VSS),.VDD(VDD),.Y(g7023),.A(I11166));
  NOT NOT1_1421(.VSS(VSS),.VDD(VDD),.Y(I7952),.A(g3664));
  NOT NOT1_1422(.VSS(VSS),.VDD(VDD),.Y(g4963),.A(I8337));
  NOT NOT1_1423(.VSS(VSS),.VDD(VDD),.Y(g10206),.A(g10178));
  NOT NOT1_1424(.VSS(VSS),.VDD(VDD),.Y(I5801),.A(g1984));
  NOT NOT1_1425(.VSS(VSS),.VDD(VDD),.Y(I7276),.A(g2861));
  NOT NOT1_1426(.VSS(VSS),.VDD(VDD),.Y(g9670),.A(I14799));
  NOT NOT1_1427(.VSS(VSS),.VDD(VDD),.Y(I16781),.A(g10893));
  NOT NOT1_1428(.VSS(VSS),.VDD(VDD),.Y(g4791),.A(I8161));
  NOT NOT1_1429(.VSS(VSS),.VDD(VDD),.Y(g7977),.A(I12779));
  NOT NOT1_1430(.VSS(VSS),.VDD(VDD),.Y(g2828),.A(I5940));
  NOT NOT1_1431(.VSS(VSS),.VDD(VDD),.Y(g6272),.A(I10075));
  NOT NOT1_1432(.VSS(VSS),.VDD(VDD),.Y(I16236),.A(g10535));
  NOT NOT1_1433(.VSS(VSS),.VDD(VDD),.Y(g3262),.A(I6432));
  NOT NOT1_1434(.VSS(VSS),.VDD(VDD),.Y(g2727),.A(g2022));
  NOT NOT1_1435(.VSS(VSS),.VDD(VDD),.Y(g3736),.A(I6924));
  NOT NOT1_1436(.VSS(VSS),.VDD(VDD),.Y(g5534),.A(g4545));
  NOT NOT1_1437(.VSS(VSS),.VDD(VDD),.Y(g5729),.A(I9279));
  NOT NOT1_1438(.VSS(VSS),.VDD(VDD),.Y(g7361),.A(I11731));
  NOT NOT1_1439(.VSS(VSS),.VDD(VDD),.Y(g10114),.A(I15350));
  NOT NOT1_1440(.VSS(VSS),.VDD(VDD),.Y(I16175),.A(g10488));
  NOT NOT1_1441(.VSS(VSS),.VDD(VDD),.Y(g9813),.A(I14948));
  NOT NOT1_1442(.VSS(VSS),.VDD(VDD),.Y(I15193),.A(g9968));
  NOT NOT1_1443(.VSS(VSS),.VDD(VDD),.Y(g6417),.A(g6136));
  NOT NOT1_1444(.VSS(VSS),.VDD(VDD),.Y(I13051),.A(g8060));
  NOT NOT1_1445(.VSS(VSS),.VDD(VDD),.Y(I15362),.A(g9987));
  NOT NOT1_1446(.VSS(VSS),.VDD(VDD),.Y(g6935),.A(I11065));
  NOT NOT1_1447(.VSS(VSS),.VDD(VDD),.Y(g11193),.A(g11112));
  NOT NOT1_1448(.VSS(VSS),.VDD(VDD),.Y(g7051),.A(I11232));
  NOT NOT1_1449(.VSS(VSS),.VDD(VDD),.Y(g10107),.A(I15341));
  NOT NOT1_1450(.VSS(VSS),.VDD(VDD),.Y(I11756),.A(g7191));
  NOT NOT1_1451(.VSS(VSS),.VDD(VDD),.Y(g2221),.A(I5198));
  NOT NOT1_1452(.VSS(VSS),.VDD(VDD),.Y(g3076),.A(I6282));
  NOT NOT1_1453(.VSS(VSS),.VDD(VDD),.Y(I13592),.A(g8362));
  NOT NOT1_1454(.VSS(VSS),.VDD(VDD),.Y(g8783),.A(g8746));
  NOT NOT1_1455(.VSS(VSS),.VDD(VDD),.Y(I15523),.A(g10058));
  NOT NOT1_1456(.VSS(VSS),.VDD(VDD),.Y(g7327),.A(I11629));
  NOT NOT1_1457(.VSS(VSS),.VDD(VDD),.Y(I12232),.A(g7072));
  NOT NOT1_1458(.VSS(VSS),.VDD(VDD),.Y(I6528),.A(g3274));
  NOT NOT1_1459(.VSS(VSS),.VDD(VDD),.Y(I16264),.A(g10557));
  NOT NOT1_1460(.VSS(VSS),.VDD(VDD),.Y(g8979),.A(I14358));
  NOT NOT1_1461(.VSS(VSS),.VDD(VDD),.Y(I16790),.A(g10900));
  NOT NOT1_1462(.VSS(VSS),.VDD(VDD),.Y(I8490),.A(g4526));
  NOT NOT1_1463(.VSS(VSS),.VDD(VDD),.Y(g4201),.A(I7420));
  NOT NOT1_1464(.VSS(VSS),.VDD(VDD),.Y(I6648),.A(g2635));
  NOT NOT1_1465(.VSS(VSS),.VDD(VDD),.Y(g8218),.A(g7826));
  NOT NOT1_1466(.VSS(VSS),.VDD(VDD),.Y(I9658),.A(g5150));
  NOT NOT1_1467(.VSS(VSS),.VDD(VDD),.Y(g8312),.A(I13320));
  NOT NOT1_1468(.VSS(VSS),.VDD(VDD),.Y(I7546),.A(g4105));
  NOT NOT1_1469(.VSS(VSS),.VDD(VDD),.Y(g6128),.A(I9829));
  NOT NOT1_1470(.VSS(VSS),.VDD(VDD),.Y(g6629),.A(I10584));
  NOT NOT1_1471(.VSS(VSS),.VDD(VDD),.Y(g5885),.A(g5361));
  NOT NOT1_1472(.VSS(VSS),.VDD(VDD),.Y(g10345),.A(I15801));
  NOT NOT1_1473(.VSS(VSS),.VDD(VDD),.Y(g7999),.A(I12825));
  NOT NOT1_1474(.VSS(VSS),.VDD(VDD),.Y(g7146),.A(I11391));
  NOT NOT1_1475(.VSS(VSS),.VDD(VDD),.Y(g5660),.A(I9141));
  NOT NOT1_1476(.VSS(VSS),.VDD(VDD),.Y(I5445),.A(g922));
  NOT NOT1_1477(.VSS(VSS),.VDD(VDD),.Y(g6330),.A(I10221));
  NOT NOT1_1478(.VSS(VSS),.VDD(VDD),.Y(g7346),.A(I11686));
  NOT NOT1_1479(.VSS(VSS),.VDD(VDD),.Y(I10162),.A(g5943));
  NOT NOT1_1480(.VSS(VSS),.VDD(VDD),.Y(g7633),.A(I12239));
  NOT NOT1_1481(.VSS(VSS),.VDD(VDD),.Y(g4049),.A(g3144));
  NOT NOT1_1482(.VSS(VSS),.VDD(VDD),.Y(g3375),.A(I6569));
  NOT NOT1_1483(.VSS(VSS),.VDD(VDD),.Y(g8001),.A(I12829));
  NOT NOT1_1484(.VSS(VSS),.VDD(VDD),.Y(I12261),.A(g7078));
  NOT NOT1_1485(.VSS(VSS),.VDD(VDD),.Y(g4449),.A(g4144));
  NOT NOT1_1486(.VSS(VSS),.VDD(VDD),.Y(g3722),.A(I6894));
  NOT NOT1_1487(.VSS(VSS),.VDD(VDD),.Y(I8456),.A(g4472));
  NOT NOT1_1488(.VSS(VSS),.VDD(VDD),.Y(g7103),.A(I11338));
  NOT NOT1_1489(.VSS(VSS),.VDD(VDD),.Y(g5903),.A(I9536));
  NOT NOT1_1490(.VSS(VSS),.VDD(VDD),.Y(g4575),.A(g3880));
  NOT NOT1_1491(.VSS(VSS),.VDD(VDD),.Y(g10848),.A(I16546));
  NOT NOT1_1492(.VSS(VSS),.VDD(VDD),.Y(g11475),.A(I17466));
  NOT NOT1_1493(.VSS(VSS),.VDD(VDD),.Y(g8293),.A(I13233));
  NOT NOT1_1494(.VSS(VSS),.VDD(VDD),.Y(g8129),.A(g8015));
  NOT NOT1_1495(.VSS(VSS),.VDD(VDD),.Y(I6010),.A(g2256));
  NOT NOT1_1496(.VSS(VSS),.VDD(VDD),.Y(g2068),.A(I4866));
  NOT NOT1_1497(.VSS(VSS),.VDD(VDD),.Y(I11152),.A(g6469));
  NOT NOT1_1498(.VSS(VSS),.VDD(VDD),.Y(g8329),.A(I13367));
  NOT NOT1_1499(.VSS(VSS),.VDD(VDD),.Y(g10141),.A(I15421));
  NOT NOT1_1500(.VSS(VSS),.VDD(VDD),.Y(g7696),.A(g7148));
  NOT NOT1_1501(.VSS(VSS),.VDD(VDD),.Y(g10804),.A(I16514));
  NOT NOT1_1502(.VSS(VSS),.VDD(VDD),.Y(g6800),.A(I10810));
  NOT NOT1_1503(.VSS(VSS),.VDD(VDD),.Y(g4098),.A(I7240));
  NOT NOT1_1504(.VSS(VSS),.VDD(VDD),.Y(g3500),.A(I6690));
  NOT NOT1_1505(.VSS(VSS),.VDD(VDD),.Y(I15437),.A(g10050));
  NOT NOT1_1506(.VSS(VSS),.VDD(VDD),.Y(I16209),.A(g10452));
  NOT NOT1_1507(.VSS(VSS),.VDD(VDD),.Y(I8851),.A(g4498));
  NOT NOT1_1508(.VSS(VSS),.VDD(VDD),.Y(I11731),.A(g7021));
  NOT NOT1_1509(.VSS(VSS),.VDD(VDD),.Y(g8828),.A(g8744));
  NOT NOT1_1510(.VSS(VSS),.VDD(VDD),.Y(g11437),.A(I17362));
  NOT NOT1_1511(.VSS(VSS),.VDD(VDD),.Y(g2677),.A(g2034));
  NOT NOT1_1512(.VSS(VSS),.VDD(VDD),.Y(g10263),.A(g10127));
  NOT NOT1_1513(.VSS(VSS),.VDD(VDD),.Y(g7753),.A(I12424));
  NOT NOT1_1514(.VSS(VSS),.VDD(VDD),.Y(I9981),.A(g5514));
  NOT NOT1_1515(.VSS(VSS),.VDD(VDD),.Y(g8727),.A(g8592));
  NOT NOT1_1516(.VSS(VSS),.VDD(VDD),.Y(g5679),.A(I9194));
  NOT NOT1_1517(.VSS(VSS),.VDD(VDD),.Y(g7508),.A(g6950));
  NOT NOT1_1518(.VSS(VSS),.VDD(VDD),.Y(g3384),.A(g3143));
  NOT NOT1_1519(.VSS(VSS),.VDD(VDD),.Y(g10332),.A(I15782));
  NOT NOT1_1520(.VSS(VSS),.VDD(VDD),.Y(g6213),.A(g5426));
  NOT NOT1_1521(.VSS(VSS),.VDD(VDD),.Y(g8592),.A(I13837));
  NOT NOT1_1522(.VSS(VSS),.VDD(VDD),.Y(g7944),.A(g7410));
  NOT NOT1_1523(.VSS(VSS),.VDD(VDD),.Y(I15347),.A(g9995));
  NOT NOT1_1524(.VSS(VSS),.VDD(VDD),.Y(g7072),.A(I11293));
  NOT NOT1_1525(.VSS(VSS),.VDD(VDD),.Y(I15253),.A(g9987));
  NOT NOT1_1526(.VSS(VSS),.VDD(VDD),.Y(g10135),.A(I15403));
  NOT NOT1_1527(.VSS(VSS),.VDD(VDD),.Y(I12445),.A(g7521));
  NOT NOT1_1528(.VSS(VSS),.VDD(VDD),.Y(g11347),.A(I17164));
  NOT NOT1_1529(.VSS(VSS),.VDD(VDD),.Y(g4896),.A(I8253));
  NOT NOT1_1530(.VSS(VSS),.VDD(VDD),.Y(I7906),.A(g3907));
  NOT NOT1_1531(.VSS(VSS),.VDD(VDD),.Y(g2349),.A(I5421));
  NOT NOT1_1532(.VSS(VSS),.VDD(VDD),.Y(g7043),.A(I11214));
  NOT NOT1_1533(.VSS(VSS),.VDD(VDD),.Y(I12499),.A(g7725));
  NOT NOT1_1534(.VSS(VSS),.VDD(VDD),.Y(I11405),.A(g6627));
  NOT NOT1_1535(.VSS(VSS),.VDD(VDD),.Y(g5288),.A(g4438));
  NOT NOT1_1536(.VSS(VSS),.VDD(VDD),.Y(g9341),.A(I14528));
  NOT NOT1_1537(.VSS(VSS),.VDD(VDD),.Y(g3424),.A(g2896));
  NOT NOT1_1538(.VSS(VSS),.VDD(VDD),.Y(I9132),.A(g4893));
  NOT NOT1_1539(.VSS(VSS),.VDD(VDD),.Y(g10361),.A(g10268));
  NOT NOT1_1540(.VSS(VSS),.VDD(VDD),.Y(g3737),.A(g2834));
  NOT NOT1_1541(.VSS(VSS),.VDD(VDD),.Y(g7443),.A(I11841));
  NOT NOT1_1542(.VSS(VSS),.VDD(VDD),.Y(I9332),.A(g4935));
  NOT NOT1_1543(.VSS(VSS),.VDD(VDD),.Y(g9525),.A(g9257));
  NOT NOT1_1544(.VSS(VSS),.VDD(VDD),.Y(I9153),.A(g5027));
  NOT NOT1_1545(.VSS(VSS),.VDD(VDD),.Y(I9680),.A(g5194));
  NOT NOT1_1546(.VSS(VSS),.VDD(VDD),.Y(I10147),.A(g5697));
  NOT NOT1_1547(.VSS(VSS),.VDD(VDD),.Y(I6343),.A(g1963));
  NOT NOT1_1548(.VSS(VSS),.VDD(VDD),.Y(I10355),.A(g6003));
  NOT NOT1_1549(.VSS(VSS),.VDD(VDD),.Y(g7116),.A(I11351));
  NOT NOT1_1550(.VSS(VSS),.VDD(VDD),.Y(g5805),.A(I9409));
  NOT NOT1_1551(.VSS(VSS),.VDD(VDD),.Y(g5916),.A(I9550));
  NOT NOT1_1552(.VSS(VSS),.VDD(VDD),.Y(g7316),.A(I11596));
  NOT NOT1_1553(.VSS(VSS),.VDD(VDD),.Y(g2198),.A(g668));
  NOT NOT1_1554(.VSS(VSS),.VDD(VDD),.Y(I6282),.A(g2231));
  NOT NOT1_1555(.VSS(VSS),.VDD(VDD),.Y(g4268),.A(I7523));
  NOT NOT1_1556(.VSS(VSS),.VDD(VDD),.Y(I7771),.A(g3418));
  NOT NOT1_1557(.VSS(VSS),.VDD(VDD),.Y(I16607),.A(g10787));
  NOT NOT1_1558(.VSS(VSS),.VDD(VDD),.Y(g2855),.A(I5989));
  NOT NOT1_1559(.VSS(VSS),.VDD(VDD),.Y(g4362),.A(I7651));
  NOT NOT1_1560(.VSS(VSS),.VDD(VDD),.Y(I11929),.A(g6901));
  NOT NOT1_1561(.VSS(VSS),.VDD(VDD),.Y(I14355),.A(g8948));
  NOT NOT1_1562(.VSS(VSS),.VDD(VDD),.Y(I12989),.A(g8043));
  NOT NOT1_1563(.VSS(VSS),.VDD(VDD),.Y(g11351),.A(I17170));
  NOT NOT1_1564(.VSS(VSS),.VDD(VDD),.Y(g3077),.A(g2213));
  NOT NOT1_1565(.VSS(VSS),.VDD(VDD),.Y(g5422),.A(g4470));
  NOT NOT1_1566(.VSS(VSS),.VDD(VDD),.Y(g7034),.A(I11191));
  NOT NOT1_1567(.VSS(VSS),.VDD(VDD),.Y(I10825),.A(g6588));
  NOT NOT1_1568(.VSS(VSS),.VDD(VDD),.Y(g4419),.A(I7763));
  NOT NOT1_1569(.VSS(VSS),.VDD(VDD),.Y(I9744),.A(g5263));
  NOT NOT1_1570(.VSS(VSS),.VDD(VDD),.Y(I12056),.A(g6929));
  NOT NOT1_1571(.VSS(VSS),.VDD(VDD),.Y(I10370),.A(g5857));
  NOT NOT1_1572(.VSS(VSS),.VDD(VDD),.Y(g6166),.A(I9893));
  NOT NOT1_1573(.VSS(VSS),.VDD(VDD),.Y(g8624),.A(g8486));
  NOT NOT1_1574(.VSS(VSS),.VDD(VDD),.Y(g3523),.A(g2971));
  NOT NOT1_1575(.VSS(VSS),.VDD(VDD),.Y(I14370),.A(g8954));
  NOT NOT1_1576(.VSS(VSS),.VDD(VDD),.Y(g8953),.A(I14312));
  NOT NOT1_1577(.VSS(VSS),.VDD(VDD),.Y(I10858),.A(g6688));
  NOT NOT1_1578(.VSS(VSS),.VDD(VDD),.Y(I13020),.A(g8049));
  NOT NOT1_1579(.VSS(VSS),.VDD(VDD),.Y(I13583),.A(g8344));
  NOT NOT1_1580(.VSS(VSS),.VDD(VDD),.Y(g4452),.A(g3365));
  NOT NOT1_1581(.VSS(VSS),.VDD(VDD),.Y(I8872),.A(g4529));
  NOT NOT1_1582(.VSS(VSS),.VDD(VDD),.Y(I15063),.A(g9699));
  NOT NOT1_1583(.VSS(VSS),.VDD(VDD),.Y(g2241),.A(g722));
  NOT NOT1_1584(.VSS(VSS),.VDD(VDD),.Y(g7147),.A(I11394));
  NOT NOT1_1585(.VSS(VSS),.VDD(VDD),.Y(g6056),.A(g5426));
  NOT NOT1_1586(.VSS(VSS),.VDD(VDD),.Y(g5947),.A(I9585));
  NOT NOT1_1587(.VSS(VSS),.VDD(VDD),.Y(g7347),.A(I11689));
  NOT NOT1_1588(.VSS(VSS),.VDD(VDD),.Y(g11063),.A(g10974));
  NOT NOT1_1589(.VSS(VSS),.VDD(VDD),.Y(I11046),.A(g6635));
  NOT NOT1_1590(.VSS(VSS),.VDD(VDD),.Y(I10996),.A(g6786));
  NOT NOT1_1591(.VSS(VSS),.VDD(VDD),.Y(I12271),.A(g7218));
  NOT NOT1_1592(.VSS(VSS),.VDD(VDD),.Y(g7681),.A(g7148));
  NOT NOT1_1593(.VSS(VSS),.VDD(VDD),.Y(g6649),.A(I10610));
  NOT NOT1_1594(.VSS(VSS),.VDD(VDD),.Y(I8989),.A(g4746));
  NOT NOT1_1595(.VSS(VSS),.VDD(VDD),.Y(g8677),.A(I13962));
  NOT NOT1_1596(.VSS(VSS),.VDD(VDD),.Y(g110),.A(I4786));
  NOT NOT1_1597(.VSS(VSS),.VDD(VDD),.Y(I10367),.A(g6234));
  NOT NOT1_1598(.VSS(VSS),.VDD(VDD),.Y(I10394),.A(g5824));
  NOT NOT1_1599(.VSS(VSS),.VDD(VDD),.Y(I9901),.A(g5557));
  NOT NOT1_1600(.VSS(VSS),.VDD(VDD),.Y(g7697),.A(g7101));
  NOT NOT1_1601(.VSS(VSS),.VDD(VDD),.Y(I14367),.A(g8953));
  NOT NOT1_1602(.VSS(VSS),.VDD(VDD),.Y(I14394),.A(g8884));
  NOT NOT1_1603(.VSS(VSS),.VDD(VDD),.Y(I16641),.A(g10864));
  NOT NOT1_1604(.VSS(VSS),.VDD(VDD),.Y(g3742),.A(I6929));
  NOT NOT1_1605(.VSS(VSS),.VDD(VDD),.Y(g7914),.A(g7651));
  NOT NOT1_1606(.VSS(VSS),.VDD(VDD),.Y(g8576),.A(I13819));
  NOT NOT1_1607(.VSS(VSS),.VDD(VDD),.Y(g2524),.A(g986));
  NOT NOT1_1608(.VSS(VSS),.VDD(VDD),.Y(g7210),.A(I11440));
  NOT NOT1_1609(.VSS(VSS),.VDD(VDD),.Y(g4728),.A(I8080));
  NOT NOT1_1610(.VSS(VSS),.VDD(VDD),.Y(I16292),.A(g10551));
  NOT NOT1_1611(.VSS(VSS),.VDD(VDD),.Y(g2644),.A(g1990));
  NOT NOT1_1612(.VSS(VSS),.VDD(VDD),.Y(g6698),.A(I10671));
  NOT NOT1_1613(.VSS(VSS),.VDD(VDD),.Y(g4730),.A(g3546));
  NOT NOT1_1614(.VSS(VSS),.VDD(VDD),.Y(g8716),.A(g8576));
  NOT NOT1_1615(.VSS(VSS),.VDD(VDD),.Y(I17546),.A(g11500));
  NOT NOT1_1616(.VSS(VSS),.VDD(VDD),.Y(g8149),.A(I13036));
  NOT NOT1_1617(.VSS(VSS),.VDD(VDD),.Y(g10947),.A(I16708));
  NOT NOT1_1618(.VSS(VSS),.VDD(VDD),.Y(g4504),.A(I7899));
  NOT NOT1_1619(.VSS(VSS),.VDD(VDD),.Y(I11357),.A(g6594));
  NOT NOT1_1620(.VSS(VSS),.VDD(VDD),.Y(g6964),.A(g6509));
  NOT NOT1_1621(.VSS(VSS),.VDD(VDD),.Y(g8349),.A(I13427));
  NOT NOT1_1622(.VSS(VSS),.VDD(VDD),.Y(g2119),.A(I5031));
  NOT NOT1_1623(.VSS(VSS),.VDD(VDD),.Y(g5095),.A(I8465));
  NOT NOT1_1624(.VSS(VSS),.VDD(VDD),.Y(g6260),.A(I10039));
  NOT NOT1_1625(.VSS(VSS),.VDD(VDD),.Y(g5037),.A(I8414));
  NOT NOT1_1626(.VSS(VSS),.VDD(VDD),.Y(I13357),.A(g8125));
  NOT NOT1_1627(.VSS(VSS),.VDD(VDD),.Y(I12199),.A(g7278));
  NOT NOT1_1628(.VSS(VSS),.VDD(VDD),.Y(g4185),.A(I7372));
  NOT NOT1_1629(.VSS(VSS),.VDD(VDD),.Y(I7244),.A(g3226));
  NOT NOT1_1630(.VSS(VSS),.VDD(VDD),.Y(g9311),.A(I14506));
  NOT NOT1_1631(.VSS(VSS),.VDD(VDD),.Y(g11422),.A(I17321));
  NOT NOT1_1632(.VSS(VSS),.VDD(VDD),.Y(I11743),.A(g7035));
  NOT NOT1_1633(.VSS(VSS),.VDD(VDD),.Y(I13105),.A(g7929));
  NOT NOT1_1634(.VSS(VSS),.VDD(VDD),.Y(g5653),.A(I9120));
  NOT NOT1_1635(.VSS(VSS),.VDD(VDD),.Y(g4385),.A(I7710));
  NOT NOT1_1636(.VSS(VSS),.VDD(VDD),.Y(g7413),.A(g7197));
  NOT NOT1_1637(.VSS(VSS),.VDD(VDD),.Y(g5102),.A(I8476));
  NOT NOT1_1638(.VSS(VSS),.VDD(VDD),.Y(g2258),.A(I5289));
  NOT NOT1_1639(.VSS(VSS),.VDD(VDD),.Y(I14319),.A(g8816));
  NOT NOT1_1640(.VSS(VSS),.VDD(VDD),.Y(g2352),.A(I5430));
  NOT NOT1_1641(.VSS(VSS),.VDD(VDD),.Y(g2818),.A(I5922));
  NOT NOT1_1642(.VSS(VSS),.VDD(VDD),.Y(I7140),.A(g2641));
  NOT NOT1_1643(.VSS(VSS),.VDD(VDD),.Y(g6063),.A(g5446));
  NOT NOT1_1644(.VSS(VSS),.VDD(VDD),.Y(I12529),.A(g7589));
  NOT NOT1_1645(.VSS(VSS),.VDD(VDD),.Y(I5940),.A(g2175));
  NOT NOT1_1646(.VSS(VSS),.VDD(VDD),.Y(g2867),.A(I6007));
  NOT NOT1_1647(.VSS(VSS),.VDD(VDD),.Y(I16635),.A(g10862));
  NOT NOT1_1648(.VSS(VSS),.VDD(VDD),.Y(g10463),.A(I15980));
  NOT NOT1_1649(.VSS(VSS),.VDD(VDD),.Y(g11208),.A(g11077));
  NOT NOT1_1650(.VSS(VSS),.VDD(VDD),.Y(g4470),.A(I7843));
  NOT NOT1_1651(.VSS(VSS),.VDD(VDD),.Y(g8198),.A(I13131));
  NOT NOT1_1652(.VSS(VSS),.VDD(VDD),.Y(g4897),.A(I8256));
  NOT NOT1_1653(.VSS(VSS),.VDD(VDD),.Y(g8747),.A(I14040));
  NOT NOT1_1654(.VSS(VSS),.VDD(VDD),.Y(I7478),.A(g3566));
  NOT NOT1_1655(.VSS(VSS),.VDD(VDD),.Y(g5719),.A(I9259));
  NOT NOT1_1656(.VSS(VSS),.VDD(VDD),.Y(g4425),.A(I7771));
  NOT NOT1_1657(.VSS(VSS),.VDD(VDD),.Y(I12843),.A(g7683));
  NOT NOT1_1658(.VSS(VSS),.VDD(VDD),.Y(I15542),.A(g10065));
  NOT NOT1_1659(.VSS(VSS),.VDD(VDD),.Y(g10972),.A(I16717));
  NOT NOT1_1660(.VSS(VSS),.VDD(VDD),.Y(g10033),.A(I15235));
  NOT NOT1_1661(.VSS(VSS),.VDD(VDD),.Y(I5388),.A(g889));
  NOT NOT1_1662(.VSS(VSS),.VDD(VDD),.Y(g10234),.A(g10188));
  NOT NOT1_1663(.VSS(VSS),.VDD(VDD),.Y(I7435),.A(g3459));
  NOT NOT1_1664(.VSS(VSS),.VDD(VDD),.Y(g7936),.A(g7712));
  NOT NOT1_1665(.VSS(VSS),.VDD(VDD),.Y(g11542),.A(g11519));
  NOT NOT1_1666(.VSS(VSS),.VDD(VDD),.Y(g11453),.A(I17416));
  NOT NOT1_1667(.VSS(VSS),.VDD(VDD),.Y(g5752),.A(I9326));
  NOT NOT1_1668(.VSS(VSS),.VDD(VDD),.Y(I6094),.A(g2110));
  NOT NOT1_1669(.VSS(VSS),.VDD(VDD),.Y(I13803),.A(g8476));
  NOT NOT1_1670(.VSS(VSS),.VDD(VDD),.Y(g3044),.A(I6256));
  NOT NOT1_1671(.VSS(VSS),.VDD(VDD),.Y(g2211),.A(g153));
  NOT NOT1_1672(.VSS(VSS),.VDD(VDD),.Y(I14540),.A(g9310));
  NOT NOT1_1673(.VSS(VSS),.VDD(VDD),.Y(g6279),.A(I10096));
  NOT NOT1_1674(.VSS(VSS),.VDD(VDD),.Y(g2186),.A(g90));
  NOT NOT1_1675(.VSS(VSS),.VDD(VDD),.Y(g7317),.A(I11599));
  NOT NOT1_1676(.VSS(VSS),.VDD(VDD),.Y(g6720),.A(I10713));
  NOT NOT1_1677(.VSS(VSS),.VDD(VDD),.Y(I8253),.A(g4637));
  NOT NOT1_1678(.VSS(VSS),.VDD(VDD),.Y(g6118),.A(I9807));
  NOT NOT1_1679(.VSS(VSS),.VDD(VDD),.Y(g3983),.A(g3222));
  NOT NOT1_1680(.VSS(VSS),.VDD(VDD),.Y(g11614),.A(I17662));
  NOT NOT1_1681(.VSS(VSS),.VDD(VDD),.Y(g7601),.A(I12153));
  NOT NOT1_1682(.VSS(VSS),.VDD(VDD),.Y(I5430),.A(g916));
  NOT NOT1_1683(.VSS(VSS),.VDD(VDD),.Y(g5265),.A(g4362));
  NOT NOT1_1684(.VSS(VSS),.VDD(VDD),.Y(g11436),.A(I17359));
  NOT NOT1_1685(.VSS(VSS),.VDD(VDD),.Y(g3862),.A(g2920));
  NOT NOT1_1686(.VSS(VSS),.VDD(VDD),.Y(g5042),.A(g4840));
  NOT NOT1_1687(.VSS(VSS),.VDD(VDD),.Y(I15320),.A(g10013));
  NOT NOT1_1688(.VSS(VSS),.VDD(VDD),.Y(g9832),.A(I14989));
  NOT NOT1_1689(.VSS(VSS),.VDD(VDD),.Y(g6652),.A(I10613));
  NOT NOT1_1690(.VSS(VSS),.VDD(VDD),.Y(g4678),.A(g3546));
  NOT NOT1_1691(.VSS(VSS),.VDD(VDD),.Y(g6057),.A(g5446));
  NOT NOT1_1692(.VSS(VSS),.VDD(VDD),.Y(g6843),.A(I10901));
  NOT NOT1_1693(.VSS(VSS),.VDD(VDD),.Y(I15530),.A(g10107));
  NOT NOT1_1694(.VSS(VSS),.VDD(VDD),.Y(g11073),.A(g10913));
  NOT NOT1_1695(.VSS(VSS),.VDD(VDD),.Y(g4331),.A(I7606));
  NOT NOT1_1696(.VSS(VSS),.VDD(VDD),.Y(g3543),.A(g3101));
  NOT NOT1_1697(.VSS(VSS),.VDD(VDD),.Y(g2170),.A(g30));
  NOT NOT1_1698(.VSS(VSS),.VDD(VDD),.Y(g2614),.A(g1994));
  NOT NOT1_1699(.VSS(VSS),.VDD(VDD),.Y(g7775),.A(I12490));
  NOT NOT1_1700(.VSS(VSS),.VDD(VDD),.Y(g11593),.A(I17633));
  NOT NOT1_1701(.VSS(VSS),.VDD(VDD),.Y(g7922),.A(I12712));
  NOT NOT1_1702(.VSS(VSS),.VDD(VDD),.Y(g2125),.A(I5053));
  NOT NOT1_1703(.VSS(VSS),.VDD(VDD),.Y(g8319),.A(I13341));
  NOT NOT1_1704(.VSS(VSS),.VDD(VDD),.Y(g11346),.A(I17161));
  NOT NOT1_1705(.VSS(VSS),.VDD(VDD),.Y(I15565),.A(g10101));
  NOT NOT1_1706(.VSS(VSS),.VDD(VDD),.Y(g2821),.A(I5929));
  NOT NOT1_1707(.VSS(VSS),.VDD(VDD),.Y(g9507),.A(g9268));
  NOT NOT1_1708(.VSS(VSS),.VDD(VDD),.Y(I15464),.A(g10094));
  NOT NOT1_1709(.VSS(VSS),.VDD(VDD),.Y(I6965),.A(g2880));
  NOT NOT1_1710(.VSS(VSS),.VDD(VDD),.Y(I10120),.A(g6248));
  NOT NOT1_1711(.VSS(VSS),.VDD(VDD),.Y(g4766),.A(g3440));
  NOT NOT1_1712(.VSS(VSS),.VDD(VDD),.Y(I11662),.A(g7033));
  NOT NOT1_1713(.VSS(VSS),.VDD(VDD),.Y(I10739),.A(g5942));
  NOT NOT1_1714(.VSS(VSS),.VDD(VDD),.Y(g4087),.A(I7220));
  NOT NOT1_1715(.VSS(VSS),.VDD(VDD),.Y(g4105),.A(I7249));
  NOT NOT1_1716(.VSS(VSS),.VDD(VDD),.Y(g8152),.A(I13043));
  NOT NOT1_1717(.VSS(VSS),.VDD(VDD),.Y(g10421),.A(g10331));
  NOT NOT1_1718(.VSS(VSS),.VDD(VDD),.Y(I16537),.A(g10721));
  NOT NOT1_1719(.VSS(VSS),.VDD(VDD),.Y(g8352),.A(I13436));
  NOT NOT1_1720(.VSS(VSS),.VDD(VDD),.Y(g4305),.A(g4013));
  NOT NOT1_1721(.VSS(VSS),.VDD(VDD),.Y(g6971),.A(g6517));
  NOT NOT1_1722(.VSS(VSS),.VDD(VDD),.Y(I13027),.A(g8051));
  NOT NOT1_1723(.VSS(VSS),.VDD(VDD),.Y(I12258),.A(g7103));
  NOT NOT1_1724(.VSS(VSS),.VDD(VDD),.Y(g3729),.A(I6907));
  NOT NOT1_1725(.VSS(VSS),.VDD(VDD),.Y(I6264),.A(g2118));
  NOT NOT1_1726(.VSS(VSS),.VDD(VDD),.Y(I16108),.A(g10383));
  NOT NOT1_1727(.VSS(VSS),.VDD(VDD),.Y(g6686),.A(I10651));
  NOT NOT1_1728(.VSS(VSS),.VDD(VDD),.Y(g10163),.A(I15485));
  NOT NOT1_1729(.VSS(VSS),.VDD(VDD),.Y(g8717),.A(I14010));
  NOT NOT1_1730(.VSS(VSS),.VDD(VDD),.Y(g11034),.A(I16763));
  NOT NOT1_1731(.VSS(VSS),.VDD(VDD),.Y(g7460),.A(g7148));
  NOT NOT1_1732(.VSS(VSS),.VDD(VDD),.Y(g7597),.A(I12133));
  NOT NOT1_1733(.VSS(VSS),.VDD(VDD),.Y(g5296),.A(g4444));
  NOT NOT1_1734(.VSS(VSS),.VDD(VDD),.Y(I11249),.A(g6541));
  NOT NOT1_1735(.VSS(VSS),.VDD(VDD),.Y(I5638),.A(g936));
  NOT NOT1_1736(.VSS(VSS),.VDD(VDD),.Y(I14645),.A(g9088));
  NOT NOT1_1737(.VSS(VSS),.VDD(VDD),.Y(I16283),.A(g10538));
  NOT NOT1_1738(.VSS(VSS),.VDD(VDD),.Y(g2083),.A(g139));
  NOT NOT1_1739(.VSS(VSS),.VDD(VDD),.Y(I6360),.A(g2261));
  NOT NOT1_1740(.VSS(VSS),.VDD(VDD),.Y(g4748),.A(g3546));
  NOT NOT1_1741(.VSS(VSS),.VDD(VDD),.Y(I16492),.A(g10773));
  NOT NOT1_1742(.VSS(VSS),.VDD(VDD),.Y(I13482),.A(g8193));
  NOT NOT1_1743(.VSS(VSS),.VDD(VDD),.Y(I5308),.A(g97));
  NOT NOT1_1744(.VSS(VSS),.VDD(VDD),.Y(I11710),.A(g7020));
  NOT NOT1_1745(.VSS(VSS),.VDD(VDD),.Y(g7784),.A(I12517));
  NOT NOT1_1746(.VSS(VSS),.VDD(VDD),.Y(I4992),.A(g1170));
  NOT NOT1_1747(.VSS(VSS),.VDD(VDD),.Y(g4755),.A(g3440));
  NOT NOT1_1748(.VSS(VSS),.VDD(VDD),.Y(g10541),.A(I16190));
  NOT NOT1_1749(.VSS(VSS),.VDD(VDD),.Y(I10698),.A(g5856));
  NOT NOT1_1750(.VSS(VSS),.VDD(VDD),.Y(g6121),.A(I9816));
  NOT NOT1_1751(.VSS(VSS),.VDD(VDD),.Y(I15409),.A(g10065));
  NOT NOT1_1752(.VSS(VSS),.VDD(VDD),.Y(I7002),.A(g2907));
  NOT NOT1_1753(.VSS(VSS),.VDD(VDD),.Y(g8186),.A(I13109));
  NOT NOT1_1754(.VSS(VSS),.VDD(VDD),.Y(g10473),.A(g10380));
  NOT NOT1_1755(.VSS(VSS),.VDD(VDD),.Y(g4226),.A(g3698));
  NOT NOT1_1756(.VSS(VSS),.VDD(VDD),.Y(I11204),.A(g6523));
  NOT NOT1_1757(.VSS(VSS),.VDD(VDD),.Y(g6670),.A(I10633));
  NOT NOT1_1758(.VSS(VSS),.VDD(VDD),.Y(I7402),.A(g4121));
  NOT NOT1_1759(.VSS(VSS),.VDD(VDD),.Y(g11409),.A(I17268));
  NOT NOT1_1760(.VSS(VSS),.VDD(VDD),.Y(I6996),.A(g2904));
  NOT NOT1_1761(.VSS(VSS),.VDD(VDD),.Y(g3946),.A(I7099));
  NOT NOT1_1762(.VSS(VSS),.VDD(VDD),.Y(I13779),.A(g8514));
  NOT NOT1_1763(.VSS(VSS),.VDD(VDD),.Y(I7236),.A(g3219));
  NOT NOT1_1764(.VSS(VSS),.VDD(VDD),.Y(I15635),.A(g10185));
  NOT NOT1_1765(.VSS(VSS),.VDD(VDD),.Y(I16982),.A(g11088));
  NOT NOT1_1766(.VSS(VSS),.VDD(VDD),.Y(g8599),.A(g8546));
  NOT NOT1_1767(.VSS(VSS),.VDD(VDD),.Y(g7995),.A(I12817));
  NOT NOT1_1768(.VSS(VSS),.VDD(VDD),.Y(g2790),.A(g2276));
  NOT NOT1_1769(.VSS(VSS),.VDD(VDD),.Y(g11408),.A(I17265));
  NOT NOT1_1770(.VSS(VSS),.VDD(VDD),.Y(g7079),.A(I11312));
  NOT NOT1_1771(.VSS(VSS),.VDD(VDD),.Y(g11635),.A(I17719));
  NOT NOT1_1772(.VSS(VSS),.VDD(VDD),.Y(I11778),.A(g7210));
  NOT NOT1_1773(.VSS(VSS),.VDD(VDD),.Y(g3903),.A(I7070));
  NOT NOT1_1774(.VSS(VSS),.VDD(VDD),.Y(g5012),.A(I8388));
  NOT NOT1_1775(.VSS(VSS),.VDD(VDD),.Y(g9100),.A(g8892));
  NOT NOT1_1776(.VSS(VSS),.VDD(VDD),.Y(g8274),.A(I13194));
  NOT NOT1_1777(.VSS(VSS),.VDD(VDD),.Y(I10427),.A(g5839));
  NOT NOT1_1778(.VSS(VSS),.VDD(VDD),.Y(g7479),.A(I11873));
  NOT NOT1_1779(.VSS(VSS),.VDD(VDD),.Y(g8426),.A(I13592));
  NOT NOT1_1780(.VSS(VSS),.VDD(VDD),.Y(g1994),.A(g794));
  NOT NOT1_1781(.VSS(VSS),.VDD(VDD),.Y(g4445),.A(I7803));
  NOT NOT1_1782(.VSS(VSS),.VDD(VDD),.Y(g6253),.A(I10018));
  NOT NOT1_1783(.VSS(VSS),.VDD(VDD),.Y(g2061),.A(g1828));
  NOT NOT1_1784(.VSS(VSS),.VDD(VDD),.Y(g2187),.A(g746));
  NOT NOT1_1785(.VSS(VSS),.VDD(VDD),.Y(g6938),.A(I11068));
  NOT NOT1_1786(.VSS(VSS),.VDD(VDD),.Y(g4173),.A(I7336));
  NOT NOT1_1787(.VSS(VSS),.VDD(VDD),.Y(g6813),.A(I10849));
  NOT NOT1_1788(.VSS(VSS),.VDD(VDD),.Y(g4373),.A(I7680));
  NOT NOT1_1789(.VSS(VSS),.VDD(VDD),.Y(I11786),.A(g7246));
  NOT NOT1_1790(.VSS(VSS),.VDD(VDD),.Y(I16796),.A(g11016));
  NOT NOT1_1791(.VSS(VSS),.VDD(VDD),.Y(g10535),.A(I16172));
  NOT NOT1_1792(.VSS(VSS),.VDD(VDD),.Y(g4491),.A(g3546));
  NOT NOT1_1793(.VSS(VSS),.VDD(VDD),.Y(g8125),.A(I12986));
  NOT NOT1_1794(.VSS(VSS),.VDD(VDD),.Y(g7190),.A(I11412));
  NOT NOT1_1795(.VSS(VSS),.VDD(VDD),.Y(g8325),.A(I13357));
  NOT NOT1_1796(.VSS(VSS),.VDD(VDD),.Y(I11647),.A(g6925));
  NOT NOT1_1797(.VSS(VSS),.VDD(VDD),.Y(g7390),.A(g6847));
  NOT NOT1_1798(.VSS(VSS),.VDD(VDD),.Y(I12878),.A(g7638));
  NOT NOT1_1799(.VSS(VSS),.VDD(VDD),.Y(g5888),.A(g5102));
  NOT NOT1_1800(.VSS(VSS),.VDD(VDD),.Y(I13945),.A(g8488));
  NOT NOT1_1801(.VSS(VSS),.VDD(VDD),.Y(I12171),.A(g6885));
  NOT NOT1_1802(.VSS(VSS),.VDD(VDD),.Y(g10121),.A(I15371));
  NOT NOT1_1803(.VSS(VSS),.VDD(VDD),.Y(g8984),.A(I14373));
  NOT NOT1_1804(.VSS(VSS),.VDD(VDD),.Y(g3436),.A(g3144));
  NOT NOT1_1805(.VSS(VSS),.VDD(VDD),.Y(g4369),.A(I7668));
  NOT NOT1_1806(.VSS(VSS),.VDD(VDD),.Y(g8280),.A(I13212));
  NOT NOT1_1807(.VSS(VSS),.VDD(VDD),.Y(I7556),.A(g4080));
  NOT NOT1_1808(.VSS(VSS),.VDD(VDD),.Y(g4602),.A(I8011));
  NOT NOT1_1809(.VSS(VSS),.VDD(VDD),.Y(g7501),.A(I11879));
  NOT NOT1_1810(.VSS(VSS),.VDD(VDD),.Y(I17450),.A(g11450));
  NOT NOT1_1811(.VSS(VSS),.VDD(VDD),.Y(g3378),.A(I6572));
  NOT NOT1_1812(.VSS(VSS),.VDD(VDD),.Y(g5787),.A(I9383));
  NOT NOT1_1813(.VSS(VSS),.VDD(VDD),.Y(I9424),.A(g4963));
  NOT NOT1_1814(.VSS(VSS),.VDD(VDD),.Y(I9795),.A(g5404));
  NOT NOT1_1815(.VSS(VSS),.VDD(VDD),.Y(I17315),.A(g11393));
  NOT NOT1_1816(.VSS(VSS),.VDD(VDD),.Y(g10344),.A(I15798));
  NOT NOT1_1817(.VSS(VSS),.VDD(VDD),.Y(I9737),.A(g5258));
  NOT NOT1_1818(.VSS(VSS),.VDD(VDD),.Y(g2904),.A(I6065));
  NOT NOT1_1819(.VSS(VSS),.VDD(VDD),.Y(g2200),.A(g92));
  NOT NOT1_1820(.VSS(VSS),.VDD(VDD),.Y(g6552),.A(g5733));
  NOT NOT1_1821(.VSS(VSS),.VDD(VDD),.Y(g7356),.A(I11716));
  NOT NOT1_1822(.VSS(VSS),.VDD(VDD),.Y(g2046),.A(g1845));
  NOT NOT1_1823(.VSS(VSS),.VDD(VDD),.Y(I17707),.A(g11619));
  NOT NOT1_1824(.VSS(VSS),.VDD(VDD),.Y(g4920),.A(I8293));
  NOT NOT1_1825(.VSS(VSS),.VDD(VDD),.Y(I5827),.A(g2271));
  NOT NOT1_1826(.VSS(VSS),.VDD(VDD),.Y(g2446),.A(g1400));
  NOT NOT1_1827(.VSS(VSS),.VDD(VDD),.Y(g4459),.A(I7820));
  NOT NOT1_1828(.VSS(VSS),.VDD(VDD),.Y(I17202),.A(g11322));
  NOT NOT1_1829(.VSS(VSS),.VDD(VDD),.Y(g3335),.A(I6520));
  NOT NOT1_1830(.VSS(VSS),.VDD(VDD),.Y(I13233),.A(g8265));
  NOT NOT1_1831(.VSS(VSS),.VDD(VDD),.Y(g8483),.A(g8332));
  NOT NOT1_1832(.VSS(VSS),.VDD(VDD),.Y(g4767),.A(I8123));
  NOT NOT1_1833(.VSS(VSS),.VDD(VDD),.Y(I7064),.A(g2984));
  NOT NOT1_1834(.VSS(VSS),.VDD(VDD),.Y(g11575),.A(g11561));
  NOT NOT1_1835(.VSS(VSS),.VDD(VDD),.Y(g2003),.A(g822));
  NOT NOT1_1836(.VSS(VSS),.VDD(VDD),.Y(g5281),.A(g4428));
  NOT NOT1_1837(.VSS(VSS),.VDD(VDD),.Y(g3382),.A(I6580));
  NOT NOT1_1838(.VSS(VSS),.VDD(VDD),.Y(I9077),.A(g4765));
  NOT NOT1_1839(.VSS(VSS),.VDD(VDD),.Y(I7899),.A(g3380));
  NOT NOT1_1840(.VSS(VSS),.VDD(VDD),.Y(g4535),.A(g3946));
  NOT NOT1_1841(.VSS(VSS),.VDD(VDD),.Y(I8358),.A(g4794));
  NOT NOT1_1842(.VSS(VSS),.VDD(VDD),.Y(I6611),.A(g2626));
  NOT NOT1_1843(.VSS(VSS),.VDD(VDD),.Y(I8506),.A(g4334));
  NOT NOT1_1844(.VSS(VSS),.VDD(VDD),.Y(g2345),.A(g1936));
  NOT NOT1_1845(.VSS(VSS),.VDD(VDD),.Y(g10173),.A(g10120));
  NOT NOT1_1846(.VSS(VSS),.VDD(VDD),.Y(I17070),.A(g11233));
  NOT NOT1_1847(.VSS(VSS),.VDD(VDD),.Y(g8106),.A(g7950));
  NOT NOT1_1848(.VSS(VSS),.VDD(VDD),.Y(g11109),.A(g10974));
  NOT NOT1_1849(.VSS(VSS),.VDD(VDD),.Y(g8306),.A(I13290));
  NOT NOT1_1850(.VSS(VSS),.VDD(VDD),.Y(g2763),.A(I5847));
  NOT NOT1_1851(.VSS(VSS),.VDD(VDD),.Y(g2191),.A(g1696));
  NOT NOT1_1852(.VSS(VSS),.VDD(VDD),.Y(g2391),.A(I5478));
  NOT NOT1_1853(.VSS(VSS),.VDD(VDD),.Y(g6586),.A(g5949));
  NOT NOT1_1854(.VSS(VSS),.VDD(VDD),.Y(I12919),.A(g8003));
  NOT NOT1_1855(.VSS(VSS),.VDD(VDD),.Y(I6799),.A(g2750));
  NOT NOT1_1856(.VSS(VSS),.VDD(VDD),.Y(I11932),.A(g6908));
  NOT NOT1_1857(.VSS(VSS),.VDD(VDD),.Y(g3749),.A(I6938));
  NOT NOT1_1858(.VSS(VSS),.VDD(VDD),.Y(g8790),.A(I14101));
  NOT NOT1_1859(.VSS(VSS),.VDD(VDD),.Y(I9205),.A(g5309));
  NOT NOT1_1860(.VSS(VSS),.VDD(VDD),.Y(g11108),.A(g10974));
  NOT NOT1_1861(.VSS(VSS),.VDD(VDD),.Y(g2695),.A(g2039));
  NOT NOT1_1862(.VSS(VSS),.VDD(VDD),.Y(g9666),.A(I14793));
  NOT NOT1_1863(.VSS(VSS),.VDD(VDD),.Y(g8061),.A(I12901));
  NOT NOT1_1864(.VSS(VSS),.VDD(VDD),.Y(g5684),.A(I9205));
  NOT NOT1_1865(.VSS(VSS),.VDD(VDD),.Y(I8275),.A(g4351));
  NOT NOT1_1866(.VSS(VSS),.VDD(VDD),.Y(I8311),.A(g4794));
  NOT NOT1_1867(.VSS(VSS),.VDD(VDD),.Y(g4415),.A(g3914));
  NOT NOT1_1868(.VSS(VSS),.VDD(VDD),.Y(g5639),.A(I9080));
  NOT NOT1_1869(.VSS(VSS),.VDD(VDD),.Y(I14127),.A(g8768));
  NOT NOT1_1870(.VSS(VSS),.VDD(VDD),.Y(I17384),.A(g11437));
  NOT NOT1_1871(.VSS(VSS),.VDD(VDD),.Y(g7810),.A(I12595));
  NOT NOT1_1872(.VSS(VSS),.VDD(VDD),.Y(g7363),.A(I11737));
  NOT NOT1_1873(.VSS(VSS),.VDD(VDD),.Y(g10134),.A(I15400));
  NOT NOT1_1874(.VSS(VSS),.VDD(VDD),.Y(I7295),.A(g3260));
  NOT NOT1_1875(.VSS(VSS),.VDD(VDD),.Y(I11961),.A(g7053));
  NOT NOT1_1876(.VSS(VSS),.VDD(VDD),.Y(I16553),.A(g10754));
  NOT NOT1_1877(.VSS(VSS),.VDD(VDD),.Y(g5109),.A(I8495));
  NOT NOT1_1878(.VSS(VSS),.VDD(VDD),.Y(g5791),.A(I9391));
  NOT NOT1_1879(.VSS(VSS),.VDD(VDD),.Y(g3798),.A(g3228));
  NOT NOT1_1880(.VSS(VSS),.VDD(VDD),.Y(I13448),.A(g8150));
  NOT NOT1_1881(.VSS(VSS),.VDD(VDD),.Y(I9099),.A(g5572));
  NOT NOT1_1882(.VSS(VSS),.VDD(VDD),.Y(g2159),.A(I5080));
  NOT NOT1_1883(.VSS(VSS),.VDD(VDD),.Y(g7432),.A(I11824));
  NOT NOT1_1884(.VSS(VSS),.VDD(VDD),.Y(I14490),.A(g8885));
  NOT NOT1_1885(.VSS(VSS),.VDD(VDD),.Y(g6141),.A(I9854));
  NOT NOT1_1886(.VSS(VSS),.VDD(VDD),.Y(g8622),.A(g8485));
  NOT NOT1_1887(.VSS(VSS),.VDD(VDD),.Y(g6570),.A(g5949));
  NOT NOT1_1888(.VSS(VSS),.VDD(VDD),.Y(g6860),.A(g6475));
  NOT NOT1_1889(.VSS(VSS),.VDD(VDD),.Y(g7053),.A(I11238));
  NOT NOT1_1890(.VSS(VSS),.VDD(VDD),.Y(I11505),.A(g6585));
  NOT NOT1_1891(.VSS(VSS),.VDD(VDD),.Y(g9351),.A(I14558));
  NOT NOT1_1892(.VSS(VSS),.VDD(VDD),.Y(I5662),.A(g563));
  NOT NOT1_1893(.VSS(VSS),.VDD(VDD),.Y(g9875),.A(I15036));
  NOT NOT1_1894(.VSS(VSS),.VDD(VDD),.Y(g8427),.A(I13595));
  NOT NOT1_1895(.VSS(VSS),.VDD(VDD),.Y(I5067),.A(g33));
  NOT NOT1_1896(.VSS(VSS),.VDD(VDD),.Y(g9530),.A(I14675));
  NOT NOT1_1897(.VSS(VSS),.VDD(VDD),.Y(g6710),.A(I10693));
  NOT NOT1_1898(.VSS(VSS),.VDD(VDD),.Y(g5808),.A(g5320));
  NOT NOT1_1899(.VSS(VSS),.VDD(VDD),.Y(I5418),.A(g907));
  NOT NOT1_1900(.VSS(VSS),.VDD(VDD),.Y(g2858),.A(I5992));
  NOT NOT1_1901(.VSS(VSS),.VDD(VDD),.Y(I12598),.A(g7628));
  NOT NOT1_1902(.VSS(VSS),.VDD(VDD),.Y(I7194),.A(g2629));
  NOT NOT1_1903(.VSS(VSS),.VDD(VDD),.Y(I14376),.A(g8959));
  NOT NOT1_1904(.VSS(VSS),.VDD(VDD),.Y(I14385),.A(g8890));
  NOT NOT1_1905(.VSS(VSS),.VDD(VDD),.Y(g4203),.A(I7426));
  NOT NOT1_1906(.VSS(VSS),.VDD(VDD),.Y(I8985),.A(g4733));
  NOT NOT1_1907(.VSS(VSS),.VDD(VDD),.Y(I13717),.A(g8354));
  NOT NOT1_1908(.VSS(VSS),.VDD(VDD),.Y(g11381),.A(I17206));
  NOT NOT1_1909(.VSS(VSS),.VDD(VDD),.Y(g4721),.A(g3546));
  NOT NOT1_1910(.VSS(VSS),.VDD(VDD),.Y(g2016),.A(g1361));
  NOT NOT1_1911(.VSS(VSS),.VDD(VDD),.Y(I13212),.A(g8195));
  NOT NOT1_1912(.VSS(VSS),.VDD(VDD),.Y(g2757),.A(I5837));
  NOT NOT1_1913(.VSS(VSS),.VDD(VDD),.Y(g8446),.A(I13636));
  NOT NOT1_1914(.VSS(VSS),.VDD(VDD),.Y(g7568),.A(I12026));
  NOT NOT1_1915(.VSS(VSS),.VDD(VDD),.Y(g5759),.A(I9341));
  NOT NOT1_1916(.VSS(VSS),.VDD(VDD),.Y(I9754),.A(g5271));
  NOT NOT1_1917(.VSS(VSS),.VDD(VDD),.Y(I10888),.A(g6333));
  NOT NOT1_1918(.VSS(VSS),.VDD(VDD),.Y(g8514),.A(I13711));
  NOT NOT1_1919(.VSS(VSS),.VDD(VDD),.Y(I6802),.A(g2751));
  NOT NOT1_1920(.VSS(VSS),.VDD(VDD),.Y(g3632),.A(I6799));
  NOT NOT1_1921(.VSS(VSS),.VDD(VDD),.Y(g3095),.A(g2482));
  NOT NOT1_1922(.VSS(VSS),.VDD(VDD),.Y(g3037),.A(g2135));
  NOT NOT1_1923(.VSS(VSS),.VDD(VDD),.Y(g8003),.A(I12835));
  NOT NOT1_1924(.VSS(VSS),.VDD(VDD),.Y(I14888),.A(g9454));
  NOT NOT1_1925(.VSS(VSS),.VDD(VDD),.Y(I16252),.A(g10515));
  NOT NOT1_1926(.VSS(VSS),.VDD(VDD),.Y(g3437),.A(I6654));
  NOT NOT1_1927(.VSS(VSS),.VDD(VDD),.Y(I12817),.A(g7692));
  NOT NOT1_1928(.VSS(VSS),.VDD(VDD),.Y(I9273),.A(g5091));
  NOT NOT1_1929(.VSS(VSS),.VDD(VDD),.Y(I10671),.A(g6045));
  NOT NOT1_1930(.VSS(VSS),.VDD(VDD),.Y(I17695),.A(g11614));
  NOT NOT1_1931(.VSS(VSS),.VDD(VDD),.Y(g3102),.A(g2482));
  NOT NOT1_1932(.VSS(VSS),.VDD(VDD),.Y(I4924),.A(g123));
  NOT NOT1_1933(.VSS(VSS),.VDD(VDD),.Y(g3208),.A(I6381));
  NOT NOT1_1934(.VSS(VSS),.VDD(VDD),.Y(I12322),.A(g7246));
  NOT NOT1_1935(.VSS(VSS),.VDD(VDD),.Y(g7912),.A(g7651));
  NOT NOT1_1936(.VSS(VSS),.VDD(VDD),.Y(g8145),.A(I13030));
  NOT NOT1_1937(.VSS(VSS),.VDD(VDD),.Y(g8345),.A(I13415));
  NOT NOT1_1938(.VSS(VSS),.VDD(VDD),.Y(g2251),.A(g731));
  NOT NOT1_1939(.VSS(VSS),.VDD(VDD),.Y(g2642),.A(g1988));
  NOT NOT1_1940(.VSS(VSS),.VDD(VDD),.Y(I12159),.A(g7243));
  NOT NOT1_1941(.VSS(VSS),.VDD(VDD),.Y(g7357),.A(I11719));
  NOT NOT1_1942(.VSS(VSS),.VDD(VDD),.Y(g2047),.A(g1857));
  NOT NOT1_1943(.VSS(VSS),.VDD(VDD),.Y(I12532),.A(g7594));
  NOT NOT1_1944(.VSS(VSS),.VDD(VDD),.Y(I12901),.A(g7984));
  NOT NOT1_1945(.VSS(VSS),.VDD(VDD),.Y(g8191),.A(I13114));
  NOT NOT1_1946(.VSS(VSS),.VDD(VDD),.Y(g10927),.A(g10827));
  NOT NOT1_1947(.VSS(VSS),.VDD(VDD),.Y(g9884),.A(I15063));
  NOT NOT1_1948(.VSS(VSS),.VDD(VDD),.Y(g6158),.A(I9883));
  NOT NOT1_1949(.VSS(VSS),.VDD(VDD),.Y(g3719),.A(g2920));
  NOT NOT1_1950(.VSS(VSS),.VDD(VDD),.Y(I12783),.A(g7590));
  NOT NOT1_1951(.VSS(VSS),.VDD(VDD),.Y(g11390),.A(I17219));
  NOT NOT1_1952(.VSS(VSS),.VDD(VDD),.Y(I13723),.A(g8359));
  NOT NOT1_1953(.VSS(VSS),.VDD(VDD),.Y(g5865),.A(I9486));
  NOT NOT1_1954(.VSS(VSS),.VDD(VDD),.Y(g8695),.A(I13978));
  NOT NOT1_1955(.VSS(VSS),.VDD(VDD),.Y(I5847),.A(g2275));
  NOT NOT1_1956(.VSS(VSS),.VDD(VDD),.Y(I6901),.A(g2818));
  NOT NOT1_1957(.VSS(VSS),.VDD(VDD),.Y(I11149),.A(g6468));
  NOT NOT1_1958(.VSS(VSS),.VDD(VDD),.Y(g2874),.A(I6022));
  NOT NOT1_1959(.VSS(VSS),.VDD(VDD),.Y(g7929),.A(g7519));
  NOT NOT1_1960(.VSS(VSS),.VDD(VDD),.Y(g3752),.A(I6947));
  NOT NOT1_1961(.VSS(VSS),.VDD(VDD),.Y(I16673),.A(g10782));
  NOT NOT1_1962(.VSS(VSS),.VDD(VDD),.Y(I11433),.A(g6424));
  NOT NOT1_1963(.VSS(VSS),.VDD(VDD),.Y(I16847),.A(g10886));
  NOT NOT1_1964(.VSS(VSS),.VDD(VDD),.Y(I11387),.A(g6672));
  NOT NOT1_1965(.VSS(VSS),.VDD(VDD),.Y(g5604),.A(I9032));
  NOT NOT1_1966(.VSS(VSS),.VDD(VDD),.Y(I13433),.A(g8181));
  NOT NOT1_1967(.VSS(VSS),.VDD(VDD),.Y(g5098),.A(g4840));
  NOT NOT1_1968(.VSS(VSS),.VDD(VDD),.Y(g2654),.A(g2012));
  NOT NOT1_1969(.VSS(VSS),.VDD(VDD),.Y(I11620),.A(g6840));
  NOT NOT1_1970(.VSS(VSS),.VDD(VDD),.Y(g4188),.A(I7381));
  NOT NOT1_1971(.VSS(VSS),.VDD(VDD),.Y(g5498),.A(I8919));
  NOT NOT1_1972(.VSS(VSS),.VDD(VDD),.Y(I9712),.A(g5230));
  NOT NOT1_1973(.VSS(VSS),.VDD(VDD),.Y(g6587),.A(g5827));
  NOT NOT1_1974(.VSS(VSS),.VDD(VDD),.Y(g4388),.A(I7719));
  NOT NOT1_1975(.VSS(VSS),.VDD(VDD),.Y(g10491),.A(I16108));
  NOT NOT1_1976(.VSS(VSS),.VDD(VDD),.Y(g10903),.A(g10809));
  NOT NOT1_1977(.VSS(VSS),.VDD(VDD),.Y(I11097),.A(g6748));
  NOT NOT1_1978(.VSS(VSS),.VDD(VDD),.Y(I5421),.A(g549));
  NOT NOT1_1979(.VSS(VSS),.VDD(VDD),.Y(g8359),.A(I13457));
  NOT NOT1_1980(.VSS(VSS),.VDD(VDD),.Y(g6111),.A(I9786));
  NOT NOT1_1981(.VSS(VSS),.VDD(VDD),.Y(g6275),.A(I10084));
  NOT NOT1_1982(.VSS(VSS),.VDD(VDD),.Y(g6311),.A(I10192));
  NOT NOT1_1983(.VSS(VSS),.VDD(VDD),.Y(g4216),.A(I7465));
  NOT NOT1_1984(.VSS(VSS),.VDD(VDD),.Y(g10604),.A(I16280));
  NOT NOT1_1985(.VSS(VSS),.VDD(VDD),.Y(g9343),.A(I14534));
  NOT NOT1_1986(.VSS(VSS),.VDD(VDD),.Y(g8858),.A(g8743));
  NOT NOT1_1987(.VSS(VSS),.VDD(VDD),.Y(g4671),.A(g3354));
  NOT NOT1_1988(.VSS(VSS),.VDD(VDD),.Y(g2880),.A(I6028));
  NOT NOT1_1989(.VSS(VSS),.VDD(VDD),.Y(g4428),.A(I7776));
  NOT NOT1_1990(.VSS(VSS),.VDD(VDD),.Y(g2537),.A(I5646));
  NOT NOT1_1991(.VSS(VSS),.VDD(VDD),.Y(I10546),.A(g5914));
  NOT NOT1_1992(.VSS(VSS),.VDD(VDD),.Y(g5896),.A(I9525));
  NOT NOT1_1993(.VSS(VSS),.VDD(VDD),.Y(g4430),.A(I7782));
  NOT NOT1_1994(.VSS(VSS),.VDD(VDD),.Y(I14546),.A(g9312));
  NOT NOT1_1995(.VSS(VSS),.VDD(VDD),.Y(I7438),.A(g3461));
  NOT NOT1_1996(.VSS(VSS),.VDD(VDD),.Y(g3164),.A(I6370));
  NOT NOT1_1997(.VSS(VSS),.VDD(VDD),.Y(g3364),.A(g3121));
  NOT NOT1_1998(.VSS(VSS),.VDD(VDD),.Y(I7009),.A(g2913));
  NOT NOT1_1999(.VSS(VSS),.VDD(VDD),.Y(I10024),.A(g5700));
  NOT NOT1_2000(.VSS(VSS),.VDD(VDD),.Y(I8204),.A(g3976));
  NOT NOT1_2001(.VSS(VSS),.VDD(VDD),.Y(I12631),.A(g7705));
  NOT NOT1_2002(.VSS(VSS),.VDD(VDD),.Y(g8115),.A(g7953));
  NOT NOT1_2003(.VSS(VSS),.VDD(VDD),.Y(g4564),.A(g3880));
  NOT NOT1_2004(.VSS(VSS),.VDD(VDD),.Y(g8251),.A(I13166));
  NOT NOT1_2005(.VSS(VSS),.VDD(VDD),.Y(g8315),.A(I13329));
  NOT NOT1_2006(.VSS(VSS),.VDD(VDD),.Y(g2612),.A(I5737));
  NOT NOT1_2007(.VSS(VSS),.VDD(VDD),.Y(I15326),.A(g10025));
  NOT NOT1_2008(.VSS(VSS),.VDD(VDD),.Y(g2017),.A(g1218));
  NOT NOT1_2009(.VSS(VSS),.VDD(VDD),.Y(g6284),.A(I10111));
  NOT NOT1_2010(.VSS(VSS),.VDD(VDD),.Y(g2243),.A(I5248));
  NOT NOT1_2011(.VSS(VSS),.VDD(VDD),.Y(g8447),.A(I13639));
  NOT NOT1_2012(.VSS(VSS),.VDD(VDD),.Y(I6580),.A(g3186));
  NOT NOT1_2013(.VSS(VSS),.VDD(VDD),.Y(g3770),.A(I6985));
  NOT NOT1_2014(.VSS(VSS),.VDD(VDD),.Y(g6239),.A(I9988));
  NOT NOT1_2015(.VSS(VSS),.VDD(VDD),.Y(g10794),.A(I16496));
  NOT NOT1_2016(.VSS(VSS),.VDD(VDD),.Y(I15536),.A(g10111));
  NOT NOT1_2017(.VSS(VSS),.VDD(VDD),.Y(g10395),.A(g10320));
  NOT NOT1_2018(.VSS(VSS),.VDD(VDD),.Y(g5419),.A(I8858));
  NOT NOT1_2019(.VSS(VSS),.VDD(VDD),.Y(g9804),.A(I14939));
  NOT NOT1_2020(.VSS(VSS),.VDD(VDD),.Y(g10262),.A(g10142));
  NOT NOT1_2021(.VSS(VSS),.VDD(VDD),.Y(g7683),.A(g7148));
  NOT NOT1_2022(.VSS(VSS),.VDD(VDD),.Y(g11040),.A(I16781));
  NOT NOT1_2023(.VSS(VSS),.VDD(VDD),.Y(g10899),.A(g10803));
  NOT NOT1_2024(.VSS(VSS),.VDD(VDD),.Y(g6591),.A(I10553));
  NOT NOT1_2025(.VSS(VSS),.VDD(VDD),.Y(I11412),.A(g6411));
  NOT NOT1_2026(.VSS(VSS),.VDD(VDD),.Y(g5052),.A(g4394));
  NOT NOT1_2027(.VSS(VSS),.VDD(VDD),.Y(I13412),.A(g8142));
  NOT NOT1_2028(.VSS(VSS),.VDD(VDD),.Y(I5101),.A(g1960));
  NOT NOT1_2029(.VSS(VSS),.VDD(VDD),.Y(g8874),.A(I14194));
  NOT NOT1_2030(.VSS(VSS),.VDD(VDD),.Y(g3532),.A(g3164));
  NOT NOT1_2031(.VSS(VSS),.VDD(VDD),.Y(g7778),.A(I12499));
  NOT NOT1_2032(.VSS(VSS),.VDD(VDD),.Y(g2234),.A(g87));
  NOT NOT1_2033(.VSS(VSS),.VDD(VDD),.Y(g6853),.A(I10917));
  NOT NOT1_2034(.VSS(VSS),.VDD(VDD),.Y(I10126),.A(g5682));
  NOT NOT1_2035(.VSS(VSS),.VDD(VDD),.Y(I10659),.A(g6038));
  NOT NOT1_2036(.VSS(VSS),.VDD(VDD),.Y(I16574),.A(g10821));
  NOT NOT1_2037(.VSS(VSS),.VDD(VDD),.Y(g2629),.A(g2001));
  NOT NOT1_2038(.VSS(VSS),.VDD(VDD),.Y(g4638),.A(g3354));
  NOT NOT1_2039(.VSS(VSS),.VDD(VDD),.Y(g2328),.A(g1882));
  NOT NOT1_2040(.VSS(VSS),.VDD(VDD),.Y(I12289),.A(g7142));
  NOT NOT1_2041(.VSS(VSS),.VDD(VDD),.Y(I6968),.A(g2881));
  NOT NOT1_2042(.VSS(VSS),.VDD(VDD),.Y(g6420),.A(I10334));
  NOT NOT1_2043(.VSS(VSS),.VDD(VDD),.Y(g11621),.A(I17681));
  NOT NOT1_2044(.VSS(VSS),.VDD(VDD),.Y(g2130),.A(I5057));
  NOT NOT1_2045(.VSS(VSS),.VDD(VDD),.Y(g10191),.A(I15551));
  NOT NOT1_2046(.VSS(VSS),.VDD(VDD),.Y(g2542),.A(g1868));
  NOT NOT1_2047(.VSS(VSS),.VDD(VDD),.Y(I8973),.A(g4488));
  NOT NOT1_2048(.VSS(VSS),.VDD(VDD),.Y(g2330),.A(g1891));
  NOT NOT1_2049(.VSS(VSS),.VDD(VDD),.Y(g7735),.A(I12384));
  NOT NOT1_2050(.VSS(VSS),.VDD(VDD),.Y(I16311),.A(g10584));
  NOT NOT1_2051(.VSS(VSS),.VDD(VDD),.Y(g4308),.A(g3863));
  NOT NOT1_2052(.VSS(VSS),.VDD(VDD),.Y(I11228),.A(g6471));
  NOT NOT1_2053(.VSS(VSS),.VDD(VDD),.Y(I17231),.A(g11303));
  NOT NOT1_2054(.VSS(VSS),.VDD(VDD),.Y(g7782),.A(I12511));
  NOT NOT1_2055(.VSS(VSS),.VDD(VDD),.Y(g6559),.A(g5758));
  NOT NOT1_2056(.VSS(VSS),.VDD(VDD),.Y(I12571),.A(g7509));
  NOT NOT1_2057(.VSS(VSS),.VDD(VDD),.Y(g3012),.A(I6247));
  NOT NOT1_2058(.VSS(VSS),.VDD(VDD),.Y(I11011),.A(g6340));
  NOT NOT1_2059(.VSS(VSS),.VDD(VDD),.Y(I5751),.A(g2296));
  NOT NOT1_2060(.VSS(VSS),.VDD(VDD),.Y(g8595),.A(I13840));
  NOT NOT1_2061(.VSS(VSS),.VDD(VDD),.Y(g6931),.A(I11055));
  NOT NOT1_2062(.VSS(VSS),.VDD(VDD),.Y(g5728),.A(I9276));
  NOT NOT1_2063(.VSS(VSS),.VDD(VDD),.Y(g5486),.A(g4395));
  NOT NOT1_2064(.VSS(VSS),.VDD(VDD),.Y(I10296),.A(g6242));
  NOT NOT1_2065(.VSS(VSS),.VDD(VDD),.Y(I11716),.A(g7026));
  NOT NOT1_2066(.VSS(VSS),.VDD(VDD),.Y(g5730),.A(I9282));
  NOT NOT1_2067(.VSS(VSS),.VDD(VDD),.Y(g5504),.A(g4419));
  NOT NOT1_2068(.VSS(VSS),.VDD(VDD),.Y(g7949),.A(g7422));
  NOT NOT1_2069(.VSS(VSS),.VDD(VDD),.Y(g4217),.A(I7468));
  NOT NOT1_2070(.VSS(VSS),.VDD(VDD),.Y(g11183),.A(I16950));
  NOT NOT1_2071(.VSS(VSS),.VDD(VDD),.Y(I8123),.A(g3630));
  NOT NOT1_2072(.VSS(VSS),.VDD(VDD),.Y(g3990),.A(g3121));
  NOT NOT1_2073(.VSS(VSS),.VDD(VDD),.Y(g2554),.A(I5672));
  NOT NOT1_2074(.VSS(VSS),.VDD(VDD),.Y(g4758),.A(g3586));
  NOT NOT1_2075(.VSS(VSS),.VDD(VDD),.Y(g4066),.A(I7191));
  NOT NOT1_2076(.VSS(VSS),.VDD(VDD),.Y(g8272),.A(I13188));
  NOT NOT1_2077(.VSS(VSS),.VDD(VDD),.Y(I16592),.A(g10781));
  NOT NOT1_2078(.VSS(VSS),.VDD(VDD),.Y(g4589),.A(I7996));
  NOT NOT1_2079(.VSS(VSS),.VDD(VDD),.Y(g5185),.A(g4682));
  NOT NOT1_2080(.VSS(VSS),.VDD(VDD),.Y(g11397),.A(I17234));
  NOT NOT1_2081(.VSS(VSS),.VDD(VDD),.Y(g5881),.A(g5361));
  NOT NOT1_2082(.VSS(VSS),.VDD(VDD),.Y(g7627),.A(I12223));
  NOT NOT1_2083(.VSS(VSS),.VDD(VDD),.Y(g9094),.A(g8892));
  NOT NOT1_2084(.VSS(VSS),.VDD(VDD),.Y(I5041),.A(g1179));
  NOT NOT1_2085(.VSS(VSS),.VDD(VDD),.Y(I9135),.A(g5198));
  NOT NOT1_2086(.VSS(VSS),.VDD(VDD),.Y(g4466),.A(I7833));
  NOT NOT1_2087(.VSS(VSS),.VDD(VDD),.Y(g1992),.A(g782));
  NOT NOT1_2088(.VSS(VSS),.VDD(VDD),.Y(g6905),.A(I11011));
  NOT NOT1_2089(.VSS(VSS),.VDD(VDD),.Y(g8978),.A(I14355));
  NOT NOT1_2090(.VSS(VSS),.VDD(VDD),.Y(I5441),.A(g919));
  NOT NOT1_2091(.VSS(VSS),.VDD(VDD),.Y(g3371),.A(g2837));
  NOT NOT1_2092(.VSS(VSS),.VDD(VDD),.Y(g11062),.A(g10937));
  NOT NOT1_2093(.VSS(VSS),.VDD(VDD),.Y(I10060),.A(g5752));
  NOT NOT1_2094(.VSS(VSS),.VDD(VDD),.Y(g2213),.A(g1110));
  NOT NOT1_2095(.VSS(VSS),.VDD(VDD),.Y(g11509),.A(I17546));
  NOT NOT1_2096(.VSS(VSS),.VDD(VDD),.Y(g7998),.A(I12822));
  NOT NOT1_2097(.VSS(VSS),.VDD(VDD),.Y(g10247),.A(I15639));
  NOT NOT1_2098(.VSS(VSS),.VDD(VDD),.Y(g4165),.A(g3164));
  NOT NOT1_2099(.VSS(VSS),.VDD(VDD),.Y(g4365),.A(g3880));
  NOT NOT1_2100(.VSS(VSS),.VDD(VDD),.Y(I13627),.A(g8326));
  NOT NOT1_2101(.VSS(VSS),.VDD(VDD),.Y(g5425),.A(g4300));
  NOT NOT1_2102(.VSS(VSS),.VDD(VDD),.Y(g10389),.A(g10307));
  NOT NOT1_2103(.VSS(VSS),.VDD(VDD),.Y(g10926),.A(g10827));
  NOT NOT1_2104(.VSS(VSS),.VDD(VDD),.Y(I10855),.A(g6685));
  NOT NOT1_2105(.VSS(VSS),.VDD(VDD),.Y(I13959),.A(g8451));
  NOT NOT1_2106(.VSS(VSS),.VDD(VDD),.Y(I13379),.A(g8133));
  NOT NOT1_2107(.VSS(VSS),.VDD(VDD),.Y(g11508),.A(I17543));
  NOT NOT1_2108(.VSS(VSS),.VDD(VDD),.Y(g4711),.A(I8061));
  NOT NOT1_2109(.VSS(VSS),.VDD(VDD),.Y(g6100),.A(I9759));
  NOT NOT1_2110(.VSS(VSS),.VDD(VDD),.Y(I11112),.A(g6445));
  NOT NOT1_2111(.VSS(VSS),.VDD(VDD),.Y(g8982),.A(I14367));
  NOT NOT1_2112(.VSS(VSS),.VDD(VDD),.Y(g11634),.A(I17716));
  NOT NOT1_2113(.VSS(VSS),.VDD(VDD),.Y(g10612),.A(I16286));
  NOT NOT1_2114(.VSS(VSS),.VDD(VDD),.Y(g6300),.A(I10159));
  NOT NOT1_2115(.VSS(VSS),.VDD(VDD),.Y(g7603),.A(I12159));
  NOT NOT1_2116(.VSS(VSS),.VDD(VDD),.Y(g4055),.A(g3144));
  NOT NOT1_2117(.VSS(VSS),.VDD(VDD),.Y(g7039),.A(I11204));
  NOT NOT1_2118(.VSS(VSS),.VDD(VDD),.Y(I9749),.A(g5266));
  NOT NOT1_2119(.VSS(VSS),.VDD(VDD),.Y(g10388),.A(g10305));
  NOT NOT1_2120(.VSS(VSS),.VDD(VDD),.Y(I8351),.A(g4794));
  NOT NOT1_2121(.VSS(VSS),.VDD(VDD),.Y(g8234),.A(g7826));
  NOT NOT1_2122(.VSS(VSS),.VDD(VDD),.Y(g2902),.A(I6061));
  NOT NOT1_2123(.VSS(VSS),.VDD(VDD),.Y(g7439),.A(I11833));
  NOT NOT1_2124(.VSS(VSS),.VDD(VDD),.Y(g8128),.A(I12993));
  NOT NOT1_2125(.VSS(VSS),.VDD(VDD),.Y(g8328),.A(I13364));
  NOT NOT1_2126(.VSS(VSS),.VDD(VDD),.Y(g7850),.A(I12647));
  NOT NOT1_2127(.VSS(VSS),.VDD(VDD),.Y(g10534),.A(I16169));
  NOT NOT1_2128(.VSS(VSS),.VDD(VDD),.Y(g10098),.A(I15332));
  NOT NOT1_2129(.VSS(VSS),.VDD(VDD),.Y(I17456),.A(g11453));
  NOT NOT1_2130(.VSS(VSS),.VDD(VDD),.Y(g4333),.A(g4144));
  NOT NOT1_2131(.VSS(VSS),.VDD(VDD),.Y(I7837),.A(g4158));
  NOT NOT1_2132(.VSS(VSS),.VDD(VDD),.Y(g8330),.A(I13370));
  NOT NOT1_2133(.VSS(VSS),.VDD(VDD),.Y(g10251),.A(g10195));
  NOT NOT1_2134(.VSS(VSS),.VDD(VDD),.Y(g10272),.A(g10168));
  NOT NOT1_2135(.VSS(VSS),.VDD(VDD),.Y(g2090),.A(I4920));
  NOT NOT1_2136(.VSS(VSS),.VDD(VDD),.Y(g4774),.A(I8136));
  NOT NOT1_2137(.VSS(VSS),.VDD(VDD),.Y(I7462),.A(g3721));
  NOT NOT1_2138(.VSS(VSS),.VDD(VDD),.Y(I9798),.A(g5415));
  NOT NOT1_2139(.VSS(VSS),.VDD(VDD),.Y(I13096),.A(g7925));
  NOT NOT1_2140(.VSS(VSS),.VDD(VDD),.Y(g2166),.A(I5101));
  NOT NOT1_2141(.VSS(VSS),.VDD(VDD),.Y(g6750),.A(I10759));
  NOT NOT1_2142(.VSS(VSS),.VDD(VDD),.Y(g9264),.A(I14477));
  NOT NOT1_2143(.VSS(VSS),.VDD(VDD),.Y(I6424),.A(g2462));
  NOT NOT1_2144(.VSS(VSS),.VDD(VDD),.Y(g7702),.A(g7079));
  NOT NOT1_2145(.VSS(VSS),.VDD(VDD),.Y(g4196),.A(I7405));
  NOT NOT1_2146(.VSS(VSS),.VDD(VDD),.Y(g5678),.A(I9191));
  NOT NOT1_2147(.VSS(VSS),.VDD(VDD),.Y(I10503),.A(g5858));
  NOT NOT1_2148(.VSS(VSS),.VDD(VDD),.Y(I16413),.A(g10663));
  NOT NOT1_2149(.VSS(VSS),.VDD(VDD),.Y(g10462),.A(I15977));
  NOT NOT1_2150(.VSS(VSS),.VDD(VDD),.Y(g4396),.A(I7735));
  NOT NOT1_2151(.VSS(VSS),.VDD(VDD),.Y(g3138),.A(I6356));
  NOT NOT1_2152(.VSS(VSS),.VDD(VDD),.Y(g8800),.A(I14123));
  NOT NOT1_2153(.VSS(VSS),.VDD(VDD),.Y(I14503),.A(g8920));
  NOT NOT1_2154(.VSS(VSS),.VDD(VDD),.Y(I8410),.A(g4283));
  NOT NOT1_2155(.VSS(VSS),.VDD(VDD),.Y(g2056),.A(I4859));
  NOT NOT1_2156(.VSS(VSS),.VDD(VDD),.Y(I16691),.A(g10788));
  NOT NOT1_2157(.VSS(VSS),.VDD(VDD),.Y(g9360),.A(I14579));
  NOT NOT1_2158(.VSS(VSS),.VDD(VDD),.Y(g3109),.A(g2482));
  NOT NOT1_2159(.VSS(VSS),.VDD(VDD),.Y(g3791),.A(I7014));
  NOT NOT1_2160(.VSS(VSS),.VDD(VDD),.Y(g2456),.A(g1397));
  NOT NOT1_2161(.VSS(VSS),.VDD(VDD),.Y(g7919),.A(g7512));
  NOT NOT1_2162(.VSS(VSS),.VDD(VDD),.Y(g10032),.A(I15232));
  NOT NOT1_2163(.VSS(VSS),.VDD(VDD),.Y(g2529),.A(I5638));
  NOT NOT1_2164(.VSS(VSS),.VDD(VDD),.Y(g2649),.A(g2005));
  NOT NOT1_2165(.VSS(VSS),.VDD(VDD),.Y(g10140),.A(I15418));
  NOT NOT1_2166(.VSS(VSS),.VDD(VDD),.Y(g4780),.A(g3440));
  NOT NOT1_2167(.VSS(VSS),.VDD(VDD),.Y(I8839),.A(g4484));
  NOT NOT1_2168(.VSS(VSS),.VDD(VDD),.Y(g6040),.A(I9655));
  NOT NOT1_2169(.VSS(VSS),.VDD(VDD),.Y(g2348),.A(I5418));
  NOT NOT1_2170(.VSS(VSS),.VDD(VDD),.Y(I6077),.A(g2349));
  NOT NOT1_2171(.VSS(VSS),.VDD(VDD),.Y(g11574),.A(g11561));
  NOT NOT1_2172(.VSS(VSS),.VDD(VDD),.Y(g11452),.A(I17413));
  NOT NOT1_2173(.VSS(VSS),.VDD(VDD),.Y(g11047),.A(I16802));
  NOT NOT1_2174(.VSS(VSS),.VDD(VDD),.Y(g5682),.A(I9199));
  NOT NOT1_2175(.VSS(VSS),.VDD(VDD),.Y(g5766),.A(I9346));
  NOT NOT1_2176(.VSS(VSS),.VDD(VDD),.Y(g5105),.A(I8487));
  NOT NOT1_2177(.VSS(VSS),.VDD(VDD),.Y(g4509),.A(I7906));
  NOT NOT1_2178(.VSS(VSS),.VDD(VDD),.Y(g6440),.A(g6150));
  NOT NOT1_2179(.VSS(VSS),.VDD(VDD),.Y(g1976),.A(g643));
  NOT NOT1_2180(.VSS(VSS),.VDD(VDD),.Y(g11205),.A(g11112));
  NOT NOT1_2181(.VSS(VSS),.VDD(VDD),.Y(I6477),.A(g2069));
  NOT NOT1_2182(.VSS(VSS),.VDD(VDD),.Y(I9632),.A(g5557));
  NOT NOT1_2183(.VSS(VSS),.VDD(VDD),.Y(g7952),.A(g7427));
  NOT NOT1_2184(.VSS(VSS),.VDD(VDD),.Y(I15311),.A(g10013));
  NOT NOT1_2185(.VSS(VSS),.VDD(VDD),.Y(g9450),.A(g9097));
  NOT NOT1_2186(.VSS(VSS),.VDD(VDD),.Y(g5305),.A(g4378));
  NOT NOT1_2187(.VSS(VSS),.VDD(VDD),.Y(g5801),.A(g5320));
  NOT NOT1_2188(.VSS(VSS),.VDD(VDD),.Y(I5734),.A(g2097));
  NOT NOT1_2189(.VSS(VSS),.VDD(VDD),.Y(I6523),.A(g2819));
  NOT NOT1_2190(.VSS(VSS),.VDD(VDD),.Y(g2155),.A(I5070));
  NOT NOT1_2191(.VSS(VSS),.VDD(VDD),.Y(I4820),.A(g865));
  NOT NOT1_2192(.VSS(VSS),.VDD(VDD),.Y(I17243),.A(g11396));
  NOT NOT1_2193(.VSS(VSS),.VDD(VDD),.Y(g2355),.A(I5435));
  NOT NOT1_2194(.VSS(VSS),.VDD(VDD),.Y(g2851),.A(I5979));
  NOT NOT1_2195(.VSS(VSS),.VDD(VDD),.Y(I7249),.A(g2833));
  NOT NOT1_2196(.VSS(VSS),.VDD(VDD),.Y(I12559),.A(g7477));
  NOT NOT1_2197(.VSS(VSS),.VDD(VDD),.Y(I14315),.A(g8815));
  NOT NOT1_2198(.VSS(VSS),.VDD(VDD),.Y(I6643),.A(g3008));
  NOT NOT1_2199(.VSS(VSS),.VDD(VDD),.Y(g8213),.A(g7826));
  NOT NOT1_2200(.VSS(VSS),.VDD(VDD),.Y(I10819),.A(g6706));
  NOT NOT1_2201(.VSS(VSS),.VDD(VDD),.Y(g11311),.A(I17100));
  NOT NOT1_2202(.VSS(VSS),.VDD(VDD),.Y(I10910),.A(g6703));
  NOT NOT1_2203(.VSS(VSS),.VDD(VDD),.Y(I12424),.A(g7635));
  NOT NOT1_2204(.VSS(VSS),.VDD(VDD),.Y(I9102),.A(g5586));
  NOT NOT1_2205(.VSS(VSS),.VDD(VDD),.Y(I9208),.A(g5047));
  NOT NOT1_2206(.VSS(VSS),.VDD(VDD),.Y(g3707),.A(g2920));
  NOT NOT1_2207(.VSS(VSS),.VDD(VDD),.Y(I9302),.A(g5576));
  NOT NOT1_2208(.VSS(VSS),.VDD(VDD),.Y(I14910),.A(g9532));
  NOT NOT1_2209(.VSS(VSS),.VDD(VDD),.Y(g7616),.A(I12196));
  NOT NOT1_2210(.VSS(VSS),.VDD(VDD),.Y(g7561),.A(I12015));
  NOT NOT1_2211(.VSS(VSS),.VDD(VDD),.Y(g4067),.A(I7194));
  NOT NOT1_2212(.VSS(VSS),.VDD(VDD),.Y(g3759),.A(I6958));
  NOT NOT1_2213(.VSS(VSS),.VDD(VDD),.Y(I8278),.A(g4495));
  NOT NOT1_2214(.VSS(VSS),.VDD(VDD),.Y(I14257),.A(g8805));
  NOT NOT1_2215(.VSS(VSS),.VDD(VDD),.Y(g5748),.A(I9320));
  NOT NOT1_2216(.VSS(VSS),.VDD(VDD),.Y(I10979),.A(g6565));
  NOT NOT1_2217(.VSS(VSS),.VDD(VDD),.Y(g2964),.A(I6193));
  NOT NOT1_2218(.VSS(VSS),.VDD(VDD),.Y(g4418),.A(I7760));
  NOT NOT1_2219(.VSS(VSS),.VDD(VDD),.Y(I9869),.A(g5405));
  NOT NOT1_2220(.VSS(VSS),.VDD(VDD),.Y(g4467),.A(g3829));
  NOT NOT1_2221(.VSS(VSS),.VDD(VDD),.Y(I15072),.A(g9713));
  NOT NOT1_2222(.VSS(VSS),.VDD(VDD),.Y(I14979),.A(g9671));
  NOT NOT1_2223(.VSS(VSS),.VDD(VDD),.Y(g4290),.A(g3586));
  NOT NOT1_2224(.VSS(VSS),.VDD(VDD),.Y(I10111),.A(g5754));
  NOT NOT1_2225(.VSS(VSS),.VDD(VDD),.Y(I14055),.A(g8650));
  NOT NOT1_2226(.VSS(VSS),.VDD(VDD),.Y(g10871),.A(I16583));
  NOT NOT1_2227(.VSS(VSS),.VDD(VDD),.Y(g11051),.A(I16814));
  NOT NOT1_2228(.VSS(VSS),.VDD(VDD),.Y(I5992),.A(g2195));
  NOT NOT1_2229(.VSS(VSS),.VDD(VDD),.Y(g7004),.A(I11143));
  NOT NOT1_2230(.VSS(VSS),.VDD(VDD),.Y(I16583),.A(g10848));
  NOT NOT1_2231(.VSS(VSS),.VDD(VDD),.Y(g11072),.A(g10913));
  NOT NOT1_2232(.VSS(VSS),.VDD(VDD),.Y(I17773),.A(g11650));
  NOT NOT1_2233(.VSS(VSS),.VDD(VDD),.Y(I15592),.A(g10163));
  NOT NOT1_2234(.VSS(VSS),.VDD(VDD),.Y(I15756),.A(g10266));
  NOT NOT1_2235(.VSS(VSS),.VDD(VDD),.Y(g7527),.A(g7148));
  NOT NOT1_2236(.VSS(VSS),.VDD(VDD),.Y(I17268),.A(g11351));
  NOT NOT1_2237(.VSS(VSS),.VDD(VDD),.Y(I6742),.A(g3326));
  NOT NOT1_2238(.VSS(VSS),.VDD(VDD),.Y(I12544),.A(g7669));
  NOT NOT1_2239(.VSS(VSS),.VDD(VDD),.Y(g4093),.A(g2965));
  NOT NOT1_2240(.VSS(VSS),.VDD(VDD),.Y(I8282),.A(g4770));
  NOT NOT1_2241(.VSS(VSS),.VDD(VDD),.Y(g6151),.A(I9872));
  NOT NOT1_2242(.VSS(VSS),.VDD(VDD),.Y(g7764),.A(I12457));
  NOT NOT1_2243(.VSS(VSS),.VDD(VDD),.Y(g4256),.A(g3664));
  NOT NOT1_2244(.VSS(VSS),.VDD(VDD),.Y(g6648),.A(I10607));
  NOT NOT1_2245(.VSS(VSS),.VDD(VDD),.Y(g9777),.A(g9474));
  NOT NOT1_2246(.VSS(VSS),.VDD(VDD),.Y(g7546),.A(I11970));
  NOT NOT1_2247(.VSS(VSS),.VDD(VDD),.Y(I5080),.A(g36));
  NOT NOT1_2248(.VSS(VSS),.VDD(VDD),.Y(I15350),.A(g10001));
  NOT NOT1_2249(.VSS(VSS),.VDD(VDD),.Y(I10384),.A(g5842));
  NOT NOT1_2250(.VSS(VSS),.VDD(VDD),.Y(g10162),.A(I15482));
  NOT NOT1_2251(.VSS(VSS),.VDD(VDD),.Y(g3715),.A(g2920));
  NOT NOT1_2252(.VSS(VSS),.VDD(VDD),.Y(I9265),.A(g5085));
  NOT NOT1_2253(.VSS(VSS),.VDD(VDD),.Y(I16787),.A(g10896));
  NOT NOT1_2254(.VSS(VSS),.VDD(VDD),.Y(g11350),.A(g11287));
  NOT NOT1_2255(.VSS(VSS),.VDD(VDD),.Y(I5713),.A(g2436));
  NOT NOT1_2256(.VSS(VSS),.VDD(VDD),.Y(I15820),.A(g10204));
  NOT NOT1_2257(.VSS(VSS),.VDD(VDD),.Y(g5091),.A(g4385));
  NOT NOT1_2258(.VSS(VSS),.VDD(VDD),.Y(g8056),.A(g7671));
  NOT NOT1_2259(.VSS(VSS),.VDD(VDD),.Y(I13317),.A(g8093));
  NOT NOT1_2260(.VSS(VSS),.VDD(VDD),.Y(I12610),.A(g7627));
  NOT NOT1_2261(.VSS(VSS),.VDD(VDD),.Y(g4181),.A(I7360));
  NOT NOT1_2262(.VSS(VSS),.VDD(VDD),.Y(I6754),.A(g2906));
  NOT NOT1_2263(.VSS(VSS),.VDD(VDD),.Y(g8529),.A(I13738));
  NOT NOT1_2264(.VSS(VSS),.VDD(VDD),.Y(I14094),.A(g8700));
  NOT NOT1_2265(.VSS(VSS),.VDD(VDD),.Y(g4381),.A(g3914));
  NOT NOT1_2266(.VSS(VSS),.VDD(VDD),.Y(g7925),.A(g7476));
  NOT NOT1_2267(.VSS(VSS),.VDD(VDD),.Y(I9786),.A(g5396));
  NOT NOT1_2268(.VSS(VSS),.VDD(VDD),.Y(g2118),.A(g1854));
  NOT NOT1_2269(.VSS(VSS),.VDD(VDD),.Y(g8348),.A(I13424));
  NOT NOT1_2270(.VSS(VSS),.VDD(VDD),.Y(I12255),.A(g7203));
  NOT NOT1_2271(.VSS(VSS),.VDD(VDD),.Y(I6273),.A(g2482));
  NOT NOT1_2272(.VSS(VSS),.VDD(VDD),.Y(g2872),.A(I6016));
  NOT NOT1_2273(.VSS(VSS),.VDD(VDD),.Y(I16105),.A(g10382));
  NOT NOT1_2274(.VSS(VSS),.VDD(VDD),.Y(g10629),.A(g10583));
  NOT NOT1_2275(.VSS(VSS),.VDD(VDD),.Y(I10150),.A(g5705));
  NOT NOT1_2276(.VSS(VSS),.VDD(VDD),.Y(g5169),.A(g4596));
  NOT NOT1_2277(.VSS(VSS),.VDD(VDD),.Y(g4197),.A(I7408));
  NOT NOT1_2278(.VSS(VSS),.VDD(VDD),.Y(I10801),.A(g6536));
  NOT NOT1_2279(.VSS(VSS),.VDD(VDD),.Y(g8155),.A(I13048));
  NOT NOT1_2280(.VSS(VSS),.VDD(VDD),.Y(g11396),.A(I17231));
  NOT NOT1_2281(.VSS(VSS),.VDD(VDD),.Y(I13002),.A(g8045));
  NOT NOT1_2282(.VSS(VSS),.VDD(VDD),.Y(g8355),.A(I13445));
  NOT NOT1_2283(.VSS(VSS),.VDD(VDD),.Y(g10220),.A(I15592));
  NOT NOT1_2284(.VSS(VSS),.VDD(VDD),.Y(g5007),.A(I8379));
  NOT NOT1_2285(.VSS(VSS),.VDD(VDD),.Y(I13057),.A(g7843));
  NOT NOT1_2286(.VSS(VSS),.VDD(VDD),.Y(g2652),.A(g2008));
  NOT NOT1_2287(.VSS(VSS),.VDD(VDD),.Y(g2057),.A(g754));
  NOT NOT1_2288(.VSS(VSS),.VDD(VDD),.Y(g10628),.A(I16307));
  NOT NOT1_2289(.VSS(VSS),.VDD(VDD),.Y(I12678),.A(g7376));
  NOT NOT1_2290(.VSS(VSS),.VDD(VDD),.Y(I13128),.A(g7976));
  NOT NOT1_2291(.VSS(VSS),.VDD(VDD),.Y(g2843),.A(I5963));
  NOT NOT1_2292(.VSS(VSS),.VDD(VDD),.Y(g10911),.A(I16685));
  NOT NOT1_2293(.VSS(VSS),.VDD(VDD),.Y(g7320),.A(I11608));
  NOT NOT1_2294(.VSS(VSS),.VDD(VDD),.Y(g2989),.A(g2135));
  NOT NOT1_2295(.VSS(VSS),.VDD(VDD),.Y(g3539),.A(g3015));
  NOT NOT1_2296(.VSS(VSS),.VDD(VDD),.Y(g4263),.A(g3586));
  NOT NOT1_2297(.VSS(VSS),.VDD(VDD),.Y(I13245),.A(g8269));
  NOT NOT1_2298(.VSS(VSS),.VDD(VDD),.Y(I11626),.A(g7042));
  NOT NOT1_2299(.VSS(VSS),.VDD(VDD),.Y(I16769),.A(g10894));
  NOT NOT1_2300(.VSS(VSS),.VDD(VDD),.Y(g5718),.A(I9256));
  NOT NOT1_2301(.VSS(VSS),.VDD(VDD),.Y(I12460),.A(g7569));
  NOT NOT1_2302(.VSS(VSS),.VDD(VDD),.Y(I12939),.A(g7977));
  NOT NOT1_2303(.VSS(VSS),.VDD(VDD),.Y(g5767),.A(I9349));
  NOT NOT1_2304(.VSS(VSS),.VDD(VDD),.Y(I15691),.A(g10233));
  NOT NOT1_2305(.VSS(VSS),.VDD(VDD),.Y(I9296),.A(g4908));
  NOT NOT1_2306(.VSS(VSS),.VDD(VDD),.Y(I10018),.A(g5862));
  NOT NOT1_2307(.VSS(VSS),.VDD(VDD),.Y(I11299),.A(g6727));
  NOT NOT1_2308(.VSS(VSS),.VDD(VDD),.Y(I13323),.A(g8203));
  NOT NOT1_2309(.VSS(VSS),.VDD(VDD),.Y(I7176),.A(g2623));
  NOT NOT1_2310(.VSS(VSS),.VDD(VDD),.Y(I5976),.A(g2186));
  NOT NOT1_2311(.VSS(VSS),.VDD(VDD),.Y(g2549),.A(g1386));
  NOT NOT1_2312(.VSS(VSS),.VDD(VDD),.Y(I6572),.A(g2853));
  NOT NOT1_2313(.VSS(VSS),.VDD(VDD),.Y(I10526),.A(g6161));
  NOT NOT1_2314(.VSS(VSS),.VDD(VDD),.Y(g8063),.A(I12907));
  NOT NOT1_2315(.VSS(VSS),.VDD(VDD),.Y(g2834),.A(I5952));
  NOT NOT1_2316(.VSS(VSS),.VDD(VDD),.Y(g2971),.A(g2046));
  NOT NOT1_2317(.VSS(VSS),.VDD(VDD),.Y(g6172),.A(I9901));
  NOT NOT1_2318(.VSS(VSS),.VDD(VDD),.Y(g6278),.A(I10093));
  NOT NOT1_2319(.VSS(VSS),.VDD(VDD),.Y(g7617),.A(I12199));
  NOT NOT1_2320(.VSS(VSS),.VDD(VDD),.Y(I7405),.A(g3861));
  NOT NOT1_2321(.VSS(VSS),.VDD(VDD),.Y(g7906),.A(I12694));
  NOT NOT1_2322(.VSS(VSS),.VDD(VDD),.Y(g7789),.A(I12532));
  NOT NOT1_2323(.VSS(VSS),.VDD(VDD),.Y(g11405),.A(I17258));
  NOT NOT1_2324(.VSS(VSS),.VDD(VDD),.Y(g5261),.A(g4640));
  NOT NOT1_2325(.VSS(VSS),.VDD(VDD),.Y(g10591),.A(I16258));
  NOT NOT1_2326(.VSS(VSS),.VDD(VDD),.Y(I6543),.A(g3186));
  NOT NOT1_2327(.VSS(VSS),.VDD(VDD),.Y(g3362),.A(I6546));
  NOT NOT1_2328(.VSS(VSS),.VDD(VDD),.Y(g3419),.A(g3104));
  NOT NOT1_2329(.VSS(VSS),.VDD(VDD),.Y(I7829),.A(g3425));
  NOT NOT1_2330(.VSS(VSS),.VDD(VDD),.Y(g6667),.A(I10630));
  NOT NOT1_2331(.VSS(VSS),.VDD(VDD),.Y(g7516),.A(g7148));
  NOT NOT1_2332(.VSS(VSS),.VDD(VDD),.Y(g4562),.A(I7973));
  NOT NOT1_2333(.VSS(VSS),.VDD(VDD),.Y(g6343),.A(I10248));
  NOT NOT1_2334(.VSS(VSS),.VDD(VDD),.Y(g10754),.A(I16439));
  NOT NOT1_2335(.VSS(VSS),.VDD(VDD),.Y(g9353),.A(I14564));
  NOT NOT1_2336(.VSS(VSS),.VDD(VDD),.Y(g3052),.A(I6264));
  NOT NOT1_2337(.VSS(VSS),.VDD(VDD),.Y(g10355),.A(I15829));
  NOT NOT1_2338(.VSS(VSS),.VDD(VDD),.Y(g5415),.A(I8848));
  NOT NOT1_2339(.VSS(VSS),.VDD(VDD),.Y(g6282),.A(I10105));
  NOT NOT1_2340(.VSS(VSS),.VDD(VDD),.Y(g7771),.A(I12478));
  NOT NOT1_2341(.VSS(VSS),.VDD(VDD),.Y(g6566),.A(g5791));
  NOT NOT1_2342(.VSS(VSS),.VDD(VDD),.Y(I11737),.A(g7027));
  NOT NOT1_2343(.VSS(VSS),.VDD(VDD),.Y(g8279),.A(I13209));
  NOT NOT1_2344(.VSS(VSS),.VDD(VDD),.Y(g2121),.A(I5041));
  NOT NOT1_2345(.VSS(VSS),.VDD(VDD),.Y(g4631),.A(g3820));
  NOT NOT1_2346(.VSS(VSS),.VDD(VDD),.Y(I12875),.A(g7638));
  NOT NOT1_2347(.VSS(VSS),.VDD(VDD),.Y(g10825),.A(I16537));
  NOT NOT1_2348(.VSS(VSS),.VDD(VDD),.Y(I10917),.A(g6732));
  NOT NOT1_2349(.VSS(VSS),.VDD(VDD),.Y(I15583),.A(g10157));
  NOT NOT1_2350(.VSS(VSS),.VDD(VDD),.Y(g9802),.A(g9490));
  NOT NOT1_2351(.VSS(VSS),.VDD(VDD),.Y(g1999),.A(g806));
  NOT NOT1_2352(.VSS(VSS),.VDD(VDD),.Y(I11232),.A(g6537));
  NOT NOT1_2353(.VSS(VSS),.VDD(VDD),.Y(g4257),.A(g3664));
  NOT NOT1_2354(.VSS(VSS),.VDD(VDD),.Y(g6134),.A(I9839));
  NOT NOT1_2355(.VSS(VSS),.VDD(VDD),.Y(g5664),.A(I9153));
  NOT NOT1_2356(.VSS(VSS),.VDD(VDD),.Y(g8318),.A(I13338));
  NOT NOT1_2357(.VSS(VSS),.VDD(VDD),.Y(g8872),.A(I14188));
  NOT NOT1_2358(.VSS(VSS),.VDD(VDD),.Y(I9706),.A(g5221));
  NOT NOT1_2359(.VSS(VSS),.VDD(VDD),.Y(g2232),.A(I5221));
  NOT NOT1_2360(.VSS(VSS),.VDD(VDD),.Y(g10172),.A(I15510));
  NOT NOT1_2361(.VSS(VSS),.VDD(VDD),.Y(g11046),.A(I16799));
  NOT NOT1_2362(.VSS(VSS),.VDD(VDD),.Y(g3086),.A(g2276));
  NOT NOT1_2363(.VSS(VSS),.VDD(VDD),.Y(g5203),.A(g4640));
  NOT NOT1_2364(.VSS(VSS),.VDD(VDD),.Y(g2253),.A(g100));
  NOT NOT1_2365(.VSS(VSS),.VDD(VDD),.Y(g3728),.A(I6904));
  NOT NOT1_2366(.VSS(VSS),.VDD(VDD),.Y(g2813),.A(I5913));
  NOT NOT1_2367(.VSS(VSS),.VDD(VDD),.Y(I9029),.A(g4781));
  NOT NOT1_2368(.VSS(VSS),.VDD(VDD),.Y(g8989),.A(I14388));
  NOT NOT1_2369(.VSS(VSS),.VDD(VDD),.Y(I14077),.A(g8758));
  NOT NOT1_2370(.VSS(VSS),.VDD(VDD),.Y(I9171),.A(g4902));
  NOT NOT1_2371(.VSS(VSS),.VDD(VDD),.Y(g6555),.A(g5740));
  NOT NOT1_2372(.VSS(VSS),.VDD(VDD),.Y(I10706),.A(g6080));
  NOT NOT1_2373(.VSS(VSS),.VDD(VDD),.Y(I9371),.A(g5075));
  NOT NOT1_2374(.VSS(VSS),.VDD(VDD),.Y(g6804),.A(I10822));
  NOT NOT1_2375(.VSS(VSS),.VDD(VDD),.Y(I15787),.A(g10269));
  NOT NOT1_2376(.VSS(VSS),.VDD(VDD),.Y(I6414),.A(g2342));
  NOT NOT1_2377(.VSS(VSS),.VDD(VDD),.Y(g3730),.A(g3015));
  NOT NOT1_2378(.VSS(VSS),.VDD(VDD),.Y(g2909),.A(I6080));
  NOT NOT1_2379(.VSS(VSS),.VDD(VDD),.Y(I9956),.A(g5485));
  NOT NOT1_2380(.VSS(VSS),.VDD(VDD),.Y(I10689),.A(g6059));
  NOT NOT1_2381(.VSS(VSS),.VDD(VDD),.Y(g3385),.A(g3121));
  NOT NOT1_2382(.VSS(VSS),.VDD(VDD),.Y(I5383),.A(g886));
  NOT NOT1_2383(.VSS(VSS),.VDD(VDD),.Y(I15302),.A(g10007));
  NOT NOT1_2384(.VSS(VSS),.VDD(VDD),.Y(g11357),.A(I17182));
  NOT NOT1_2385(.VSS(VSS),.VDD(VDD),.Y(g7991),.A(I12809));
  NOT NOT1_2386(.VSS(VSS),.VDD(VDD),.Y(I6513),.A(g2812));
  NOT NOT1_2387(.VSS(VSS),.VDD(VDD),.Y(g2606),.A(I5719));
  NOT NOT1_2388(.VSS(VSS),.VDD(VDD),.Y(g10319),.A(g10270));
  NOT NOT1_2389(.VSS(VSS),.VDD(VDD),.Y(g4441),.A(g3914));
  NOT NOT1_2390(.VSS(VSS),.VDD(VDD),.Y(g6113),.A(I9792));
  NOT NOT1_2391(.VSS(VSS),.VDD(VDD),.Y(g6313),.A(I10198));
  NOT NOT1_2392(.VSS(VSS),.VDD(VDD),.Y(g7078),.A(I11309));
  NOT NOT1_2393(.VSS(VSS),.VDD(VDD),.Y(g7340),.A(I11668));
  NOT NOT1_2394(.VSS(VSS),.VDD(VDD),.Y(I10102),.A(g5730));
  NOT NOT1_2395(.VSS(VSS),.VDD(VDD),.Y(I16778),.A(g10891));
  NOT NOT1_2396(.VSS(VSS),.VDD(VDD),.Y(I13831),.A(g8560));
  NOT NOT1_2397(.VSS(VSS),.VDD(VDD),.Y(g10318),.A(I15752));
  NOT NOT1_2398(.VSS(VSS),.VDD(VDD),.Y(I8050),.A(g4089));
  NOT NOT1_2399(.VSS(VSS),.VDD(VDD),.Y(I13445),.A(g8149));
  NOT NOT1_2400(.VSS(VSS),.VDD(VDD),.Y(I5588),.A(g1203));
  NOT NOT1_2401(.VSS(VSS),.VDD(VDD),.Y(g8121),.A(I12978));
  NOT NOT1_2402(.VSS(VSS),.VDD(VDD),.Y(g10227),.A(I15601));
  NOT NOT1_2403(.VSS(VSS),.VDD(VDD),.Y(g7907),.A(g7664));
  NOT NOT1_2404(.VSS(VSS),.VDD(VDD),.Y(I6436),.A(g2351));
  NOT NOT1_2405(.VSS(VSS),.VDD(VDD),.Y(I6679),.A(g2902));
  NOT NOT1_2406(.VSS(VSS),.VDD(VDD),.Y(g8321),.A(I13347));
  NOT NOT1_2407(.VSS(VSS),.VDD(VDD),.Y(g4673),.A(g4013));
  NOT NOT1_2408(.VSS(VSS),.VDD(VDD),.Y(g6202),.A(g5426));
  NOT NOT1_2409(.VSS(VSS),.VDD(VDD),.Y(g8670),.A(g8551));
  NOT NOT1_2410(.VSS(VSS),.VDD(VDD),.Y(g5689),.A(I9216));
  NOT NOT1_2411(.VSS(VSS),.VDD(VDD),.Y(I8996),.A(g4757));
  NOT NOT1_2412(.VSS(VSS),.VDD(VDD),.Y(I9684),.A(g5426));
  NOT NOT1_2413(.VSS(VSS),.VDD(VDD),.Y(g7035),.A(I11194));
  NOT NOT1_2414(.VSS(VSS),.VDD(VDD),.Y(I15768),.A(g10249));
  NOT NOT1_2415(.VSS(VSS),.VDD(VDD),.Y(I9138),.A(g5210));
  NOT NOT1_2416(.VSS(VSS),.VDD(VDD),.Y(I9639),.A(g5126));
  NOT NOT1_2417(.VSS(VSS),.VDD(VDD),.Y(g7959),.A(I12751));
  NOT NOT1_2418(.VSS(VSS),.VDD(VDD),.Y(I10066),.A(g5778));
  NOT NOT1_2419(.VSS(VSS),.VDD(VDD),.Y(I9338),.A(g5576));
  NOT NOT1_2420(.VSS(VSS),.VDD(VDD),.Y(I10231),.A(g6111));
  NOT NOT1_2421(.VSS(VSS),.VDD(VDD),.Y(g8625),.A(g8487));
  NOT NOT1_2422(.VSS(VSS),.VDD(VDD),.Y(g7082),.A(I11315));
  NOT NOT1_2423(.VSS(VSS),.VDD(VDD),.Y(g2586),.A(g1972));
  NOT NOT1_2424(.VSS(VSS),.VDD(VDD),.Y(g5216),.A(g4445));
  NOT NOT1_2425(.VSS(VSS),.VDD(VDD),.Y(g10540),.A(I16187));
  NOT NOT1_2426(.VSS(VSS),.VDD(VDD),.Y(I17410),.A(g11419));
  NOT NOT1_2427(.VSS(VSS),.VDD(VDD),.Y(g6094),.A(I9749));
  NOT NOT1_2428(.VSS(VSS),.VDD(VDD),.Y(I11498),.A(g6578));
  NOT NOT1_2429(.VSS(VSS),.VDD(VDD),.Y(I12595),.A(g7706));
  NOT NOT1_2430(.VSS(VSS),.VDD(VDD),.Y(I16647),.A(g10866));
  NOT NOT1_2431(.VSS(VSS),.VDD(VDD),.Y(g10058),.A(I15281));
  NOT NOT1_2432(.VSS(VSS),.VDD(VDD),.Y(I16356),.A(g10597));
  NOT NOT1_2433(.VSS(VSS),.VDD(VDD),.Y(g4669),.A(g4013));
  NOT NOT1_2434(.VSS(VSS),.VDD(VDD),.Y(I8724),.A(g4791));
  NOT NOT1_2435(.VSS(VSS),.VDD(VDD),.Y(g6567),.A(I10495));
  NOT NOT1_2436(.VSS(VSS),.VDD(VDD),.Y(g5671),.A(I9174));
  NOT NOT1_2437(.VSS(VSS),.VDD(VDD),.Y(g4368),.A(I7665));
  NOT NOT1_2438(.VSS(VSS),.VDD(VDD),.Y(I11989),.A(g6919));
  NOT NOT1_2439(.VSS(VSS),.VDD(VDD),.Y(I17666),.A(g11603));
  NOT NOT1_2440(.VSS(VSS),.VDD(VDD),.Y(I10885),.A(g6332));
  NOT NOT1_2441(.VSS(VSS),.VDD(VDD),.Y(I8379),.A(g4231));
  NOT NOT1_2442(.VSS(VSS),.VDD(VDD),.Y(g3331),.A(I6510));
  NOT NOT1_2443(.VSS(VSS),.VDD(VDD),.Y(g10203),.A(g10177));
  NOT NOT1_2444(.VSS(VSS),.VDD(VDD),.Y(I14876),.A(g9526));
  NOT NOT1_2445(.VSS(VSS),.VDD(VDD),.Y(I11611),.A(g6913));
  NOT NOT1_2446(.VSS(VSS),.VDD(VDD),.Y(g7656),.A(I12265));
  NOT NOT1_2447(.VSS(VSS),.VDD(VDD),.Y(g4772),.A(g3440));
  NOT NOT1_2448(.VSS(VSS),.VDD(VDD),.Y(g3406),.A(I6611));
  NOT NOT1_2449(.VSS(VSS),.VDD(VDD),.Y(I11722),.A(g7034));
  NOT NOT1_2450(.VSS(VSS),.VDD(VDD),.Y(I7399),.A(g4113));
  NOT NOT1_2451(.VSS(VSS),.VDD(VDD),.Y(g10044),.A(I15263));
  NOT NOT1_2452(.VSS(VSS),.VDD(VDD),.Y(g3635),.A(I6812));
  NOT NOT1_2453(.VSS(VSS),.VDD(VDD),.Y(I6022),.A(g2258));
  NOT NOT1_2454(.VSS(VSS),.VDD(VDD),.Y(g4458),.A(I7817));
  NOT NOT1_2455(.VSS(VSS),.VDD(VDD),.Y(g2570),.A(g207));
  NOT NOT1_2456(.VSS(VSS),.VDD(VDD),.Y(g2860),.A(I5998));
  NOT NOT1_2457(.VSS(VSS),.VDD(VDD),.Y(g2341),.A(I5403));
  NOT NOT1_2458(.VSS(VSS),.VDD(VDD),.Y(g9262),.A(I14473));
  NOT NOT1_2459(.VSS(VSS),.VDD(VDD),.Y(g3682),.A(g2920));
  NOT NOT1_2460(.VSS(VSS),.VDD(VDD),.Y(g6593),.A(I10557));
  NOT NOT1_2461(.VSS(VSS),.VDD(VDD),.Y(I9759),.A(g5344));
  NOT NOT1_2462(.VSS(VSS),.VDD(VDD),.Y(g8519),.A(I13726));
  NOT NOT1_2463(.VSS(VSS),.VDD(VDD),.Y(g3105),.A(g2482));
  NOT NOT1_2464(.VSS(VSS),.VDD(VDD),.Y(g7915),.A(g7473));
  NOT NOT1_2465(.VSS(VSS),.VDD(VDD),.Y(g3305),.A(I6474));
  NOT NOT1_2466(.VSS(VSS),.VDD(VDD),.Y(g10281),.A(g10162));
  NOT NOT1_2467(.VSS(VSS),.VDD(VDD),.Y(g98),.A(I4783));
  NOT NOT1_2468(.VSS(VSS),.VDD(VDD),.Y(g2645),.A(g1991));
  NOT NOT1_2469(.VSS(VSS),.VDD(VDD),.Y(I8835),.A(g4791));
  NOT NOT1_2470(.VSS(VSS),.VDD(VDD),.Y(g5826),.A(I9440));
  NOT NOT1_2471(.VSS(VSS),.VDD(VDD),.Y(I12418),.A(g7568));
  NOT NOT1_2472(.VSS(VSS),.VDD(VDD),.Y(I12822),.A(g7677));
  NOT NOT1_2473(.VSS(VSS),.VDD(VDD),.Y(g10902),.A(I16660));
  NOT NOT1_2474(.VSS(VSS),.VDD(VDD),.Y(g10377),.A(I15855));
  NOT NOT1_2475(.VSS(VSS),.VDD(VDD),.Y(g8606),.A(g8481));
  NOT NOT1_2476(.VSS(VSS),.VDD(VDD),.Y(g7214),.A(I11450));
  NOT NOT1_2477(.VSS(VSS),.VDD(VDD),.Y(I6947),.A(g2860));
  NOT NOT1_2478(.VSS(VSS),.VDD(VDD),.Y(g10120),.A(I15368));
  NOT NOT1_2479(.VSS(VSS),.VDD(VDD),.Y(g4011),.A(I7151));
  NOT NOT1_2480(.VSS(VSS),.VDD(VDD),.Y(g9076),.A(g8892));
  NOT NOT1_2481(.VSS(VSS),.VDD(VDD),.Y(g5741),.A(I9305));
  NOT NOT1_2482(.VSS(VSS),.VDD(VDD),.Y(g3748),.A(g2971));
  NOT NOT1_2483(.VSS(VSS),.VDD(VDD),.Y(g4411),.A(I7743));
  NOT NOT1_2484(.VSS(VSS),.VDD(VDD),.Y(g4734),.A(g3586));
  NOT NOT1_2485(.VSS(VSS),.VDD(VDD),.Y(I11342),.A(g6686));
  NOT NOT1_2486(.VSS(VSS),.VDD(VDD),.Y(g9889),.A(I15072));
  NOT NOT1_2487(.VSS(VSS),.VDD(VDD),.Y(g7110),.A(I11345));
  NOT NOT1_2488(.VSS(VSS),.VDD(VDD),.Y(g6264),.A(I10051));
  NOT NOT1_2489(.VSS(VSS),.VDD(VDD),.Y(g7310),.A(I11578));
  NOT NOT1_2490(.VSS(VSS),.VDD(VDD),.Y(I6560),.A(g2845));
  NOT NOT1_2491(.VSS(VSS),.VDD(VDD),.Y(I7291),.A(g3212));
  NOT NOT1_2492(.VSS(VSS),.VDD(VDD),.Y(I8611),.A(g4562));
  NOT NOT1_2493(.VSS(VSS),.VDD(VDD),.Y(I10456),.A(g5844));
  NOT NOT1_2494(.VSS(VSS),.VDD(VDD),.Y(I15482),.A(g10115));
  NOT NOT1_2495(.VSS(VSS),.VDD(VDD),.Y(g5638),.A(I9077));
  NOT NOT1_2496(.VSS(VSS),.VDD(VDD),.Y(g3226),.A(I6403));
  NOT NOT1_2497(.VSS(VSS),.VDD(VDD),.Y(g6933),.A(I11061));
  NOT NOT1_2498(.VSS(VSS),.VDD(VDD),.Y(g7663),.A(I12282));
  NOT NOT1_2499(.VSS(VSS),.VDD(VDD),.Y(I11650),.A(g6938));
  NOT NOT1_2500(.VSS(VSS),.VDD(VDD),.Y(g10699),.A(I16376));
  NOT NOT1_2501(.VSS(VSS),.VDD(VDD),.Y(g2607),.A(I5722));
  NOT NOT1_2502(.VSS(VSS),.VDD(VDD),.Y(I12853),.A(g7638));
  NOT NOT1_2503(.VSS(VSS),.VDD(VDD),.Y(I16897),.A(g10947));
  NOT NOT1_2504(.VSS(VSS),.VDD(VDD),.Y(I5240),.A(g64));
  NOT NOT1_2505(.VSS(VSS),.VDD(VDD),.Y(g2962),.A(I6183));
  NOT NOT1_2506(.VSS(VSS),.VDD(VDD),.Y(g6521),.A(I10437));
  NOT NOT1_2507(.VSS(VSS),.VDD(VDD),.Y(I17084),.A(g11249));
  NOT NOT1_2508(.VSS(VSS),.VDD(VDD),.Y(g4474),.A(g3820));
  NOT NOT1_2509(.VSS(VSS),.VDD(VDD),.Y(g10290),.A(I15694));
  NOT NOT1_2510(.VSS(VSS),.VDD(VDD),.Y(g2158),.A(I5077));
  NOT NOT1_2511(.VSS(VSS),.VDD(VDD),.Y(g6050),.A(I9677));
  NOT NOT1_2512(.VSS(VSS),.VDD(VDD),.Y(g6641),.A(I10598));
  NOT NOT1_2513(.VSS(VSS),.VDD(VDD),.Y(I11198),.A(g6521));
  NOT NOT1_2514(.VSS(VSS),.VDD(VDD),.Y(I9498),.A(g5081));
  NOT NOT1_2515(.VSS(VSS),.VDD(VDD),.Y(I12589),.A(g7571));
  NOT NOT1_2516(.VSS(VSS),.VDD(VDD),.Y(g10698),.A(I16373));
  NOT NOT1_2517(.VSS(VSS),.VDD(VDD),.Y(g2506),.A(g636));
  NOT NOT1_2518(.VSS(VSS),.VDD(VDD),.Y(g6450),.A(I10378));
  NOT NOT1_2519(.VSS(VSS),.VDD(VDD),.Y(I6037),.A(g2560));
  NOT NOT1_2520(.VSS(VSS),.VDD(VDD),.Y(I17321),.A(g11348));
  NOT NOT1_2521(.VSS(VSS),.VDD(VDD),.Y(g5883),.A(g5309));
  NOT NOT1_2522(.VSS(VSS),.VDD(VDD),.Y(I10314),.A(g6251));
  NOT NOT1_2523(.VSS(VSS),.VDD(VDD),.Y(g7402),.A(g6860));
  NOT NOT1_2524(.VSS(VSS),.VDD(VDD),.Y(I6495),.A(g2076));
  NOT NOT1_2525(.VSS(VSS),.VDD(VDD),.Y(I9833),.A(g5197));
  NOT NOT1_2526(.VSS(VSS),.VDD(VDD),.Y(I17179),.A(g11307));
  NOT NOT1_2527(.VSS(VSS),.VDD(VDD),.Y(I11528),.A(g6796));
  NOT NOT1_2528(.VSS(VSS),.VDD(VDD),.Y(I6102),.A(g2240));
  NOT NOT1_2529(.VSS(VSS),.VDD(VDD),.Y(I16717),.A(g10779));
  NOT NOT1_2530(.VSS(VSS),.VDD(VDD),.Y(I17531),.A(g11488));
  NOT NOT1_2531(.VSS(VSS),.VDD(VDD),.Y(I7694),.A(g3742));
  NOT NOT1_2532(.VSS(VSS),.VDD(VDD),.Y(I11330),.A(g6571));
  NOT NOT1_2533(.VSS(VSS),.VDD(VDD),.Y(I6302),.A(g2243));
  NOT NOT1_2534(.VSS(VSS),.VDD(VDD),.Y(g3373),.A(I6565));
  NOT NOT1_2535(.VSS(VSS),.VDD(VDD),.Y(I15778),.A(g10255));
  NOT NOT1_2536(.VSS(VSS),.VDD(VDD),.Y(g7762),.A(I12451));
  NOT NOT1_2537(.VSS(VSS),.VDD(VDD),.Y(g3491),.A(g2669));
  NOT NOT1_2538(.VSS(VSS),.VDD(VDD),.Y(g4080),.A(g2903));
  NOT NOT1_2539(.VSS(VSS),.VDD(VDD),.Y(I5116),.A(g40));
  NOT NOT1_2540(.VSS(VSS),.VDD(VDD),.Y(g11081),.A(I16856));
  NOT NOT1_2541(.VSS(VSS),.VDD(VDD),.Y(I7852),.A(g3438));
  NOT NOT1_2542(.VSS(VSS),.VDD(VDD),.Y(I7923),.A(g3394));
  NOT NOT1_2543(.VSS(VSS),.VDD(VDD),.Y(g5758),.A(I9338));
  NOT NOT1_2544(.VSS(VSS),.VDD(VDD),.Y(g8141),.A(I13020));
  NOT NOT1_2545(.VSS(VSS),.VDD(VDD),.Y(g8570),.A(I13803));
  NOT NOT1_2546(.VSS(VSS),.VDD(VDD),.Y(g5066),.A(I8436));
  NOT NOT1_2547(.VSS(VSS),.VDD(VDD),.Y(g5589),.A(I9001));
  NOT NOT1_2548(.VSS(VSS),.VDD(VDD),.Y(g6724),.A(I10719));
  NOT NOT1_2549(.VSS(VSS),.VDD(VDD),.Y(g8341),.A(I13403));
  NOT NOT1_2550(.VSS(VSS),.VDD(VDD),.Y(I10054),.A(g5728));
  NOT NOT1_2551(.VSS(VSS),.VDD(VDD),.Y(g2275),.A(g757));
  NOT NOT1_2552(.VSS(VSS),.VDD(VDD),.Y(I9539),.A(g5354));
  NOT NOT1_2553(.VSS(VSS),.VDD(VDD),.Y(I9896),.A(g5295));
  NOT NOT1_2554(.VSS(VSS),.VDD(VDD),.Y(g4713),.A(g3546));
  NOT NOT1_2555(.VSS(VSS),.VDD(VDD),.Y(I10243),.A(g5918));
  NOT NOT1_2556(.VSS(VSS),.VDD(VDD),.Y(I11132),.A(g6451));
  NOT NOT1_2557(.VSS(VSS),.VDD(VDD),.Y(I11869),.A(g6894));
  NOT NOT1_2558(.VSS(VSS),.VDD(VDD),.Y(g7877),.A(g7479));
  NOT NOT1_2559(.VSS(VSS),.VDD(VDD),.Y(I7701),.A(g3513));
  NOT NOT1_2560(.VSS(VSS),.VDD(VDD),.Y(g3369),.A(I6557));
  NOT NOT1_2561(.VSS(VSS),.VDD(VDD),.Y(I5565),.A(g1713));
  NOT NOT1_2562(.VSS(VSS),.VDD(VDD),.Y(g3007),.A(I6240));
  NOT NOT1_2563(.VSS(VSS),.VDD(VDD),.Y(g9339),.A(I14522));
  NOT NOT1_2564(.VSS(VSS),.VDD(VDD),.Y(I15356),.A(g10013));
  NOT NOT1_2565(.VSS(VSS),.VDD(VDD),.Y(g7657),.A(I12268));
  NOT NOT1_2566(.VSS(VSS),.VDD(VDD),.Y(g6878),.A(I10966));
  NOT NOT1_2567(.VSS(VSS),.VDD(VDD),.Y(I15826),.A(g10205));
  NOT NOT1_2568(.VSS(VSS),.VDD(VDD),.Y(I6917),.A(g2832));
  NOT NOT1_2569(.VSS(VSS),.VDD(VDD),.Y(I15380),.A(g10098));
  NOT NOT1_2570(.VSS(VSS),.VDD(VDD),.Y(I4894),.A(g258));
  NOT NOT1_2571(.VSS(VSS),.VDD(VDD),.Y(g2174),.A(g31));
  NOT NOT1_2572(.VSS(VSS),.VDD(VDD),.Y(g3459),.A(I6661));
  NOT NOT1_2573(.VSS(VSS),.VDD(VDD),.Y(g6289),.A(I10126));
  NOT NOT1_2574(.VSS(VSS),.VDD(VDD),.Y(g9024),.A(I14409));
  NOT NOT1_2575(.VSS(VSS),.VDD(VDD),.Y(g2374),.A(g591));
  NOT NOT1_2576(.VSS(VSS),.VDD(VDD),.Y(I12616),.A(g7534));
  NOT NOT1_2577(.VSS(VSS),.VDD(VDD),.Y(I9162),.A(g5035));
  NOT NOT1_2578(.VSS(VSS),.VDD(VDD),.Y(g7556),.A(I11992));
  NOT NOT1_2579(.VSS(VSS),.VDD(VDD),.Y(I9268),.A(g5305));
  NOT NOT1_2580(.VSS(VSS),.VDD(VDD),.Y(I16723),.A(g10851));
  NOT NOT1_2581(.VSS(VSS),.VDD(VDD),.Y(g3767),.A(I6976));
  NOT NOT1_2582(.VSS(VSS),.VDD(VDD),.Y(g10547),.A(I16206));
  NOT NOT1_2583(.VSS(VSS),.VDD(VDD),.Y(g9424),.A(g9076));
  NOT NOT1_2584(.VSS(VSS),.VDD(VDD),.Y(g10895),.A(I16647));
  NOT NOT1_2585(.VSS(VSS),.VDD(VDD),.Y(I7886),.A(g4076));
  NOT NOT1_2586(.VSS(VSS),.VDD(VDD),.Y(I9362),.A(g5013));
  NOT NOT1_2587(.VSS(VSS),.VDD(VDD),.Y(g6835),.A(I10885));
  NOT NOT1_2588(.VSS(VSS),.VDD(VDD),.Y(g2985),.A(I6217));
  NOT NOT1_2589(.VSS(VSS),.VDD(VDD),.Y(g9809),.A(I14944));
  NOT NOT1_2590(.VSS(VSS),.VDD(VDD),.Y(g5827),.A(I9443));
  NOT NOT1_2591(.VSS(VSS),.VDD(VDD),.Y(g6882),.A(I10974));
  NOT NOT1_2592(.VSS(VSS),.VDD(VDD),.Y(g7928),.A(g7508));
  NOT NOT1_2593(.VSS(VSS),.VDD(VDD),.Y(I10156),.A(g6100));
  NOT NOT1_2594(.VSS(VSS),.VDD(VDD),.Y(I10655),.A(g6036));
  NOT NOT1_2595(.VSS(VSS),.VDD(VDD),.Y(I15672),.A(g10132));
  NOT NOT1_2596(.VSS(VSS),.VDD(VDD),.Y(g3582),.A(g3164));
  NOT NOT1_2597(.VSS(VSS),.VDD(VDD),.Y(I16387),.A(g10629));
  NOT NOT1_2598(.VSS(VSS),.VDD(VDD),.Y(I17334),.A(g11360));
  NOT NOT1_2599(.VSS(VSS),.VDD(VDD),.Y(g6271),.A(I10072));
  NOT NOT1_2600(.VSS(VSS),.VDD(VDD),.Y(I11225),.A(g6534));
  NOT NOT1_2601(.VSS(VSS),.VDD(VDD),.Y(g10226),.A(I15598));
  NOT NOT1_2602(.VSS(VSS),.VDD(VDD),.Y(I9452),.A(g5085));
  NOT NOT1_2603(.VSS(VSS),.VDD(VDD),.Y(g11182),.A(I16947));
  NOT NOT1_2604(.VSS(VSS),.VDD(VDD),.Y(g11651),.A(I17755));
  NOT NOT1_2605(.VSS(VSS),.VDD(VDD),.Y(g7064),.A(I11269));
  NOT NOT1_2606(.VSS(VSS),.VDD(VDD),.Y(I5210),.A(g58));
  NOT NOT1_2607(.VSS(VSS),.VDD(VDD),.Y(g2239),.A(I5240));
  NOT NOT1_2608(.VSS(VSS),.VDD(VDD),.Y(I10180),.A(g6107));
  NOT NOT1_2609(.VSS(VSS),.VDD(VDD),.Y(g9672),.A(I14805));
  NOT NOT1_2610(.VSS(VSS),.VDD(VDD),.Y(I13708),.A(g8337));
  NOT NOT1_2611(.VSS(VSS),.VDD(VDD),.Y(g5774),.A(I9362));
  NOT NOT1_2612(.VSS(VSS),.VDD(VDD),.Y(g7899),.A(I12683));
  NOT NOT1_2613(.VSS(VSS),.VDD(VDD),.Y(g3793),.A(g2593));
  NOT NOT1_2614(.VSS(VSS),.VDD(VDD),.Y(g7464),.A(I11858));
  NOT NOT1_2615(.VSS(VSS),.VDD(VDD),.Y(I12053),.A(g6928));
  NOT NOT1_2616(.VSS(VSS),.VDD(VDD),.Y(g8358),.A(I13454));
  NOT NOT1_2617(.VSS(VSS),.VDD(VDD),.Y(I12809),.A(g7686));
  NOT NOT1_2618(.VSS(VSS),.VDD(VDD),.Y(g7785),.A(I12520));
  NOT NOT1_2619(.VSS(VSS),.VDD(VDD),.Y(I16811),.A(g10908));
  NOT NOT1_2620(.VSS(VSS),.VDD(VDD),.Y(g10551),.A(I16214));
  NOT NOT1_2621(.VSS(VSS),.VDD(VDD),.Y(I6233),.A(g2299));
  NOT NOT1_2622(.VSS(VSS),.VDD(VDD),.Y(g2832),.A(I5946));
  NOT NOT1_2623(.VSS(VSS),.VDD(VDD),.Y(I12466),.A(g7585));
  NOT NOT1_2624(.VSS(VSS),.VDD(VDD),.Y(g3415),.A(g3121));
  NOT NOT1_2625(.VSS(VSS),.VDD(VDD),.Y(g3227),.A(I6406));
  NOT NOT1_2626(.VSS(VSS),.VDD(VDD),.Y(I7825),.A(g3414));
  NOT NOT1_2627(.VSS(VSS),.VDD(VDD),.Y(g6799),.A(I10807));
  NOT NOT1_2628(.VSS(VSS),.VDD(VDD),.Y(g2853),.A(g2171));
  NOT NOT1_2629(.VSS(VSS),.VDD(VDD),.Y(I11043),.A(g6412));
  NOT NOT1_2630(.VSS(VSS),.VDD(VDD),.Y(I6454),.A(g2368));
  NOT NOT1_2631(.VSS(VSS),.VDD(VDD),.Y(I13043),.A(g8055));
  NOT NOT1_2632(.VSS(VSS),.VDD(VDD),.Y(I17216),.A(g11291));
  NOT NOT1_2633(.VSS(VSS),.VDD(VDD),.Y(g2420),.A(g237));
  NOT NOT1_2634(.VSS(VSS),.VDD(VDD),.Y(g6674),.A(I10639));
  NOT NOT1_2635(.VSS(VSS),.VDD(VDD),.Y(I9486),.A(g5066));
  NOT NOT1_2636(.VSS(VSS),.VDD(VDD),.Y(g11513),.A(I17558));
  NOT NOT1_2637(.VSS(VSS),.VDD(VDD),.Y(I12177),.A(g7259));
  NOT NOT1_2638(.VSS(VSS),.VDD(VDD),.Y(g10127),.A(I15383));
  NOT NOT1_2639(.VSS(VSS),.VDD(VDD),.Y(g3664),.A(g3209));
  NOT NOT1_2640(.VSS(VSS),.VDD(VDD),.Y(g8275),.A(I13197));
  NOT NOT1_2641(.VSS(VSS),.VDD(VDD),.Y(g2507),.A(I5584));
  NOT NOT1_2642(.VSS(VSS),.VDD(VDD),.Y(g8311),.A(I13317));
  NOT NOT1_2643(.VSS(VSS),.VDD(VDD),.Y(g3246),.A(g2482));
  NOT NOT1_2644(.VSS(VSS),.VDD(VDD),.Y(I15448),.A(g10056));
  NOT NOT1_2645(.VSS(VSS),.VDD(VDD),.Y(g5509),.A(g4739));
  NOT NOT1_2646(.VSS(VSS),.VDD(VDD),.Y(g4326),.A(g3863));
  NOT NOT1_2647(.VSS(VSS),.VDD(VDD),.Y(I14694),.A(g9259));
  NOT NOT1_2648(.VSS(VSS),.VDD(VDD),.Y(I7408),.A(g4125));
  NOT NOT1_2649(.VSS(VSS),.VDD(VDD),.Y(g7237),.A(I11477));
  NOT NOT1_2650(.VSS(VSS),.VDD(VDD),.Y(g10490),.A(I16105));
  NOT NOT1_2651(.VSS(VSS),.VDD(VDD),.Y(I9185),.A(g4915));
  NOT NOT1_2652(.VSS(VSS),.VDD(VDD),.Y(I7336),.A(g3997));
  NOT NOT1_2653(.VSS(VSS),.VDD(VDD),.Y(g3721),.A(I6891));
  NOT NOT1_2654(.VSS(VSS),.VDD(VDD),.Y(g11505),.A(I17534));
  NOT NOT1_2655(.VSS(VSS),.VDD(VDD),.Y(I11602),.A(g6833));
  NOT NOT1_2656(.VSS(VSS),.VDD(VDD),.Y(I11810),.A(g7246));
  NOT NOT1_2657(.VSS(VSS),.VDD(VDD),.Y(g11404),.A(I17255));
  NOT NOT1_2658(.VSS(VSS),.VDD(VDD),.Y(g6132),.A(I9833));
  NOT NOT1_2659(.VSS(VSS),.VDD(VDD),.Y(g5662),.A(I9147));
  NOT NOT1_2660(.VSS(VSS),.VDD(VDD),.Y(I6553),.A(g3186));
  NOT NOT1_2661(.VSS(VSS),.VDD(VDD),.Y(I4850),.A(g1958));
  NOT NOT1_2662(.VSS(VSS),.VDD(VDD),.Y(g7844),.A(I12631));
  NOT NOT1_2663(.VSS(VSS),.VDD(VDD),.Y(I17543),.A(g11499));
  NOT NOT1_2664(.VSS(VSS),.VDD(VDD),.Y(I11068),.A(g6426));
  NOT NOT1_2665(.VSS(VSS),.VDD(VDD),.Y(I13068),.A(g7906));
  NOT NOT1_2666(.VSS(VSS),.VDD(VDD),.Y(g6680),.A(I10643));
  NOT NOT1_2667(.VSS(VSS),.VDD(VDD),.Y(g6209),.A(I9956));
  NOT NOT1_2668(.VSS(VSS),.VDD(VDD),.Y(g8985),.A(I14376));
  NOT NOT1_2669(.VSS(VSS),.VDD(VDD),.Y(I11879),.A(g6893));
  NOT NOT1_2670(.VSS(VSS),.VDD(VDD),.Y(g5994),.A(I9612));
  NOT NOT1_2671(.VSS(VSS),.VDD(VDD),.Y(g10889),.A(I16629));
  NOT NOT1_2672(.VSS(VSS),.VDD(VDD),.Y(I16850),.A(g10905));
  NOT NOT1_2673(.VSS(VSS),.VDD(VDD),.Y(I11970),.A(g6918));
  NOT NOT1_2674(.VSS(VSS),.VDD(VDD),.Y(g7394),.A(I11778));
  NOT NOT1_2675(.VSS(VSS),.VDD(VDD),.Y(I10557),.A(g6197));
  NOT NOT1_2676(.VSS(VSS),.VDD(VDD),.Y(g10354),.A(I15826));
  NOT NOT1_2677(.VSS(VSS),.VDD(VDD),.Y(g2905),.A(I6068));
  NOT NOT1_2678(.VSS(VSS),.VDD(VDD),.Y(g7089),.A(I11322));
  NOT NOT1_2679(.VSS(VSS),.VDD(VDD),.Y(g7731),.A(I12376));
  NOT NOT1_2680(.VSS(VSS),.VDD(VDD),.Y(g10888),.A(I16626));
  NOT NOT1_2681(.VSS(VSS),.VDD(VDD),.Y(g6802),.A(I10816));
  NOT NOT1_2682(.VSS(VSS),.VDD(VDD),.Y(g8239),.A(g7826));
  NOT NOT1_2683(.VSS(VSS),.VDD(VDD),.Y(g4183),.A(I7366));
  NOT NOT1_2684(.VSS(VSS),.VDD(VDD),.Y(g9273),.A(I14490));
  NOT NOT1_2685(.VSS(VSS),.VDD(VDD),.Y(g4608),.A(g3829));
  NOT NOT1_2686(.VSS(VSS),.VDD(VDD),.Y(g5816),.A(I9424));
  NOT NOT1_2687(.VSS(VSS),.VDD(VDD),.Y(I5922),.A(g2170));
  NOT NOT1_2688(.VSS(VSS),.VDD(VDD),.Y(I7465),.A(g3726));
  NOT NOT1_2689(.VSS(VSS),.VDD(VDD),.Y(g7966),.A(I12762));
  NOT NOT1_2690(.VSS(VSS),.VDD(VDD),.Y(g2100),.A(I4948));
  NOT NOT1_2691(.VSS(VSS),.VDD(VDD),.Y(I10278),.A(g5815));
  NOT NOT1_2692(.VSS(VSS),.VDD(VDD),.Y(g3940),.A(g2920));
  NOT NOT1_2693(.VSS(VSS),.VDD(VDD),.Y(g6558),.A(I10484));
  NOT NOT1_2694(.VSS(VSS),.VDD(VDD),.Y(I12009),.A(g6915));
  NOT NOT1_2695(.VSS(VSS),.VDD(VDD),.Y(I6888),.A(g2960));
  NOT NOT1_2696(.VSS(VSS),.VDD(VDD),.Y(I8262),.A(g4636));
  NOT NOT1_2697(.VSS(VSS),.VDD(VDD),.Y(I11967),.A(g6911));
  NOT NOT1_2698(.VSS(VSS),.VDD(VDD),.Y(g8020),.A(I12862));
  NOT NOT1_2699(.VSS(VSS),.VDD(VDD),.Y(I10286),.A(g6237));
  NOT NOT1_2700(.VSS(VSS),.VDD(VDD),.Y(g8420),.A(I13574));
  NOT NOT1_2701(.VSS(VSS),.VDD(VDD),.Y(I5060),.A(g1191));
  NOT NOT1_2702(.VSS(VSS),.VDD(VDD),.Y(g10931),.A(g10827));
  NOT NOT1_2703(.VSS(VSS),.VDD(VDD),.Y(g3388),.A(I6590));
  NOT NOT1_2704(.VSS(VSS),.VDD(VDD),.Y(I10039),.A(g5718));
  NOT NOT1_2705(.VSS(VSS),.VDD(VDD),.Y(I14306),.A(g8812));
  NOT NOT1_2706(.VSS(VSS),.VDD(VDD),.Y(I11459),.A(g6488));
  NOT NOT1_2707(.VSS(VSS),.VDD(VDD),.Y(g11433),.A(I17350));
  NOT NOT1_2708(.VSS(VSS),.VDD(VDD),.Y(g9572),.A(I14709));
  NOT NOT1_2709(.VSS(VSS),.VDD(VDD),.Y(g5685),.A(I9208));
  NOT NOT1_2710(.VSS(VSS),.VDD(VDD),.Y(g5197),.A(I8611));
  NOT NOT1_2711(.VSS(VSS),.VDD(VDD),.Y(g5700),.A(I9237));
  NOT NOT1_2712(.VSS(VSS),.VDD(VDD),.Y(g8794),.A(I14109));
  NOT NOT1_2713(.VSS(VSS),.VDD(VDD),.Y(g5397),.A(I8835));
  NOT NOT1_2714(.VSS(VSS),.VDD(VDD),.Y(g2750),.A(I5818));
  NOT NOT1_2715(.VSS(VSS),.VDD(VDD),.Y(I8889),.A(g4553));
  NOT NOT1_2716(.VSS(VSS),.VDD(VDD),.Y(g11620),.A(I17678));
  NOT NOT1_2717(.VSS(VSS),.VDD(VDD),.Y(g10190),.A(I15548));
  NOT NOT1_2718(.VSS(VSS),.VDD(VDD),.Y(I8476),.A(g4577));
  NOT NOT1_2719(.VSS(VSS),.VDD(VDD),.Y(g4361),.A(I7648));
  NOT NOT1_2720(.VSS(VSS),.VDD(VDD),.Y(I9766),.A(g5348));
  NOT NOT1_2721(.VSS(VSS),.VDD(VDD),.Y(I15811),.A(g10200));
  NOT NOT1_2722(.VSS(VSS),.VDD(VDD),.Y(g3428),.A(I6639));
  NOT NOT1_2723(.VSS(VSS),.VDD(VDD),.Y(I7096),.A(g3186));
  NOT NOT1_2724(.VSS(VSS),.VDD(VDD),.Y(I12454),.A(g7544));
  NOT NOT1_2725(.VSS(VSS),.VDD(VDD),.Y(I9087),.A(g5113));
  NOT NOT1_2726(.VSS(VSS),.VDD(VDD),.Y(I9105),.A(g5589));
  NOT NOT1_2727(.VSS(VSS),.VDD(VDD),.Y(I9305),.A(g4970));
  NOT NOT1_2728(.VSS(VSS),.VDD(VDD),.Y(I9801),.A(g5416));
  NOT NOT1_2729(.VSS(VSS),.VDD(VDD),.Y(g3430),.A(I6643));
  NOT NOT1_2730(.VSS(VSS),.VDD(VDD),.Y(g7814),.A(I12607));
  NOT NOT1_2731(.VSS(VSS),.VDD(VDD),.Y(I12712),.A(g7441));
  NOT NOT1_2732(.VSS(VSS),.VDD(VDD),.Y(g11646),.A(I17742));
  NOT NOT1_2733(.VSS(VSS),.VDD(VDD),.Y(g4051),.A(I7166));
  NOT NOT1_2734(.VSS(VSS),.VDD(VDD),.Y(I10601),.A(g5996));
  NOT NOT1_2735(.VSS(VSS),.VDD(VDD),.Y(I13010),.A(g8047));
  NOT NOT1_2736(.VSS(VSS),.VDD(VDD),.Y(g11343),.A(I17152));
  NOT NOT1_2737(.VSS(VSS),.VDD(VDD),.Y(I13918),.A(g8451));
  NOT NOT1_2738(.VSS(VSS),.VDD(VDD),.Y(I16379),.A(g10598));
  NOT NOT1_2739(.VSS(VSS),.VDD(VDD),.Y(g4127),.A(I7276));
  NOT NOT1_2740(.VSS(VSS),.VDD(VDD),.Y(g4451),.A(g3638));
  NOT NOT1_2741(.VSS(VSS),.VDD(VDD),.Y(I15971),.A(g10408));
  NOT NOT1_2742(.VSS(VSS),.VDD(VDD),.Y(g4327),.A(I7600));
  NOT NOT1_2743(.VSS(VSS),.VDD(VDD),.Y(I17265),.A(g11352));
  NOT NOT1_2744(.VSS(VSS),.VDD(VDD),.Y(g7350),.A(I11698));
  NOT NOT1_2745(.VSS(VSS),.VDD(VDD),.Y(g2040),.A(g1786));
  NOT NOT1_2746(.VSS(VSS),.VDD(VDD),.Y(g6574),.A(I10514));
  NOT NOT1_2747(.VSS(VSS),.VDD(VDD),.Y(I12907),.A(g7959));
  NOT NOT1_2748(.VSS(VSS),.VDD(VDD),.Y(I5995),.A(g2196));
  NOT NOT1_2749(.VSS(VSS),.VDD(VDD),.Y(I11079),.A(g6649));
  NOT NOT1_2750(.VSS(VSS),.VDD(VDD),.Y(g10546),.A(I16203));
  NOT NOT1_2751(.VSS(VSS),.VDD(VDD),.Y(g7038),.A(I11201));
  NOT NOT1_2752(.VSS(VSS),.VDD(VDD),.Y(I11444),.A(g6653));
  NOT NOT1_2753(.VSS(VSS),.VDD(VDD),.Y(I17416),.A(g11420));
  NOT NOT1_2754(.VSS(VSS),.VDD(VDD),.Y(g10211),.A(I15583));
  NOT NOT1_2755(.VSS(VSS),.VDD(VDD),.Y(g9534),.A(I14687));
  NOT NOT1_2756(.VSS(VSS),.VDD(VDD),.Y(g9961),.A(I15162));
  NOT NOT1_2757(.VSS(VSS),.VDD(VDD),.Y(g6714),.A(g5867));
  NOT NOT1_2758(.VSS(VSS),.VDD(VDD),.Y(g7438),.A(g7232));
  NOT NOT1_2759(.VSS(VSS),.VDD(VDD),.Y(g7773),.A(I12484));
  NOT NOT1_2760(.VSS(VSS),.VDD(VDD),.Y(I11599),.A(g6832));
  NOT NOT1_2761(.VSS(VSS),.VDD(VDD),.Y(g7009),.A(I11152));
  NOT NOT1_2762(.VSS(VSS),.VDD(VDD),.Y(g11369),.A(I17194));
  NOT NOT1_2763(.VSS(VSS),.VDD(VDD),.Y(g2123),.A(I5047));
  NOT NOT1_2764(.VSS(VSS),.VDD(VDD),.Y(I6639),.A(g2632));
  NOT NOT1_2765(.VSS(VSS),.VDD(VDD),.Y(g4346),.A(I7625));
  NOT NOT1_2766(.VSS(VSS),.VDD(VDD),.Y(g8515),.A(I13714));
  NOT NOT1_2767(.VSS(VSS),.VDD(VDD),.Y(g10088),.A(I15317));
  NOT NOT1_2768(.VSS(VSS),.VDD(VDD),.Y(I8285),.A(g4771));
  NOT NOT1_2769(.VSS(VSS),.VDD(VDD),.Y(I10937),.A(g6552));
  NOT NOT1_2770(.VSS(VSS),.VDD(VDD),.Y(I12239),.A(g7073));
  NOT NOT1_2771(.VSS(VSS),.VDD(VDD),.Y(I5840),.A(g2432));
  NOT NOT1_2772(.VSS(VSS),.VDD(VDD),.Y(I15368),.A(g9990));
  NOT NOT1_2773(.VSS(VSS),.VDD(VDD),.Y(I17510),.A(g11481));
  NOT NOT1_2774(.VSS(VSS),.VDD(VDD),.Y(I16742),.A(g10857));
  NOT NOT1_2775(.VSS(VSS),.VDD(VDD),.Y(g8100),.A(g7947));
  NOT NOT1_2776(.VSS(VSS),.VDD(VDD),.Y(I16944),.A(g11079));
  NOT NOT1_2777(.VSS(VSS),.VDD(VDD),.Y(g3910),.A(g3015));
  NOT NOT1_2778(.VSS(VSS),.VDD(VDD),.Y(I13086),.A(g7924));
  NOT NOT1_2779(.VSS(VSS),.VDD(VDD),.Y(g7769),.A(I12472));
  NOT NOT1_2780(.VSS(VSS),.VDD(VDD),.Y(I15412),.A(g10075));
  NOT NOT1_2781(.VSS(VSS),.VDD(VDD),.Y(g3638),.A(I6821));
  NOT NOT1_2782(.VSS(VSS),.VDD(VDD),.Y(I8139),.A(g3681));
  NOT NOT1_2783(.VSS(VSS),.VDD(VDD),.Y(g7212),.A(I11444));
  NOT NOT1_2784(.VSS(VSS),.VDD(VDD),.Y(g5723),.A(I9265));
  NOT NOT1_2785(.VSS(VSS),.VDD(VDD),.Y(I14884),.A(g9454));
  NOT NOT1_2786(.VSS(VSS),.VDD(VDD),.Y(g11412),.A(I17277));
  NOT NOT1_2787(.VSS(VSS),.VDD(VDD),.Y(I11817),.A(g7246));
  NOT NOT1_2788(.VSS(VSS),.VDD(VDD),.Y(I10168),.A(g5982));
  NOT NOT1_2789(.VSS(VSS),.VDD(VDD),.Y(g5101),.A(I8473));
  NOT NOT1_2790(.VSS(VSS),.VDD(VDD),.Y(g5817),.A(I9427));
  NOT NOT1_2791(.VSS(VSS),.VDD(VDD),.Y(I11322),.A(g6652));
  NOT NOT1_2792(.VSS(VSS),.VDD(VDD),.Y(g7918),.A(g7505));
  NOT NOT1_2793(.VSS(VSS),.VDD(VDD),.Y(g5301),.A(g4373));
  NOT NOT1_2794(.VSS(VSS),.VDD(VDD),.Y(g7967),.A(I12765));
  NOT NOT1_2795(.VSS(VSS),.VDD(VDD),.Y(g6262),.A(I10045));
  NOT NOT1_2796(.VSS(VSS),.VDD(VDD),.Y(I15229),.A(g9968));
  NOT NOT1_2797(.VSS(VSS),.VDD(VDD),.Y(g2351),.A(I5427));
  NOT NOT1_2798(.VSS(VSS),.VDD(VDD),.Y(I11159),.A(g6478));
  NOT NOT1_2799(.VSS(VSS),.VDD(VDD),.Y(g10700),.A(I16379));
  NOT NOT1_2800(.VSS(VSS),.VDD(VDD),.Y(g2648),.A(I5765));
  NOT NOT1_2801(.VSS(VSS),.VDD(VDD),.Y(I9491),.A(g5072));
  NOT NOT1_2802(.VSS(VSS),.VDD(VDD),.Y(g10126),.A(I15380));
  NOT NOT1_2803(.VSS(VSS),.VDD(VDD),.Y(I8024),.A(g4117));
  NOT NOT1_2804(.VSS(VSS),.VDD(VDD),.Y(I11901),.A(g6897));
  NOT NOT1_2805(.VSS(VSS),.VDD(VDD),.Y(I16802),.A(g10902));
  NOT NOT1_2806(.VSS(VSS),.VDD(VDD),.Y(g2530),.A(I5641));
  NOT NOT1_2807(.VSS(VSS),.VDD(VDD),.Y(g6736),.A(I10739));
  NOT NOT1_2808(.VSS(VSS),.VDD(VDD),.Y(I13125),.A(g7975));
  NOT NOT1_2809(.VSS(VSS),.VDD(VDD),.Y(g8750),.A(I14045));
  NOT NOT1_2810(.VSS(VSS),.VDD(VDD),.Y(I10666),.A(g6042));
  NOT NOT1_2811(.VSS(VSS),.VDD(VDD),.Y(g4508),.A(g3946));
  NOT NOT1_2812(.VSS(VSS),.VDD(VDD),.Y(g10250),.A(g10136));
  NOT NOT1_2813(.VSS(VSS),.VDD(VDD),.Y(g2655),.A(g2013));
  NOT NOT1_2814(.VSS(VSS),.VDD(VDD),.Y(g4944),.A(g4430));
  NOT NOT1_2815(.VSS(VSS),.VDD(VDD),.Y(g4240),.A(g3664));
  NOT NOT1_2816(.VSS(VSS),.VDD(VDD),.Y(I11783),.A(g7246));
  NOT NOT1_2817(.VSS(VSS),.VDD(VDD),.Y(I16793),.A(g11014));
  NOT NOT1_2818(.VSS(VSS),.VDD(VDD),.Y(I7342),.A(g4011));
  NOT NOT1_2819(.VSS(VSS),.VDD(VDD),.Y(I9602),.A(g5013));
  NOT NOT1_2820(.VSS(VSS),.VDD(VDD),.Y(g4472),.A(I7847));
  NOT NOT1_2821(.VSS(VSS),.VDD(VDD),.Y(I10015),.A(g5641));
  NOT NOT1_2822(.VSS(VSS),.VDD(VDD),.Y(I5704),.A(g2056));
  NOT NOT1_2823(.VSS(VSS),.VDD(VDD),.Y(g7993),.A(I12813));
  NOT NOT1_2824(.VSS(VSS),.VDD(VDD),.Y(I7255),.A(g3227));
  NOT NOT1_2825(.VSS(VSS),.VDD(VDD),.Y(g6076),.A(I9717));
  NOT NOT1_2826(.VSS(VSS),.VDD(VDD),.Y(I4906),.A(g119));
  NOT NOT1_2827(.VSS(VSS),.VDD(VDD),.Y(I11656),.A(g7122));
  NOT NOT1_2828(.VSS(VSS),.VDD(VDD),.Y(I6049),.A(g2219));
  NOT NOT1_2829(.VSS(VSS),.VDD(VDD),.Y(g5751),.A(I9323));
  NOT NOT1_2830(.VSS(VSS),.VDD(VDD),.Y(g3758),.A(I6955));
  NOT NOT1_2831(.VSS(VSS),.VDD(VDD),.Y(g3066),.A(g2135));
  NOT NOT1_2832(.VSS(VSS),.VDD(VDD),.Y(I8231),.A(g4170));
  NOT NOT1_2833(.VSS(VSS),.VDD(VDD),.Y(g4443),.A(g3359));
  NOT NOT1_2834(.VSS(VSS),.VDD(VDD),.Y(g10296),.A(I15708));
  NOT NOT1_2835(.VSS(VSS),.VDD(VDD),.Y(g8440),.A(I13618));
  NOT NOT1_2836(.VSS(VSS),.VDD(VDD),.Y(I11680),.A(g7064));
  NOT NOT1_2837(.VSS(VSS),.VDD(VDD),.Y(g8969),.A(I14340));
  NOT NOT1_2838(.VSS(VSS),.VDD(VDD),.Y(I17116),.A(g11229));
  NOT NOT1_2839(.VSS(VSS),.VDD(VDD),.Y(g2410),.A(g1453));
  NOT NOT1_2840(.VSS(VSS),.VDD(VDD),.Y(g9679),.A(g9452));
  NOT NOT1_2841(.VSS(VSS),.VDD(VDD),.Y(I7726),.A(g3378));
  NOT NOT1_2842(.VSS(VSS),.VDD(VDD),.Y(g6175),.A(g5320));
  NOT NOT1_2843(.VSS(VSS),.VDD(VDD),.Y(g4116),.A(I7260));
  NOT NOT1_2844(.VSS(VSS),.VDD(VDD),.Y(I7154),.A(g2617));
  NOT NOT1_2845(.VSS(VSS),.VDD(VDD),.Y(g8323),.A(I13351));
  NOT NOT1_2846(.VSS(VSS),.VDD(VDD),.Y(g6871),.A(g6724));
  NOT NOT1_2847(.VSS(VSS),.VDD(VDD),.Y(g2884),.A(I6040));
  NOT NOT1_2848(.VSS(VSS),.VDD(VDD),.Y(I7354),.A(g4066));
  NOT NOT1_2849(.VSS(VSS),.VDD(VDD),.Y(g2839),.A(I5957));
  NOT NOT1_2850(.VSS(VSS),.VDD(VDD),.Y(g3365),.A(I6553));
  NOT NOT1_2851(.VSS(VSS),.VDD(VDD),.Y(g3861),.A(I7054));
  NOT NOT1_2852(.VSS(VSS),.VDD(VDD),.Y(I6498),.A(g2958));
  NOT NOT1_2853(.VSS(VSS),.VDD(VDD),.Y(I17746),.A(g11643));
  NOT NOT1_2854(.VSS(VSS),.VDD(VDD),.Y(g3055),.A(g2135));
  NOT NOT1_2855(.VSS(VSS),.VDD(VDD),.Y(I5053),.A(g1188));
  NOT NOT1_2856(.VSS(VSS),.VDD(VDD),.Y(I15959),.A(g10402));
  NOT NOT1_2857(.VSS(VSS),.VDD(VDD),.Y(g6285),.A(I10114));
  NOT NOT1_2858(.VSS(VSS),.VDD(VDD),.Y(g11627),.A(I17695));
  NOT NOT1_2859(.VSS(VSS),.VDD(VDD),.Y(g7921),.A(g7463));
  NOT NOT1_2860(.VSS(VSS),.VDD(VDD),.Y(g10197),.A(I15565));
  NOT NOT1_2861(.VSS(VSS),.VDD(VDD),.Y(g5673),.A(I9180));
  NOT NOT1_2862(.VSS(VSS),.VDD(VDD),.Y(g4347),.A(g3880));
  NOT NOT1_2863(.VSS(VSS),.VDD(VDD),.Y(I8551),.A(g4342));
  NOT NOT1_2864(.VSS(VSS),.VDD(VDD),.Y(I10084),.A(g5742));
  NOT NOT1_2865(.VSS(VSS),.VDD(VDD),.Y(g2172),.A(g43));
  NOT NOT1_2866(.VSS(VSS),.VDD(VDD),.Y(g3333),.A(g2779));
  NOT NOT1_2867(.VSS(VSS),.VDD(VDD),.Y(I9415),.A(g5047));
  NOT NOT1_2868(.VSS(VSS),.VDD(VDD),.Y(g11112),.A(I16897));
  NOT NOT1_2869(.VSS(VSS),.VDD(VDD),.Y(I17237),.A(g11394));
  NOT NOT1_2870(.VSS(VSS),.VDD(VDD),.Y(g4681),.A(g3546));
  NOT NOT1_2871(.VSS(VSS),.VDD(VDD),.Y(g10870),.A(I16580));
  NOT NOT1_2872(.VSS(VSS),.VDD(VDD),.Y(g11050),.A(I16811));
  NOT NOT1_2873(.VSS(VSS),.VDD(VDD),.Y(I8499),.A(g4330));
  NOT NOT1_2874(.VSS(VSS),.VDD(VDD),.Y(I12577),.A(g7532));
  NOT NOT1_2875(.VSS(VSS),.VDD(VDD),.Y(g8151),.A(g8036));
  NOT NOT1_2876(.VSS(VSS),.VDD(VDD),.Y(g10527),.A(g10462));
  NOT NOT1_2877(.VSS(VSS),.VDD(VDD),.Y(g3774),.A(I6999));
  NOT NOT1_2878(.VSS(VSS),.VDD(VDD),.Y(g8351),.A(I13433));
  NOT NOT1_2879(.VSS(VSS),.VDD(VDD),.Y(I17340),.A(g11366));
  NOT NOT1_2880(.VSS(VSS),.VDD(VDD),.Y(g4533),.A(I7938));
  NOT NOT1_2881(.VSS(VSS),.VDD(VDD),.Y(I13017),.A(g7848));
  NOT NOT1_2882(.VSS(VSS),.VDD(VDD),.Y(I13364),.A(g8221));
  NOT NOT1_2883(.VSS(VSS),.VDD(VDD),.Y(I15386),.A(g10101));
  NOT NOT1_2884(.VSS(VSS),.VDD(VDD),.Y(g6184),.A(I9915));
  NOT NOT1_2885(.VSS(VSS),.VDD(VDD),.Y(g2235),.A(g96));
  NOT NOT1_2886(.VSS(VSS),.VDD(VDD),.Y(g2343),.A(g1927));
  NOT NOT1_2887(.VSS(VSS),.VDD(VDD),.Y(I12439),.A(g7663));
  NOT NOT1_2888(.VSS(VSS),.VDD(VDD),.Y(g5669),.A(I9168));
  NOT NOT1_2889(.VSS(VSS),.VDD(VDD),.Y(I10531),.A(g6169));
  NOT NOT1_2890(.VSS(VSS),.VDD(VDD),.Y(I17684),.A(g11609));
  NOT NOT1_2891(.VSS(VSS),.VDD(VDD),.Y(g6339),.A(I10240));
  NOT NOT1_2892(.VSS(VSS),.VDD(VDD),.Y(I14179),.A(g8785));
  NOT NOT1_2893(.VSS(VSS),.VDD(VDD),.Y(g4210),.A(I7447));
  NOT NOT1_2894(.VSS(VSS),.VDD(VDD),.Y(I14531),.A(g9273));
  NOT NOT1_2895(.VSS(VSS),.VDD(VDD),.Y(I7112),.A(g3186));
  NOT NOT1_2896(.VSS(VSS),.VDD(VDD),.Y(I17142),.A(g11301));
  NOT NOT1_2897(.VSS(VSS),.VDD(VDD),.Y(g11096),.A(I16879));
  NOT NOT1_2898(.VSS(VSS),.VDD(VDD),.Y(g7620),.A(I12208));
  NOT NOT1_2899(.VSS(VSS),.VDD(VDD),.Y(g4596),.A(I8007));
  NOT NOT1_2900(.VSS(VSS),.VDD(VDD),.Y(g3538),.A(I6726));
  NOT NOT1_2901(.VSS(VSS),.VDD(VDD),.Y(I6019),.A(g2554));
  NOT NOT1_2902(.VSS(VSS),.VDD(VDD),.Y(g4013),.A(I7157));
  NOT NOT1_2903(.VSS(VSS),.VDD(VDD),.Y(g6424),.A(g6140));
  NOT NOT1_2904(.VSS(VSS),.VDD(VDD),.Y(I16626),.A(g10859));
  NOT NOT1_2905(.VSS(VSS),.VDD(VDD),.Y(I10186),.A(g6110));
  NOT NOT1_2906(.VSS(VSS),.VDD(VDD),.Y(g6737),.A(g6016));
  NOT NOT1_2907(.VSS(VSS),.VDD(VDD),.Y(g10867),.A(I16571));
  NOT NOT1_2908(.VSS(VSS),.VDD(VDD),.Y(g2334),.A(I5388));
  NOT NOT1_2909(.VSS(VSS),.VDD(VDD),.Y(g10894),.A(I16644));
  NOT NOT1_2910(.VSS(VSS),.VDD(VDD),.Y(g6809),.A(I10837));
  NOT NOT1_2911(.VSS(VSS),.VDD(VDD),.Y(I10685),.A(g6054));
  NOT NOT1_2912(.VSS(VSS),.VDD(VDD),.Y(g5743),.A(I9311));
  NOT NOT1_2913(.VSS(VSS),.VDD(VDD),.Y(g4413),.A(I7749));
  NOT NOT1_2914(.VSS(VSS),.VDD(VDD),.Y(g5890),.A(g5361));
  NOT NOT1_2915(.VSS(VSS),.VDD(VDD),.Y(I11289),.A(g6508));
  NOT NOT1_2916(.VSS(VSS),.VDD(VDD),.Y(I6052),.A(g2220));
  NOT NOT1_2917(.VSS(VSS),.VDD(VDD),.Y(g2548),.A(I5667));
  NOT NOT1_2918(.VSS(VSS),.VDD(VDD),.Y(I14373),.A(g8956));
  NOT NOT1_2919(.VSS(VSS),.VDD(VDD),.Y(I11309),.A(g6531));
  NOT NOT1_2920(.VSS(VSS),.VDD(VDD),.Y(I5929),.A(g2225));
  NOT NOT1_2921(.VSS(VSS),.VDD(VDD),.Y(I13023),.A(g8050));
  NOT NOT1_2922(.VSS(VSS),.VDD(VDD),.Y(g8884),.A(I14224));
  NOT NOT1_2923(.VSS(VSS),.VDD(VDD),.Y(I16298),.A(g10553));
  NOT NOT1_2924(.VSS(VSS),.VDD(VDD),.Y(I13224),.A(g8261));
  NOT NOT1_2925(.VSS(VSS),.VDD(VDD),.Y(g7788),.A(I12529));
  NOT NOT1_2926(.VSS(VSS),.VDD(VDD),.Y(g6077),.A(I9720));
  NOT NOT1_2927(.VSS(VSS),.VDD(VDD),.Y(g11429),.A(I17340));
  NOT NOT1_2928(.VSS(VSS),.VDD(VDD),.Y(g5011),.A(I8385));
  NOT NOT1_2929(.VSS(VSS),.VDD(VDD),.Y(I16775),.A(g10889));
  NOT NOT1_2930(.VSS(VSS),.VDD(VDD),.Y(g3067),.A(I6273));
  NOT NOT1_2931(.VSS(VSS),.VDD(VDD),.Y(I13571),.A(g8355));
  NOT NOT1_2932(.VSS(VSS),.VDD(VDD),.Y(g10315),.A(g10243));
  NOT NOT1_2933(.VSS(VSS),.VDD(VDD),.Y(g5856),.A(g5245));
  NOT NOT1_2934(.VSS(VSS),.VDD(VDD),.Y(g5734),.A(I9290));
  NOT NOT1_2935(.VSS(VSS),.VDD(VDD),.Y(g10819),.A(I16525));
  NOT NOT1_2936(.VSS(VSS),.VDD(VDD),.Y(g11428),.A(I17337));
  NOT NOT1_2937(.VSS(VSS),.VDD(VDD),.Y(g10910),.A(I16682));
  NOT NOT1_2938(.VSS(VSS),.VDD(VDD),.Y(g3290),.A(I6461));
  NOT NOT1_2939(.VSS(VSS),.VDD(VDD),.Y(I17362),.A(g11376));
  NOT NOT1_2940(.VSS(VSS),.VDD(VDD),.Y(g10202),.A(g10171));
  NOT NOT1_2941(.VSS(VSS),.VDD(VDD),.Y(I10334),.A(g6003));
  NOT NOT1_2942(.VSS(VSS),.VDD(VDD),.Y(g10257),.A(g10197));
  NOT NOT1_2943(.VSS(VSS),.VDD(VDD),.Y(g4317),.A(I7586));
  NOT NOT1_2944(.VSS(VSS),.VDD(VDD),.Y(g8278),.A(I13206));
  NOT NOT1_2945(.VSS(VSS),.VDD(VDD),.Y(I4876),.A(g580));
  NOT NOT1_2946(.VSS(VSS),.VDD(VDD),.Y(g3093),.A(I6299));
  NOT NOT1_2947(.VSS(VSS),.VDD(VDD),.Y(g1998),.A(g802));
  NOT NOT1_2948(.VSS(VSS),.VDD(VDD),.Y(g5474),.A(I8889));
  NOT NOT1_2949(.VSS(VSS),.VDD(VDD),.Y(g10111),.A(I15347));
  NOT NOT1_2950(.VSS(VSS),.VDD(VDD),.Y(g7192),.A(g6742));
  NOT NOT1_2951(.VSS(VSS),.VDD(VDD),.Y(g5992),.A(I9608));
  NOT NOT1_2952(.VSS(VSS),.VDD(VDD),.Y(g7085),.A(I11318));
  NOT NOT1_2953(.VSS(VSS),.VDD(VDD),.Y(g3256),.A(I6424));
  NOT NOT1_2954(.VSS(VSS),.VDD(VDD),.Y(I7746),.A(g3763));
  NOT NOT1_2955(.VSS(VSS),.VDD(VDD),.Y(g6634),.A(I10589));
  NOT NOT1_2956(.VSS(VSS),.VDD(VDD),.Y(I9188),.A(g4908));
  NOT NOT1_2957(.VSS(VSS),.VDD(VDD),.Y(I10762),.A(g6127));
  NOT NOT1_2958(.VSS(VSS),.VDD(VDD),.Y(g8667),.A(I13952));
  NOT NOT1_2959(.VSS(VSS),.VDD(VDD),.Y(g3816),.A(g3228));
  NOT NOT1_2960(.VSS(VSS),.VDD(VDD),.Y(g8143),.A(g8029));
  NOT NOT1_2961(.VSS(VSS),.VDD(VDD),.Y(I13816),.A(g8559));
  NOT NOT1_2962(.VSS(VSS),.VDD(VDD),.Y(I15548),.A(g10083));
  NOT NOT1_2963(.VSS(VSS),.VDD(VDD),.Y(I6504),.A(g3214));
  NOT NOT1_2964(.VSS(VSS),.VDD(VDD),.Y(I9388),.A(g5576));
  NOT NOT1_2965(.VSS(VSS),.VDD(VDD),.Y(g8235),.A(g7967));
  NOT NOT1_2966(.VSS(VSS),.VDD(VDD),.Y(g8343),.A(I13409));
  NOT NOT1_2967(.VSS(VSS),.VDD(VDD),.Y(g6742),.A(g5830));
  NOT NOT1_2968(.VSS(VSS),.VDD(VDD),.Y(g11548),.A(g11519));
  NOT NOT1_2969(.VSS(VSS),.VDD(VDD),.Y(g6104),.A(I9769));
  NOT NOT1_2970(.VSS(VSS),.VDD(VDD),.Y(I14964),.A(g9762));
  NOT NOT1_2971(.VSS(VSS),.VDD(VDD),.Y(g10590),.A(I16255));
  NOT NOT1_2972(.VSS(VSS),.VDD(VDD),.Y(I9216),.A(g4935));
  NOT NOT1_2973(.VSS(VSS),.VDD(VDD),.Y(I6385),.A(g2260));
  NOT NOT1_2974(.VSS(VSS),.VDD(VDD),.Y(g6304),.A(I10171));
  NOT NOT1_2975(.VSS(VSS),.VDD(VDD),.Y(I16856),.A(g10909));
  NOT NOT1_2976(.VSS(VSS),.VDD(VDD),.Y(g8566),.A(I13791));
  NOT NOT1_2977(.VSS(VSS),.VDD(VDD),.Y(g6499),.A(g5867));
  NOT NOT1_2978(.VSS(VSS),.VDD(VDD),.Y(I16261),.A(g10556));
  NOT NOT1_2979(.VSS(VSS),.VDD(VDD),.Y(g2202),.A(g148));
  NOT NOT1_2980(.VSS(VSS),.VDD(VDD),.Y(g11504),.A(I17531));
  NOT NOT1_2981(.VSS(VSS),.VDD(VDD),.Y(g8988),.A(I14385));
  NOT NOT1_2982(.VSS(VSS),.VDD(VDD),.Y(g4775),.A(I8139));
  NOT NOT1_2983(.VSS(VSS),.VDD(VDD),.Y(I11752),.A(g7032));
  NOT NOT1_2984(.VSS(VSS),.VDD(VDD),.Y(g8134),.A(I13005));
  NOT NOT1_2985(.VSS(VSS),.VDD(VDD),.Y(g7941),.A(g7406));
  NOT NOT1_2986(.VSS(VSS),.VDD(VDD),.Y(I15317),.A(g10025));
  NOT NOT1_2987(.VSS(VSS),.VDD(VDD),.Y(I6025),.A(g2259));
  NOT NOT1_2988(.VSS(VSS),.VDD(VDD),.Y(g2908),.A(I6077));
  NOT NOT1_2989(.VSS(VSS),.VDD(VDD),.Y(g8334),.A(I13382));
  NOT NOT1_2990(.VSS(VSS),.VDD(VDD),.Y(g9265),.A(g8892));
  NOT NOT1_2991(.VSS(VSS),.VDD(VDD),.Y(g6926),.A(I11046));
  NOT NOT1_2992(.VSS(VSS),.VDD(VDD),.Y(g2094),.A(I4924));
  NOT NOT1_2993(.VSS(VSS),.VDD(VDD),.Y(I12415),.A(g7631));
  NOT NOT1_2994(.VSS(VSS),.VDD(VDD),.Y(g11317),.A(I17112));
  NOT NOT1_2995(.VSS(VSS),.VDD(VDD),.Y(g10094),.A(I15329));
  NOT NOT1_2996(.VSS(VSS),.VDD(VDD),.Y(g3397),.A(g2896));
  NOT NOT1_2997(.VSS(VSS),.VDD(VDD),.Y(g8548),.A(g8390));
  NOT NOT1_2998(.VSS(VSS),.VDD(VDD),.Y(g2518),.A(g590));
  NOT NOT1_2999(.VSS(VSS),.VDD(VDD),.Y(g4060),.A(g3144));
  NOT NOT1_3000(.VSS(VSS),.VDD(VDD),.Y(g4460),.A(g3820));
  NOT NOT1_3001(.VSS(VSS),.VDD(VDD),.Y(I9564),.A(g5109));
  NOT NOT1_3002(.VSS(VSS),.VDD(VDD),.Y(I7468),.A(g3697));
  NOT NOT1_3003(.VSS(VSS),.VDD(VDD),.Y(g6273),.A(I10078));
  NOT NOT1_3004(.VSS(VSS),.VDD(VDD),.Y(I8885),.A(g4548));
  NOT NOT1_3005(.VSS(VSS),.VDD(VDD),.Y(g8804),.A(I14133));
  NOT NOT1_3006(.VSS(VSS),.VDD(VDD),.Y(I14543),.A(g9311));
  NOT NOT1_3007(.VSS(VSS),.VDD(VDD),.Y(I8414),.A(g4293));
  NOT NOT1_3008(.VSS(VSS),.VDD(VDD),.Y(g10150),.A(I15448));
  NOT NOT1_3009(.VSS(VSS),.VDD(VDD),.Y(g10801),.A(I16507));
  NOT NOT1_3010(.VSS(VSS),.VDD(VDD),.Y(I9826),.A(g5390));
  NOT NOT1_3011(.VSS(VSS),.VDD(VDD),.Y(I10117),.A(g6241));
  NOT NOT1_3012(.VSS(VSS),.VDD(VDD),.Y(g7708),.A(I12339));
  NOT NOT1_3013(.VSS(VSS),.VDD(VDD),.Y(I13669),.A(g8294));
  NOT NOT1_3014(.VSS(VSS),.VDD(VDD),.Y(g10735),.A(I16416));
  NOT NOT1_3015(.VSS(VSS),.VDD(VDD),.Y(g10877),.A(I16601));
  NOT NOT1_3016(.VSS(VSS),.VDD(VDD),.Y(g11057),.A(g10937));
  NOT NOT1_3017(.VSS(VSS),.VDD(VDD),.Y(g7520),.A(I11898));
  NOT NOT1_3018(.VSS(VSS),.VDD(VDD),.Y(g8792),.A(I14105));
  NOT NOT1_3019(.VSS(VSS),.VDD(VDD),.Y(I17347),.A(g11373));
  NOT NOT1_3020(.VSS(VSS),.VDD(VDD),.Y(I7677),.A(g3735));
  NOT NOT1_3021(.VSS(VSS),.VDD(VDD),.Y(I11668),.A(g7043));
  NOT NOT1_3022(.VSS(VSS),.VDD(VDD),.Y(g6044),.A(I9665));
  NOT NOT1_3023(.VSS(VSS),.VDD(VDD),.Y(g2593),.A(g1973));
  NOT NOT1_3024(.VSS(VSS),.VDD(VDD),.Y(g7031),.A(g6413));
  NOT NOT1_3025(.VSS(VSS),.VDD(VDD),.Y(g4739),.A(g4117));
  NOT NOT1_3026(.VSS(VSS),.VDD(VDD),.Y(I8903),.A(g4561));
  NOT NOT1_3027(.VSS(VSS),.VDD(VDD),.Y(g6444),.A(g6158));
  NOT NOT1_3028(.VSS(VSS),.VDD(VDD),.Y(g11245),.A(g11112));
  NOT NOT1_3029(.VSS(VSS),.VDD(VDD),.Y(g7431),.A(I11821));
  NOT NOT1_3030(.VSS(VSS),.VDD(VDD),.Y(I15323),.A(g10019));
  NOT NOT1_3031(.VSS(VSS),.VDD(VDD),.Y(g6269),.A(I10066));
  NOT NOT1_3032(.VSS(VSS),.VDD(VDD),.Y(I15299),.A(g9995));
  NOT NOT1_3033(.VSS(VSS),.VDD(VDD),.Y(g7812),.A(I12601));
  NOT NOT1_3034(.VSS(VSS),.VDD(VDD),.Y(g11626),.A(I17692));
  NOT NOT1_3035(.VSS(VSS),.VDD(VDD),.Y(g9770),.A(g9432));
  NOT NOT1_3036(.VSS(VSS),.VDD(VDD),.Y(g10196),.A(I15562));
  NOT NOT1_3037(.VSS(VSS),.VDD(VDD),.Y(I11489),.A(g6569));
  NOT NOT1_3038(.VSS(VSS),.VDD(VDD),.Y(g10695),.A(I16366));
  NOT NOT1_3039(.VSS(VSS),.VDD(VDD),.Y(g5688),.A(I9213));
  NOT NOT1_3040(.VSS(VSS),.VDD(VDD),.Y(g11323),.A(I17124));
  NOT NOT1_3041(.VSS(VSS),.VDD(VDD),.Y(I13489),.A(g8233));
  NOT NOT1_3042(.VSS(VSS),.VDD(VDD),.Y(g2965),.A(I6196));
  NOT NOT1_3043(.VSS(VSS),.VDD(VDD),.Y(I6406),.A(g2339));
  NOT NOT1_3044(.VSS(VSS),.VDD(VDD),.Y(I5475),.A(g1289));
  NOT NOT1_3045(.VSS(VSS),.VDD(VDD),.Y(I7716),.A(g3751));
  NOT NOT1_3046(.VSS(VSS),.VDD(VDD),.Y(g6572),.A(g5805));
  NOT NOT1_3047(.VSS(VSS),.VDD(VDD),.Y(g6862),.A(g6720));
  NOT NOT1_3048(.VSS(VSS),.VDD(VDD),.Y(g7376),.A(I11756));
  NOT NOT1_3049(.VSS(VSS),.VDD(VDD),.Y(I5949),.A(g2540));
  NOT NOT1_3050(.VSS(VSS),.VDD(VDD),.Y(g10526),.A(g10460));
  NOT NOT1_3051(.VSS(VSS),.VDD(VDD),.Y(g8313),.A(I13323));
  NOT NOT1_3052(.VSS(VSS),.VDD(VDD),.Y(I12484),.A(g7580));
  NOT NOT1_3053(.VSS(VSS),.VDD(VDD),.Y(I14242),.A(g8787));
  NOT NOT1_3054(.VSS(VSS),.VDD(VDD),.Y(I9108),.A(g5593));
  NOT NOT1_3055(.VSS(VSS),.VDD(VDD),.Y(I15775),.A(g10253));
  NOT NOT1_3056(.VSS(VSS),.VDD(VDD),.Y(I13424),.A(g8200));
  NOT NOT1_3057(.VSS(VSS),.VDD(VDD),.Y(g4479),.A(I7858));
  NOT NOT1_3058(.VSS(VSS),.VDD(VDD),.Y(g9532),.A(I14681));
  NOT NOT1_3059(.VSS(VSS),.VDD(VDD),.Y(I9308),.A(g5494));
  NOT NOT1_3060(.VSS(VSS),.VDD(VDD),.Y(g6712),.A(g5984));
  NOT NOT1_3061(.VSS(VSS),.VDD(VDD),.Y(I8036),.A(g3820));
  NOT NOT1_3062(.VSS(VSS),.VDD(VDD),.Y(g4294),.A(g3664));
  NOT NOT1_3063(.VSS(VSS),.VDD(VDD),.Y(I10123),.A(g5676));
  NOT NOT1_3064(.VSS(VSS),.VDD(VDD),.Y(g6543),.A(g5888));
  NOT NOT1_3065(.VSS(VSS),.VDD(VDD),.Y(g4840),.A(I8199));
  NOT NOT1_3066(.VSS(VSS),.VDD(VDD),.Y(I8436),.A(g4462));
  NOT NOT1_3067(.VSS(VSS),.VDD(VDD),.Y(g9553),.A(I14694));
  NOT NOT1_3068(.VSS(VSS),.VDD(VDD),.Y(I5292),.A(g76));
  NOT NOT1_3069(.VSS(VSS),.VDD(VDD),.Y(I9883),.A(g5557));
  NOT NOT1_3070(.VSS(VSS),.VDD(VDD),.Y(I14123),.A(g8767));
  NOT NOT1_3071(.VSS(VSS),.VDD(VDD),.Y(g3723),.A(g3071));
  NOT NOT1_3072(.VSS(VSS),.VDD(VDD),.Y(g7765),.A(I12460));
  NOT NOT1_3073(.VSS(VSS),.VDD(VDD),.Y(g7286),.A(I11534));
  NOT NOT1_3074(.VSS(VSS),.VDD(VDD),.Y(g4190),.A(I7387));
  NOT NOT1_3075(.VSS(VSS),.VDD(VDD),.Y(I5998),.A(g2197));
  NOT NOT1_3076(.VSS(VSS),.VDD(VDD),.Y(g4390),.A(g3914));
  NOT NOT1_3077(.VSS(VSS),.VDD(VDD),.Y(I10807),.A(g6396));
  NOT NOT1_3078(.VSS(VSS),.VDD(VDD),.Y(g10457),.A(I15962));
  NOT NOT1_3079(.VSS(VSS),.VDD(VDD),.Y(g3817),.A(I7043));
  NOT NOT1_3080(.VSS(VSS),.VDD(VDD),.Y(g7911),.A(g7664));
  NOT NOT1_3081(.VSS(VSS),.VDD(VDD),.Y(I5646),.A(g940));
  NOT NOT1_3082(.VSS(VSS),.VDD(VDD),.Y(I10974),.A(g6563));
  NOT NOT1_3083(.VSS(VSS),.VDD(VDD),.Y(g8094),.A(g7987));
  NOT NOT1_3084(.VSS(VSS),.VDD(VDD),.Y(g2050),.A(g1861));
  NOT NOT1_3085(.VSS(VSS),.VDD(VDD),.Y(g2641),.A(g1987));
  NOT NOT1_3086(.VSS(VSS),.VDD(VDD),.Y(I8831),.A(g4480));
  NOT NOT1_3087(.VSS(VSS),.VDD(VDD),.Y(I15232),.A(g9974));
  NOT NOT1_3088(.VSS(VSS),.VDD(VDD),.Y(I10639),.A(g5830));
  NOT NOT1_3089(.VSS(VSS),.VDD(VDD),.Y(I17516),.A(g11483));
  NOT NOT1_3090(.VSS(VSS),.VDD(VDD),.Y(g2450),.A(g1351));
  NOT NOT1_3091(.VSS(VSS),.VDD(VDD),.Y(I16432),.A(g10702));
  NOT NOT1_3092(.VSS(VSS),.VDD(VDD),.Y(g4501),.A(g3946));
  NOT NOT1_3093(.VSS(VSS),.VDD(VDD),.Y(g8518),.A(I13723));
  NOT NOT1_3094(.VSS(VSS),.VDD(VDD),.Y(g6729),.A(I10724));
  NOT NOT1_3095(.VSS(VSS),.VDD(VDD),.Y(g6961),.A(I11115));
  NOT NOT1_3096(.VSS(VSS),.VDD(VDD),.Y(g8567),.A(I13794));
  NOT NOT1_3097(.VSS(VSS),.VDD(VDD),.Y(I10293),.A(g5863));
  NOT NOT1_3098(.VSS(VSS),.VDD(VDD),.Y(g4156),.A(I7295));
  NOT NOT1_3099(.VSS(VSS),.VDD(VDD),.Y(I11713),.A(g7023));
  NOT NOT1_3100(.VSS(VSS),.VDD(VDD),.Y(g7733),.A(I12380));
  NOT NOT1_3101(.VSS(VSS),.VDD(VDD),.Y(I5850),.A(g2273));
  NOT NOT1_3102(.VSS(VSS),.VDD(VDD),.Y(g7270),.A(I11515));
  NOT NOT1_3103(.VSS(VSS),.VDD(VDD),.Y(g9990),.A(I15190));
  NOT NOT1_3104(.VSS(VSS),.VDD(VDD),.Y(g6927),.A(I11049));
  NOT NOT1_3105(.VSS(VSS),.VDD(VDD),.Y(g3751),.A(I6944));
  NOT NOT1_3106(.VSS(VSS),.VDD(VDD),.Y(I9165),.A(g5037));
  NOT NOT1_3107(.VSS(VSS),.VDD(VDD),.Y(I16461),.A(g10735));
  NOT NOT1_3108(.VSS(VSS),.VDD(VDD),.Y(I9571),.A(g5509));
  NOT NOT1_3109(.VSS(VSS),.VDD(VDD),.Y(I9365),.A(g5392));
  NOT NOT1_3110(.VSS(VSS),.VDD(VDD),.Y(g7610),.A(I12180));
  NOT NOT1_3111(.VSS(VSS),.VDD(VDD),.Y(g2179),.A(g89));
  NOT NOT1_3112(.VSS(VSS),.VDD(VDD),.Y(g4942),.A(I8308));
  NOT NOT1_3113(.VSS(VSS),.VDD(VDD),.Y(g9029),.A(I14424));
  NOT NOT1_3114(.VSS(VSS),.VDD(VDD),.Y(g6014),.A(g5309));
  NOT NOT1_3115(.VSS(VSS),.VDD(VDD),.Y(g7073),.A(I11296));
  NOT NOT1_3116(.VSS(VSS),.VDD(VDD),.Y(I12799),.A(g7556));
  NOT NOT1_3117(.VSS(VSS),.VDD(VDD),.Y(g7796),.A(I12553));
  NOT NOT1_3118(.VSS(VSS),.VDD(VDD),.Y(I12813),.A(g7688));
  NOT NOT1_3119(.VSS(VSS),.VDD(VDD),.Y(g6885),.A(I10979));
  NOT NOT1_3120(.VSS(VSS),.VDD(VDD),.Y(g9429),.A(g9082));
  NOT NOT1_3121(.VSS(VSS),.VDD(VDD),.Y(g22),.A(I4777));
  NOT NOT1_3122(.VSS(VSS),.VDD(VDD),.Y(g7473),.A(g7148));
  NOT NOT1_3123(.VSS(VSS),.VDD(VDD),.Y(I10391),.A(g5838));
  NOT NOT1_3124(.VSS(VSS),.VDD(VDD),.Y(I17209),.A(g11289));
  NOT NOT1_3125(.VSS(VSS),.VDD(VDD),.Y(g6660),.A(I10623));
  NOT NOT1_3126(.VSS(VSS),.VDD(VDD),.Y(I11255),.A(g6547));
  NOT NOT1_3127(.VSS(VSS),.VDD(VDD),.Y(g10256),.A(g10140));
  NOT NOT1_3128(.VSS(VSS),.VDD(VDD),.Y(I6173),.A(g2125));
  NOT NOT1_3129(.VSS(VSS),.VDD(VDD),.Y(g11512),.A(I17555));
  NOT NOT1_3130(.VSS(VSS),.VDD(VDD),.Y(I13255),.A(g8270));
  NOT NOT1_3131(.VSS(VSS),.VDD(VDD),.Y(I14391),.A(g8928));
  NOT NOT1_3132(.VSS(VSS),.VDD(VDD),.Y(I16650),.A(g10776));
  NOT NOT1_3133(.VSS(VSS),.VDD(VDD),.Y(I6373),.A(g2024));
  NOT NOT1_3134(.VSS(VSS),.VDD(VDD),.Y(I6091),.A(g2270));
  NOT NOT1_3135(.VSS(VSS),.VDD(VDD),.Y(g5183),.A(g4640));
  NOT NOT1_3136(.VSS(VSS),.VDD(VDD),.Y(g7124),.A(I11363));
  NOT NOT1_3137(.VSS(VSS),.VDD(VDD),.Y(g7980),.A(I12786));
  NOT NOT1_3138(.VSS(VSS),.VDD(VDD),.Y(g7324),.A(I11620));
  NOT NOT1_3139(.VSS(VSS),.VDD(VDD),.Y(g10280),.A(g10160));
  NOT NOT1_3140(.VSS(VSS),.VDD(VDD),.Y(g6903),.A(I11005));
  NOT NOT1_3141(.VSS(VSS),.VDD(VDD),.Y(g2777),.A(g2276));
  NOT NOT1_3142(.VSS(VSS),.VDD(VDD),.Y(I5919),.A(g2530));
  NOT NOT1_3143(.VSS(VSS),.VDD(VDD),.Y(I11188),.A(g6513));
  NOT NOT1_3144(.VSS(VSS),.VDD(VDD),.Y(g7069),.A(I11286));
  NOT NOT1_3145(.VSS(VSS),.VDD(VDD),.Y(I12805),.A(g7684));
  NOT NOT1_3146(.VSS(VSS),.VDD(VDD),.Y(I13188),.A(g8171));
  NOT NOT1_3147(.VSS(VSS),.VDD(VDD),.Y(g5779),.A(I9371));
  NOT NOT1_3148(.VSS(VSS),.VDD(VDD),.Y(I13678),.A(g8306));
  NOT NOT1_3149(.VSS(VSS),.VDD(VDD),.Y(I14579),.A(g9272));
  NOT NOT1_3150(.VSS(VSS),.VDD(VDD),.Y(g4954),.A(g4509));
  NOT NOT1_3151(.VSS(VSS),.VDD(VDD),.Y(g4250),.A(g3698));
  NOT NOT1_3152(.VSS(VSS),.VDD(VDD),.Y(g4163),.A(I7308));
  NOT NOT1_3153(.VSS(VSS),.VDD(VDD),.Y(I5952),.A(g2506));
  NOT NOT1_3154(.VSS(VSS),.VDD(VDD),.Y(g2882),.A(I6034));
  NOT NOT1_3155(.VSS(VSS),.VDD(VDD),.Y(g7540),.A(I11956));
  NOT NOT1_3156(.VSS(VSS),.VDD(VDD),.Y(g8160),.A(I13057));
  NOT NOT1_3157(.VSS(VSS),.VDD(VDD),.Y(g4363),.A(I7654));
  NOT NOT1_3158(.VSS(VSS),.VDD(VDD),.Y(I11686),.A(g7039));
  NOT NOT1_3159(.VSS(VSS),.VDD(VDD),.Y(I16528),.A(g10732));
  NOT NOT1_3160(.VSS(VSS),.VDD(VDD),.Y(I7577),.A(g4124));
  NOT NOT1_3161(.VSS(VSS),.VDD(VDD),.Y(I5276),.A(g1411));
  NOT NOT1_3162(.VSS(VSS),.VDD(VDD),.Y(g8360),.A(I13460));
  NOT NOT1_3163(.VSS(VSS),.VDD(VDD),.Y(I16843),.A(g10898));
  NOT NOT1_3164(.VSS(VSS),.VDD(VDD),.Y(I6007),.A(g2199));
  NOT NOT1_3165(.VSS(VSS),.VDD(VDD),.Y(g5423),.A(g4300));
  NOT NOT1_3166(.VSS(VSS),.VDD(VDD),.Y(I13460),.A(g8155));
  NOT NOT1_3167(.VSS(VSS),.VDD(VDD),.Y(I17453),.A(g11451));
  NOT NOT1_3168(.VSS(VSS),.VDD(VDD),.Y(I11383),.A(g6385));
  NOT NOT1_3169(.VSS(VSS),.VDD(VDD),.Y(g2271),.A(g877));
  NOT NOT1_3170(.VSS(VSS),.VDD(VDD),.Y(g7377),.A(I11759));
  NOT NOT1_3171(.VSS(VSS),.VDD(VDD),.Y(g7206),.A(I11436));
  NOT NOT1_3172(.VSS(VSS),.VDD(VDD),.Y(g10157),.A(I15467));
  NOT NOT1_3173(.VSS(VSS),.VDD(VDD),.Y(g11445),.A(I17384));
  NOT NOT1_3174(.VSS(VSS),.VDD(VDD),.Y(g6036),.A(I9647));
  NOT NOT1_3175(.VSS(VSS),.VDD(VDD),.Y(I5561),.A(g869));
  NOT NOT1_3176(.VSS(VSS),.VDD(VDD),.Y(I13030),.A(g8052));
  NOT NOT1_3177(.VSS(VSS),.VDD(VDD),.Y(g2611),.A(I5734));
  NOT NOT1_3178(.VSS(VSS),.VDD(VDD),.Y(g4453),.A(I7810));
  NOT NOT1_3179(.VSS(VSS),.VDD(VDD),.Y(g8450),.A(I13648));
  NOT NOT1_3180(.VSS(VSS),.VDD(VDD),.Y(g6178),.A(g4977));
  NOT NOT1_3181(.VSS(VSS),.VDD(VDD),.Y(I6767),.A(g2914));
  NOT NOT1_3182(.VSS(VSS),.VDD(VDD),.Y(g11499),.A(I17516));
  NOT NOT1_3183(.VSS(VSS),.VDD(VDD),.Y(I8495),.A(g4325));
  NOT NOT1_3184(.VSS(VSS),.VDD(VDD),.Y(g3368),.A(g3138));
  NOT NOT1_3185(.VSS(VSS),.VDD(VDD),.Y(g9745),.A(g9454));
  NOT NOT1_3186(.VSS(VSS),.VDD(VDD),.Y(I11065),.A(g6750));
  NOT NOT1_3187(.VSS(VSS),.VDD(VDD),.Y(I6535),.A(g2826));
  NOT NOT1_3188(.VSS(VSS),.VDD(VDD),.Y(g1987),.A(g762));
  NOT NOT1_3189(.VSS(VSS),.VDD(VDD),.Y(g9338),.A(I14519));
  NOT NOT1_3190(.VSS(VSS),.VDD(VDD),.Y(g7287),.A(I11537));
  NOT NOT1_3191(.VSS(VSS),.VDD(VDD),.Y(g2799),.A(g2276));
  NOT NOT1_3192(.VSS(VSS),.VDD(VDD),.Y(g11498),.A(I17513));
  NOT NOT1_3193(.VSS(VSS),.VDD(VDD),.Y(I5986),.A(g2194));
  NOT NOT1_3194(.VSS(VSS),.VDD(VDD),.Y(g6135),.A(I9842));
  NOT NOT1_3195(.VSS(VSS),.VDD(VDD),.Y(g5665),.A(I9156));
  NOT NOT1_3196(.VSS(VSS),.VDD(VDD),.Y(g9109),.A(I14452));
  NOT NOT1_3197(.VSS(VSS),.VDD(VDD),.Y(g6335),.A(I10228));
  NOT NOT1_3198(.VSS(VSS),.VDD(VDD),.Y(I15989),.A(g10417));
  NOT NOT1_3199(.VSS(VSS),.VDD(VDD),.Y(g9309),.A(g8892));
  NOT NOT1_3200(.VSS(VSS),.VDD(VDD),.Y(g3531),.A(g2971));
  NOT NOT1_3201(.VSS(VSS),.VDD(VDD),.Y(I8869),.A(g4421));
  NOT NOT1_3202(.VSS(VSS),.VDD(VDD),.Y(g5127),.A(I8535));
  NOT NOT1_3203(.VSS(VSS),.VDD(VDD),.Y(g3458),.A(g3144));
  NOT NOT1_3204(.VSS(VSS),.VDD(VDD),.Y(g6182),.A(g5446));
  NOT NOT1_3205(.VSS(VSS),.VDD(VDD),.Y(g6288),.A(I10123));
  NOT NOT1_3206(.VSS(VSS),.VDD(VDD),.Y(I17274),.A(g11389));
  NOT NOT1_3207(.VSS(VSS),.VDD(VDD),.Y(g6382),.A(I10278));
  NOT NOT1_3208(.VSS(VSS),.VDD(VDD),.Y(I9662),.A(g5319));
  NOT NOT1_3209(.VSS(VSS),.VDD(VDD),.Y(g8179),.A(I13086));
  NOT NOT1_3210(.VSS(VSS),.VDD(VDD),.Y(g7849),.A(I12644));
  NOT NOT1_3211(.VSS(VSS),.VDD(VDD),.Y(g10876),.A(I16598));
  NOT NOT1_3212(.VSS(VSS),.VDD(VDD),.Y(g10885),.A(g10809));
  NOT NOT1_3213(.VSS(VSS),.VDD(VDD),.Y(g11056),.A(g10950));
  NOT NOT1_3214(.VSS(VSS),.VDD(VDD),.Y(g3743),.A(I6932));
  NOT NOT1_3215(.VSS(VSS),.VDD(VDD),.Y(g8379),.A(I13485));
  NOT NOT1_3216(.VSS(VSS),.VDD(VDD),.Y(g4912),.A(I8282));
  NOT NOT1_3217(.VSS(VSS),.VDD(VDD),.Y(I14116),.A(g8766));
  NOT NOT1_3218(.VSS(VSS),.VDD(VDD),.Y(g2997),.A(g2135));
  NOT NOT1_3219(.VSS(VSS),.VDD(VDD),.Y(g11611),.A(I17657));
  NOT NOT1_3220(.VSS(VSS),.VDD(VDD),.Y(I12400),.A(g7537));
  NOT NOT1_3221(.VSS(VSS),.VDD(VDD),.Y(g2541),.A(I5658));
  NOT NOT1_3222(.VSS(VSS),.VDD(VDD),.Y(g11080),.A(I16853));
  NOT NOT1_3223(.VSS(VSS),.VDD(VDD),.Y(I7426),.A(g3334));
  NOT NOT1_3224(.VSS(VSS),.VDD(VDD),.Y(I9290),.A(g5052));
  NOT NOT1_3225(.VSS(VSS),.VDD(VDD),.Y(g5146),.A(g4596));
  NOT NOT1_3226(.VSS(VSS),.VDD(VDD),.Y(g10854),.A(g10708));
  NOT NOT1_3227(.VSS(VSS),.VDD(VDD),.Y(g6805),.A(I10825));
  NOT NOT1_3228(.VSS(VSS),.VDD(VDD),.Y(g5633),.A(g4388));
  NOT NOT1_3229(.VSS(VSS),.VDD(VDD),.Y(g3505),.A(I6694));
  NOT NOT1_3230(.VSS(VSS),.VDD(VDD),.Y(g7781),.A(I12508));
  NOT NOT1_3231(.VSS(VSS),.VDD(VDD),.Y(I5970),.A(g2185));
  NOT NOT1_3232(.VSS(VSS),.VDD(VDD),.Y(g6749),.A(I10756));
  NOT NOT1_3233(.VSS(VSS),.VDD(VDD),.Y(I16708),.A(g10822));
  NOT NOT1_3234(.VSS(VSS),.VDD(VDD),.Y(g2238),.A(I5237));
  NOT NOT1_3235(.VSS(VSS),.VDD(VDD),.Y(g11432),.A(I17347));
  NOT NOT1_3236(.VSS(VSS),.VDD(VDD),.Y(I13837),.A(g8488));
  NOT NOT1_3237(.VSS(VSS),.VDD(VDD),.Y(g3411),.A(I6616));
  NOT NOT1_3238(.VSS(VSS),.VDD(VDD),.Y(I9093),.A(g5397));
  NOT NOT1_3239(.VSS(VSS),.VDD(VDD),.Y(g7900),.A(g7712));
  NOT NOT1_3240(.VSS(VSS),.VDD(VDD),.Y(I16258),.A(g10555));
  NOT NOT1_3241(.VSS(VSS),.VDD(VDD),.Y(I4948),.A(g586));
  NOT NOT1_3242(.VSS(VSS),.VDD(VDD),.Y(g2209),.A(g93));
  NOT NOT1_3243(.VSS(VSS),.VDD(VDD),.Y(g7797),.A(I12556));
  NOT NOT1_3244(.VSS(VSS),.VDD(VDD),.Y(I9256),.A(g5078));
  NOT NOT1_3245(.VSS(VSS),.VDD(VDD),.Y(I8265),.A(g4602));
  NOT NOT1_3246(.VSS(VSS),.VDD(VDD),.Y(I9816),.A(g5576));
  NOT NOT1_3247(.VSS(VSS),.VDD(VDD),.Y(g5696),.A(I9229));
  NOT NOT1_3248(.VSS(VSS),.VDD(VDD),.Y(I15461),.A(g10074));
  NOT NOT1_3249(.VSS(VSS),.VDD(VDD),.Y(g6947),.A(I11085));
  NOT NOT1_3250(.VSS(VSS),.VDD(VDD),.Y(I7984),.A(g3621));
  NOT NOT1_3251(.VSS(VSS),.VDD(VDD),.Y(I5224),.A(g61));
  NOT NOT1_3252(.VSS(VSS),.VDD(VDD),.Y(I7280),.A(g3208));
  NOT NOT1_3253(.VSS(VSS),.VDD(VDD),.Y(I10237),.A(g6120));
  NOT NOT1_3254(.VSS(VSS),.VDD(VDD),.Y(g6798),.A(I10804));
  NOT NOT1_3255(.VSS(VSS),.VDD(VDD),.Y(I8442),.A(g4464));
  NOT NOT1_3256(.VSS(VSS),.VDD(VDD),.Y(I12538),.A(g7658));
  NOT NOT1_3257(.VSS(VSS),.VDD(VDD),.Y(g8271),.A(I13185));
  NOT NOT1_3258(.VSS(VSS),.VDD(VDD),.Y(g2802),.A(g2276));
  NOT NOT1_3259(.VSS(VSS),.VDD(VDD),.Y(g11342),.A(I17149));
  NOT NOT1_3260(.VSS(VSS),.VDD(VDD),.Y(I10340),.A(g6205));
  NOT NOT1_3261(.VSS(VSS),.VDD(VDD),.Y(g1991),.A(g778));
  NOT NOT1_3262(.VSS(VSS),.VDD(VDD),.Y(I5120),.A(g622));
  NOT NOT1_3263(.VSS(VSS),.VDD(VDD),.Y(g3474),.A(I6679));
  NOT NOT1_3264(.VSS(VSS),.VDD(VDD),.Y(g9449),.A(g9094));
  NOT NOT1_3265(.VSS(VSS),.VDD(VDD),.Y(g6560),.A(g5759));
  NOT NOT1_3266(.VSS(VSS),.VDD(VDD),.Y(I14340),.A(g8820));
  NOT NOT1_3267(.VSS(VSS),.VDD(VDD),.Y(g5753),.A(I9329));
  NOT NOT1_3268(.VSS(VSS),.VDD(VDD),.Y(I8164),.A(g3566));
  NOT NOT1_3269(.VSS(VSS),.VDD(VDD),.Y(I15736),.A(g10258));
  NOT NOT1_3270(.VSS(VSS),.VDD(VDD),.Y(g10456),.A(I15959));
  NOT NOT1_3271(.VSS(VSS),.VDD(VDD),.Y(g5508),.A(I8929));
  NOT NOT1_3272(.VSS(VSS),.VDD(VDD),.Y(g11199),.A(g11112));
  NOT NOT1_3273(.VSS(VSS),.VDD(VDD),.Y(I14684),.A(g9124));
  NOT NOT1_3274(.VSS(VSS),.VDD(VDD),.Y(g11650),.A(I17752));
  NOT NOT1_3275(.VSS(VSS),.VDD(VDD),.Y(g7144),.A(I11387));
  NOT NOT1_3276(.VSS(VSS),.VDD(VDD),.Y(I11617),.A(g6839));
  NOT NOT1_3277(.VSS(VSS),.VDD(VDD),.Y(g7344),.A(I11680));
  NOT NOT1_3278(.VSS(VSS),.VDD(VDD),.Y(g5072),.A(I8442));
  NOT NOT1_3279(.VSS(VSS),.VDD(VDD),.Y(I7636),.A(g3330));
  NOT NOT1_3280(.VSS(VSS),.VDD(VDD),.Y(I13915),.A(g8451));
  NOT NOT1_3281(.VSS(VSS),.VDD(VDD),.Y(g5472),.A(I8885));
  NOT NOT1_3282(.VSS(VSS),.VDD(VDD),.Y(g8981),.A(I14364));
  NOT NOT1_3283(.VSS(VSS),.VDD(VDD),.Y(I9421),.A(g5063));
  NOT NOT1_3284(.VSS(VSS),.VDD(VDD),.Y(g8674),.A(I13959));
  NOT NOT1_3285(.VSS(VSS),.VDD(VDD),.Y(I5789),.A(g2162));
  NOT NOT1_3286(.VSS(VSS),.VDD(VDD),.Y(g5043),.A(g4840));
  NOT NOT1_3287(.VSS(VSS),.VDD(VDD),.Y(I11201),.A(g6522));
  NOT NOT1_3288(.VSS(VSS),.VDD(VDD),.Y(g10314),.A(I15744));
  NOT NOT1_3289(.VSS(VSS),.VDD(VDD),.Y(g7259),.A(I11494));
  NOT NOT1_3290(.VSS(VSS),.VDD(VDD),.Y(g5443),.A(I8872));
  NOT NOT1_3291(.VSS(VSS),.VDD(VDD),.Y(g6208),.A(I9953));
  NOT NOT1_3292(.VSS(VSS),.VDD(VDD),.Y(I7790),.A(g3782));
  NOT NOT1_3293(.VSS(VSS),.VDD(VDD),.Y(I16879),.A(g10936));
  NOT NOT1_3294(.VSS(VSS),.VDD(VDD),.Y(g6302),.A(I10165));
  NOT NOT1_3295(.VSS(VSS),.VDD(VDD),.Y(g10307),.A(I15729));
  NOT NOT1_3296(.VSS(VSS),.VDD(VDD),.Y(I15365),.A(g10025));
  NOT NOT1_3297(.VSS(VSS),.VDD(VDD),.Y(I7061),.A(g3050));
  NOT NOT1_3298(.VSS(VSS),.VDD(VDD),.Y(g6579),.A(g5949));
  NOT NOT1_3299(.VSS(VSS),.VDD(VDD),.Y(g5116),.A(g4682));
  NOT NOT1_3300(.VSS(VSS),.VDD(VDD),.Y(g6869),.A(I10949));
  NOT NOT1_3301(.VSS(VSS),.VDD(VDD),.Y(g7852),.A(g7479));
  NOT NOT1_3302(.VSS(VSS),.VDD(VDD),.Y(g7923),.A(g7527));
  NOT NOT1_3303(.VSS(VSS),.VDD(VDD),.Y(I17164),.A(g11320));
  NOT NOT1_3304(.VSS(VSS),.VDD(VDD),.Y(I7387),.A(g4083));
  NOT NOT1_3305(.VSS(VSS),.VDD(VDD),.Y(g10596),.A(I16269));
  NOT NOT1_3306(.VSS(VSS),.VDD(VDD),.Y(I11467),.A(g6488));
  NOT NOT1_3307(.VSS(VSS),.VDD(VDD),.Y(I11494),.A(g6574));
  NOT NOT1_3308(.VSS(VSS),.VDD(VDD),.Y(I13595),.A(g8339));
  NOT NOT1_3309(.VSS(VSS),.VDD(VDD),.Y(g8132),.A(I12999));
  NOT NOT1_3310(.VSS(VSS),.VDD(VDD),.Y(g6719),.A(I10710));
  NOT NOT1_3311(.VSS(VSS),.VDD(VDD),.Y(I12235),.A(g7082));
  NOT NOT1_3312(.VSS(VSS),.VDD(VDD),.Y(g8332),.A(I13376));
  NOT NOT1_3313(.VSS(VSS),.VDD(VDD),.Y(g10243),.A(I15635));
  NOT NOT1_3314(.VSS(VSS),.VDD(VDD),.Y(I11623),.A(g6841));
  NOT NOT1_3315(.VSS(VSS),.VDD(VDD),.Y(I12683),.A(g7387));
  NOT NOT1_3316(.VSS(VSS),.VDD(VDD),.Y(I6388),.A(g2329));
  NOT NOT1_3317(.VSS(VSS),.VDD(VDD),.Y(g8680),.A(I13965));
  NOT NOT1_3318(.VSS(VSS),.VDD(VDD),.Y(g10431),.A(g10328));
  NOT NOT1_3319(.VSS(VSS),.VDD(VDD),.Y(I11037),.A(g6629));
  NOT NOT1_3320(.VSS(VSS),.VDD(VDD),.Y(g8353),.A(I13439));
  NOT NOT1_3321(.VSS(VSS),.VDD(VDD),.Y(I14130),.A(g8769));
  NOT NOT1_3322(.VSS(VSS),.VDD(VDD),.Y(I10362),.A(g6224));
  NOT NOT1_3323(.VSS(VSS),.VDD(VDD),.Y(g2864),.A(g2298));
  NOT NOT1_3324(.VSS(VSS),.VDD(VDD),.Y(I10165),.A(g5948));
  NOT NOT1_3325(.VSS(VSS),.VDD(VDD),.Y(I13782),.A(g8515));
  NOT NOT1_3326(.VSS(VSS),.VDD(VDD),.Y(g6917),.A(I11029));
  NOT NOT1_3327(.VSS(VSS),.VDD(VDD),.Y(g4894),.A(I8247));
  NOT NOT1_3328(.VSS(VSS),.VDD(VDD),.Y(I6028),.A(g2208));
  NOT NOT1_3329(.VSS(VSS),.VDD(VDD),.Y(g10269),.A(g10154));
  NOT NOT1_3330(.VSS(VSS),.VDD(VDD),.Y(g8802),.A(I14127));
  NOT NOT1_3331(.VSS(VSS),.VDD(VDD),.Y(I6671),.A(g2757));
  NOT NOT1_3332(.VSS(VSS),.VDD(VDD),.Y(I6428),.A(g2348));
  NOT NOT1_3333(.VSS(VSS),.VDD(VDD),.Y(g7886),.A(g7479));
  NOT NOT1_3334(.VSS(VSS),.VDD(VDD),.Y(g4735),.A(g3546));
  NOT NOT1_3335(.VSS(VSS),.VDD(VDD),.Y(I17327),.A(g11349));
  NOT NOT1_3336(.VSS(VSS),.VDD(VDD),.Y(g6265),.A(I10054));
  NOT NOT1_3337(.VSS(VSS),.VDD(VDD),.Y(g3976),.A(I7109));
  NOT NOT1_3338(.VSS(VSS),.VDD(VDD),.Y(I6247),.A(g2462));
  NOT NOT1_3339(.VSS(VSS),.VDD(VDD),.Y(g4782),.A(g4089));
  NOT NOT1_3340(.VSS(VSS),.VDD(VDD),.Y(I11155),.A(g6470));
  NOT NOT1_3341(.VSS(VSS),.VDD(VDD),.Y(g10156),.A(I15464));
  NOT NOT1_3342(.VSS(VSS),.VDD(VDD),.Y(I15708),.A(g10241));
  NOT NOT1_3343(.VSS(VSS),.VDD(VDD),.Y(I17537),.A(g11497));
  NOT NOT1_3344(.VSS(VSS),.VDD(VDD),.Y(I13418),.A(g8145));
  NOT NOT1_3345(.VSS(VSS),.VDD(VDD),.Y(I13822),.A(g8488));
  NOT NOT1_3346(.VSS(VSS),.VDD(VDD),.Y(g5697),.A(I9232));
  NOT NOT1_3347(.VSS(VSS),.VDD(VDD),.Y(I10006),.A(g5633));
  NOT NOT1_3348(.VSS(VSS),.VDD(VDD),.Y(g6442),.A(I10362));
  NOT NOT1_3349(.VSS(VSS),.VDD(VDD),.Y(g9452),.A(I14645));
  NOT NOT1_3350(.VSS(VSS),.VDD(VDD),.Y(g7314),.A(I11590));
  NOT NOT1_3351(.VSS(VSS),.VDD(VDD),.Y(g5210),.A(I8631));
  NOT NOT1_3352(.VSS(VSS),.VDD(VDD),.Y(I17108),.A(g11225));
  NOT NOT1_3353(.VSS(VSS),.VDD(VDD),.Y(g11471),.A(I17450));
  NOT NOT1_3354(.VSS(VSS),.VDD(VDD),.Y(I7345),.A(g4050));
  NOT NOT1_3355(.VSS(VSS),.VDD(VDD),.Y(I16458),.A(g10734));
  NOT NOT1_3356(.VSS(VSS),.VDD(VDD),.Y(I8429),.A(g4458));
  NOT NOT1_3357(.VSS(VSS),.VDD(VDD),.Y(I9605),.A(g5620));
  NOT NOT1_3358(.VSS(VSS),.VDD(VDD),.Y(g4475),.A(I7852));
  NOT NOT1_3359(.VSS(VSS),.VDD(VDD),.Y(g5596),.A(I9020));
  NOT NOT1_3360(.VSS(VSS),.VDD(VDD),.Y(g6164),.A(g5426));
  NOT NOT1_3361(.VSS(VSS),.VDD(VDD),.Y(I7763),.A(g3769));
  NOT NOT1_3362(.VSS(VSS),.VDD(VDD),.Y(I7191),.A(g2646));
  NOT NOT1_3363(.VSS(VSS),.VDD(VDD),.Y(g10734),.A(I16413));
  NOT NOT1_3364(.VSS(VSS),.VDD(VDD),.Y(I10437),.A(g5755));
  NOT NOT1_3365(.VSS(VSS),.VDD(VDD),.Y(g10335),.A(I15787));
  NOT NOT1_3366(.VSS(VSS),.VDD(VDD),.Y(g7650),.A(I12261));
  NOT NOT1_3367(.VSS(VSS),.VDD(VDD),.Y(g3326),.A(I6495));
  NOT NOT1_3368(.VSS(VSS),.VDD(VDD),.Y(I15244),.A(g10031));
  NOT NOT1_3369(.VSS(VSS),.VDD(VDD),.Y(g4292),.A(g3863));
  NOT NOT1_3370(.VSS(VSS),.VDD(VDD),.Y(g10930),.A(g10827));
  NOT NOT1_3371(.VSS(VSS),.VDD(VDD),.Y(g11043),.A(I16790));
  NOT NOT1_3372(.VSS(VSS),.VDD(VDD),.Y(g6454),.A(I10388));
  NOT NOT1_3373(.VSS(VSS),.VDD(VDD),.Y(g11244),.A(g11112));
  NOT NOT1_3374(.VSS(VSS),.VDD(VDD),.Y(g4526),.A(I7931));
  NOT NOT1_3375(.VSS(VSS),.VDD(VDD),.Y(I5478),.A(g1212));
  NOT NOT1_3376(.VSS(VSS),.VDD(VDD),.Y(g6296),.A(I10147));
  NOT NOT1_3377(.VSS(VSS),.VDD(VDD),.Y(I11194),.A(g6515));
  NOT NOT1_3378(.VSS(VSS),.VDD(VDD),.Y(g3760),.A(g3003));
  NOT NOT1_3379(.VSS(VSS),.VDD(VDD),.Y(g7008),.A(I11149));
  NOT NOT1_3380(.VSS(VSS),.VDD(VDD),.Y(I13194),.A(g8140));
  NOT NOT1_3381(.VSS(VSS),.VDD(VDD),.Y(I13589),.A(g8361));
  NOT NOT1_3382(.VSS(VSS),.VDD(VDD),.Y(g2623),.A(g1999));
  NOT NOT1_3383(.VSS(VSS),.VDD(VDD),.Y(I17381),.A(g11436));
  NOT NOT1_3384(.VSS(VSS),.VDD(VDD),.Y(I7536),.A(g4098));
  NOT NOT1_3385(.VSS(VSS),.VDD(VDD),.Y(I9585),.A(g5241));
  NOT NOT1_3386(.VSS(VSS),.VDD(VDD),.Y(g2076),.A(I4886));
  NOT NOT1_3387(.VSS(VSS),.VDD(VDD),.Y(g10131),.A(I15395));
  NOT NOT1_3388(.VSS(VSS),.VDD(VDD),.Y(g2889),.A(I6049));
  NOT NOT1_3389(.VSS(VSS),.VDD(VDD),.Y(I11524),.A(g6593));
  NOT NOT1_3390(.VSS(VSS),.VDD(VDD),.Y(I16598),.A(g10804));
  NOT NOT1_3391(.VSS(VSS),.VDD(VDD),.Y(g11069),.A(g10974));
  NOT NOT1_3392(.VSS(VSS),.VDD(VDD),.Y(g4084),.A(g3119));
  NOT NOT1_3393(.VSS(VSS),.VDD(VDD),.Y(I11836),.A(g7220));
  NOT NOT1_3394(.VSS(VSS),.VDD(VDD),.Y(I5435),.A(g18));
  NOT NOT1_3395(.VSS(VSS),.VDD(VDD),.Y(g4603),.A(g3829));
  NOT NOT1_3396(.VSS(VSS),.VDD(VDD),.Y(g5936),.A(I9564));
  NOT NOT1_3397(.VSS(VSS),.VDD(VDD),.Y(g7336),.A(I11656));
  NOT NOT1_3398(.VSS(VSS),.VDD(VDD),.Y(g8600),.A(g8475));
  NOT NOT1_3399(.VSS(VSS),.VDD(VDD),.Y(I15068),.A(g9710));
  NOT NOT1_3400(.VSS(VSS),.VDD(VDD),.Y(g7768),.A(I12469));
  NOT NOT1_3401(.VSS(VSS),.VDD(VDD),.Y(g4439),.A(I7793));
  NOT NOT1_3402(.VSS(VSS),.VDD(VDD),.Y(g11657),.A(I17773));
  NOT NOT1_3403(.VSS(VSS),.VDD(VDD),.Y(g5117),.A(g4682));
  NOT NOT1_3404(.VSS(VSS),.VDD(VDD),.Y(g6553),.A(I10477));
  NOT NOT1_3405(.VSS(VSS),.VDD(VDD),.Y(g8714),.A(I14005));
  NOT NOT1_3406(.VSS(VSS),.VDD(VDD),.Y(g11068),.A(g10974));
  NOT NOT1_3407(.VSS(VSS),.VDD(VDD),.Y(I7858),.A(g3631));
  NOT NOT1_3408(.VSS(VSS),.VDD(VDD),.Y(I11477),.A(g6488));
  NOT NOT1_3409(.VSS(VSS),.VDD(VDD),.Y(g7594),.A(I12120));
  NOT NOT1_3410(.VSS(VSS),.VDD(VDD),.Y(g10487),.A(I16098));
  NOT NOT1_3411(.VSS(VSS),.VDD(VDD),.Y(g7972),.A(I12770));
  NOT NOT1_3412(.VSS(VSS),.VDD(VDD),.Y(g2175),.A(g44));
  NOT NOT1_3413(.VSS(VSS),.VDD(VDD),.Y(I11119),.A(g6461));
  NOT NOT1_3414(.VSS(VSS),.VDD(VDD),.Y(g9025),.A(I14412));
  NOT NOT1_3415(.VSS(VSS),.VDD(VDD),.Y(g2871),.A(I6013));
  NOT NOT1_3416(.VSS(VSS),.VDD(VDD),.Y(g10619),.A(I16292));
  NOT NOT1_3417(.VSS(VSS),.VDD(VDD),.Y(I12759),.A(g7702));
  NOT NOT1_3418(.VSS(VSS),.VDD(VDD),.Y(I7757),.A(g3767));
  NOT NOT1_3419(.VSS(VSS),.VDD(VDD),.Y(I16817),.A(g10912));
  NOT NOT1_3420(.VSS(VSS),.VDD(VDD),.Y(I9673),.A(g5182));
  NOT NOT1_3421(.VSS(VSS),.VDD(VDD),.Y(I14236),.A(g8802));
  NOT NOT1_3422(.VSS(VSS),.VDD(VDD),.Y(g7806),.A(I12583));
  NOT NOT1_3423(.VSS(VSS),.VDD(VDD),.Y(I10952),.A(g6556));
  NOT NOT1_3424(.VSS(VSS),.VDD(VDD),.Y(g3220),.A(I6398));
  NOT NOT1_3425(.VSS(VSS),.VDD(VDD),.Y(I8109),.A(g3622));
  NOT NOT1_3426(.VSS(VSS),.VDD(VDD),.Y(g2651),.A(g2007));
  NOT NOT1_3427(.VSS(VSS),.VDD(VDD),.Y(I6217),.A(g2302));
  NOT NOT1_3428(.VSS(VSS),.VDD(VDD),.Y(g4583),.A(g3880));
  NOT NOT1_3429(.VSS(VSS),.VDD(VDD),.Y(g6412),.A(I10322));
  NOT NOT1_3430(.VSS(VSS),.VDD(VDD),.Y(I17390),.A(g11430));
  NOT NOT1_3431(.VSS(VSS),.VDD(VDD),.Y(g10279),.A(g10158));
  NOT NOT1_3432(.VSS(VSS),.VDD(VDD),.Y(g7065),.A(I11272));
  NOT NOT1_3433(.VSS(VSS),.VDD(VDD),.Y(I7315),.A(g2891));
  NOT NOT1_3434(.VSS(VSS),.VDD(VDD),.Y(g6389),.A(I10289));
  NOT NOT1_3435(.VSS(VSS),.VDD(VDD),.Y(I7642),.A(g3440));
  NOT NOT1_3436(.VSS(VSS),.VDD(VDD),.Y(I9168),.A(g5040));
  NOT NOT1_3437(.VSS(VSS),.VDD(VDD),.Y(g6706),.A(I10685));
  NOT NOT1_3438(.VSS(VSS),.VDD(VDD),.Y(I9669),.A(g5426));
  NOT NOT1_3439(.VSS(VSS),.VDD(VDD),.Y(g7887),.A(g7693));
  NOT NOT1_3440(.VSS(VSS),.VDD(VDD),.Y(g7122),.A(I11357));
  NOT NOT1_3441(.VSS(VSS),.VDD(VDD),.Y(I15792),.A(g10279));
  NOT NOT1_3442(.VSS(VSS),.VDD(VDD),.Y(I9368),.A(g5288));
  NOT NOT1_3443(.VSS(VSS),.VDD(VDD),.Y(g7322),.A(I11614));
  NOT NOT1_3444(.VSS(VSS),.VDD(VDD),.Y(g4919),.A(I8290));
  NOT NOT1_3445(.VSS(VSS),.VDD(VDD),.Y(I10063),.A(g5766));
  NOT NOT1_3446(.VSS(VSS),.VDD(VDD),.Y(g6990),.A(I11132));
  NOT NOT1_3447(.VSS(VSS),.VDD(VDD),.Y(I7447),.A(g3694));
  NOT NOT1_3448(.VSS(VSS),.VDD(VDD),.Y(g10278),.A(g10182));
  NOT NOT1_3449(.VSS(VSS),.VDD(VDD),.Y(g3977),.A(I7112));
  NOT NOT1_3450(.VSS(VSS),.VDD(VDD),.Y(I6861),.A(g2942));
  NOT NOT1_3451(.VSS(VSS),.VDD(VDD),.Y(g6888),.A(I10984));
  NOT NOT1_3452(.VSS(VSS),.VDD(VDD),.Y(I16656),.A(g10791));
  NOT NOT1_3453(.VSS(VSS),.VDD(VDD),.Y(I9531),.A(g5004));
  NOT NOT1_3454(.VSS(VSS),.VDD(VDD),.Y(g6171),.A(g5446));
  NOT NOT1_3455(.VSS(VSS),.VDD(VDD),.Y(g2184),.A(g1806));
  NOT NOT1_3456(.VSS(VSS),.VDD(VDD),.Y(I16295),.A(g10552));
  NOT NOT1_3457(.VSS(VSS),.VDD(VDD),.Y(I9458),.A(g5091));
  NOT NOT1_3458(.VSS(VSS),.VDD(VDD),.Y(g3161),.A(I6367));
  NOT NOT1_3459(.VSS(VSS),.VDD(VDD),.Y(I11704),.A(g7008));
  NOT NOT1_3460(.VSS(VSS),.VDD(VDD),.Y(I12849),.A(g7632));
  NOT NOT1_3461(.VSS(VSS),.VDD(VDD),.Y(I6055),.A(g2569));
  NOT NOT1_3462(.VSS(VSS),.VDD(VDD),.Y(I17522),.A(g11485));
  NOT NOT1_3463(.VSS(VSS),.VDD(VDD),.Y(g2339),.A(I5399));
  NOT NOT1_3464(.VSS(VSS),.VDD(VDD),.Y(g7033),.A(I11188));
  NOT NOT1_3465(.VSS(VSS),.VDD(VDD),.Y(g10039),.A(I15244));
  NOT NOT1_3466(.VSS(VSS),.VDD(VDD),.Y(I10873),.A(g6331));
  NOT NOT1_3467(.VSS(VSS),.VDD(VDD),.Y(g6956),.A(I11106));
  NOT NOT1_3468(.VSS(VSS),.VDD(VDD),.Y(g5597),.A(I9023));
  NOT NOT1_3469(.VSS(VSS),.VDD(VDD),.Y(I14873),.A(g9525));
  NOT NOT1_3470(.VSS(VSS),.VDD(VDD),.Y(I7654),.A(g3728));
  NOT NOT1_3471(.VSS(VSS),.VDD(VDD),.Y(I13809),.A(g8480));
  NOT NOT1_3472(.VSS(VSS),.VDD(VDD),.Y(I6133),.A(g2253));
  NOT NOT1_3473(.VSS(VSS),.VDD(VDD),.Y(g3051),.A(g2135));
  NOT NOT1_3474(.VSS(VSS),.VDD(VDD),.Y(g2838),.A(g2165));
  NOT NOT1_3475(.VSS(VSS),.VDD(VDD),.Y(g8076),.A(I12930));
  NOT NOT1_3476(.VSS(VSS),.VDD(VDD),.Y(g2024),.A(g1718));
  NOT NOT1_3477(.VSS(VSS),.VDD(VDD),.Y(I15458),.A(g10069));
  NOT NOT1_3478(.VSS(VSS),.VDD(VDD),.Y(I13466),.A(g8160));
  NOT NOT1_3479(.VSS(VSS),.VDD(VDD),.Y(I9505),.A(g5088));
  NOT NOT1_3480(.VSS(VSS),.VDD(VDD),.Y(g6281),.A(I10102));
  NOT NOT1_3481(.VSS(VSS),.VDD(VDD),.Y(g8476),.A(I13674));
  NOT NOT1_3482(.VSS(VSS),.VDD(VDD),.Y(g3327),.A(I6498));
  NOT NOT1_3483(.VSS(VSS),.VDD(VDD),.Y(g2424),.A(g1690));
  NOT NOT1_3484(.VSS(VSS),.VDD(VDD),.Y(I8449),.A(g4469));
  NOT NOT1_3485(.VSS(VSS),.VDD(VDD),.Y(I12652),.A(g7458));
  NOT NOT1_3486(.VSS(VSS),.VDD(VDD),.Y(g9766),.A(g9432));
  NOT NOT1_3487(.VSS(VSS),.VDD(VDD),.Y(g2809),.A(I5909));
  NOT NOT1_3488(.VSS(VSS),.VDD(VDD),.Y(g5784),.A(I9380));
  NOT NOT1_3489(.VSS(VSS),.VDD(VDD),.Y(g4004),.A(I7140));
  NOT NOT1_3490(.VSS(VSS),.VDD(VDD),.Y(I9734),.A(g5257));
  NOT NOT1_3491(.VSS(VSS),.VDD(VDD),.Y(I13036),.A(g8053));
  NOT NOT1_3492(.VSS(VSS),.VDD(VDD),.Y(I5002),.A(g1173));
  NOT NOT1_3493(.VSS(VSS),.VDD(VDD),.Y(I8865),.A(g4518));
  NOT NOT1_3494(.VSS(VSS),.VDD(VDD),.Y(g7550),.A(g6974));
  NOT NOT1_3495(.VSS(VSS),.VDD(VDD),.Y(g6297),.A(I10150));
  NOT NOT1_3496(.VSS(VSS),.VDD(VDD),.Y(I11560),.A(g7037));
  NOT NOT1_3497(.VSS(VSS),.VDD(VDD),.Y(g10187),.A(I15539));
  NOT NOT1_3498(.VSS(VSS),.VDD(VDD),.Y(I6196),.A(g2462));
  NOT NOT1_3499(.VSS(VSS),.VDD(VDD),.Y(I5824),.A(g2502));
  NOT NOT1_3500(.VSS(VSS),.VDD(VDD),.Y(g7845),.A(I12634));
  NOT NOT1_3501(.VSS(VSS),.VDD(VDD),.Y(I10834),.A(g6715));
  NOT NOT1_3502(.VSS(VSS),.VDD(VDD),.Y(g8871),.A(I14185));
  NOT NOT1_3503(.VSS(VSS),.VDD(VDD),.Y(g8375),.A(I13475));
  NOT NOT1_3504(.VSS(VSS),.VDD(VDD),.Y(I15545),.A(g10075));
  NOT NOT1_3505(.VSS(VSS),.VDD(VDD),.Y(g3633),.A(I6802));
  NOT NOT1_3506(.VSS(VSS),.VDD(VDD),.Y(I15079),.A(g9745));
  NOT NOT1_3507(.VSS(VSS),.VDD(VDD),.Y(I8098),.A(g3583));
  NOT NOT1_3508(.VSS(VSS),.VDD(VDD),.Y(g2077),.A(g219));
  NOT NOT1_3509(.VSS(VSS),.VDD(VDD),.Y(g2231),.A(I5218));
  NOT NOT1_3510(.VSS(VSS),.VDD(VDD),.Y(g7195),.A(I11417));
  NOT NOT1_3511(.VSS(VSS),.VDD(VDD),.Y(g11545),.A(g11519));
  NOT NOT1_3512(.VSS(VSS),.VDD(VDD),.Y(g11079),.A(I16850));
  NOT NOT1_3513(.VSS(VSS),.VDD(VDD),.Y(g11444),.A(I17381));
  NOT NOT1_3514(.VSS(VSS),.VDD(VDD),.Y(g5937),.A(I9567));
  NOT NOT1_3515(.VSS(VSS),.VDD(VDD),.Y(g7395),.A(g6941));
  NOT NOT1_3516(.VSS(VSS),.VDD(VDD),.Y(I13642),.A(g8378));
  NOT NOT1_3517(.VSS(VSS),.VDD(VDD),.Y(g7337),.A(I11659));
  NOT NOT1_3518(.VSS(VSS),.VDD(VDD),.Y(g3103),.A(g2391));
  NOT NOT1_3519(.VSS(VSS),.VDD(VDD),.Y(I9074),.A(g4764));
  NOT NOT1_3520(.VSS(VSS),.VDD(VDD),.Y(g7913),.A(g7467));
  NOT NOT1_3521(.VSS(VSS),.VDD(VDD),.Y(I6538),.A(g2827));
  NOT NOT1_3522(.VSS(VSS),.VDD(VDD),.Y(g2523),.A(I5632));
  NOT NOT1_3523(.VSS(VSS),.VDD(VDD),.Y(I7272),.A(g3253));
  NOT NOT1_3524(.VSS(VSS),.VDD(VDD),.Y(g2643),.A(g1989));
  NOT NOT1_3525(.VSS(VSS),.VDD(VDD),.Y(I9992),.A(g5633));
  NOT NOT1_3526(.VSS(VSS),.VDD(VDD),.Y(g10143),.A(I15427));
  NOT NOT1_3527(.VSS(VSS),.VDD(VDD),.Y(g5668),.A(I9165));
  NOT NOT1_3528(.VSS(VSS),.VDD(VDD),.Y(g11078),.A(I16847));
  NOT NOT1_3529(.VSS(VSS),.VDD(VDD),.Y(g6338),.A(I10237));
  NOT NOT1_3530(.VSS(VSS),.VDD(VDD),.Y(I15598),.A(g10170));
  NOT NOT1_3531(.VSS(VSS),.VDD(VDD),.Y(I10021),.A(g5692));
  NOT NOT1_3532(.VSS(VSS),.VDD(VDD),.Y(g5840),.A(g5320));
  NOT NOT1_3533(.VSS(VSS),.VDD(VDD),.Y(g4970),.A(g4411));
  NOT NOT1_3534(.VSS(VSS),.VDD(VDD),.Y(g8500),.A(I13695));
  NOT NOT1_3535(.VSS(VSS),.VDD(VDD),.Y(I7612),.A(g3817));
  NOT NOT1_3536(.VSS(VSS),.VDD(VDD),.Y(g11598),.A(I17642));
  NOT NOT1_3537(.VSS(VSS),.VDD(VDD),.Y(I7017),.A(g3068));
  NOT NOT1_3538(.VSS(VSS),.VDD(VDD),.Y(g6109),.A(g5052));
  NOT NOT1_3539(.VSS(VSS),.VDD(VDD),.Y(I12406),.A(g7464));
  NOT NOT1_3540(.VSS(VSS),.VDD(VDD),.Y(g6309),.A(I10186));
  NOT NOT1_3541(.VSS(VSS),.VDD(VDD),.Y(g11086),.A(I16867));
  NOT NOT1_3542(.VSS(VSS),.VDD(VDD),.Y(g7807),.A(I12586));
  NOT NOT1_3543(.VSS(VSS),.VDD(VDD),.Y(I7417),.A(g4160));
  NOT NOT1_3544(.VSS(VSS),.VDD(VDD),.Y(g3732),.A(I6914));
  NOT NOT1_3545(.VSS(VSS),.VDD(VDD),.Y(I17252),.A(g11343));
  NOT NOT1_3546(.VSS(VSS),.VDD(VDD),.Y(g10169),.A(I15503));
  NOT NOT1_3547(.VSS(VSS),.VDD(VDD),.Y(I7935),.A(g3440));
  NOT NOT1_3548(.VSS(VSS),.VDD(VDD),.Y(I9080),.A(g4775));
  NOT NOT1_3549(.VSS(VSS),.VDD(VDD),.Y(g8184),.A(I13105));
  NOT NOT1_3550(.VSS(VSS),.VDD(VDD),.Y(g10884),.A(g10809));
  NOT NOT1_3551(.VSS(VSS),.VDD(VDD),.Y(g6808),.A(I10834));
  NOT NOT1_3552(.VSS(VSS),.VDD(VDD),.Y(I15817),.A(g10199));
  NOT NOT1_3553(.VSS(VSS),.VDD(VDD),.Y(I9863),.A(g5557));
  NOT NOT1_3554(.VSS(VSS),.VDD(VDD),.Y(g8139),.A(g8025));
  NOT NOT1_3555(.VSS(VSS),.VDD(VDD),.Y(I16289),.A(g10541));
  NOT NOT1_3556(.VSS(VSS),.VDD(VDD),.Y(g8339),.A(I13397));
  NOT NOT1_3557(.VSS(VSS),.VDD(VDD),.Y(g2742),.A(I5798));
  NOT NOT1_3558(.VSS(VSS),.VDD(VDD),.Y(g3944),.A(g2920));
  NOT NOT1_3559(.VSS(VSS),.VDD(VDD),.Y(g10168),.A(I15500));
  NOT NOT1_3560(.VSS(VSS),.VDD(VDD),.Y(I10607),.A(g5763));
  NOT NOT1_3561(.VSS(VSS),.VDD(VDD),.Y(g6707),.A(g5949));
  NOT NOT1_3562(.VSS(VSS),.VDD(VDD),.Y(I13630),.A(g8334));
  NOT NOT1_3563(.VSS(VSS),.VDD(VDD),.Y(g2304),.A(I5348));
  NOT NOT1_3564(.VSS(VSS),.VDD(VDD),.Y(g11322),.A(I17121));
  NOT NOT1_3565(.VSS(VSS),.VDD(VDD),.Y(g9091),.A(g8892));
  NOT NOT1_3566(.VSS(VSS),.VDD(VDD),.Y(g4320),.A(g4013));
  NOT NOT1_3567(.VSS(VSS),.VDD(VDD),.Y(I15977),.A(g10411));
  NOT NOT1_3568(.VSS(VSS),.VDD(VDD),.Y(g11159),.A(g10950));
  NOT NOT1_3569(.VSS(VSS),.VDD(VDD),.Y(I10274),.A(g5811));
  NOT NOT1_3570(.VSS(VSS),.VDD(VDD),.Y(I11166),.A(g6480));
  NOT NOT1_3571(.VSS(VSS),.VDD(VDD),.Y(I11665),.A(g7038));
  NOT NOT1_3572(.VSS(VSS),.VDD(VDD),.Y(I16571),.A(g10819));
  NOT NOT1_3573(.VSS(VSS),.VDD(VDD),.Y(I13166),.A(g8009));
  NOT NOT1_3574(.VSS(VSS),.VDD(VDD),.Y(I7330),.A(g3761));
  NOT NOT1_3575(.VSS(VSS),.VDD(VDD),.Y(I8268),.A(g4674));
  NOT NOT1_3576(.VSS(VSS),.VDD(VDD),.Y(g8424),.A(I13586));
  NOT NOT1_3577(.VSS(VSS),.VDD(VDD),.Y(I5064),.A(g1690));
  NOT NOT1_3578(.VSS(VSS),.VDD(VDD),.Y(g8795),.A(I14112));
  NOT NOT1_3579(.VSS(VSS),.VDD(VDD),.Y(g10217),.A(I15589));
  NOT NOT1_3580(.VSS(VSS),.VDD(VDD),.Y(g7142),.A(I11383));
  NOT NOT1_3581(.VSS(VSS),.VDD(VDD),.Y(I6256),.A(g2462));
  NOT NOT1_3582(.VSS(VSS),.VDD(VDD),.Y(g4277),.A(g3688));
  NOT NOT1_3583(.VSS(VSS),.VDD(VDD),.Y(g6201),.A(I9938));
  NOT NOT1_3584(.VSS(VSS),.VDD(VDD),.Y(g7342),.A(I11674));
  NOT NOT1_3585(.VSS(VSS),.VDD(VDD),.Y(I11008),.A(g6795));
  NOT NOT1_3586(.VSS(VSS),.VDD(VDD),.Y(g6957),.A(I11109));
  NOT NOT1_3587(.VSS(VSS),.VDD(VDD),.Y(I15353),.A(g10007));
  NOT NOT1_3588(.VSS(VSS),.VDD(VDD),.Y(g2754),.A(I5830));
  NOT NOT1_3589(.VSS(VSS),.VDD(VDD),.Y(g4906),.A(I8275));
  NOT NOT1_3590(.VSS(VSS),.VDD(VDD),.Y(g7815),.A(I12610));
  NOT NOT1_3591(.VSS(VSS),.VDD(VDD),.Y(g11656),.A(I17770));
  NOT NOT1_3592(.VSS(VSS),.VDD(VDD),.Y(g4789),.A(g3337));
  NOT NOT1_3593(.VSS(VSS),.VDD(VDD),.Y(I7800),.A(g3791));
  NOT NOT1_3594(.VSS(VSS),.VDD(VDD),.Y(g10486),.A(I16095));
  NOT NOT1_3595(.VSS(VSS),.VDD(VDD),.Y(g11353),.A(I17176));
  NOT NOT1_3596(.VSS(VSS),.VDD(VDD),.Y(g8077),.A(I12933));
  NOT NOT1_3597(.VSS(VSS),.VDD(VDD),.Y(I15823),.A(g10201));
  NOT NOT1_3598(.VSS(VSS),.VDD(VDD),.Y(g6449),.A(g6172));
  NOT NOT1_3599(.VSS(VSS),.VDD(VDD),.Y(I13485),.A(g8194));
  NOT NOT1_3600(.VSS(VSS),.VDD(VDD),.Y(g2273),.A(g881));
  NOT NOT1_3601(.VSS(VSS),.VDD(VDD),.Y(g8477),.A(g8317));
  NOT NOT1_3602(.VSS(VSS),.VDD(VDD),.Y(g6575),.A(g5949));
  NOT NOT1_3603(.VSS(VSS),.VDD(VDD),.Y(g7692),.A(g7148));
  NOT NOT1_3604(.VSS(VSS),.VDD(VDD),.Y(I12613),.A(g7525));
  NOT NOT1_3605(.VSS(VSS),.VDD(VDD),.Y(g8523),.A(I13732));
  NOT NOT1_3606(.VSS(VSS),.VDD(VDD),.Y(I6381),.A(g2257));
  NOT NOT1_3607(.VSS(VSS),.VDD(VDD),.Y(g9767),.A(I14914));
  NOT NOT1_3608(.VSS(VSS),.VDD(VDD),.Y(g7097),.A(I11330));
  NOT NOT1_3609(.VSS(VSS),.VDD(VDD),.Y(I9688),.A(g5201));
  NOT NOT1_3610(.VSS(VSS),.VDD(VDD),.Y(g7726),.A(I12363));
  NOT NOT1_3611(.VSS(VSS),.VDD(VDD),.Y(I9857),.A(g5269));
  NOT NOT1_3612(.VSS(VSS),.VDD(VDD),.Y(I13454),.A(g8183));
  NOT NOT1_3613(.VSS(VSS),.VDD(VDD),.Y(g2613),.A(I5740));
  NOT NOT1_3614(.VSS(VSS),.VDD(VDD),.Y(g7497),.A(g7148));
  NOT NOT1_3615(.VSS(VSS),.VDD(VDD),.Y(g9535),.A(I14690));
  NOT NOT1_3616(.VSS(VSS),.VDD(VDD),.Y(g6715),.A(I10702));
  NOT NOT1_3617(.VSS(VSS),.VDD(VDD),.Y(g2044),.A(I4850));
  NOT NOT1_3618(.VSS(VSS),.VDD(VDD),.Y(g7354),.A(I11710));
  NOT NOT1_3619(.VSS(VSS),.VDD(VDD),.Y(g10580),.A(g10530));
  NOT NOT1_3620(.VSS(VSS),.VDD(VDD),.Y(I10153),.A(g5947));
  NOT NOT1_3621(.VSS(VSS),.VDD(VDD),.Y(g2444),.A(g876));
  NOT NOT1_3622(.VSS(VSS),.VDD(VDD),.Y(I5237),.A(g1107));
  NOT NOT1_3623(.VSS(VSS),.VDD(VDD),.Y(g5032),.A(I8403));
  NOT NOT1_3624(.VSS(VSS),.VDD(VDD),.Y(g2269),.A(I5308));
  NOT NOT1_3625(.VSS(VSS),.VDD(VDD),.Y(g10223),.A(I15595));
  NOT NOT1_3626(.VSS(VSS),.VDD(VDD),.Y(I7213),.A(g2635));
  NOT NOT1_3627(.VSS(VSS),.VDD(VDD),.Y(g9261),.A(g8892));
  NOT NOT1_3628(.VSS(VSS),.VDD(VDD),.Y(I6421),.A(g2346));
  NOT NOT1_3629(.VSS(VSS),.VDD(VDD),.Y(g4299),.A(g4144));
  NOT NOT1_3630(.VSS(VSS),.VDD(VDD),.Y(I14409),.A(g8938));
  NOT NOT1_3631(.VSS(VSS),.VDD(VDD),.Y(I12463),.A(g7579));
  NOT NOT1_3632(.VSS(VSS),.VDD(VDD),.Y(g3697),.A(I6856));
  NOT NOT1_3633(.VSS(VSS),.VDD(VDD),.Y(g8099),.A(g7990));
  NOT NOT1_3634(.VSS(VSS),.VDD(VDD),.Y(I8385),.A(g4238));
  NOT NOT1_3635(.VSS(VSS),.VDD(VDD),.Y(I14136),.A(g8775));
  NOT NOT1_3636(.VSS(VSS),.VDD(VDD),.Y(g8304),.A(I13280));
  NOT NOT1_3637(.VSS(VSS),.VDD(VDD),.Y(g3914),.A(g3015));
  NOT NOT1_3638(.VSS(VSS),.VDD(VDD),.Y(I9126),.A(g4891));
  NOT NOT1_3639(.VSS(VSS),.VDD(VDD),.Y(I13239),.A(g8266));
  NOT NOT1_3640(.VSS(VSS),.VDD(VDD),.Y(g10110),.A(I15344));
  NOT NOT1_3641(.VSS(VSS),.VDD(VDD),.Y(g11631),.A(I17707));
  NOT NOT1_3642(.VSS(VSS),.VDD(VDD),.Y(I9326),.A(g5320));
  NOT NOT1_3643(.VSS(VSS),.VDD(VDD),.Y(g2543),.A(I5662));
  NOT NOT1_3644(.VSS(VSS),.VDD(VDD),.Y(g6584),.A(I10538));
  NOT NOT1_3645(.VSS(VSS),.VDD(VDD),.Y(g11017),.A(I16742));
  NOT NOT1_3646(.VSS(VSS),.VDD(VDD),.Y(g6539),.A(I10461));
  NOT NOT1_3647(.VSS(VSS),.VDD(VDD),.Y(g6896),.A(I10996));
  NOT NOT1_3648(.VSS(VSS),.VDD(VDD),.Y(g5568),.A(I8985));
  NOT NOT1_3649(.VSS(VSS),.VDD(VDD),.Y(g10321),.A(I15759));
  NOT NOT1_3650(.VSS(VSS),.VDD(VDD),.Y(I5089),.A(g1854));
  NOT NOT1_3651(.VSS(VSS),.VDD(VDD),.Y(I5731),.A(g2089));
  NOT NOT1_3652(.VSS(VSS),.VDD(VDD),.Y(I11238),.A(g6543));
  NOT NOT1_3653(.VSS(VSS),.VDD(VDD),.Y(I17213),.A(g11290));
  NOT NOT1_3654(.VSS(VSS),.VDD(VDD),.Y(g7783),.A(I12514));
  NOT NOT1_3655(.VSS(VSS),.VDD(VDD),.Y(g10179),.A(g10041));
  NOT NOT1_3656(.VSS(VSS),.VDD(VDD),.Y(g10531),.A(g10471));
  NOT NOT1_3657(.VSS(VSS),.VDD(VDD),.Y(g7979),.A(I12783));
  NOT NOT1_3658(.VSS(VSS),.VDD(VDD),.Y(g3413),.A(g2896));
  NOT NOT1_3659(.VSS(VSS),.VDD(VDD),.Y(g5912),.A(I9544));
  NOT NOT1_3660(.VSS(VSS),.VDD(VDD),.Y(g7312),.A(I11584));
  NOT NOT1_3661(.VSS(VSS),.VDD(VDD),.Y(I7166),.A(g2620));
  NOT NOT1_3662(.VSS(VSS),.VDD(VDD),.Y(I5966),.A(g2541));
  NOT NOT1_3663(.VSS(VSS),.VDD(VDD),.Y(g10178),.A(I15526));
  NOT NOT1_3664(.VSS(VSS),.VDD(VDD),.Y(I7366),.A(g4012));
  NOT NOT1_3665(.VSS(VSS),.VDD(VDD),.Y(g4738),.A(g3440));
  NOT NOT1_3666(.VSS(VSS),.VDD(VDD),.Y(I13941),.A(g8488));
  NOT NOT1_3667(.VSS(VSS),.VDD(VDD),.Y(I13382),.A(g8134));
  NOT NOT1_3668(.VSS(VSS),.VDD(VDD),.Y(g6268),.A(I10063));
  NOT NOT1_3669(.VSS(VSS),.VDD(VDD),.Y(I11519),.A(g6591));
  NOT NOT1_3670(.VSS(VSS),.VDD(VDD),.Y(I11176),.A(g6501));
  NOT NOT1_3671(.VSS(VSS),.VDD(VDD),.Y(g10186),.A(I15536));
  NOT NOT1_3672(.VSS(VSS),.VDD(VDD),.Y(g7001),.A(I11140));
  NOT NOT1_3673(.VSS(VSS),.VDD(VDD),.Y(g8273),.A(I13191));
  NOT NOT1_3674(.VSS(VSS),.VDD(VDD),.Y(g10676),.A(g10570));
  NOT NOT1_3675(.VSS(VSS),.VDD(VDD),.Y(g6419),.A(I10331));
  NOT NOT1_3676(.VSS(VSS),.VDD(VDD),.Y(I10891),.A(g6334));
  NOT NOT1_3677(.VSS(VSS),.VDD(VDD),.Y(I13185),.A(g8192));
  NOT NOT1_3678(.VSS(VSS),.VDD(VDD),.Y(g11289),.A(I17070));
  NOT NOT1_3679(.VSS(VSS),.VDD(VDD),.Y(I7456),.A(g3716));
  NOT NOT1_3680(.VSS(VSS),.VDD(VDD),.Y(g1993),.A(g786));
  NOT NOT1_3681(.VSS(VSS),.VDD(VDD),.Y(g3820),.A(I7048));
  NOT NOT1_3682(.VSS(VSS),.VDD(VDD),.Y(g7676),.A(I12303));
  NOT NOT1_3683(.VSS(VSS),.VDD(VDD),.Y(g4140),.A(I7284));
  NOT NOT1_3684(.VSS(VSS),.VDD(VDD),.Y(g6052),.A(g5426));
  NOT NOT1_3685(.VSS(VSS),.VDD(VDD),.Y(g11309),.A(I17096));
  NOT NOT1_3686(.VSS(VSS),.VDD(VDD),.Y(g4078),.A(I7205));
  NOT NOT1_3687(.VSS(VSS),.VDD(VDD),.Y(I12514),.A(g7735));
  NOT NOT1_3688(.VSS(VSS),.VDD(VDD),.Y(g8613),.A(g8484));
  NOT NOT1_3689(.VSS(VSS),.VDD(VDD),.Y(I16525),.A(g10719));
  NOT NOT1_3690(.VSS(VSS),.VDD(VDD),.Y(I7348),.A(g4056));
  NOT NOT1_3691(.VSS(VSS),.VDD(VDD),.Y(g6452),.A(I10384));
  NOT NOT1_3692(.VSS(VSS),.VDD(VDD),.Y(I9383),.A(g5296));
  NOT NOT1_3693(.VSS(VSS),.VDD(VDD),.Y(I9608),.A(g5127));
  NOT NOT1_3694(.VSS(VSS),.VDD(VDD),.Y(I15308),.A(g10019));
  NOT NOT1_3695(.VSS(VSS),.VDD(VDD),.Y(g7329),.A(I11635));
  NOT NOT1_3696(.VSS(VSS),.VDD(VDD),.Y(g4478),.A(g3820));
  NOT NOT1_3697(.VSS(VSS),.VDD(VDD),.Y(g7761),.A(I12448));
  NOT NOT1_3698(.VSS(VSS),.VDD(VDD),.Y(g2014),.A(g1104));
  NOT NOT1_3699(.VSS(VSS),.VDD(VDD),.Y(g4907),.A(I8278));
  NOT NOT1_3700(.VSS(VSS),.VDD(VDD),.Y(g8444),.A(I13630));
  NOT NOT1_3701(.VSS(VSS),.VDD(VDD),.Y(g2885),.A(I6043));
  NOT NOT1_3702(.VSS(VSS),.VDD(VDD),.Y(I9779),.A(g5391));
  NOT NOT1_3703(.VSS(VSS),.VDD(VDD),.Y(g2946),.A(I6133));
  NOT NOT1_3704(.VSS(VSS),.VDD(VDD),.Y(g4435),.A(g3914));
  NOT NOT1_3705(.VSS(VSS),.VDD(VDD),.Y(I9023),.A(g4727));
  NOT NOT1_3706(.VSS(VSS),.VDD(VDD),.Y(g8983),.A(I14370));
  NOT NOT1_3707(.VSS(VSS),.VDD(VDD),.Y(g4082),.A(I7213));
  NOT NOT1_3708(.VSS(VSS),.VDD(VDD),.Y(I12421),.A(g7634));
  NOT NOT1_3709(.VSS(VSS),.VDD(VDD),.Y(I8406),.A(g4274));
  NOT NOT1_3710(.VSS(VSS),.VDD(VDD),.Y(I5254),.A(g1700));
  NOT NOT1_3711(.VSS(VSS),.VDD(VDD),.Y(I14109),.A(g8765));
  NOT NOT1_3712(.VSS(VSS),.VDD(VDD),.Y(g8572),.A(I13809));
  NOT NOT1_3713(.VSS(VSS),.VDD(VDD),.Y(g7727),.A(I12366));
  NOT NOT1_3714(.VSS(VSS),.VDD(VDD),.Y(I7964),.A(g3433));
  NOT NOT1_3715(.VSS(VSS),.VDD(VDD),.Y(g2903),.A(g2166));
  NOT NOT1_3716(.VSS(VSS),.VDD(VDD),.Y(I7260),.A(g2844));
  NOT NOT1_3717(.VSS(VSS),.VDD(VDD),.Y(I14537),.A(g9308));
  NOT NOT1_3718(.VSS(VSS),.VDD(VDD),.Y(I10108),.A(g5743));
  NOT NOT1_3719(.VSS(VSS),.VDD(VDD),.Y(g6086),.A(I9737));
  NOT NOT1_3720(.VSS(VSS),.VDD(VDD),.Y(g8712),.A(g8680));
  NOT NOT1_3721(.VSS(VSS),.VDD(VDD),.Y(g11495),.A(I17500));
  NOT NOT1_3722(.VSS(VSS),.VDD(VDD),.Y(I12012),.A(g6916));
  NOT NOT1_3723(.VSS(VSS),.VDD(VDD),.Y(I9588),.A(g5114));
  NOT NOT1_3724(.VSS(VSS),.VDD(VDD),.Y(g7746),.A(I12403));
  NOT NOT1_3725(.VSS(VSS),.VDD(VDD),.Y(I8487),.A(g4526));
  NOT NOT1_3726(.VSS(VSS),.VDD(VDD),.Y(I5438),.A(g18));
  NOT NOT1_3727(.VSS(VSS),.VDD(VDD),.Y(g3775),.A(I7002));
  NOT NOT1_3728(.VSS(VSS),.VDD(VDD),.Y(g7221),.A(I11459));
  NOT NOT1_3729(.VSS(VSS),.VDD(VDD),.Y(I17350),.A(g11377));
  NOT NOT1_3730(.VSS(VSS),.VDD(VDD),.Y(I14303),.A(g8811));
  NOT NOT1_3731(.VSS(VSS),.VDD(VDD),.Y(g6385),.A(g6119));
  NOT NOT1_3732(.VSS(VSS),.VDD(VDD),.Y(g6881),.A(I10971));
  NOT NOT1_3733(.VSS(VSS),.VDD(VDD),.Y(I12541),.A(g7662));
  NOT NOT1_3734(.VSS(VSS),.VDD(VDD),.Y(g7703),.A(g7085));
  NOT NOT1_3735(.VSS(VSS),.VDD(VDD),.Y(I9665),.A(g5174));
  NOT NOT1_3736(.VSS(VSS),.VDD(VDD),.Y(I15752),.A(g10264));
  NOT NOT1_3737(.VSS(VSS),.VDD(VDD),.Y(g4915),.A(g4413));
  NOT NOT1_3738(.VSS(VSS),.VDD(VDD),.Y(g2178),.A(g45));
  NOT NOT1_3739(.VSS(VSS),.VDD(VDD),.Y(g2436),.A(I5525));
  NOT NOT1_3740(.VSS(VSS),.VDD(VDD),.Y(I15374),.A(g10007));
  NOT NOT1_3741(.VSS(VSS),.VDD(VDD),.Y(g9028),.A(I14421));
  NOT NOT1_3742(.VSS(VSS),.VDD(VDD),.Y(g8729),.A(g8595));
  NOT NOT1_3743(.VSS(VSS),.VDD(VDD),.Y(g8961),.A(I14330));
  NOT NOT1_3744(.VSS(VSS),.VDD(VDD),.Y(I4900),.A(g583));
  NOT NOT1_3745(.VSS(VSS),.VDD(VDD),.Y(I11501),.A(g6581));
  NOT NOT1_3746(.VSS(VSS),.VDD(VDD),.Y(I16610),.A(g10792));
  NOT NOT1_3747(.VSS(VSS),.VDD(VDD),.Y(g9671),.A(I14802));
  NOT NOT1_3748(.VSS(VSS),.VDD(VDD),.Y(I17152),.A(g11308));
  NOT NOT1_3749(.VSS(VSS),.VDD(VDD),.Y(g3060),.A(g2135));
  NOT NOT1_3750(.VSS(VSS),.VDD(VDD),.Y(I13729),.A(g8290));
  NOT NOT1_3751(.VSS(VSS),.VDD(VDD),.Y(I13577),.A(g8330));
  NOT NOT1_3752(.VSS(VSS),.VDD(VDD),.Y(I10381),.A(g5847));
  NOT NOT1_3753(.VSS(VSS),.VDD(VDD),.Y(g4214),.A(I7459));
  NOT NOT1_3754(.VSS(VSS),.VDD(VDD),.Y(I16255),.A(g10554));
  NOT NOT1_3755(.VSS(VSS),.VDD(VDD),.Y(I14982),.A(g9672));
  NOT NOT1_3756(.VSS(VSS),.VDD(VDD),.Y(g6425),.A(g6141));
  NOT NOT1_3757(.VSS(VSS),.VDD(VDD),.Y(I11728),.A(g7010));
  NOT NOT1_3758(.VSS(VSS),.VDD(VDD),.Y(g11643),.A(I17733));
  NOT NOT1_3759(.VSS(VSS),.VDD(VDD),.Y(g2135),.A(I5064));
  NOT NOT1_3760(.VSS(VSS),.VDD(VDD),.Y(I16679),.A(g10784));
  NOT NOT1_3761(.VSS(VSS),.VDD(VDD),.Y(g2335),.A(I5391));
  NOT NOT1_3762(.VSS(VSS),.VDD(VDD),.Y(g5683),.A(I9202));
  NOT NOT1_3763(.VSS(VSS),.VDD(VDD),.Y(I13439),.A(g8187));
  NOT NOT1_3764(.VSS(VSS),.VDD(VDD),.Y(I9346),.A(g5281));
  NOT NOT1_3765(.VSS(VSS),.VDD(VDD),.Y(I7118),.A(g2979));
  NOT NOT1_3766(.VSS(VSS),.VDD(VDD),.Y(g4310),.A(I7577));
  NOT NOT1_3767(.VSS(VSS),.VDD(VDD),.Y(g2382),.A(g599));
  NOT NOT1_3768(.VSS(VSS),.VDD(VDD),.Y(I7318),.A(g3266));
  NOT NOT1_3769(.VSS(VSS),.VDD(VDD),.Y(I12829),.A(g7680));
  NOT NOT1_3770(.VSS(VSS),.VDD(VDD),.Y(I16124),.A(g10396));
  NOT NOT1_3771(.VSS(VSS),.VDD(VDD),.Y(g10909),.A(I16679));
  NOT NOT1_3772(.VSS(VSS),.VDD(VDD),.Y(I12535),.A(g7656));
  NOT NOT1_3773(.VSS(VSS),.VDD(VDD),.Y(g5778),.A(I9368));
  NOT NOT1_3774(.VSS(VSS),.VDD(VDD),.Y(I10174),.A(g5994));
  NOT NOT1_3775(.VSS(VSS),.VDD(VDD),.Y(I15669),.A(g10194));
  NOT NOT1_3776(.VSS(VSS),.VDD(VDD),.Y(g10543),.A(I16196));
  NOT NOT1_3777(.VSS(VSS),.VDD(VDD),.Y(g3784),.A(g2586));
  NOT NOT1_3778(.VSS(VSS),.VDD(VDD),.Y(I17413),.A(g11425));
  NOT NOT1_3779(.VSS(VSS),.VDD(VDD),.Y(g5894),.A(g5361));
  NOT NOT1_3780(.VSS(VSS),.VDD(VDD),.Y(g9826),.A(I14979));
  NOT NOT1_3781(.VSS(VSS),.VDD(VDD),.Y(g10117),.A(I15359));
  NOT NOT1_3782(.VSS(VSS),.VDD(VDD),.Y(g8660),.A(I13945));
  NOT NOT1_3783(.VSS(VSS),.VDD(VDD),.Y(g8946),.A(I14295));
  NOT NOT1_3784(.VSS(VSS),.VDD(VDD),.Y(g10908),.A(I16676));
  NOT NOT1_3785(.VSS(VSS),.VDD(VDD),.Y(g2916),.A(I6097));
  NOT NOT1_3786(.VSS(VSS),.VDD(VDD),.Y(I7843),.A(g3440));
  NOT NOT1_3787(.VSS(VSS),.VDD(VDD),.Y(g2022),.A(g1346));
  NOT NOT1_3788(.VSS(VSS),.VDD(VDD),.Y(g5735),.A(I9293));
  NOT NOT1_3789(.VSS(VSS),.VDD(VDD),.Y(I15392),.A(g10104));
  NOT NOT1_3790(.VSS(VSS),.VDD(VDD),.Y(g7677),.A(g7148));
  NOT NOT1_3791(.VSS(VSS),.VDD(VDD),.Y(g2749),.A(I5815));
  NOT NOT1_3792(.VSS(VSS),.VDD(VDD),.Y(g3995),.A(g3121));
  NOT NOT1_3793(.VSS(VSS),.VDD(VDD),.Y(g3937),.A(I7086));
  NOT NOT1_3794(.VSS(VSS),.VDD(VDD),.Y(I10840),.A(g6719));
  NOT NOT1_3795(.VSS(VSS),.VDD(VDD),.Y(g9741),.A(I14888));
  NOT NOT1_3796(.VSS(VSS),.VDD(VDD),.Y(g4002),.A(g3121));
  NOT NOT1_3797(.VSS(VSS),.VDD(VDD),.Y(I7393),.A(g4096));
  NOT NOT1_3798(.VSS(VSS),.VDD(VDD),.Y(I16938),.A(g11086));
  NOT NOT1_3799(.VSS(VSS),.VDD(VDD),.Y(I6531),.A(g3186));
  NOT NOT1_3800(.VSS(VSS),.VDD(VDD),.Y(I11348),.A(g6695));
  NOT NOT1_3801(.VSS(VSS),.VDD(VDD),.Y(I12344),.A(g7062));
  NOT NOT1_3802(.VSS(VSS),.VDD(VDD),.Y(I13083),.A(g7921));
  NOT NOT1_3803(.VSS(VSS),.VDD(VDD),.Y(g3479),.A(g2655));
  NOT NOT1_3804(.VSS(VSS),.VDD(VDD),.Y(g11195),.A(g11112));
  NOT NOT1_3805(.VSS(VSS),.VDD(VDD),.Y(g11489),.A(I17482));
  NOT NOT1_3806(.VSS(VSS),.VDD(VDD),.Y(g6131),.A(g5548));
  NOT NOT1_3807(.VSS(VSS),.VDD(VDD),.Y(g5661),.A(I9144));
  NOT NOT1_3808(.VSS(VSS),.VDD(VDD),.Y(g10747),.A(I16432));
  NOT NOT1_3809(.VSS(VSS),.VDD(VDD),.Y(I15559),.A(g10094));
  NOT NOT1_3810(.VSS(VSS),.VDD(VDD),.Y(g5075),.A(g4439));
  NOT NOT1_3811(.VSS(VSS),.VDD(VDD),.Y(g8513),.A(I13708));
  NOT NOT1_3812(.VSS(VSS),.VDD(VDD),.Y(I15488),.A(g10116));
  NOT NOT1_3813(.VSS(VSS),.VDD(VDD),.Y(I15424),.A(g10080));
  NOT NOT1_3814(.VSS(VSS),.VDD(VDD),.Y(g6406),.A(I10314));
  NOT NOT1_3815(.VSS(VSS),.VDD(VDD),.Y(g10242),.A(I15632));
  NOT NOT1_3816(.VSS(VSS),.VDD(VDD),.Y(I8007),.A(g3829));
  NOT NOT1_3817(.VSS(VSS),.VDD(VDD),.Y(g5475),.A(I8892));
  NOT NOT1_3818(.VSS(VSS),.VDD(VDD),.Y(g4762),.A(I8116));
  NOT NOT1_3819(.VSS(VSS),.VDD(VDD),.Y(g2798),.A(g2449));
  NOT NOT1_3820(.VSS(VSS),.VDD(VDD),.Y(g5949),.A(I9591));
  NOT NOT1_3821(.VSS(VSS),.VDD(VDD),.Y(g7349),.A(I11695));
  NOT NOT1_3822(.VSS(VSS),.VDD(VDD),.Y(I10192),.A(g6115));
  NOT NOT1_3823(.VSS(VSS),.VDD(VDD),.Y(g11424),.A(I17327));
  NOT NOT1_3824(.VSS(VSS),.VDD(VDD),.Y(I9240),.A(g5069));
  NOT NOT1_3825(.VSS(VSS),.VDD(VDD),.Y(g6635),.A(I10592));
  NOT NOT1_3826(.VSS(VSS),.VDD(VDD),.Y(I11566),.A(g6820));
  NOT NOT1_3827(.VSS(VSS),.VDD(VDD),.Y(g11016),.A(I16739));
  NOT NOT1_3828(.VSS(VSS),.VDD(VDD),.Y(g9108),.A(I14449));
  NOT NOT1_3829(.VSS(VSS),.VDD(VDD),.Y(g3390),.A(g3161));
  NOT NOT1_3830(.VSS(VSS),.VDD(VDD),.Y(g9308),.A(I14499));
  NOT NOT1_3831(.VSS(VSS),.VDD(VDD),.Y(g8036),.A(I12878));
  NOT NOT1_3832(.VSS(VSS),.VDD(VDD),.Y(g2560),.A(I5684));
  NOT NOT1_3833(.VSS(VSS),.VDD(VDD),.Y(g5627),.A(g4840));
  NOT NOT1_3834(.VSS(VSS),.VDD(VDD),.Y(g8436),.A(I13606));
  NOT NOT1_3835(.VSS(VSS),.VDD(VDD),.Y(g8178),.A(I13083));
  NOT NOT1_3836(.VSS(VSS),.VDD(VDD),.Y(g6801),.A(I10813));
  NOT NOT1_3837(.VSS(VSS),.VDD(VDD),.Y(g6305),.A(I10174));
  NOT NOT1_3838(.VSS(VSS),.VDD(VDD),.Y(I6856),.A(g3318));
  NOT NOT1_3839(.VSS(VSS),.VDD(VDD),.Y(g4590),.A(I7999));
  NOT NOT1_3840(.VSS(VSS),.VDD(VDD),.Y(g7848),.A(I12641));
  NOT NOT1_3841(.VSS(VSS),.VDD(VDD),.Y(g5292),.A(g4445));
  NOT NOT1_3842(.VSS(VSS),.VDD(VDD),.Y(I10663),.A(g6040));
  NOT NOT1_3843(.VSS(VSS),.VDD(VDD),.Y(g8378),.A(I13482));
  NOT NOT1_3844(.VSS(VSS),.VDD(VDD),.Y(g9883),.A(I15060));
  NOT NOT1_3845(.VSS(VSS),.VDD(VDD),.Y(I9043),.A(g4786));
  NOT NOT1_3846(.VSS(VSS),.VDD(VDD),.Y(g3501),.A(g3077));
  NOT NOT1_3847(.VSS(VSS),.VDD(VDD),.Y(I14522),.A(g9108));
  NOT NOT1_3848(.VSS(VSS),.VDD(VDD),.Y(I8535),.A(g4340));
  NOT NOT1_3849(.VSS(VSS),.VDD(VDD),.Y(I9443),.A(g5557));
  NOT NOT1_3850(.VSS(VSS),.VDD(VDD),.Y(g7747),.A(I12406));
  NOT NOT1_3851(.VSS(VSS),.VDD(VDD),.Y(g5998),.A(I9620));
  NOT NOT1_3852(.VSS(VSS),.VDD(VDD),.Y(g5646),.A(I9099));
  NOT NOT1_3853(.VSS(VSS),.VDD(VDD),.Y(g10974),.A(I16723));
  NOT NOT1_3854(.VSS(VSS),.VDD(VDD),.Y(g8335),.A(I13385));
  NOT NOT1_3855(.VSS(VSS),.VDD(VDD),.Y(g2873),.A(I6019));
  NOT NOT1_3856(.VSS(VSS),.VDD(VDD),.Y(g6748),.A(I10753));
  NOT NOT1_3857(.VSS(VSS),.VDD(VDD),.Y(g2632),.A(g2002));
  NOT NOT1_3858(.VSS(VSS),.VDD(VDD),.Y(I6074),.A(g2228));
  NOT NOT1_3859(.VSS(VSS),.VDD(VDD),.Y(g2095),.A(g143));
  NOT NOT1_3860(.VSS(VSS),.VDD(VDD),.Y(I11653),.A(g6954));
  NOT NOT1_3861(.VSS(VSS),.VDD(VDD),.Y(g2037),.A(g1771));
  NOT NOT1_3862(.VSS(VSS),.VDD(VDD),.Y(g8182),.A(I13099));
  NOT NOT1_3863(.VSS(VSS),.VDD(VDD),.Y(I4886),.A(g257));
  NOT NOT1_3864(.VSS(VSS),.VDD(VDD),.Y(g4222),.A(g3638));
  NOT NOT1_3865(.VSS(VSS),.VDD(VDD),.Y(g5603),.A(I9029));
  NOT NOT1_3866(.VSS(VSS),.VDD(VDD),.Y(I6474),.A(g2297));
  NOT NOT1_3867(.VSS(VSS),.VDD(VDD),.Y(I7625),.A(g4164));
  NOT NOT1_3868(.VSS(VSS),.VDD(VDD),.Y(g5039),.A(I8418));
  NOT NOT1_3869(.VSS(VSS),.VDD(VDD),.Y(I4951),.A(g262));
  NOT NOT1_3870(.VSS(VSS),.VDD(VDD),.Y(g10293),.A(I15701));
  NOT NOT1_3871(.VSS(VSS),.VDD(VDD),.Y(g2653),.A(g2011));
  NOT NOT1_3872(.VSS(VSS),.VDD(VDD),.Y(g2208),.A(g84));
  NOT NOT1_3873(.VSS(VSS),.VDD(VDD),.Y(g2302),.A(g29));
  NOT NOT1_3874(.VSS(VSS),.VDD(VDD),.Y(I12029),.A(g6922));
  NOT NOT1_3875(.VSS(VSS),.VDD(VDD),.Y(g5850),.A(g5320));
  NOT NOT1_3876(.VSS(VSS),.VDD(VDD),.Y(g6226),.A(I9973));
  NOT NOT1_3877(.VSS(VSS),.VDD(VDD),.Y(I10553),.A(g6192));
  NOT NOT1_3878(.VSS(VSS),.VDD(VDD),.Y(g3704),.A(I6861));
  NOT NOT1_3879(.VSS(VSS),.VDD(VDD),.Y(g8805),.A(I14136));
  NOT NOT1_3880(.VSS(VSS),.VDD(VDD),.Y(g10265),.A(g10143));
  NOT NOT1_3881(.VSS(VSS),.VDD(VDD),.Y(g2579),.A(g1969));
  NOT NOT1_3882(.VSS(VSS),.VDD(VDD),.Y(I5837),.A(g2507));
  NOT NOT1_3883(.VSS(VSS),.VDD(VDD),.Y(I7938),.A(g3406));
  NOT NOT1_3884(.VSS(VSS),.VDD(VDD),.Y(I9147),.A(g5011));
  NOT NOT1_3885(.VSS(VSS),.VDD(VDD),.Y(I13636),.A(g8357));
  NOT NOT1_3886(.VSS(VSS),.VDD(VDD),.Y(g8422),.A(I13580));
  NOT NOT1_3887(.VSS(VSS),.VDD(VDD),.Y(I10949),.A(g6747));
  NOT NOT1_3888(.VSS(VSS),.VDD(VDD),.Y(I17302),.A(g11391));
  NOT NOT1_3889(.VSS(VSS),.VDD(VDD),.Y(g4899),.A(I8262));
  NOT NOT1_3890(.VSS(VSS),.VDD(VDD),.Y(I11333),.A(g6670));
  NOT NOT1_3891(.VSS(VSS),.VDD(VDD),.Y(I13415),.A(g8144));
  NOT NOT1_3892(.VSS(VSS),.VDD(VDD),.Y(g4464),.A(I7829));
  NOT NOT1_3893(.VSS(VSS),.VDD(VDD),.Y(g2719),.A(g2043));
  NOT NOT1_3894(.VSS(VSS),.VDD(VDD),.Y(g9448),.A(g9091));
  NOT NOT1_3895(.VSS(VSS),.VDD(VDD),.Y(I7909),.A(g3387));
  NOT NOT1_3896(.VSS(VSS),.VDD(VDD),.Y(I6080),.A(g2108));
  NOT NOT1_3897(.VSS(VSS),.VDD(VDD),.Y(I14326),.A(g8818));
  NOT NOT1_3898(.VSS(VSS),.VDD(VDD),.Y(g4785),.A(g3337));
  NOT NOT1_3899(.VSS(VSS),.VDD(VDD),.Y(g11042),.A(I16787));
  NOT NOT1_3900(.VSS(VSS),.VDD(VDD),.Y(g10391),.A(g10313));
  NOT NOT1_3901(.VSS(VSS),.VDD(VDD),.Y(I6480),.A(g2462));
  NOT NOT1_3902(.VSS(VSS),.VDD(VDD),.Y(g5702),.A(I9243));
  NOT NOT1_3903(.VSS(VSS),.VDD(VDD),.Y(g6445),.A(I10367));
  NOT NOT1_3904(.VSS(VSS),.VDD(VDD),.Y(g2752),.A(I5824));
  NOT NOT1_3905(.VSS(VSS),.VDD(VDD),.Y(I14040),.A(g8649));
  NOT NOT1_3906(.VSS(VSS),.VDD(VDD),.Y(I14948),.A(g9555));
  NOT NOT1_3907(.VSS(VSS),.VDD(VDD),.Y(g9827),.A(I14982));
  NOT NOT1_3908(.VSS(VSS),.VDD(VDD),.Y(g6091),.A(I9744));
  NOT NOT1_3909(.VSS(VSS),.VDD(VDD),.Y(I10702),.A(g6071));
  NOT NOT1_3910(.VSS(VSS),.VDD(VDD),.Y(g3810),.A(g3228));
  NOT NOT1_3911(.VSS(VSS),.VDD(VDD),.Y(g3363),.A(I6549));
  NOT NOT1_3912(.VSS(VSS),.VDD(VDD),.Y(I10904),.A(g6558));
  NOT NOT1_3913(.VSS(VSS),.VDD(VDD),.Y(g8798),.A(I14119));
  NOT NOT1_3914(.VSS(VSS),.VDD(VDD),.Y(g7119),.A(I11354));
  NOT NOT1_3915(.VSS(VSS),.VDD(VDD),.Y(g7319),.A(I11605));
  NOT NOT1_3916(.VSS(VSS),.VDD(VDD),.Y(g3432),.A(g3144));
  NOT NOT1_3917(.VSS(VSS),.VDD(VDD),.Y(I6569),.A(g3186));
  NOT NOT1_3918(.VSS(VSS),.VDD(VDD),.Y(g10579),.A(g10528));
  NOT NOT1_3919(.VSS(VSS),.VDD(VDD),.Y(g4563),.A(g3946));
  NOT NOT1_3920(.VSS(VSS),.VDD(VDD),.Y(g9774),.A(g9474));
  NOT NOT1_3921(.VSS(VSS),.VDD(VDD),.Y(I7606),.A(g4166));
  NOT NOT1_3922(.VSS(VSS),.VDD(VDD),.Y(g8560),.A(I13773));
  NOT NOT1_3923(.VSS(VSS),.VDD(VDD),.Y(I14252),.A(g8783));
  NOT NOT1_3924(.VSS(VSS),.VDD(VDD),.Y(g6169),.A(I9896));
  NOT NOT1_3925(.VSS(VSS),.VDD(VDD),.Y(I15383),.A(g10107));
  NOT NOT1_3926(.VSS(VSS),.VDD(VDD),.Y(I16277),.A(g10536));
  NOT NOT1_3927(.VSS(VSS),.VDD(VDD),.Y(g6283),.A(I10108));
  NOT NOT1_3928(.VSS(VSS),.VDD(VDD),.Y(g7352),.A(I11704));
  NOT NOT1_3929(.VSS(VSS),.VDD(VDD),.Y(g2042),.A(g1796));
  NOT NOT1_3930(.VSS(VSS),.VDD(VDD),.Y(g4295),.A(I7556));
  NOT NOT1_3931(.VSS(VSS),.VDD(VDD),.Y(g10578),.A(g10527));
  NOT NOT1_3932(.VSS(VSS),.VDD(VDD),.Y(I9013),.A(g4767));
  NOT NOT1_3933(.VSS(VSS),.VDD(VDD),.Y(g4237),.A(g4013));
  NOT NOT1_3934(.VSS(VSS),.VDD(VDD),.Y(g6407),.A(I10317));
  NOT NOT1_3935(.VSS(VSS),.VDD(VDD),.Y(I14564),.A(g9026));
  NOT NOT1_3936(.VSS(VSS),.VDD(VDD),.Y(g6920),.A(I11034));
  NOT NOT1_3937(.VSS(VSS),.VDD(VDD),.Y(g6578),.A(I10526));
  NOT NOT1_3938(.VSS(VSS),.VDD(VDD),.Y(g6868),.A(I10946));
  NOT NOT1_3939(.VSS(VSS),.VDD(VDD),.Y(g5616),.A(I9046));
  NOT NOT1_3940(.VSS(VSS),.VDD(VDD),.Y(I16595),.A(g10783));
  NOT NOT1_3941(.VSS(VSS),.VDD(VDD),.Y(g8873),.A(I14191));
  NOT NOT1_3942(.VSS(VSS),.VDD(VDD),.Y(g8632),.A(I13915));
  NOT NOT1_3943(.VSS(VSS),.VDD(VDD),.Y(g8095),.A(g7942));
  NOT NOT1_3944(.VSS(VSS),.VDD(VDD),.Y(g2164),.A(I5095));
  NOT NOT1_3945(.VSS(VSS),.VDD(VDD),.Y(g6718),.A(g5949));
  NOT NOT1_3946(.VSS(VSS),.VDD(VDD),.Y(g2364),.A(g611));
  NOT NOT1_3947(.VSS(VSS),.VDD(VDD),.Y(g2233),.A(I5224));
  NOT NOT1_3948(.VSS(VSS),.VDD(VDD),.Y(g9780),.A(g9474));
  NOT NOT1_3949(.VSS(VSS),.VDD(VDD),.Y(g4194),.A(I7399));
  NOT NOT1_3950(.VSS(VSS),.VDD(VDD),.Y(I16623),.A(g10858));
  NOT NOT1_3951(.VSS(VSS),.VDD(VDD),.Y(g8437),.A(I13609));
  NOT NOT1_3952(.VSS(VSS),.VDD(VDD),.Y(I10183),.A(g6108));
  NOT NOT1_3953(.VSS(VSS),.VDD(VDD),.Y(I7586),.A(g4127));
  NOT NOT1_3954(.VSS(VSS),.VDD(VDD),.Y(g11065),.A(g10974));
  NOT NOT1_3955(.VSS(VSS),.VDD(VDD),.Y(g4394),.A(I7729));
  NOT NOT1_3956(.VSS(VSS),.VDD(VDD),.Y(I5192),.A(g55));
  NOT NOT1_3957(.VSS(VSS),.VDD(VDD),.Y(I6976),.A(g2884));
  NOT NOT1_3958(.VSS(VSS),.VDD(VDD),.Y(g2054),.A(g1864));
  NOT NOT1_3959(.VSS(VSS),.VDD(VDD),.Y(g6582),.A(g5949));
  NOT NOT1_3960(.VSS(VSS),.VDD(VDD),.Y(I13609),.A(g8312));
  NOT NOT1_3961(.VSS(VSS),.VDD(VDD),.Y(I14397),.A(g8888));
  NOT NOT1_3962(.VSS(VSS),.VDD(VDD),.Y(g7386),.A(I11767));
  NOT NOT1_3963(.VSS(VSS),.VDD(VDD),.Y(g4731),.A(I8085));
  NOT NOT1_3964(.VSS(VSS),.VDD(VDD),.Y(I11312),.A(g6488));
  NOT NOT1_3965(.VSS(VSS),.VDD(VDD),.Y(g5647),.A(I9102));
  NOT NOT1_3966(.VSS(VSS),.VDD(VDD),.Y(g2454),.A(I5549));
  NOT NOT1_3967(.VSS(VSS),.VDD(VDD),.Y(g8579),.A(I13822));
  NOT NOT1_3968(.VSS(VSS),.VDD(VDD),.Y(g8869),.A(I14179));
  NOT NOT1_3969(.VSS(VSS),.VDD(VDD),.Y(g7975),.A(I12773));
  NOT NOT1_3970(.VSS(VSS),.VDD(VDD),.Y(I13200),.A(g8251));
  NOT NOT1_3971(.VSS(VSS),.VDD(VDD),.Y(g6261),.A(I10042));
  NOT NOT1_3972(.VSS(VSS),.VDD(VDD),.Y(I11608),.A(g6903));
  NOT NOT1_3973(.VSS(VSS),.VDD(VDD),.Y(g2296),.A(I5332));
  NOT NOT1_3974(.VSS(VSS),.VDD(VDD),.Y(I11115),.A(g6462));
  NOT NOT1_3975(.VSS(VSS),.VDD(VDD),.Y(I12604),.A(g7630));
  NOT NOT1_3976(.VSS(VSS),.VDD(VDD),.Y(g10116),.A(I15356));
  NOT NOT1_3977(.VSS(VSS),.VDD(VDD),.Y(I9117),.A(g5615));
  NOT NOT1_3978(.VSS(VSS),.VDD(VDD),.Y(g6793),.A(I10795));
  NOT NOT1_3979(.VSS(VSS),.VDD(VDD),.Y(g8719),.A(g8579));
  NOT NOT1_3980(.VSS(VSS),.VDD(VDD),.Y(g4557),.A(g3946));
  NOT NOT1_3981(.VSS(VSS),.VDD(VDD),.Y(I9317),.A(g5576));
  NOT NOT1_3982(.VSS(VSS),.VDD(VDD),.Y(g2725),.A(g2018));
  NOT NOT1_3983(.VSS(VSS),.VDD(VDD),.Y(g1974),.A(g627));
  NOT NOT1_3984(.VSS(VSS),.VDD(VDD),.Y(I14509),.A(g8926));
  NOT NOT1_3985(.VSS(VSS),.VDD(VDD),.Y(g5546),.A(I8973));
  NOT NOT1_3986(.VSS(VSS),.VDD(VDD),.Y(g7026),.A(I11173));
  NOT NOT1_3987(.VSS(VSS),.VDD(VDD),.Y(I5854),.A(g2523));
  NOT NOT1_3988(.VSS(VSS),.VDD(VDD),.Y(I8388),.A(g4239));
  NOT NOT1_3989(.VSS(VSS),.VDD(VDD),.Y(g4966),.A(I8340));
  NOT NOT1_3990(.VSS(VSS),.VDD(VDD),.Y(I12770),.A(g7638));
  NOT NOT1_3991(.VSS(VSS),.VDD(VDD),.Y(I14933),.A(g9454));
  NOT NOT1_3992(.VSS(VSS),.VDD(VDD),.Y(g7426),.A(I11814));
  NOT NOT1_3993(.VSS(VSS),.VDD(VDD),.Y(g9994),.A(I15196));
  NOT NOT1_3994(.VSS(VSS),.VDD(VDD),.Y(g9290),.A(I14494));
  NOT NOT1_3995(.VSS(VSS),.VDD(VDD),.Y(I11921),.A(g6904));
  NOT NOT1_3996(.VSS(VSS),.VDD(VDD),.Y(I17662),.A(g11602));
  NOT NOT1_3997(.VSS(VSS),.VDD(VDD),.Y(I12981),.A(g8041));
  NOT NOT1_3998(.VSS(VSS),.VDD(VDD),.Y(g8752),.A(g8635));
  NOT NOT1_3999(.VSS(VSS),.VDD(VDD),.Y(g6227),.A(g5446));
  NOT NOT1_4000(.VSS(VSS),.VDD(VDD),.Y(g10041),.A(I15250));
  NOT NOT1_4001(.VSS(VSS),.VDD(VDD),.Y(g5503),.A(g4515));
  NOT NOT1_4002(.VSS(VSS),.VDD(VDD),.Y(I7710),.A(g3749));
  NOT NOT1_4003(.VSS(VSS),.VDD(VDD),.Y(g7614),.A(I12190));
  NOT NOT1_4004(.VSS(VSS),.VDD(VDD),.Y(g10275),.A(I15669));
  NOT NOT1_4005(.VSS(VSS),.VDD(VDD),.Y(g4242),.A(g3664));
  NOT NOT1_4006(.VSS(VSS),.VDD(VDD),.Y(g10493),.A(I16114));
  NOT NOT1_4007(.VSS(VSS),.VDD(VDD),.Y(g7325),.A(I11623));
  NOT NOT1_4008(.VSS(VSS),.VDD(VDD),.Y(I17249),.A(g11342));
  NOT NOT1_4009(.VSS(VSS),.VDD(VDD),.Y(g4948),.A(I8315));
  NOT NOT1_4010(.VSS(VSS),.VDD(VDD),.Y(I7691),.A(g3363));
  NOT NOT1_4011(.VSS(VSS),.VDD(VDD),.Y(g9816),.A(g9490));
  NOT NOT1_4012(.VSS(VSS),.VDD(VDD),.Y(I17482),.A(g11479));
  NOT NOT1_4013(.VSS(VSS),.VDD(VDD),.Y(g10465),.A(I15986));
  NOT NOT1_4014(.VSS(VSS),.VDD(VDD),.Y(g1980),.A(g646));
  NOT NOT1_4015(.VSS(VSS),.VDD(VDD),.Y(I8247),.A(g4615));
  NOT NOT1_4016(.VSS(VSS),.VDD(VDD),.Y(g7984),.A(I12796));
  NOT NOT1_4017(.VSS(VSS),.VDD(VDD),.Y(g2012),.A(g981));
  NOT NOT1_4018(.VSS(VSS),.VDD(VDD),.Y(g11160),.A(g10950));
  NOT NOT1_4019(.VSS(VSS),.VDD(VDD),.Y(g8442),.A(I13624));
  NOT NOT1_4020(.VSS(VSS),.VDD(VDD),.Y(I17710),.A(g11620));
  NOT NOT1_4021(.VSS(VSS),.VDD(VDD),.Y(g6203),.A(g5446));
  NOT NOT1_4022(.VSS(VSS),.VDD(VDD),.Y(I17552),.A(g11502));
  NOT NOT1_4023(.VSS(VSS),.VDD(VDD),.Y(I16853),.A(g10907));
  NOT NOT1_4024(.VSS(VSS),.VDD(VDD),.Y(I9581),.A(g5111));
  NOT NOT1_4025(.VSS(VSS),.VDD(VDD),.Y(g10035),.A(I15241));
  NOT NOT1_4026(.VSS(VSS),.VDD(VDD),.Y(g5120),.A(I8520));
  NOT NOT1_4027(.VSS(VSS),.VDD(VDD),.Y(I5031),.A(g928));
  NOT NOT1_4028(.VSS(VSS),.VDD(VDD),.Y(g5320),.A(g4418));
  NOT NOT1_4029(.VSS(VSS),.VDD(VDD),.Y(g4254),.A(g4013));
  NOT NOT1_4030(.VSS(VSS),.VDD(VDD),.Y(I16589),.A(g10820));
  NOT NOT1_4031(.VSS(VSS),.VDD(VDD),.Y(I11674),.A(g7051));
  NOT NOT1_4032(.VSS(VSS),.VDD(VDD),.Y(g10806),.A(I16518));
  NOT NOT1_4033(.VSS(VSS),.VDD(VDD),.Y(g7544),.A(I11964));
  NOT NOT1_4034(.VSS(VSS),.VDD(VDD),.Y(g8164),.A(g7872));
  NOT NOT1_4035(.VSS(VSS),.VDD(VDD),.Y(I13674),.A(g8304));
  NOT NOT1_4036(.VSS(VSS),.VDD(VDD),.Y(I15470),.A(g10111));
  NOT NOT1_4037(.VSS(VSS),.VDD(VDD),.Y(I5812),.A(g2090));
  NOT NOT1_4038(.VSS(VSS),.VDD(VDD),.Y(g8233),.A(g7872));
  NOT NOT1_4039(.VSS(VSS),.VDD(VDD),.Y(g11617),.A(I17669));
  NOT NOT1_4040(.VSS(VSS),.VDD(VDD),.Y(I6183),.A(g2131));
  NOT NOT1_4041(.VSS(VSS),.VDD(VDD),.Y(g11470),.A(I17447));
  NOT NOT1_4042(.VSS(VSS),.VDD(VDD),.Y(I7659),.A(g3731));
  NOT NOT1_4043(.VSS(VSS),.VDD(VDD),.Y(g10142),.A(I15424));
  NOT NOT1_4044(.VSS(VSS),.VDD(VDD),.Y(g2888),.A(I6046));
  NOT NOT1_4045(.VSS(VSS),.VDD(VDD),.Y(I6924),.A(g2843));
  NOT NOT1_4046(.VSS(VSS),.VDD(VDD),.Y(g7636),.A(I12248));
  NOT NOT1_4047(.VSS(VSS),.VDD(VDD),.Y(I6220),.A(g883));
  NOT NOT1_4048(.VSS(VSS),.VDD(VDD),.Y(I4891),.A(g582));
  NOT NOT1_4049(.VSS(VSS),.VDD(VDD),.Y(g2171),.A(I5116));
  NOT NOT1_4050(.VSS(VSS),.VDD(VDD),.Y(g4438),.A(I7790));
  NOT NOT1_4051(.VSS(VSS),.VDD(VDD),.Y(I14452),.A(g8922));
  NOT NOT1_4052(.VSS(VSS),.VDD(VDD),.Y(g4773),.A(I8133));
  NOT NOT1_4053(.VSS(VSS),.VDD(VDD),.Y(g7306),.A(I11566));
  NOT NOT1_4054(.VSS(VSS),.VDD(VDD),.Y(I13732),.A(g8291));
  NOT NOT1_4055(.VSS(VSS),.VDD(VDD),.Y(g8296),.A(I13242));
  NOT NOT1_4056(.VSS(VSS),.VDD(VDD),.Y(g2956),.A(I6159));
  NOT NOT1_4057(.VSS(VSS),.VDD(VDD),.Y(I15075),.A(g9761));
  NOT NOT1_4058(.VSS(VSS),.VDD(VDD),.Y(g8725),.A(g8589));
  NOT NOT1_4059(.VSS(VSS),.VDD(VDD),.Y(g7790),.A(I12535));
  NOT NOT1_4060(.VSS(VSS),.VDD(VDD),.Y(g9263),.A(g8892));
  NOT NOT1_4061(.VSS(VSS),.VDD(VDD),.Y(g3683),.A(I6844));
  NOT NOT1_4062(.VSS(VSS),.VDD(VDD),.Y(g11075),.A(g10937));
  NOT NOT1_4063(.VSS(VSS),.VDD(VDD),.Y(I5765),.A(g2004));
  NOT NOT1_4064(.VSS(VSS),.VDD(VDD),.Y(I15595),.A(g10165));
  NOT NOT1_4065(.VSS(VSS),.VDD(VDD),.Y(I15467),.A(g10079));
  NOT NOT1_4066(.VSS(VSS),.VDD(VDD),.Y(I15494),.A(g10117));
  NOT NOT1_4067(.VSS(VSS),.VDD(VDD),.Y(I17356),.A(g11384));
  NOT NOT1_4068(.VSS(VSS),.VDD(VDD),.Y(g8532),.A(I13741));
  NOT NOT1_4069(.VSS(VSS),.VDD(VDD),.Y(I8308),.A(g4443));
  NOT NOT1_4070(.VSS(VSS),.VDD(VDD),.Y(g7187),.A(I11405));
  NOT NOT1_4071(.VSS(VSS),.VDD(VDD),.Y(I7311),.A(g2803));
  NOT NOT1_4072(.VSS(VSS),.VDD(VDD),.Y(g4769),.A(g3586));
  NOT NOT1_4073(.VSS(VSS),.VDD(VDD),.Y(g5987),.A(I9605));
  NOT NOT1_4074(.VSS(VSS),.VDD(VDD),.Y(I11692),.A(g7048));
  NOT NOT1_4075(.VSS(VSS),.VDD(VDD),.Y(g7387),.A(I11770));
  NOT NOT1_4076(.VSS(VSS),.VDD(VDD),.Y(g11467),.A(I17438));
  NOT NOT1_4077(.VSS(VSS),.VDD(VDD),.Y(I9995),.A(g5536));
  NOT NOT1_4078(.VSS(VSS),.VDD(VDD),.Y(I12832),.A(g7681));
  NOT NOT1_4079(.VSS(VSS),.VDD(VDD),.Y(I4859),.A(g578));
  NOT NOT1_4080(.VSS(VSS),.VDD(VDD),.Y(I10051),.A(g5702));
  NOT NOT1_4081(.VSS(VSS),.VDD(VDD),.Y(I10072),.A(g5719));
  NOT NOT1_4082(.VSS(VSS),.VDD(VDD),.Y(g4212),.A(I7453));
  NOT NOT1_4083(.VSS(VSS),.VDD(VDD),.Y(I9479),.A(g4954));
  NOT NOT1_4084(.VSS(VSS),.VDD(VDD),.Y(g6689),.A(g5830));
  NOT NOT1_4085(.VSS(VSS),.VDD(VDD),.Y(g10130),.A(I15392));
  NOT NOT1_4086(.VSS(VSS),.VDD(VDD),.Y(g7756),.A(I12433));
  NOT NOT1_4087(.VSS(VSS),.VDD(VDD),.Y(g2297),.A(g865));
  NOT NOT1_4088(.VSS(VSS),.VDD(VDD),.Y(g11623),.A(I17687));
  NOT NOT1_4089(.VSS(VSS),.VDD(VDD),.Y(g6388),.A(I10286));
  NOT NOT1_4090(.VSS(VSS),.VDD(VDD),.Y(g10193),.A(g10057));
  NOT NOT1_4091(.VSS(VSS),.VDD(VDD),.Y(I16616),.A(g10796));
  NOT NOT1_4092(.VSS(VSS),.VDD(VDD),.Y(g11037),.A(I16772));
  NOT NOT1_4093(.VSS(VSS),.VDD(VDD),.Y(I10592),.A(g5865));
  NOT NOT1_4094(.VSS(VSS),.VDD(VDD),.Y(g5299),.A(g4393));
  NOT NOT1_4095(.VSS(VSS),.VDD(VDD),.Y(I10756),.A(g5810));
  NOT NOT1_4096(.VSS(VSS),.VDD(VDD),.Y(I15782),.A(g10259));
  NOT NOT1_4097(.VSS(VSS),.VDD(VDD),.Y(g7622),.A(g7067));
  NOT NOT1_4098(.VSS(VSS),.VDD(VDD),.Y(g3735),.A(I6921));
  NOT NOT1_4099(.VSS(VSS),.VDD(VDD),.Y(g7027),.A(I11176));
  NOT NOT1_4100(.VSS(VSS),.VDD(VDD),.Y(g7427),.A(I11817));
  NOT NOT1_4101(.VSS(VSS),.VDD(VDD),.Y(I17182),.A(g11309));
  NOT NOT1_4102(.VSS(VSS),.VDD(VDD),.Y(g10165),.A(I15491));
  NOT NOT1_4103(.VSS(VSS),.VDD(VDD),.Y(I13400),.A(g8236));
  NOT NOT1_4104(.VSS(VSS),.VDD(VDD),.Y(g10523),.A(g10456));
  NOT NOT1_4105(.VSS(VSS),.VDD(VDD),.Y(I17672),.A(g11605));
  NOT NOT1_4106(.VSS(VSS),.VDD(VDD),.Y(g3782),.A(I7006));
  NOT NOT1_4107(.VSS(VSS),.VDD(VDD),.Y(I13013),.A(g8048));
  NOT NOT1_4108(.VSS(VSS),.VDD(VDD),.Y(g5892),.A(I9519));
  NOT NOT1_4109(.VSS(VSS),.VDD(VDD),.Y(I11214),.A(g6528));
  NOT NOT1_4110(.VSS(VSS),.VDD(VDD),.Y(g7904),.A(I12690));
  NOT NOT1_4111(.VSS(VSS),.VDD(VDD),.Y(g11419),.A(I17312));
  NOT NOT1_4112(.VSS(VSS),.VDD(VDD),.Y(g2745),.A(I5809));
  NOT NOT1_4113(.VSS(VSS),.VDD(VDD),.Y(g2639),.A(I5754));
  NOT NOT1_4114(.VSS(VSS),.VDD(VDD),.Y(g6030),.A(I9639));
  NOT NOT1_4115(.VSS(VSS),.VDD(VDD),.Y(g2338),.A(g1909));
  NOT NOT1_4116(.VSS(VSS),.VDD(VDD),.Y(g11352),.A(I17173));
  NOT NOT1_4117(.VSS(VSS),.VDD(VDD),.Y(I15418),.A(g10083));
  NOT NOT1_4118(.VSS(VSS),.VDD(VDD),.Y(I5073),.A(g34));
  NOT NOT1_4119(.VSS(VSS),.VDD(VDD),.Y(I13329),.A(g8116));
  NOT NOT1_4120(.VSS(VSS),.VDD(VDD),.Y(I11207),.A(g6524));
  NOT NOT1_4121(.VSS(VSS),.VDD(VDD),.Y(g7446),.A(g7148));
  NOT NOT1_4122(.VSS(VSS),.VDD(VDD),.Y(g3475),.A(g3056));
  NOT NOT1_4123(.VSS(VSS),.VDD(VDD),.Y(I6999),.A(g2905));
  NOT NOT1_4124(.VSS(VSS),.VDD(VDD),.Y(g11155),.A(g10950));
  NOT NOT1_4125(.VSS(VSS),.VDD(VDD),.Y(I7284),.A(g3255));
  NOT NOT1_4126(.VSS(VSS),.VDD(VDD),.Y(I15266),.A(g10001));
  NOT NOT1_4127(.VSS(VSS),.VDD(VDD),.Y(g8990),.A(I14391));
  NOT NOT1_4128(.VSS(VSS),.VDD(VDD),.Y(I9156),.A(g5032));
  NOT NOT1_4129(.VSS(VSS),.VDD(VDD),.Y(I12099),.A(g7258));
  NOT NOT1_4130(.VSS(VSS),.VDD(VDD),.Y(I11005),.A(g6386));
  NOT NOT1_4131(.VSS(VSS),.VDD(VDD),.Y(I12388),.A(g7219));
  NOT NOT1_4132(.VSS(VSS),.VDD(VDD),.Y(I17331),.A(g11357));
  NOT NOT1_4133(.VSS(VSS),.VDD(VDD),.Y(I13005),.A(g8046));
  NOT NOT1_4134(.VSS(VSS),.VDD(VDD),.Y(g8888),.A(I14232));
  NOT NOT1_4135(.VSS(VSS),.VDD(VDD),.Y(g7403),.A(I11783));
  NOT NOT1_4136(.VSS(VSS),.VDD(VDD),.Y(g3627),.A(I6784));
  NOT NOT1_4137(.VSS(VSS),.VDD(VDD),.Y(g4822),.A(g3706));
  NOT NOT1_4138(.VSS(VSS),.VDD(VDD),.Y(g8029),.A(I12871));
  NOT NOT1_4139(.VSS(VSS),.VDD(VDD),.Y(g6564),.A(g5784));
  NOT NOT1_4140(.VSS(VSS),.VDD(VDD),.Y(I16808),.A(g10906));
  NOT NOT1_4141(.VSS(VSS),.VDD(VDD),.Y(g8171),.A(I13068));
  NOT NOT1_4142(.VSS(VSS),.VDD(VDD),.Y(g7345),.A(I11683));
  NOT NOT1_4143(.VSS(VSS),.VDD(VDD),.Y(I17513),.A(g11482));
  NOT NOT1_4144(.VSS(VSS),.VDD(VDD),.Y(I8711),.A(g4530));
  NOT NOT1_4145(.VSS(VSS),.VDD(VDD),.Y(g2808),.A(g2156));
  NOT NOT1_4146(.VSS(VSS),.VDD(VDD),.Y(g3292),.A(g2373));
  NOT NOT1_4147(.VSS(VSS),.VDD(VDD),.Y(I10846),.A(g6729));
  NOT NOT1_4148(.VSS(VSS),.VDD(VDD),.Y(g8787),.A(I14094));
  NOT NOT1_4149(.VSS(VSS),.VDD(VDD),.Y(I12251),.A(g7076));
  NOT NOT1_4150(.VSS(VSS),.VDD(VDD),.Y(g7763),.A(I12454));
  NOT NOT1_4151(.VSS(VSS),.VDD(VDD),.Y(I16101),.A(g10381));
  NOT NOT1_4152(.VSS(VSS),.VDD(VDD),.Y(g8956),.A(I14319));
  NOT NOT1_4153(.VSS(VSS),.VDD(VDD),.Y(g2707),.A(g2041));
  NOT NOT1_4154(.VSS(VSS),.VDD(VDD),.Y(I8827),.A(g4477));
  NOT NOT1_4155(.VSS(VSS),.VDD(VDD),.Y(g10437),.A(g10333));
  NOT NOT1_4156(.VSS(VSS),.VDD(VDD),.Y(I8133),.A(g3632));
  NOT NOT1_4157(.VSS(VSS),.VDD(VDD),.Y(g2759),.A(I5843));
  NOT NOT1_4158(.VSS(VSS),.VDD(VDD),.Y(I8333),.A(g4456));
  NOT NOT1_4159(.VSS(VSS),.VDD(VDD),.Y(I7420),.A(g4167));
  NOT NOT1_4160(.VSS(VSS),.VDD(VDD),.Y(g7637),.A(I12251));
  NOT NOT1_4161(.VSS(VSS),.VDD(VDD),.Y(I15589),.A(g10161));
  NOT NOT1_4162(.VSS(VSS),.VDD(VDD),.Y(g5078),.A(g4372));
  NOT NOT1_4163(.VSS(VSS),.VDD(VDD),.Y(g3039),.A(g2310));
  NOT NOT1_4164(.VSS(VSS),.VDD(VDD),.Y(g2201),.A(g102));
  NOT NOT1_4165(.VSS(VSS),.VDD(VDD),.Y(g3439),.A(g3144));
  NOT NOT1_4166(.VSS(VSS),.VDD(VDD),.Y(g7107),.A(I11342));
  NOT NOT1_4167(.VSS(VSS),.VDD(VDD),.Y(I7559),.A(g4116));
  NOT NOT1_4168(.VSS(VSS),.VDD(VDD),.Y(g7307),.A(I11569));
  NOT NOT1_4169(.VSS(VSS),.VDD(VDD),.Y(I12032),.A(g6923));
  NOT NOT1_4170(.VSS(VSS),.VDD(VDD),.Y(g8297),.A(I13245));
  NOT NOT1_4171(.VSS(VSS),.VDD(VDD),.Y(g10347),.A(I15807));
  NOT NOT1_4172(.VSS(VSS),.VDD(VDD),.Y(g5035),.A(I8410));
  NOT NOT1_4173(.VSS(VSS),.VDD(VDD),.Y(I6944),.A(g2859));
  NOT NOT1_4174(.VSS(VSS),.VDD(VDD),.Y(I8396),.A(g4255));
  NOT NOT1_4175(.VSS(VSS),.VDD(VDD),.Y(g10253),.A(g10138));
  NOT NOT1_4176(.VSS(VSS),.VDD(VDD),.Y(I6240),.A(g878));
  NOT NOT1_4177(.VSS(VSS),.VDD(VDD),.Y(I7931),.A(g3624));
  NOT NOT1_4178(.VSS(VSS),.VDD(VDD),.Y(g7359),.A(I11725));
  NOT NOT1_4179(.VSS(VSS),.VDD(VDD),.Y(g6108),.A(I9779));
  NOT NOT1_4180(.VSS(VSS),.VDD(VDD),.Y(g6308),.A(I10183));
  NOT NOT1_4181(.VSS(VSS),.VDD(VDD),.Y(I9810),.A(g5576));
  NOT NOT1_4182(.VSS(VSS),.VDD(VDD),.Y(g5082),.A(g4840));
  NOT NOT1_4183(.VSS(VSS),.VDD(VDD),.Y(g2449),.A(g790));
  NOT NOT1_4184(.VSS(VSS),.VDD(VDD),.Y(I9032),.A(g4732));
  NOT NOT1_4185(.VSS(VSS),.VDD(VDD),.Y(I11100),.A(g6442));
  NOT NOT1_4186(.VSS(VSS),.VDD(VDD),.Y(g5482),.A(I8903));
  NOT NOT1_4187(.VSS(VSS),.VDD(VDD),.Y(I14405),.A(g8937));
  NOT NOT1_4188(.VSS(VSS),.VDD(VDD),.Y(g10600),.A(I16277));
  NOT NOT1_4189(.VSS(VSS),.VDD(VDD),.Y(g11401),.A(I17246));
  NOT NOT1_4190(.VSS(VSS),.VDD(VDD),.Y(g10781),.A(I16475));
  NOT NOT1_4191(.VSS(VSS),.VDD(VDD),.Y(I4783),.A(g873));
  NOT NOT1_4192(.VSS(VSS),.VDD(VDD),.Y(I6043),.A(g2267));
  NOT NOT1_4193(.VSS(VSS),.VDD(VDD),.Y(I9053),.A(g4752));
  NOT NOT1_4194(.VSS(VSS),.VDD(VDD),.Y(g8684),.A(I13969));
  NOT NOT1_4195(.VSS(VSS),.VDD(VDD),.Y(g3583),.A(I6742));
  NOT NOT1_4196(.VSS(VSS),.VDD(VDD),.Y(g4895),.A(I8250));
  NOT NOT1_4197(.VSS(VSS),.VDD(VDD),.Y(g5876),.A(g5361));
  NOT NOT1_4198(.VSS(VSS),.VDD(VDD),.Y(g8138),.A(I13013));
  NOT NOT1_4199(.VSS(VSS),.VDD(VDD),.Y(I6443),.A(g2363));
  NOT NOT1_4200(.VSS(VSS),.VDD(VDD),.Y(I11235),.A(g6538));
  NOT NOT1_4201(.VSS(VSS),.VDD(VDD),.Y(g8338),.A(I13394));
  NOT NOT1_4202(.VSS(VSS),.VDD(VDD),.Y(g10236),.A(g10190));
  NOT NOT1_4203(.VSS(VSS),.VDD(VDD),.Y(g7757),.A(I12436));
  NOT NOT1_4204(.VSS(VSS),.VDD(VDD),.Y(g2604),.A(I5713));
  NOT NOT1_4205(.VSS(VSS),.VDD(VDD),.Y(g4062),.A(I7185));
  NOT NOT1_4206(.VSS(VSS),.VDD(VDD),.Y(g2098),.A(I4938));
  NOT NOT1_4207(.VSS(VSS),.VDD(VDD),.Y(I11683),.A(g7069));
  NOT NOT1_4208(.VSS(VSS),.VDD(VDD),.Y(g5656),.A(I9129));
  NOT NOT1_4209(.VSS(VSS),.VDD(VDD),.Y(g7416),.A(I11800));
  NOT NOT1_4210(.VSS(VSS),.VDD(VDD),.Y(g4620),.A(I8031));
  NOT NOT1_4211(.VSS(VSS),.VDD(VDD),.Y(g10351),.A(I15817));
  NOT NOT1_4212(.VSS(VSS),.VDD(VDD),.Y(g4462),.A(I7825));
  NOT NOT1_4213(.VSS(VSS),.VDD(VDD),.Y(I15864),.A(g10339));
  NOT NOT1_4214(.VSS(VSS),.VDD(VDD),.Y(I5399),.A(g895));
  NOT NOT1_4215(.VSS(VSS),.VDD(VDD),.Y(g6589),.A(I10549));
  NOT NOT1_4216(.VSS(VSS),.VDD(VDD),.Y(I12871),.A(g7638));
  NOT NOT1_4217(.VSS(VSS),.VDD(VDD),.Y(g10175),.A(I15517));
  NOT NOT1_4218(.VSS(VSS),.VDD(VDD),.Y(g10821),.A(I16531));
  NOT NOT1_4219(.VSS(VSS),.VDD(VDD),.Y(I7630),.A(g3524));
  NOT NOT1_4220(.VSS(VSS),.VDD(VDD),.Y(I15749),.A(g10263));
  NOT NOT1_4221(.VSS(VSS),.VDD(VDD),.Y(g2833),.A(I5949));
  NOT NOT1_4222(.VSS(VSS),.VDD(VDD),.Y(I6034),.A(g2210));
  NOT NOT1_4223(.VSS(VSS),.VDD(VDD),.Y(g7522),.A(I11904));
  NOT NOT1_4224(.VSS(VSS),.VDD(VDD),.Y(I8418),.A(g4794));
  NOT NOT1_4225(.VSS(VSS),.VDD(VDD),.Y(g7811),.A(I12598));
  NOT NOT1_4226(.VSS(VSS),.VDD(VDD),.Y(g7315),.A(I11593));
  NOT NOT1_4227(.VSS(VSS),.VDD(VDD),.Y(g11616),.A(I17666));
  NOT NOT1_4228(.VSS(VSS),.VDD(VDD),.Y(I17149),.A(g11306));
  NOT NOT1_4229(.VSS(VSS),.VDD(VDD),.Y(I6565),.A(g2614));
  NOT NOT1_4230(.VSS(VSS),.VDD(VDD),.Y(g7047),.A(I11222));
  NOT NOT1_4231(.VSS(VSS),.VDD(VDD),.Y(I7300),.A(g2883));
  NOT NOT1_4232(.VSS(VSS),.VDD(VDD),.Y(g11313),.A(I17104));
  NOT NOT1_4233(.VSS(VSS),.VDD(VDD),.Y(I12360),.A(g7183));
  NOT NOT1_4234(.VSS(VSS),.VDD(VDD),.Y(I8290),.A(g4778));
  NOT NOT1_4235(.VSS(VSS),.VDD(VDD),.Y(g10063),.A(I15287));
  NOT NOT1_4236(.VSS(VSS),.VDD(VDD),.Y(I17387),.A(g11438));
  NOT NOT1_4237(.VSS(VSS),.VDD(VDD),.Y(g8707),.A(g8671));
  NOT NOT1_4238(.VSS(VSS),.VDD(VDD),.Y(g6165),.A(g5446));
  NOT NOT1_4239(.VSS(VSS),.VDD(VDD),.Y(g10264),.A(g10128));
  NOT NOT1_4240(.VSS(VSS),.VDD(VDD),.Y(g6571),.A(I10503));
  NOT NOT1_4241(.VSS(VSS),.VDD(VDD),.Y(g6365),.A(I10274));
  NOT NOT1_4242(.VSS(VSS),.VDD(VDD),.Y(g6861),.A(I10941));
  NOT NOT1_4243(.VSS(VSS),.VDD(VDD),.Y(g5214),.A(g4640));
  NOT NOT1_4244(.VSS(VSS),.VDD(VDD),.Y(g10137),.A(I15409));
  NOT NOT1_4245(.VSS(VSS),.VDD(VDD),.Y(g6048),.A(I9673));
  NOT NOT1_4246(.VSS(VSS),.VDD(VDD),.Y(I11515),.A(g6589));
  NOT NOT1_4247(.VSS(VSS),.VDD(VDD),.Y(g9772),.A(g9432));
  NOT NOT1_4248(.VSS(VSS),.VDD(VDD),.Y(I11882),.A(g6895));
  NOT NOT1_4249(.VSS(VSS),.VDD(VDD),.Y(I5510),.A(g588));
  NOT NOT1_4250(.VSS(VSS),.VDD(VDD),.Y(g2539),.A(I5652));
  NOT NOT1_4251(.VSS(VSS),.VDD(VDD),.Y(g2896),.A(g2356));
  NOT NOT1_4252(.VSS(VSS),.VDD(VDD),.Y(I6347),.A(g2462));
  NOT NOT1_4253(.VSS(VSS),.VDD(VDD),.Y(I15704),.A(g10238));
  NOT NOT1_4254(.VSS(VSS),.VDD(VDD),.Y(I5245),.A(g925));
  NOT NOT1_4255(.VSS(VSS),.VDD(VDD),.Y(g6448),.A(I10374));
  NOT NOT1_4256(.VSS(VSS),.VDD(VDD),.Y(g9531),.A(I14678));
  NOT NOT1_4257(.VSS(VSS),.VDD(VDD),.Y(I15305),.A(g10001));
  NOT NOT1_4258(.VSS(VSS),.VDD(VDD),.Y(g6711),.A(g5949));
  NOT NOT1_4259(.VSS(VSS),.VDD(VDD),.Y(g6055),.A(I9688));
  NOT NOT1_4260(.VSS(VSS),.VDD(VDD),.Y(I12162),.A(g7146));
  NOT NOT1_4261(.VSS(VSS),.VDD(VDD),.Y(I17104),.A(g11223));
  NOT NOT1_4262(.VSS(VSS),.VDD(VDD),.Y(g10873),.A(I16589));
  NOT NOT1_4263(.VSS(VSS),.VDD(VDD),.Y(g11053),.A(g10950));
  NOT NOT1_4264(.VSS(VSS),.VDD(VDD),.Y(I8256),.A(g4711));
  NOT NOT1_4265(.VSS(VSS),.VDD(VDD),.Y(g9890),.A(I15075));
  NOT NOT1_4266(.VSS(VSS),.VDD(VDD),.Y(I10282),.A(g6163));
  NOT NOT1_4267(.VSS(VSS),.VDD(VDD),.Y(g3404),.A(g3121));
  NOT NOT1_4268(.VSS(VSS),.VDD(VDD),.Y(g6133),.A(I9836));
  NOT NOT1_4269(.VSS(VSS),.VDD(VDD),.Y(g11466),.A(I17435));
  NOT NOT1_4270(.VSS(VSS),.VDD(VDD),.Y(g5663),.A(I9150));
  NOT NOT1_4271(.VSS(VSS),.VDD(VDD),.Y(I10302),.A(g6179));
  NOT NOT1_4272(.VSS(VSS),.VDD(VDD),.Y(I6914),.A(g2828));
  NOT NOT1_4273(.VSS(VSS),.VDD(VDD),.Y(g9505),.A(g9052));
  NOT NOT1_4274(.VSS(VSS),.VDD(VDD),.Y(g2162),.A(I5089));
  NOT NOT1_4275(.VSS(VSS),.VDD(VDD),.Y(I7973),.A(g3437));
  NOT NOT1_4276(.VSS(VSS),.VDD(VDD),.Y(I15036),.A(g9721));
  NOT NOT1_4277(.VSS(VSS),.VDD(VDD),.Y(g2268),.A(g654));
  NOT NOT1_4278(.VSS(VSS),.VDD(VDD),.Y(g8449),.A(I13645));
  NOT NOT1_4279(.VSS(VSS),.VDD(VDD),.Y(g4192),.A(I7393));
  NOT NOT1_4280(.VSS(VSS),.VDD(VDD),.Y(I10105),.A(g5736));
  NOT NOT1_4281(.VSS(VSS),.VDD(VDD),.Y(g4298),.A(g4130));
  NOT NOT1_4282(.VSS(VSS),.VDD(VDD),.Y(g3764),.A(I6971));
  NOT NOT1_4283(.VSS(VSS),.VDD(VDD),.Y(I12451),.A(g7538));
  NOT NOT1_4284(.VSS(VSS),.VDD(VDD),.Y(g6846),.A(I10910));
  NOT NOT1_4285(.VSS(VSS),.VDD(VDD),.Y(g11036),.A(I16769));
  NOT NOT1_4286(.VSS(VSS),.VDD(VDD),.Y(I12472),.A(g7539));
  NOT NOT1_4287(.VSS(VSS),.VDD(VDD),.Y(g8575),.A(I13816));
  NOT NOT1_4288(.VSS(VSS),.VDD(VDD),.Y(g3546),.A(g3307));
  NOT NOT1_4289(.VSS(VSS),.VDD(VDD),.Y(I14105),.A(g8776));
  NOT NOT1_4290(.VSS(VSS),.VDD(VDD),.Y(g4485),.A(g3546));
  NOT NOT1_4291(.VSS(VSS),.VDD(VDD),.Y(I6013),.A(g2200));
  NOT NOT1_4292(.VSS(VSS),.VDD(VDD),.Y(g5402),.A(I8842));
  NOT NOT1_4293(.VSS(VSS),.VDD(VDD),.Y(g6196),.A(g5446));
  NOT NOT1_4294(.VSS(VSS),.VDD(VDD),.Y(g7880),.A(g7479));
  NOT NOT1_4295(.VSS(VSS),.VDD(VDD),.Y(g6396),.A(I10296));
  NOT NOT1_4296(.VSS(VSS),.VDD(VDD),.Y(g7595),.A(I12123));
  NOT NOT1_4297(.VSS(VSS),.VDD(VDD),.Y(g6803),.A(I10819));
  NOT NOT1_4298(.VSS(VSS),.VDD(VDD),.Y(g7537),.A(I11947));
  NOT NOT1_4299(.VSS(VSS),.VDD(VDD),.Y(g5236),.A(g4361));
  NOT NOT1_4300(.VSS(VSS),.VDD(VDD),.Y(I17368),.A(g11423));
  NOT NOT1_4301(.VSS(VSS),.VDD(VDD),.Y(g8604),.A(g8479));
  NOT NOT1_4302(.VSS(VSS),.VDD(VDD),.Y(g10208),.A(I15580));
  NOT NOT1_4303(.VSS(VSS),.VDD(VDD),.Y(I16239),.A(g10525));
  NOT NOT1_4304(.VSS(VSS),.VDD(VDD),.Y(g11642),.A(I17730));
  NOT NOT1_4305(.VSS(VSS),.VDD(VDD),.Y(g8498),.A(g8353));
  NOT NOT1_4306(.VSS(VSS),.VDD(VDD),.Y(I11584),.A(g6827));
  NOT NOT1_4307(.VSS(VSS),.VDD(VDD),.Y(g1972),.A(g461));
  NOT NOT1_4308(.VSS(VSS),.VDD(VDD),.Y(I8421),.A(g4309));
  NOT NOT1_4309(.VSS(VSS),.VDD(VDD),.Y(g9474),.A(g9331));
  NOT NOT1_4310(.VSS(VSS),.VDD(VDD),.Y(g7272),.A(I11519));
  NOT NOT1_4311(.VSS(VSS),.VDD(VDD),.Y(I13206),.A(g8197));
  NOT NOT1_4312(.VSS(VSS),.VDD(VDD),.Y(g10542),.A(I16193));
  NOT NOT1_4313(.VSS(VSS),.VDD(VDD),.Y(g6509),.A(I10427));
  NOT NOT1_4314(.VSS(VSS),.VDD(VDD),.Y(g11064),.A(g10974));
  NOT NOT1_4315(.VSS(VSS),.VDD(VDD),.Y(I15733),.A(g10257));
  NOT NOT1_4316(.VSS(VSS),.VDD(VDD),.Y(g7612),.A(I12186));
  NOT NOT1_4317(.VSS(VSS),.VDD(VDD),.Y(g7243),.A(I11483));
  NOT NOT1_4318(.VSS(VSS),.VDD(VDD),.Y(g2086),.A(I4906));
  NOT NOT1_4319(.VSS(VSS),.VDD(VDD),.Y(I11759),.A(g7244));
  NOT NOT1_4320(.VSS(VSS),.VDD(VDD),.Y(I11725),.A(g7040));
  NOT NOT1_4321(.VSS(VSS),.VDD(VDD),.Y(I12776),.A(g7586));
  NOT NOT1_4322(.VSS(VSS),.VDD(VDD),.Y(g5657),.A(I9132));
  NOT NOT1_4323(.VSS(VSS),.VDD(VDD),.Y(g10913),.A(I16691));
  NOT NOT1_4324(.VSS(VSS),.VDD(VDD),.Y(I16941),.A(g11076));
  NOT NOT1_4325(.VSS(VSS),.VDD(VDD),.Y(g2728),.A(g2025));
  NOT NOT1_4326(.VSS(VSS),.VDD(VDD),.Y(I13114),.A(g7930));
  NOT NOT1_4327(.VSS(VSS),.VDD(VDD),.Y(g6418),.A(g6137));
  NOT NOT1_4328(.VSS(VSS),.VDD(VDD),.Y(I11082),.A(g6749));
  NOT NOT1_4329(.VSS(VSS),.VDD(VDD),.Y(g7982),.A(I12790));
  NOT NOT1_4330(.VSS(VSS),.VDD(VDD),.Y(g4520),.A(I7923));
  NOT NOT1_4331(.VSS(VSS),.VDD(VDD),.Y(g5222),.A(g4640));
  NOT NOT1_4332(.VSS(VSS),.VDD(VDD),.Y(I17228),.A(g11300));
  NOT NOT1_4333(.VSS(VSS),.VDD(VDD),.Y(g11630),.A(I17704));
  NOT NOT1_4334(.VSS(VSS),.VDD(VDD),.Y(g2185),.A(g46));
  NOT NOT1_4335(.VSS(VSS),.VDD(VDD),.Y(g4219),.A(g3635));
  NOT NOT1_4336(.VSS(VSS),.VDD(VDD),.Y(g6290),.A(I10129));
  NOT NOT1_4337(.VSS(VSS),.VDD(VDD),.Y(I7151),.A(g2642));
  NOT NOT1_4338(.VSS(VSS),.VDD(VDD),.Y(g2881),.A(I6031));
  NOT NOT1_4339(.VSS(VSS),.VDD(VDD),.Y(I7351),.A(g4061));
  NOT NOT1_4340(.VSS(VSS),.VDD(VDD),.Y(I16518),.A(g10718));
  NOT NOT1_4341(.VSS(VSS),.VDD(VDD),.Y(I6601),.A(g3186));
  NOT NOT1_4342(.VSS(VSS),.VDD(VDD),.Y(I7648),.A(g3727));
  NOT NOT1_4343(.VSS(VSS),.VDD(VDD),.Y(I12825),.A(g7696));
  NOT NOT1_4344(.VSS(VSS),.VDD(VDD),.Y(g10320),.A(I15756));
  NOT NOT1_4345(.VSS(VSS),.VDD(VDD),.Y(g10905),.A(I16667));
  NOT NOT1_4346(.VSS(VSS),.VDD(VDD),.Y(g7629),.A(I12229));
  NOT NOT1_4347(.VSS(VSS),.VDD(VDD),.Y(I15665),.A(g10193));
  NOT NOT1_4348(.VSS(VSS),.VDD(VDD),.Y(g7328),.A(I11632));
  NOT NOT1_4349(.VSS(VSS),.VDD(VDD),.Y(g2070),.A(g213));
  NOT NOT1_4350(.VSS(VSS),.VDD(VDD),.Y(g10530),.A(g10466));
  NOT NOT1_4351(.VSS(VSS),.VDD(VDD),.Y(g3906),.A(g3015));
  NOT NOT1_4352(.VSS(VSS),.VDD(VDD),.Y(I17716),.A(g11622));
  NOT NOT1_4353(.VSS(VSS),.VDD(VDD),.Y(g7330),.A(I11638));
  NOT NOT1_4354(.VSS(VSS),.VDD(VDD),.Y(g10593),.A(I16264));
  NOT NOT1_4355(.VSS(VSS),.VDD(VDD),.Y(I4866),.A(g579));
  NOT NOT1_4356(.VSS(VSS),.VDD(VDD),.Y(g8362),.A(I13466));
  NOT NOT1_4357(.VSS(VSS),.VDD(VDD),.Y(I13744),.A(g8297));
  NOT NOT1_4358(.VSS(VSS),.VDD(VDD),.Y(g2025),.A(g1696));
  NOT NOT1_4359(.VSS(VSS),.VDD(VDD),.Y(I11345),.A(g6692));
  NOT NOT1_4360(.VSS(VSS),.VDD(VDD),.Y(g10346),.A(I15804));
  NOT NOT1_4361(.VSS(VSS),.VDD(VDD),.Y(I8631),.A(g4425));
  NOT NOT1_4362(.VSS(VSS),.VDD(VDD),.Y(g5899),.A(g5361));
  NOT NOT1_4363(.VSS(VSS),.VDD(VDD),.Y(g8419),.A(I13571));
  NOT NOT1_4364(.VSS(VSS),.VDD(VDD),.Y(g4958),.A(I8328));
  NOT NOT1_4365(.VSS(VSS),.VDD(VDD),.Y(g6256),.A(I10027));
  NOT NOT1_4366(.VSS(VSS),.VDD(VDD),.Y(g4176),.A(I7345));
  NOT NOT1_4367(.VSS(VSS),.VDD(VDD),.Y(g6816),.A(I10858));
  NOT NOT1_4368(.VSS(VSS),.VDD(VDD),.Y(g10122),.A(I15374));
  NOT NOT1_4369(.VSS(VSS),.VDD(VDD),.Y(g4376),.A(I7691));
  NOT NOT1_4370(.VSS(VSS),.VDD(VDD),.Y(g4005),.A(I7143));
  NOT NOT1_4371(.VSS(VSS),.VDD(VDD),.Y(g10464),.A(I15983));
  NOT NOT1_4372(.VSS(VSS),.VDD(VDD),.Y(I10027),.A(g5751));
  NOT NOT1_4373(.VSS(VSS),.VDD(VDD),.Y(I15476),.A(g10114));
  NOT NOT1_4374(.VSS(VSS),.VDD(VDD),.Y(I15485),.A(g10092));
  NOT NOT1_4375(.VSS(VSS),.VDD(VDD),.Y(g7800),.A(I12565));
  NOT NOT1_4376(.VSS(VSS),.VDD(VDD),.Y(g10034),.A(I15238));
  NOT NOT1_4377(.VSS(VSS),.VDD(VDD),.Y(g6181),.A(g5426));
  NOT NOT1_4378(.VSS(VSS),.VDD(VDD),.Y(I11804),.A(g7190));
  NOT NOT1_4379(.VSS(VSS),.VDD(VDD),.Y(I14249),.A(g8804));
  NOT NOT1_4380(.VSS(VSS),.VDD(VDD),.Y(g11454),.A(I17419));
  NOT NOT1_4381(.VSS(VSS),.VDD(VDD),.Y(g6847),.A(g6482));
  NOT NOT1_4382(.VSS(VSS),.VDD(VDD),.Y(g10292),.A(I15698));
  NOT NOT1_4383(.VSS(VSS),.VDD(VDD),.Y(I9475),.A(g5445));
  NOT NOT1_4384(.VSS(VSS),.VDD(VDD),.Y(I10248),.A(g6125));
  NOT NOT1_4385(.VSS(VSS),.VDD(VDD),.Y(g6685),.A(I10648));
  NOT NOT1_4386(.VSS(VSS),.VDD(VDD),.Y(g6197),.A(I9930));
  NOT NOT1_4387(.VSS(VSS),.VDD(VDD),.Y(g6700),.A(g5949));
  NOT NOT1_4388(.VSS(VSS),.VDD(VDD),.Y(I17112),.A(g11227));
  NOT NOT1_4389(.VSS(VSS),.VDD(VDD),.Y(I10710),.A(g6088));
  NOT NOT1_4390(.VSS(VSS),.VDD(VDD),.Y(g6397),.A(I10299));
  NOT NOT1_4391(.VSS(VSS),.VDD(VDD),.Y(I10003),.A(g4908));
  NOT NOT1_4392(.VSS(VSS),.VDD(VDD),.Y(g7213),.A(I11447));
  NOT NOT1_4393(.VSS(VSS),.VDD(VDD),.Y(I10204),.A(g6031));
  NOT NOT1_4394(.VSS(VSS),.VDD(VDD),.Y(I14552),.A(g9264));
  NOT NOT1_4395(.VSS(VSS),.VDD(VDD),.Y(I5336),.A(g1700));
  NOT NOT1_4396(.VSS(VSS),.VDD(VDD),.Y(g2131),.A(I5060));
  NOT NOT1_4397(.VSS(VSS),.VDD(VDD),.Y(g8486),.A(g8348));
  NOT NOT1_4398(.VSS(VSS),.VDD(VDD),.Y(I6784),.A(g2742));
  NOT NOT1_4399(.VSS(VSS),.VDD(VDD),.Y(g2006),.A(g932));
  NOT NOT1_4400(.VSS(VSS),.VDD(VDD),.Y(g2331),.A(g658));
  NOT NOT1_4401(.VSS(VSS),.VDD(VDD),.Y(I16577),.A(g10825));
  NOT NOT1_4402(.VSS(VSS),.VDD(VDD),.Y(g4733),.A(I8089));
  NOT NOT1_4403(.VSS(VSS),.VDD(VDD),.Y(g2406),.A(g1365));
  NOT NOT1_4404(.VSS(VSS),.VDD(VDD),.Y(g5844),.A(I9461));
  NOT NOT1_4405(.VSS(VSS),.VDD(VDD),.Y(I13332),.A(g8206));
  NOT NOT1_4406(.VSS(VSS),.VDD(VDD),.Y(g6263),.A(I10048));
  NOT NOT1_4407(.VSS(VSS),.VDD(VDD),.Y(g4270),.A(g4013));
  NOT NOT1_4408(.VSS(VSS),.VDD(VDD),.Y(I11135),.A(g6679));
  NOT NOT1_4409(.VSS(VSS),.VDD(VDD),.Y(I7372),.A(g4057));
  NOT NOT1_4410(.VSS(VSS),.VDD(VDD),.Y(g10136),.A(I15406));
  NOT NOT1_4411(.VSS(VSS),.VDD(VDD),.Y(g2635),.A(g2003));
  NOT NOT1_4412(.VSS(VSS),.VDD(VDD),.Y(I16439),.A(g10702));
  NOT NOT1_4413(.VSS(VSS),.VDD(VDD),.Y(I17742),.A(g11636));
  NOT NOT1_4414(.VSS(VSS),.VDD(VDD),.Y(I12318),.A(g6862));
  NOT NOT1_4415(.VSS(VSS),.VDD(VDD),.Y(g11074),.A(g10901));
  NOT NOT1_4416(.VSS(VSS),.VDD(VDD),.Y(g6950),.A(I11094));
  NOT NOT1_4417(.VSS(VSS),.VDD(VDD),.Y(g11239),.A(g11112));
  NOT NOT1_4418(.VSS(VSS),.VDD(VDD),.Y(I10081),.A(g5735));
  NOT NOT1_4419(.VSS(VSS),.VDD(VDD),.Y(I17096),.A(g11219));
  NOT NOT1_4420(.VSS(VSS),.VDD(VDD),.Y(g4225),.A(I7478));
  NOT NOT1_4421(.VSS(VSS),.VDD(VDD),.Y(I15238),.A(g9974));
  NOT NOT1_4422(.VSS(VSS),.VDD(VDD),.Y(g2087),.A(g225));
  NOT NOT1_4423(.VSS(VSS),.VDD(VDD),.Y(g11594),.A(I17636));
  NOT NOT1_4424(.VSS(VSS),.VDD(VDD),.Y(g3945),.A(I7096));
  NOT NOT1_4425(.VSS(VSS),.VDD(VDD),.Y(I7143),.A(g2614));
  NOT NOT1_4426(.VSS(VSS),.VDD(VDD),.Y(I5943),.A(g2233));
  NOT NOT1_4427(.VSS(VSS),.VDD(VDD),.Y(g2801),.A(g2117));
  NOT NOT1_4428(.VSS(VSS),.VDD(VDD),.Y(g5089),.A(g4840));
  NOT NOT1_4429(.VSS(VSS),.VDD(VDD),.Y(I13406),.A(g8179));
  NOT NOT1_4430(.VSS(VSS),.VDD(VDD),.Y(I9084),.A(g4886));
  NOT NOT1_4431(.VSS(VSS),.VDD(VDD),.Y(g3738),.A(g3062));
  NOT NOT1_4432(.VSS(VSS),.VDD(VDD),.Y(I13962),.A(g8451));
  NOT NOT1_4433(.VSS(VSS),.VDD(VDD),.Y(I14786),.A(g9266));
  NOT NOT1_4434(.VSS(VSS),.VDD(VDD),.Y(g7512),.A(g7148));
  NOT NOT1_4435(.VSS(VSS),.VDD(VDD),.Y(g8025),.A(I12867));
  NOT NOT1_4436(.VSS(VSS),.VDD(VDD),.Y(g9760),.A(g9454));
  NOT NOT1_4437(.VSS(VSS),.VDD(VDD),.Y(I6294),.A(g2238));
  NOT NOT1_4438(.VSS(VSS),.VDD(VDD),.Y(I17681),.A(g11608));
  NOT NOT1_4439(.VSS(VSS),.VDD(VDD),.Y(g8425),.A(I13589));
  NOT NOT1_4440(.VSS(VSS),.VDD(VDD),.Y(g3709),.A(I6870));
  NOT NOT1_4441(.VSS(VSS),.VDD(VDD),.Y(g4124),.A(I7269));
  NOT NOT1_4442(.VSS(VSS),.VDD(VDD),.Y(g4324),.A(g4144));
  NOT NOT1_4443(.VSS(VSS),.VDD(VDD),.Y(g2748),.A(I5812));
  NOT NOT1_4444(.VSS(VSS),.VDD(VDD),.Y(g6562),.A(g5774));
  NOT NOT1_4445(.VSS(VSS),.VDD(VDD),.Y(g7366),.A(I11746));
  NOT NOT1_4446(.VSS(VSS),.VDD(VDD),.Y(g10164),.A(I15488));
  NOT NOT1_4447(.VSS(VSS),.VDD(VDD),.Y(I11833),.A(g7077));
  NOT NOT1_4448(.VSS(VSS),.VDD(VDD),.Y(I11049),.A(g6635));
  NOT NOT1_4449(.VSS(VSS),.VDD(VDD),.Y(I15675),.A(g10133));
  NOT NOT1_4450(.VSS(VSS),.VDD(VDD),.Y(g4469),.A(I7840));
  NOT NOT1_4451(.VSS(VSS),.VDD(VDD),.Y(g5705),.A(I9248));
  NOT NOT1_4452(.VSS(VSS),.VDD(VDD),.Y(g5471),.A(g4370));
  NOT NOT1_4453(.VSS(VSS),.VDD(VDD),.Y(g2755),.A(I5833));
  NOT NOT1_4454(.VSS(VSS),.VDD(VDD),.Y(g11185),.A(I16956));
  NOT NOT1_4455(.VSS(VSS),.VDD(VDD),.Y(g7056),.A(I11249));
  NOT NOT1_4456(.VSS(VSS),.VDD(VDD),.Y(I17730),.A(g11638));
  NOT NOT1_4457(.VSS(VSS),.VDD(VDD),.Y(g3907),.A(I7076));
  NOT NOT1_4458(.VSS(VSS),.VDD(VDD),.Y(g10891),.A(I16635));
  NOT NOT1_4459(.VSS(VSS),.VDD(VDD),.Y(g2226),.A(g86));
  NOT NOT1_4460(.VSS(VSS),.VDD(VDD),.Y(I6501),.A(g2578));
  NOT NOT1_4461(.VSS(VSS),.VDD(VDD),.Y(I10090),.A(g5767));
  NOT NOT1_4462(.VSS(VSS),.VDD(VDD),.Y(g6723),.A(I10716));
  NOT NOT1_4463(.VSS(VSS),.VDD(VDD),.Y(I13048),.A(g8059));
  NOT NOT1_4464(.VSS(VSS),.VDD(VDD),.Y(g6257),.A(I10030));
  NOT NOT1_4465(.VSS(VSS),.VDD(VDD),.Y(I14090),.A(g8771));
  NOT NOT1_4466(.VSS(VSS),.VDD(VDD),.Y(g11518),.A(I17563));
  NOT NOT1_4467(.VSS(VSS),.VDD(VDD),.Y(g4177),.A(I7348));
  NOT NOT1_4468(.VSS(VSS),.VDD(VDD),.Y(I6156),.A(g2119));
  NOT NOT1_4469(.VSS(VSS),.VDD(VDD),.Y(g6101),.A(I9762));
  NOT NOT1_4470(.VSS(VSS),.VDD(VDD),.Y(g7148),.A(I11397));
  NOT NOT1_4471(.VSS(VSS),.VDD(VDD),.Y(g6817),.A(I10861));
  NOT NOT1_4472(.VSS(VSS),.VDD(VDD),.Y(g7649),.A(I12258));
  NOT NOT1_4473(.VSS(VSS),.VDD(VDD),.Y(g5948),.A(I9588));
  NOT NOT1_4474(.VSS(VSS),.VDD(VDD),.Y(g6301),.A(I10162));
  NOT NOT1_4475(.VSS(VSS),.VDD(VDD),.Y(g7348),.A(I11692));
  NOT NOT1_4476(.VSS(VSS),.VDD(VDD),.Y(I6356),.A(g2459));
  NOT NOT1_4477(.VSS(VSS),.VDD(VDD),.Y(g4377),.A(I7694));
  NOT NOT1_4478(.VSS(VSS),.VDD(VDD),.Y(g4206),.A(I7435));
  NOT NOT1_4479(.VSS(VSS),.VDD(VDD),.Y(I10651),.A(g6035));
  NOT NOT1_4480(.VSS(VSS),.VDD(VDD),.Y(g3517),.A(I6702));
  NOT NOT1_4481(.VSS(VSS),.VDD(VDD),.Y(g10575),.A(g10523));
  NOT NOT1_4482(.VSS(VSS),.VDD(VDD),.Y(I14182),.A(g8788));
  NOT NOT1_4483(.VSS(VSS),.VDD(VDD),.Y(I14672),.A(g9261));
  NOT NOT1_4484(.VSS(VSS),.VDD(VDD),.Y(g7355),.A(I11713));
  NOT NOT1_4485(.VSS(VSS),.VDD(VDD),.Y(g2045),.A(g1811));
  NOT NOT1_4486(.VSS(VSS),.VDD(VDD),.Y(g7851),.A(g7479));
  NOT NOT1_4487(.VSS(VSS),.VDD(VDD),.Y(I17549),.A(g11501));
  NOT NOT1_4488(.VSS(VSS),.VDD(VDD),.Y(g3876),.A(I7061));
  NOT NOT1_4489(.VSS(VSS),.VDD(VDD),.Y(g8131),.A(g8020));
  NOT NOT1_4490(.VSS(VSS),.VDD(VDD),.Y(g10327),.A(I15771));
  NOT NOT1_4491(.VSS(VSS),.VDD(VDD),.Y(g8331),.A(I13373));
  NOT NOT1_4492(.VSS(VSS),.VDD(VDD),.Y(g2173),.A(I5120));
  NOT NOT1_4493(.VSS(VSS),.VDD(VDD),.Y(I12120),.A(g7106));
  NOT NOT1_4494(.VSS(VSS),.VDD(VDD),.Y(g2373),.A(g471));
  NOT NOT1_4495(.VSS(VSS),.VDD(VDD),.Y(g4287),.A(I7546));
  NOT NOT1_4496(.VSS(VSS),.VDD(VDD),.Y(I9276),.A(g5241));
  NOT NOT1_4497(.VSS(VSS),.VDD(VDD),.Y(g10537),.A(I16178));
  NOT NOT1_4498(.VSS(VSS),.VDD(VDD),.Y(I10331),.A(g6198));
  NOT NOT1_4499(.VSS(VSS),.VDD(VDD),.Y(g7964),.A(g7651));
  NOT NOT1_4500(.VSS(VSS),.VDD(VDD),.Y(g8635),.A(I13918));
  NOT NOT1_4501(.VSS(VSS),.VDD(VDD),.Y(g6751),.A(I10762));
  NOT NOT1_4502(.VSS(VSS),.VDD(VDD),.Y(I12562),.A(g7377));
  NOT NOT1_4503(.VSS(VSS),.VDD(VDD),.Y(I8011),.A(g3820));
  NOT NOT1_4504(.VSS(VSS),.VDD(VDD),.Y(I11947),.A(g6905));
  NOT NOT1_4505(.VSS(VSS),.VDD(VDD),.Y(g8105),.A(g7992));
  NOT NOT1_4506(.VSS(VSS),.VDD(VDD),.Y(g2169),.A(g42));
  NOT NOT1_4507(.VSS(VSS),.VDD(VDD),.Y(I5395),.A(g892));
  NOT NOT1_4508(.VSS(VSS),.VDD(VDD),.Y(I14449),.A(g8973));
  NOT NOT1_4509(.VSS(VSS),.VDD(VDD),.Y(g10283),.A(g10166));
  NOT NOT1_4510(.VSS(VSS),.VDD(VDD),.Y(g2369),.A(g617));
  NOT NOT1_4511(.VSS(VSS),.VDD(VDD),.Y(I5913),.A(g2169));
  NOT NOT1_4512(.VSS(VSS),.VDD(VDD),.Y(I11106),.A(g6667));
  NOT NOT1_4513(.VSS(VSS),.VDD(VDD),.Y(g8487),.A(g8350));
  NOT NOT1_4514(.VSS(VSS),.VDD(VDD),.Y(g2602),.A(I5707));
  NOT NOT1_4515(.VSS(VSS),.VDD(VDD),.Y(I11605),.A(g6834));
  NOT NOT1_4516(.VSS(VSS),.VDD(VDD),.Y(g4199),.A(I7414));
  NOT NOT1_4517(.VSS(VSS),.VDD(VDD),.Y(g6585),.A(I10541));
  NOT NOT1_4518(.VSS(VSS),.VDD(VDD),.Y(g2007),.A(g936));
  NOT NOT1_4519(.VSS(VSS),.VDD(VDD),.Y(g5773),.A(I9359));
  NOT NOT1_4520(.VSS(VSS),.VDD(VDD),.Y(g10492),.A(I16111));
  NOT NOT1_4521(.VSS(VSS),.VDD(VDD),.Y(g4399),.A(g3638));
  NOT NOT1_4522(.VSS(VSS),.VDD(VDD),.Y(g7463),.A(g6921));
  NOT NOT1_4523(.VSS(VSS),.VDD(VDD),.Y(g2407),.A(g197));
  NOT NOT1_4524(.VSS(VSS),.VDD(VDD),.Y(I6163),.A(g2547));
  NOT NOT1_4525(.VSS(VSS),.VDD(VDD),.Y(g2920),.A(g2462));
  NOT NOT1_4526(.VSS(VSS),.VDD(VDD),.Y(I14961),.A(g9769));
  NOT NOT1_4527(.VSS(VSS),.VDD(VDD),.Y(g2578),.A(g1962));
  NOT NOT1_4528(.VSS(VSS),.VDD(VDD),.Y(g2868),.A(I6010));
  NOT NOT1_4529(.VSS(VSS),.VDD(VDD),.Y(g3214),.A(I6391));
  NOT NOT1_4530(.VSS(VSS),.VDD(VDD),.Y(g4781),.A(I8147));
  NOT NOT1_4531(.VSS(VSS),.VDD(VDD),.Y(g6041),.A(I9658));
  NOT NOT1_4532(.VSS(VSS),.VDD(VDD),.Y(I6363),.A(g2459));
  NOT NOT1_4533(.VSS(VSS),.VDD(VDD),.Y(I7202),.A(g2647));
  NOT NOT1_4534(.VSS(VSS),.VDD(VDD),.Y(I15729),.A(g10254));
  NOT NOT1_4535(.VSS(VSS),.VDD(VDD),.Y(I13812),.A(g8519));
  NOT NOT1_4536(.VSS(VSS),.VDD(VDD),.Y(I9647),.A(g5148));
  NOT NOT1_4537(.VSS(VSS),.VDD(VDD),.Y(g4898),.A(I8259));
  NOT NOT1_4538(.VSS(VSS),.VDD(VDD),.Y(g6441),.A(g6151));
  NOT NOT1_4539(.VSS(VSS),.VDD(VDD),.Y(I13463),.A(g8156));
  NOT NOT1_4540(.VSS(VSS),.VDD(VDD),.Y(g9451),.A(I14642));
  NOT NOT1_4541(.VSS(VSS),.VDD(VDD),.Y(g4900),.A(I8265));
  NOT NOT1_4542(.VSS(VSS),.VDD(VDD),.Y(I6432),.A(g2350));
  NOT NOT1_4543(.VSS(VSS),.VDD(VDD),.Y(g11501),.A(I17522));
  NOT NOT1_4544(.VSS(VSS),.VDD(VDD),.Y(g3110),.A(g2482));
  NOT NOT1_4545(.VSS(VSS),.VDD(VDD),.Y(g11577),.A(I17613));
  NOT NOT1_4546(.VSS(VSS),.VDD(VDD),.Y(g7279),.A(g6382));
  NOT NOT1_4547(.VSS(VSS),.VDD(VDD),.Y(g5836),.A(g5320));
  NOT NOT1_4548(.VSS(VSS),.VDD(VDD),.Y(g4510),.A(I7909));
  NOT NOT1_4549(.VSS(VSS),.VDD(VDD),.Y(g11439),.A(I17368));
  NOT NOT1_4550(.VSS(VSS),.VDD(VDD),.Y(g3663),.A(I6832));
  NOT NOT1_4551(.VSS(VSS),.VDD(VDD),.Y(I12427),.A(g7636));
  NOT NOT1_4552(.VSS(VSS),.VDD(VDD),.Y(g10091),.A(I15320));
  NOT NOT1_4553(.VSS(VSS),.VDD(VDD),.Y(g9346),.A(I14543));
  NOT NOT1_4554(.VSS(VSS),.VDD(VDD),.Y(I12366),.A(g7134));
  NOT NOT1_4555(.VSS(VSS),.VDD(VDD),.Y(g2261),.A(g1713));
  NOT NOT1_4556(.VSS(VSS),.VDD(VDD),.Y(g7619),.A(I12205));
  NOT NOT1_4557(.VSS(VSS),.VDD(VDD),.Y(g7318),.A(I11602));
  NOT NOT1_4558(.VSS(VSS),.VDD(VDD),.Y(g2793),.A(g2276));
  NOT NOT1_4559(.VSS(VSS),.VDD(VDD),.Y(g4291),.A(g4013));
  NOT NOT1_4560(.VSS(VSS),.VDD(VDD),.Y(g7872),.A(I12655));
  NOT NOT1_4561(.VSS(VSS),.VDD(VDD),.Y(g11438),.A(I17365));
  NOT NOT1_4562(.VSS(VSS),.VDD(VDD),.Y(g10174),.A(I15514));
  NOT NOT1_4563(.VSS(VSS),.VDD(VDD),.Y(g10796),.A(I16500));
  NOT NOT1_4564(.VSS(VSS),.VDD(VDD),.Y(I16664),.A(g10795));
  NOT NOT1_4565(.VSS(VSS),.VDD(VDD),.Y(g9103),.A(g8892));
  NOT NOT1_4566(.VSS(VSS),.VDD(VDD),.Y(I8080),.A(g3538));
  NOT NOT1_4567(.VSS(VSS),.VDD(VDD),.Y(g2015),.A(g1107));
  NOT NOT1_4568(.VSS(VSS),.VDD(VDD),.Y(g6368),.A(g5987));
  NOT NOT1_4569(.VSS(VSS),.VDD(VDD),.Y(g8445),.A(I13633));
  NOT NOT1_4570(.VSS(VSS),.VDD(VDD),.Y(I7776),.A(g3773));
  NOT NOT1_4571(.VSS(VSS),.VDD(VDD),.Y(g7057),.A(I11252));
  NOT NOT1_4572(.VSS(VSS),.VDD(VDD),.Y(g2227),.A(g95));
  NOT NOT1_4573(.VSS(VSS),.VDD(VDD),.Y(g4344),.A(g3946));
  NOT NOT1_4574(.VSS(VSS),.VDD(VDD),.Y(I5142),.A(g639));
  NOT NOT1_4575(.VSS(VSS),.VDD(VDD),.Y(I7593),.A(g4142));
  NOT NOT1_4576(.VSS(VSS),.VDD(VDD),.Y(I5248),.A(g1110));
  NOT NOT1_4577(.VSS(VSS),.VDD(VDD),.Y(g7989),.A(I12805));
  NOT NOT1_4578(.VSS(VSS),.VDD(VDD),.Y(I9224),.A(g5063));
  NOT NOT1_4579(.VSS(VSS),.VDD(VDD),.Y(I15284),.A(g10034));
  NOT NOT1_4580(.VSS(VSS),.VDD(VDD),.Y(g3762),.A(I6965));
  NOT NOT1_4581(.VSS(VSS),.VDD(VDD),.Y(I12403),.A(g7611));
  NOT NOT1_4582(.VSS(VSS),.VDD(VDD),.Y(I12547),.A(g7673));
  NOT NOT1_4583(.VSS(VSS),.VDD(VDD),.Y(g4207),.A(I7438));
  NOT NOT1_4584(.VSS(VSS),.VDD(VDD),.Y(g11083),.A(g10913));
  NOT NOT1_4585(.VSS(VSS),.VDD(VDD),.Y(g11348),.A(g11276));
  NOT NOT1_4586(.VSS(VSS),.VDD(VDD),.Y(g10390),.A(g10309));
  NOT NOT1_4587(.VSS(VSS),.VDD(VDD),.Y(I16484),.A(g10770));
  NOT NOT1_4588(.VSS(VSS),.VDD(VDD),.Y(g9732),.A(I14873));
  NOT NOT1_4589(.VSS(VSS),.VDD(VDD),.Y(I5815),.A(g1994));
  NOT NOT1_4590(.VSS(VSS),.VDD(VDD),.Y(I9120),.A(g5218));
  NOT NOT1_4591(.VSS(VSS),.VDD(VDD),.Y(g11284),.A(g11208));
  NOT NOT1_4592(.VSS(VSS),.VDD(VDD),.Y(I9320),.A(g5013));
  NOT NOT1_4593(.VSS(VSS),.VDD(VDD),.Y(g2246),.A(g1810));
  NOT NOT1_4594(.VSS(VSS),.VDD(VDD),.Y(g5822),.A(g5320));
  NOT NOT1_4595(.VSS(VSS),.VDD(VDD),.Y(g4819),.A(g3354));
  NOT NOT1_4596(.VSS(VSS),.VDD(VDD),.Y(g3877),.A(I7064));
  NOT NOT1_4597(.VSS(VSS),.VDD(VDD),.Y(g9508),.A(g9271));
  NOT NOT1_4598(.VSS(VSS),.VDD(VDD),.Y(I12226),.A(g7066));
  NOT NOT1_4599(.VSS(VSS),.VDD(VDD),.Y(g8007),.A(I12843));
  NOT NOT1_4600(.VSS(VSS),.VDD(VDD),.Y(I7264),.A(g3252));
  NOT NOT1_4601(.VSS(VSS),.VDD(VDD),.Y(g11622),.A(I17684));
  NOT NOT1_4602(.VSS(VSS),.VDD(VDD),.Y(g2203),.A(g677));
  NOT NOT1_4603(.VSS(VSS),.VDD(VDD),.Y(g7686),.A(g7148));
  NOT NOT1_4604(.VSS(VSS),.VDD(VDD),.Y(g10192),.A(I15554));
  NOT NOT1_4605(.VSS(VSS),.VDD(VDD),.Y(I10620),.A(g5884));
  NOT NOT1_4606(.VSS(VSS),.VDD(VDD),.Y(I5497),.A(g587));
  NOT NOT1_4607(.VSS(VSS),.VDD(VDD),.Y(I6929),.A(g2846));
  NOT NOT1_4608(.VSS(VSS),.VDD(VDD),.Y(I12481),.A(g7570));
  NOT NOT1_4609(.VSS(VSS),.VDD(VDD),.Y(I13421),.A(g8200));
  NOT NOT1_4610(.VSS(VSS),.VDD(VDD),.Y(I16200),.A(g10494));
  NOT NOT1_4611(.VSS(VSS),.VDD(VDD),.Y(g8868),.A(I14176));
  NOT NOT1_4612(.VSS(VSS),.VDD(VDD),.Y(I5960),.A(g2239));
  NOT NOT1_4613(.VSS(VSS),.VDD(VDD),.Y(I7360),.A(g4081));
  NOT NOT1_4614(.VSS(VSS),.VDD(VDD),.Y(I14097),.A(g8773));
  NOT NOT1_4615(.VSS(VSS),.VDD(VDD),.Y(I9617),.A(g5405));
  NOT NOT1_4616(.VSS(VSS),.VDD(VDD),.Y(g6856),.A(I10924));
  NOT NOT1_4617(.VSS(VSS),.VDD(VDD),.Y(g6411),.A(g6135));
  NOT NOT1_4618(.VSS(VSS),.VDD(VDD),.Y(g6734),.A(I10733));
  NOT NOT1_4619(.VSS(VSS),.VDD(VDD),.Y(I9789),.A(g5401));
  NOT NOT1_4620(.VSS(VSS),.VDD(VDD),.Y(I10343),.A(g6003));
  NOT NOT1_4621(.VSS(VSS),.VDD(VDD),.Y(g8535),.A(I13744));
  NOT NOT1_4622(.VSS(VSS),.VDD(VDD),.Y(I7450),.A(g3704));
  NOT NOT1_4623(.VSS(VSS),.VDD(VDD),.Y(I10971),.A(g6344));
  NOT NOT1_4624(.VSS(VSS),.VDD(VDD),.Y(g7321),.A(I11611));
  NOT NOT1_4625(.VSS(VSS),.VDD(VDD),.Y(g8582),.A(I13825));
  NOT NOT1_4626(.VSS(VSS),.VDD(VDD),.Y(g7670),.A(I12289));
  NOT NOT1_4627(.VSS(VSS),.VDD(VDD),.Y(I17261),.A(g11346));
  NOT NOT1_4628(.VSS(VSS),.VDD(VDD),.Y(g4215),.A(I7462));
  NOT NOT1_4629(.VSS(VSS),.VDD(VDD),.Y(I7996),.A(g3462));
  NOT NOT1_4630(.VSS(VSS),.VDD(VDD),.Y(g11653),.A(I17761));
  NOT NOT1_4631(.VSS(VSS),.VDD(VDD),.Y(g2502),.A(I5579));
  NOT NOT1_4632(.VSS(VSS),.VDD(VDD),.Y(g4886),.A(I8231));
  NOT NOT1_4633(.VSS(VSS),.VDD(VDD),.Y(g4951),.A(I8320));
  NOT NOT1_4634(.VSS(VSS),.VDD(VDD),.Y(I16799),.A(g11017));
  NOT NOT1_4635(.VSS(VSS),.VDD(VDD),.Y(g7232),.A(I11472));
  NOT NOT1_4636(.VSS(VSS),.VDD(VDD),.Y(I12490),.A(g7637));
  NOT NOT1_4637(.VSS(VSS),.VDD(VDD),.Y(g10553),.A(I16220));
  NOT NOT1_4638(.VSS(VSS),.VDD(VDD),.Y(g8015),.A(I12857));
  NOT NOT1_4639(.VSS(VSS),.VDD(VDD),.Y(I15415),.A(g10075));
  NOT NOT1_4640(.VSS(VSS),.VDD(VDD),.Y(g5895),.A(g5361));
  NOT NOT1_4641(.VSS(VSS),.VDD(VDD),.Y(g7938),.A(g7403));
  NOT NOT1_4642(.VSS(VSS),.VDD(VDD),.Y(I8126),.A(g3662));
  NOT NOT1_4643(.VSS(VSS),.VDD(VDD),.Y(g7813),.A(I12604));
  NOT NOT1_4644(.VSS(VSS),.VDD(VDD),.Y(I5979),.A(g2543));
  NOT NOT1_4645(.VSS(VSS),.VDD(VDD),.Y(g4314),.A(g4013));
  NOT NOT1_4646(.VSS(VSS),.VDD(VDD),.Y(I5218),.A(g1104));
  NOT NOT1_4647(.VSS(VSS),.VDD(VDD),.Y(g5062),.A(g4840));
  NOT NOT1_4648(.VSS(VSS),.VDD(VDD),.Y(I13788),.A(g8517));
  NOT NOT1_4649(.VSS(VSS),.VDD(VDD),.Y(g9347),.A(I14546));
  NOT NOT1_4650(.VSS(VSS),.VDD(VDD),.Y(I12376),.A(g7195));
  NOT NOT1_4651(.VSS(VSS),.VDD(VDD),.Y(g10326),.A(I15768));
  NOT NOT1_4652(.VSS(VSS),.VDD(VDD),.Y(g5620),.A(g4417));
  NOT NOT1_4653(.VSS(VSS),.VDD(VDD),.Y(g7909),.A(g7664));
  NOT NOT1_4654(.VSS(VSS),.VDD(VDD),.Y(g2689),.A(g2038));
  NOT NOT1_4655(.VSS(VSS),.VDD(VDD),.Y(I12103),.A(g6859));
  NOT NOT1_4656(.VSS(VSS),.VDD(VDD),.Y(I11829),.A(g7213));
  NOT NOT1_4657(.VSS(VSS),.VDD(VDD),.Y(g6863),.A(g6740));
  NOT NOT1_4658(.VSS(VSS),.VDD(VDD),.Y(I16184),.A(g10484));
  NOT NOT1_4659(.VSS(VSS),.VDD(VDD),.Y(I16805),.A(g10904));
  NOT NOT1_4660(.VSS(VSS),.VDD(VDD),.Y(g10536),.A(I16175));
  NOT NOT1_4661(.VSS(VSS),.VDD(VDD),.Y(g8664),.A(I13949));
  NOT NOT1_4662(.VSS(VSS),.VDD(VDD),.Y(g10040),.A(I15247));
  NOT NOT1_4663(.VSS(VSS),.VDD(VDD),.Y(I10412),.A(g5821));
  NOT NOT1_4664(.VSS(VSS),.VDD(VDD),.Y(I12354),.A(g7143));
  NOT NOT1_4665(.VSS(VSS),.VDD(VDD),.Y(g2216),.A(g41));
  NOT NOT1_4666(.VSS(VSS),.VDD(VDD),.Y(g9533),.A(I14684));
  NOT NOT1_4667(.VSS(VSS),.VDD(VDD),.Y(g6713),.A(I10698));
  NOT NOT1_4668(.VSS(VSS),.VDD(VDD),.Y(I14412),.A(g8939));
  NOT NOT1_4669(.VSS(VSS),.VDD(VDD),.Y(g7519),.A(g6956));
  NOT NOT1_4670(.VSS(VSS),.VDD(VDD),.Y(I13828),.A(g8488));
  NOT NOT1_4671(.VSS(VSS),.VDD(VDD),.Y(g10904),.A(I16664));
  NOT NOT1_4672(.VSS(VSS),.VDD(VDD),.Y(g2028),.A(g1703));
  NOT NOT1_4673(.VSS(VSS),.VDD(VDD),.Y(I14133),.A(g8772));
  NOT NOT1_4674(.VSS(VSS),.VDD(VDD),.Y(g10252),.A(g10137));
  NOT NOT1_4675(.VSS(VSS),.VDD(VDD),.Y(g8721),.A(g8582));
  NOT NOT1_4676(.VSS(VSS),.VDD(VDD),.Y(g6569),.A(I10499));
  NOT NOT1_4677(.VSS(VSS),.VDD(VDD),.Y(g10621),.A(I16298));
  NOT NOT1_4678(.VSS(VSS),.VDD(VDD),.Y(g7606),.A(I12168));
  NOT NOT1_4679(.VSS(VSS),.VDD(VDD),.Y(I6894),.A(g2813));
  NOT NOT1_4680(.VSS(VSS),.VDD(VDD),.Y(I13344),.A(g8121));
  NOT NOT1_4681(.VSS(VSS),.VDD(VDD),.Y(I10228),.A(g6113));
  NOT NOT1_4682(.VSS(VSS),.VDD(VDD),.Y(g2247),.A(I5258));
  NOT NOT1_4683(.VSS(VSS),.VDD(VDD),.Y(I14228),.A(g8797));
  NOT NOT1_4684(.VSS(VSS),.VDD(VDD),.Y(g4336),.A(g4130));
  NOT NOT1_4685(.VSS(VSS),.VDD(VDD),.Y(g3394),.A(I6598));
  NOT NOT1_4686(.VSS(VSS),.VDD(VDD),.Y(I5830),.A(g2067));
  NOT NOT1_4687(.VSS(VSS),.VDD(VDD),.Y(g2564),.A(g1814));
  NOT NOT1_4688(.VSS(VSS),.VDD(VDD),.Y(g7687),.A(I12318));
  NOT NOT1_4689(.VSS(VSS),.VDD(VDD),.Y(g4768),.A(I8126));
  NOT NOT1_4690(.VSS(VSS),.VDD(VDD),.Y(g11576),.A(I17610));
  NOT NOT1_4691(.VSS(VSS),.VDD(VDD),.Y(I10716),.A(g6093));
  NOT NOT1_4692(.VSS(VSS),.VDD(VDD),.Y(I13682),.A(g8310));
  NOT NOT1_4693(.VSS(VSS),.VDD(VDD),.Y(g3731),.A(I6911));
  NOT NOT1_4694(.VSS(VSS),.VDD(VDD),.Y(I15554),.A(g10088));
  NOT NOT1_4695(.VSS(VSS),.VDD(VDD),.Y(g2826),.A(g2163));
  NOT NOT1_4696(.VSS(VSS),.VDD(VDD),.Y(I6661),.A(g2752));
  NOT NOT1_4697(.VSS(VSS),.VDD(VDD),.Y(g6688),.A(I10655));
  NOT NOT1_4698(.VSS(VSS),.VDD(VDD),.Y(I11173),.A(g6500));
  NOT NOT1_4699(.VSS(VSS),.VDD(VDD),.Y(g10183),.A(g10042));
  NOT NOT1_4700(.VSS(VSS),.VDD(VDD),.Y(g6857),.A(I10927));
  NOT NOT1_4701(.VSS(VSS),.VDD(VDD),.Y(g5192),.A(g4640));
  NOT NOT1_4702(.VSS(VSS),.VDD(VDD),.Y(g5085),.A(g4377));
  NOT NOT1_4703(.VSS(VSS),.VDD(VDD),.Y(I5221),.A(g1407));
  NOT NOT1_4704(.VSS(VSS),.VDD(VDD),.Y(g9820),.A(I14961));
  NOT NOT1_4705(.VSS(VSS),.VDD(VDD),.Y(g4943),.A(I8311));
  NOT NOT1_4706(.VSS(VSS),.VDD(VDD),.Y(I12190),.A(g7268));
  NOT NOT1_4707(.VSS(VSS),.VDD(VDD),.Y(I7674),.A(g3352));
  NOT NOT1_4708(.VSS(VSS),.VDD(VDD),.Y(g11200),.A(g11112));
  NOT NOT1_4709(.VSS(VSS),.VDD(VDD),.Y(g10062),.A(I15284));
  NOT NOT1_4710(.VSS(VSS),.VDD(VDD),.Y(g3705),.A(g3113));
  NOT NOT1_4711(.VSS(VSS),.VDD(VDD),.Y(I16214),.A(g10500));
  NOT NOT1_4712(.VSS(VSS),.VDD(VDD),.Y(I17271),.A(g11388));
  NOT NOT1_4713(.VSS(VSS),.VDD(VDD),.Y(I12520),.A(g7415));
  NOT NOT1_4714(.VSS(VSS),.VDD(VDD),.Y(g2638),.A(I5751));
  NOT NOT1_4715(.VSS(VSS),.VDD(VDD),.Y(g4065),.A(g2794));
  NOT NOT1_4716(.VSS(VSS),.VDD(VDD),.Y(I8161),.A(g3637));
  NOT NOT1_4717(.VSS(VSS),.VDD(VDD),.Y(g4887),.A(I8234));
  NOT NOT1_4718(.VSS(VSS),.VDD(VDD),.Y(g4228),.A(g3914));
  NOT NOT1_4719(.VSS(VSS),.VDD(VDD),.Y(g4322),.A(I7593));
  NOT NOT1_4720(.VSS(VSS),.VDD(VDD),.Y(g7570),.A(I12032));
  NOT NOT1_4721(.VSS(VSS),.VDD(VDD),.Y(g2108),.A(I4992));
  NOT NOT1_4722(.VSS(VSS),.VDD(VDD),.Y(g5941),.A(I9571));
  NOT NOT1_4723(.VSS(VSS),.VDD(VDD),.Y(I14379),.A(g8961));
  NOT NOT1_4724(.VSS(VSS),.VDD(VDD),.Y(g2609),.A(I5728));
  NOT NOT1_4725(.VSS(VSS),.VDD(VDD),.Y(g4934),.A(g4243));
  NOT NOT1_4726(.VSS(VSS),.VDD(VDD),.Y(g7341),.A(I11671));
  NOT NOT1_4727(.VSS(VSS),.VDD(VDD),.Y(I11029),.A(g6485));
  NOT NOT1_4728(.VSS(VSS),.VDD(VDD),.Y(g10851),.A(I16553));
  NOT NOT1_4729(.VSS(VSS),.VDD(VDD),.Y(g10872),.A(I16586));
  NOT NOT1_4730(.VSS(VSS),.VDD(VDD),.Y(g11052),.A(I16817));
  NOT NOT1_4731(.VSS(VSS),.VDD(VDD),.Y(I5932),.A(g2539));
  NOT NOT1_4732(.VSS(VSS),.VDD(VDD),.Y(I10958),.A(g6559));
  NOT NOT1_4733(.VSS(VSS),.VDD(VDD),.Y(g6400),.A(I10308));
  NOT NOT1_4734(.VSS(VSS),.VDD(VDD),.Y(I14112),.A(g8777));
  NOT NOT1_4735(.VSS(VSS),.VDD(VDD),.Y(I10378),.A(g6244));
  NOT NOT1_4736(.VSS(VSS),.VDD(VDD),.Y(g7525),.A(I11921));
  NOT NOT1_4737(.VSS(VSS),.VDD(VDD),.Y(I7680),.A(g3736));
  NOT NOT1_4738(.VSS(VSS),.VDD(VDD),.Y(I14958),.A(g9767));
  NOT NOT1_4739(.VSS(VSS),.VDD(VDD),.Y(g2883),.A(I6037));
  NOT NOT1_4740(.VSS(VSS),.VDD(VDD),.Y(g8671),.A(I13956));
  NOT NOT1_4741(.VSS(VSS),.VDD(VDD),.Y(I6484),.A(g2073));
  NOT NOT1_4742(.VSS(VSS),.VDD(VDD),.Y(I6439),.A(g2352));
  NOT NOT1_4743(.VSS(VSS),.VDD(VDD),.Y(I9915),.A(g5304));
  NOT NOT1_4744(.VSS(VSS),.VDD(VDD),.Y(g3254),.A(g2322));
  NOT NOT1_4745(.VSS(VSS),.VDD(VDD),.Y(g9775),.A(g9474));
  NOT NOT1_4746(.VSS(VSS),.VDD(VDD),.Y(I17736),.A(g11640));
  NOT NOT1_4747(.VSS(VSS),.VDD(VDD),.Y(I15798),.A(g10281));
  NOT NOT1_4748(.VSS(VSS),.VDD(VDD),.Y(g3814),.A(g3228));
  NOT NOT1_4749(.VSS(VSS),.VDD(VDD),.Y(g5708),.A(I9253));
  NOT NOT1_4750(.VSS(VSS),.VDD(VDD),.Y(I10096),.A(g5794));
  NOT NOT1_4751(.VSS(VSS),.VDD(VDD),.Y(g2217),.A(I5192));
  NOT NOT1_4752(.VSS(VSS),.VDD(VDD),.Y(g2758),.A(I5840));
  NOT NOT1_4753(.VSS(VSS),.VDD(VDD),.Y(g5520),.A(I8943));
  NOT NOT1_4754(.VSS(VSS),.VDD(VDD),.Y(I14944),.A(g9454));
  NOT NOT1_4755(.VSS(VSS),.VDD(VDD),.Y(I17198),.A(g11319));
  NOT NOT1_4756(.VSS(VSS),.VDD(VDD),.Y(I15184),.A(g9974));
  NOT NOT1_4757(.VSS(VSS),.VDD(VDD),.Y(g4096),.A(I7236));
  NOT NOT1_4758(.VSS(VSS),.VDD(VDD),.Y(g8564),.A(I13785));
  NOT NOT1_4759(.VSS(VSS),.VDD(VDD),.Y(g3038),.A(g1982));
  NOT NOT1_4760(.VSS(VSS),.VDD(VDD),.Y(g4496),.A(I7889));
  NOT NOT1_4761(.VSS(VSS),.VDD(VDD),.Y(I8303),.A(g4784));
  NOT NOT1_4762(.VSS(VSS),.VDD(VDD),.Y(g11184),.A(I16953));
  NOT NOT1_4763(.VSS(VSS),.VDD(VDD),.Y(g5252),.A(g4640));
  NOT NOT1_4764(.VSS(VSS),.VDD(VDD),.Y(g7607),.A(I12171));
  NOT NOT1_4765(.VSS(VSS),.VDD(VDD),.Y(I17528),.A(g11487));
  NOT NOT1_4766(.VSS(VSS),.VDD(VDD),.Y(I6702),.A(g2801));
  NOT NOT1_4767(.VSS(VSS),.VDD(VDD),.Y(g3773),.A(I6996));
  NOT NOT1_4768(.VSS(VSS),.VDD(VDD),.Y(g5812),.A(g5320));
  NOT NOT1_4769(.VSS(VSS),.VDD(VDD),.Y(g3009),.A(g2135));
  NOT NOT1_4770(.VSS(VSS),.VDD(VDD),.Y(I14681),.A(g9110));
  NOT NOT1_4771(.VSS(VSS),.VDD(VDD),.Y(g2165),.A(I5098));
  NOT NOT1_4772(.VSS(VSS),.VDD(VDD),.Y(g6183),.A(g5320));
  NOT NOT1_4773(.VSS(VSS),.VDD(VDD),.Y(g2571),.A(g1822));
  NOT NOT1_4774(.VSS(VSS),.VDD(VDD),.Y(g7659),.A(I12274));
  NOT NOT1_4775(.VSS(VSS),.VDD(VDD),.Y(g2861),.A(I6001));
  NOT NOT1_4776(.VSS(VSS),.VDD(VDD),.Y(g7358),.A(I11722));
  NOT NOT1_4777(.VSS(VSS),.VDD(VDD),.Y(g4195),.A(I7402));
  NOT NOT1_4778(.VSS(VSS),.VDD(VDD),.Y(g5176),.A(g4682));
  NOT NOT1_4779(.VSS(VSS),.VDD(VDD),.Y(g6220),.A(g5446));
  NOT NOT1_4780(.VSS(VSS),.VDD(VDD),.Y(I5716),.A(g2068));
  NOT NOT1_4781(.VSS(VSS),.VDD(VDD),.Y(g10574),.A(I16239));
  NOT NOT1_4782(.VSS(VSS),.VDD(VDD),.Y(I17764),.A(g11651));
  NOT NOT1_4783(.VSS(VSS),.VDD(VDD),.Y(I5149),.A(g1453));
  NOT NOT1_4784(.VSS(VSS),.VDD(VDD),.Y(g4395),.A(I7732));
  NOT NOT1_4785(.VSS(VSS),.VDD(VDD),.Y(g10047),.A(I15266));
  NOT NOT1_4786(.VSS(VSS),.VDD(VDD),.Y(g4337),.A(g4144));
  NOT NOT1_4787(.VSS(VSS),.VDD(VDD),.Y(g4913),.A(I8285));
  NOT NOT1_4788(.VSS(VSS),.VDD(VDD),.Y(I17365),.A(g11380));
  NOT NOT1_4789(.VSS(VSS),.VDD(VDD),.Y(I14802),.A(g9666));
  NOT NOT1_4790(.VSS(VSS),.VDD(VDD),.Y(g10205),.A(g10176));
  NOT NOT1_4791(.VSS(VSS),.VDD(VDD),.Y(g2055),.A(g1950));
  NOT NOT1_4792(.VSS(VSS),.VDD(VDD),.Y(g3769),.A(I6982));
  NOT NOT1_4793(.VSS(VSS),.VDD(VDD),.Y(g10912),.A(I16688));
  NOT NOT1_4794(.VSS(VSS),.VDD(VDD),.Y(g10311),.A(g10242));
  NOT NOT1_4795(.VSS(VSS),.VDD(VDD),.Y(g2455),.A(g826));
  NOT NOT1_4796(.VSS(VSS),.VDD(VDD),.Y(g9739),.A(I14884));
  NOT NOT1_4797(.VSS(VSS),.VDD(VDD),.Y(g2827),.A(g2164));
  NOT NOT1_4798(.VSS(VSS),.VDD(VDD),.Y(I6952),.A(g2867));
  NOT NOT1_4799(.VSS(VSS),.VDD(VDD),.Y(I14793),.A(g9269));
  NOT NOT1_4800(.VSS(VSS),.VDD(VDD),.Y(g3212),.A(I6385));
  NOT NOT1_4801(.VSS(VSS),.VDD(VDD),.Y(I9402),.A(g5107));
  NOT NOT1_4802(.VSS(VSS),.VDD(VDD),.Y(I12339),.A(g7054));
  NOT NOT1_4803(.VSS(VSS),.VDD(VDD),.Y(I8240),.A(g4380));
  NOT NOT1_4804(.VSS(VSS),.VDD(VDD),.Y(g1975),.A(g622));
  NOT NOT1_4805(.VSS(VSS),.VDD(VDD),.Y(I5198),.A(g143));
  NOT NOT1_4806(.VSS(VSS),.VDD(VDD),.Y(I12296),.A(g7236));
  NOT NOT1_4807(.VSS(VSS),.VDD(VDD),.Y(g7311),.A(I11581));
  NOT NOT1_4808(.VSS(VSS),.VDD(VDD),.Y(g2774),.A(g2276));
  NOT NOT1_4809(.VSS(VSS),.VDD(VDD),.Y(I6616),.A(g3186));
  NOT NOT1_4810(.VSS(VSS),.VDD(VDD),.Y(g3967),.A(g3247));
  NOT NOT1_4811(.VSS(VSS),.VDD(VDD),.Y(I17161),.A(g11314));
  NOT NOT1_4812(.VSS(VSS),.VDD(VDD),.Y(g6588),.A(I10546));
  NOT NOT1_4813(.VSS(VSS),.VDD(VDD),.Y(I4935),.A(g585));
  NOT NOT1_4814(.VSS(VSS),.VDD(VDD),.Y(I12644),.A(g7729));
  NOT NOT1_4815(.VSS(VSS),.VDD(VDD),.Y(g2846),.A(I5970));
  NOT NOT1_4816(.VSS(VSS),.VDD(VDD),.Y(I9762),.A(g5276));
  NOT NOT1_4817(.VSS(VSS),.VDD(VDD),.Y(I10549),.A(g6184));
  NOT NOT1_4818(.VSS(VSS),.VDD(VDD),.Y(g9079),.A(g8892));
  NOT NOT1_4819(.VSS(VSS),.VDD(VDD),.Y(I13648),.A(g8376));
  NOT NOT1_4820(.VSS(VSS),.VDD(VDD),.Y(g10051),.A(I15272));
  NOT NOT1_4821(.VSS(VSS),.VDD(VDD),.Y(I14690),.A(g9150));
  NOT NOT1_4822(.VSS(VSS),.VDD(VDD),.Y(g6161),.A(I9886));
  NOT NOT1_4823(.VSS(VSS),.VDD(VDD),.Y(I14549),.A(g9262));
  NOT NOT1_4824(.VSS(VSS),.VDD(VDD),.Y(g7615),.A(I12193));
  NOT NOT1_4825(.VSS(VSS),.VDD(VDD),.Y(g6361),.A(g5867));
  NOT NOT1_4826(.VSS(VSS),.VDD(VDD),.Y(g2196),.A(g91));
  NOT NOT1_4827(.VSS(VSS),.VDD(VDD),.Y(g4266),.A(g3688));
  NOT NOT1_4828(.VSS(VSS),.VDD(VDD),.Y(I7600),.A(g4159));
  NOT NOT1_4829(.VSS(VSS),.VDD(VDD),.Y(g9668),.A(g9490));
  NOT NOT1_4830(.VSS(VSS),.VDD(VDD),.Y(g2396),.A(g1389));
  NOT NOT1_4831(.VSS(VSS),.VDD(VDD),.Y(g10592),.A(I16261));
  NOT NOT1_4832(.VSS(VSS),.VDD(VDD),.Y(I15400),.A(g10069));
  NOT NOT1_4833(.VSS(VSS),.VDD(VDD),.Y(g2803),.A(g2154));
  NOT NOT1_4834(.VSS(VSS),.VDD(VDD),.Y(g5733),.A(I9287));
  NOT NOT1_4835(.VSS(VSS),.VDD(VDD),.Y(I17225),.A(g11298));
  NOT NOT1_4836(.VSS(VSS),.VDD(VDD),.Y(g11400),.A(I17243));
  NOT NOT1_4837(.VSS(VSS),.VDD(VDD),.Y(g6051),.A(I9680));
  NOT NOT1_4838(.VSS(VSS),.VDD(VDD),.Y(I11770),.A(g7202));
  NOT NOT1_4839(.VSS(VSS),.VDD(VDD),.Y(g5270),.A(g4367));
  NOT NOT1_4840(.VSS(VSS),.VDD(VDD),.Y(g7374),.A(I11752));
  NOT NOT1_4841(.VSS(VSS),.VDD(VDD),.Y(I11563),.A(g6819));
  NOT NOT1_4842(.VSS(VSS),.VDD(VDD),.Y(I8116),.A(g3627));
  NOT NOT1_4843(.VSS(VSS),.VDD(VDD),.Y(g6127),.A(I9826));
  NOT NOT1_4844(.VSS(VSS),.VDD(VDD),.Y(g6451),.A(I10381));
  NOT NOT1_4845(.VSS(VSS),.VDD(VDD),.Y(g8758),.A(I14055));
  NOT NOT1_4846(.VSS(VSS),.VDD(VDD),.Y(g8066),.A(I12916));
  NOT NOT1_4847(.VSS(VSS),.VDD(VDD),.Y(g8589),.A(I13834));
  NOT NOT1_4848(.VSS(VSS),.VDD(VDD),.Y(I15329),.A(g9995));
  NOT NOT1_4849(.VSS(VSS),.VDD(VDD),.Y(g7985),.A(I12799));
  NOT NOT1_4850(.VSS(VSS),.VDD(VDD),.Y(I17258),.A(g11345));
  NOT NOT1_4851(.VSS(VSS),.VDD(VDD),.Y(g4142),.A(I7288));
  NOT NOT1_4852(.VSS(VSS),.VDD(VDD),.Y(g2509),.A(I5588));
  NOT NOT1_4853(.VSS(VSS),.VDD(VDD),.Y(I16407),.A(g10696));
  NOT NOT1_4854(.VSS(VSS),.VDD(VDD),.Y(I15539),.A(g10069));
  NOT NOT1_4855(.VSS(VSS),.VDD(VDD),.Y(I6546),.A(g2987));
  NOT NOT1_4856(.VSS(VSS),.VDD(VDD),.Y(g5073),.A(g4840));
  NOT NOT1_4857(.VSS(VSS),.VDD(VDD),.Y(g10350),.A(I15814));
  NOT NOT1_4858(.VSS(VSS),.VDD(VDD),.Y(g11207),.A(I16982));
  NOT NOT1_4859(.VSS(VSS),.VDD(VDD),.Y(g1984),.A(g758));
  NOT NOT1_4860(.VSS(VSS),.VDD(VDD),.Y(I10317),.A(g6003));
  NOT NOT1_4861(.VSS(VSS),.VDD(VDD),.Y(g7284),.A(I11528));
  NOT NOT1_4862(.VSS(VSS),.VDD(VDD),.Y(g11539),.A(g11519));
  NOT NOT1_4863(.VSS(VSS),.VDD(VDD),.Y(g6146),.A(I9863));
  NOT NOT1_4864(.VSS(VSS),.VDD(VDD),.Y(g10820),.A(I16528));
  NOT NOT1_4865(.VSS(VSS),.VDD(VDD),.Y(g4081),.A(I7210));
  NOT NOT1_4866(.VSS(VSS),.VDD(VDD),.Y(g7545),.A(I11967));
  NOT NOT1_4867(.VSS(VSS),.VDD(VDD),.Y(g9356),.A(I14573));
  NOT NOT1_4868(.VSS(VSS),.VDD(VDD),.Y(g8571),.A(I13806));
  NOT NOT1_4869(.VSS(VSS),.VDD(VDD),.Y(I8147),.A(g3633));
  NOT NOT1_4870(.VSS(VSS),.VDD(VDD),.Y(g2662),.A(g2014));
  NOT NOT1_4871(.VSS(VSS),.VDD(VDD),.Y(g5124),.A(g4596));
  NOT NOT1_4872(.VSS(VSS),.VDD(VDD),.Y(g2018),.A(g1336));
  NOT NOT1_4873(.VSS(VSS),.VDD(VDD),.Y(g5980),.A(I9594));
  NOT NOT1_4874(.VSS(VSS),.VDD(VDD),.Y(g2067),.A(g108));
  NOT NOT1_4875(.VSS(VSS),.VDD(VDD),.Y(g7380),.A(g7279));
  NOT NOT1_4876(.VSS(VSS),.VDD(VDD),.Y(g8448),.A(I13642));
  NOT NOT1_4877(.VSS(VSS),.VDD(VDD),.Y(g6103),.A(I9766));
  NOT NOT1_4878(.VSS(VSS),.VDD(VDD),.Y(I10129),.A(g5688));
  NOT NOT1_4879(.VSS(VSS),.VDD(VDD),.Y(I9930),.A(g5317));
  NOT NOT1_4880(.VSS(VSS),.VDD(VDD),.Y(I11767),.A(g7201));
  NOT NOT1_4881(.VSS(VSS),.VDD(VDD),.Y(I11794),.A(g7188));
  NOT NOT1_4882(.VSS(VSS),.VDD(VDD),.Y(g8711),.A(g8677));
  NOT NOT1_4883(.VSS(VSS),.VDD(VDD),.Y(g7591),.A(I12103));
  NOT NOT1_4884(.VSS(VSS),.VDD(VDD),.Y(g6303),.A(I10168));
  NOT NOT1_4885(.VSS(VSS),.VDD(VDD),.Y(g2418),.A(I5497));
  NOT NOT1_4886(.VSS(VSS),.VDD(VDD),.Y(I11845),.A(g6869));
  NOT NOT1_4887(.VSS(VSS),.VDD(VDD),.Y(g5069),.A(g4368));
  NOT NOT1_4888(.VSS(VSS),.VDD(VDD),.Y(I13794),.A(g8472));
  NOT NOT1_4889(.VSS(VSS),.VDD(VDD),.Y(I10057),.A(g5741));
  NOT NOT1_4890(.VSS(VSS),.VDD(VDD),.Y(g4726),.A(g3546));
  NOT NOT1_4891(.VSS(VSS),.VDD(VDD),.Y(g2994),.A(g2057));
  NOT NOT1_4892(.VSS(VSS),.VDD(VDD),.Y(g5469),.A(I8880));
  NOT NOT1_4893(.VSS(VSS),.VDD(VDD),.Y(g7853),.A(I12652));
  NOT NOT1_4894(.VSS(VSS),.VDD(VDD),.Y(g4354),.A(I7639));
  NOT NOT1_4895(.VSS(VSS),.VDD(VDD),.Y(I5258),.A(g67));
  NOT NOT1_4896(.VSS(VSS),.VDD(VDD),.Y(g7020),.A(I11159));
  NOT NOT1_4897(.VSS(VSS),.VDD(VDD),.Y(I5818),.A(g2098));
  NOT NOT1_4898(.VSS(VSS),.VDD(VDD),.Y(g8133),.A(I13002));
  NOT NOT1_4899(.VSS(VSS),.VDD(VDD),.Y(g8333),.A(I13379));
  NOT NOT1_4900(.VSS(VSS),.VDD(VDD),.Y(g7420),.A(I11804));
  NOT NOT1_4901(.VSS(VSS),.VDD(VDD),.Y(I15241),.A(g10013));
  NOT NOT1_4902(.VSS(VSS),.VDD(VDD),.Y(I11898),.A(g6896));
  NOT NOT1_4903(.VSS(VSS),.VDD(VDD),.Y(g5177),.A(g4596));
  NOT NOT1_4904(.VSS(VSS),.VDD(VDD),.Y(g6732),.A(I10729));
  NOT NOT1_4905(.VSS(VSS),.VDD(VDD),.Y(I12867),.A(g7638));
  NOT NOT1_4906(.VSS(VSS),.VDD(VDD),.Y(I17657),.A(g11598));
  NOT NOT1_4907(.VSS(VSS),.VDD(VDD),.Y(I13633),.A(g8346));
  NOT NOT1_4908(.VSS(VSS),.VDD(VDD),.Y(g11241),.A(g11112));
  NOT NOT1_4909(.VSS(VSS),.VDD(VDD),.Y(I16206),.A(g10453));
  NOT NOT1_4910(.VSS(VSS),.VDD(VDD),.Y(I10299),.A(g6243));
  NOT NOT1_4911(.VSS(VSS),.VDD(VDD),.Y(g2256),.A(I5279));
  NOT NOT1_4912(.VSS(VSS),.VDD(VDD),.Y(I11191),.A(g6514));
  NOT NOT1_4913(.VSS(VSS),.VDD(VDD),.Y(I11719),.A(g7029));
  NOT NOT1_4914(.VSS(VSS),.VDD(VDD),.Y(g7559),.A(I12009));
  NOT NOT1_4915(.VSS(VSS),.VDD(VDD),.Y(I14323),.A(g8817));
  NOT NOT1_4916(.VSS(VSS),.VDD(VDD),.Y(g10691),.A(I16360));
  NOT NOT1_4917(.VSS(VSS),.VDD(VDD),.Y(g7794),.A(I12547));
  NOT NOT1_4918(.VSS(VSS),.VDD(VDD),.Y(I7076),.A(g2985));
  NOT NOT1_4919(.VSS(VSS),.VDD(VDD),.Y(I13191),.A(g8132));
  NOT NOT1_4920(.VSS(VSS),.VDD(VDD),.Y(I14299),.A(g8810));
  NOT NOT1_4921(.VSS(VSS),.VDD(VDD),.Y(I7889),.A(g3373));
  NOT NOT1_4922(.VSS(VSS),.VDD(VDD),.Y(g8196),.A(I13125));
  NOT NOT1_4923(.VSS(VSS),.VDD(VDD),.Y(g6944),.A(I11082));
  NOT NOT1_4924(.VSS(VSS),.VDD(VDD),.Y(g8803),.A(I14130));
  NOT NOT1_4925(.VSS(VSS),.VDD(VDD),.Y(I6277),.A(g1206));
  NOT NOT1_4926(.VSS(VSS),.VDD(VDD),.Y(g6072),.A(g4977));
  NOT NOT1_4927(.VSS(VSS),.VDD(VDD),.Y(I15771),.A(g10250));
  NOT NOT1_4928(.VSS(VSS),.VDD(VDD),.Y(I9237),.A(g5205));
  NOT NOT1_4929(.VSS(VSS),.VDD(VDD),.Y(I17337),.A(g11363));
  NOT NOT1_4930(.VSS(VSS),.VDD(VDD),.Y(g2181),.A(I5142));
  NOT NOT1_4931(.VSS(VSS),.VDD(VDD),.Y(g8538),.A(I13747));
  NOT NOT1_4932(.VSS(VSS),.VDD(VDD),.Y(g2381),.A(g1368));
  NOT NOT1_4933(.VSS(VSS),.VDD(VDD),.Y(g9432),.A(g9313));
  NOT NOT1_4934(.VSS(VSS),.VDD(VDD),.Y(I15235),.A(g9968));
  NOT NOT1_4935(.VSS(VSS),.VDD(VDD),.Y(I6789),.A(g2748));
  NOT NOT1_4936(.VSS(VSS),.VDD(VDD),.Y(I16114),.A(g10387));
  NOT NOT1_4937(.VSS(VSS),.VDD(VDD),.Y(g4783),.A(g3829));
  NOT NOT1_4938(.VSS(VSS),.VDD(VDD),.Y(g6043),.A(I9662));
  NOT NOT1_4939(.VSS(VSS),.VDD(VDD),.Y(I12910),.A(g7922));
  NOT NOT1_4940(.VSS(VSS),.VDD(VDD),.Y(I7375),.A(g4062));
  NOT NOT1_4941(.VSS(VSS),.VDD(VDD),.Y(g2847),.A(I5973));
  NOT NOT1_4942(.VSS(VSS),.VDD(VDD),.Y(g8780),.A(I14077));
  NOT NOT1_4943(.VSS(VSS),.VDD(VDD),.Y(g6443),.A(g6157));
  NOT NOT1_4944(.VSS(VSS),.VDD(VDD),.Y(I12202),.A(g6983));
  NOT NOT1_4945(.VSS(VSS),.VDD(VDD),.Y(g8509),.A(g8366));
  NOT NOT1_4946(.VSS(VSS),.VDD(VDD),.Y(g9453),.A(g9100));
  NOT NOT1_4947(.VSS(VSS),.VDD(VDD),.Y(g4112),.A(g2994));
  NOT NOT1_4948(.VSS(VSS),.VDD(VDD),.Y(g7905),.A(g7450));
  NOT NOT1_4949(.VSS(VSS),.VDD(VDD),.Y(g2197),.A(g101));
  NOT NOT1_4950(.VSS(VSS),.VDD(VDD),.Y(I7651),.A(g3332));
  NOT NOT1_4951(.VSS(VSS),.VDD(VDD),.Y(g4312),.A(g4144));
  NOT NOT1_4952(.VSS(VSS),.VDD(VDD),.Y(I8820),.A(g4473));
  NOT NOT1_4953(.VSS(VSS),.VDD(VDD),.Y(I11440),.A(g6577));
  NOT NOT1_4954(.VSS(VSS),.VDD(VDD),.Y(g10929),.A(g10827));
  NOT NOT1_4955(.VSS(VSS),.VDD(VDD),.Y(I12496),.A(g7724));
  NOT NOT1_4956(.VSS(VSS),.VDD(VDD),.Y(g2021),.A(g1341));
  NOT NOT1_4957(.VSS(VSS),.VDD(VDD),.Y(I9194),.A(g5236));
  NOT NOT1_4958(.VSS(VSS),.VDD(VDD),.Y(g7628),.A(I12226));
  NOT NOT1_4959(.VSS(VSS),.VDD(VDD),.Y(I9394),.A(g5195));
  NOT NOT1_4960(.VSS(VSS),.VDD(VDD),.Y(g6116),.A(I9801));
  NOT NOT1_4961(.VSS(VSS),.VDD(VDD),.Y(g2421),.A(g1374));
  NOT NOT1_4962(.VSS(VSS),.VDD(VDD),.Y(g7630),.A(I12232));
  NOT NOT1_4963(.VSS(VSS),.VDD(VDD),.Y(g4001),.A(g3200));
  NOT NOT1_4964(.VSS(VSS),.VDD(VDD),.Y(I12978),.A(g8040));
  NOT NOT1_4965(.VSS(VSS),.VDD(VDD),.Y(I14232),.A(g8800));
  NOT NOT1_4966(.VSS(VSS),.VDD(VDD),.Y(g10928),.A(g10827));
  NOT NOT1_4967(.VSS(VSS),.VDD(VDD),.Y(g8067),.A(I12919));
  NOT NOT1_4968(.VSS(VSS),.VDD(VDD),.Y(I9731),.A(g5255));
  NOT NOT1_4969(.VSS(VSS),.VDD(VDD),.Y(g5898),.A(g5361));
  NOT NOT1_4970(.VSS(VSS),.VDD(VDD),.Y(g8418),.A(I13568));
  NOT NOT1_4971(.VSS(VSS),.VDD(VDD),.Y(g6434),.A(I10352));
  NOT NOT1_4972(.VSS(VSS),.VDD(VDD),.Y(g4676),.A(g3354));
  NOT NOT1_4973(.VSS(VSS),.VDD(VDD),.Y(g5900),.A(I9531));
  NOT NOT1_4974(.VSS(VSS),.VDD(VDD),.Y(g6565),.A(g5790));
  NOT NOT1_4975(.VSS(VSS),.VDD(VDD),.Y(I5821),.A(g2101));
  NOT NOT1_4976(.VSS(VSS),.VDD(VDD),.Y(I6299),.A(g2242));
  NOT NOT1_4977(.VSS(VSS),.VDD(VDD),.Y(I11926),.A(g6900));
  NOT NOT1_4978(.VSS(VSS),.VDD(VDD),.Y(g8290),.A(I13224));
  NOT NOT1_4979(.VSS(VSS),.VDD(VDD),.Y(I12986),.A(g8042));
  NOT NOT1_4980(.VSS(VSS),.VDD(VDD),.Y(g4129),.A(I7280));
  NOT NOT1_4981(.VSS(VSS),.VDD(VDD),.Y(g5797),.A(I9399));
  NOT NOT1_4982(.VSS(VSS),.VDD(VDD),.Y(g4329),.A(g4144));
  NOT NOT1_4983(.VSS(VSS),.VDD(VDD),.Y(I14697),.A(g9260));
  NOT NOT1_4984(.VSS(VSS),.VDD(VDD),.Y(g4761),.A(g3440));
  NOT NOT1_4985(.VSS(VSS),.VDD(VDD),.Y(g11515),.A(g11490));
  NOT NOT1_4986(.VSS(VSS),.VDD(VDD),.Y(I7384),.A(g4082));
  NOT NOT1_4987(.VSS(VSS),.VDD(VDD),.Y(I13612),.A(g8325));
  NOT NOT1_4988(.VSS(VSS),.VDD(VDD),.Y(g5245),.A(g4369));
  NOT NOT1_4989(.VSS(VSS),.VDD(VDD),.Y(I7339),.A(g4004));
  NOT NOT1_4990(.VSS(VSS),.VDD(VDD),.Y(I13099),.A(g7927));
  NOT NOT1_4991(.VSS(VSS),.VDD(VDD),.Y(I12384),.A(g7212));
  NOT NOT1_4992(.VSS(VSS),.VDD(VDD),.Y(g8093),.A(I12948));
  NOT NOT1_4993(.VSS(VSS),.VDD(VDD),.Y(I13388),.A(g8230));
  NOT NOT1_4994(.VSS(VSS),.VDD(VDD),.Y(g6681),.A(g5830));
  NOT NOT1_4995(.VSS(VSS),.VDD(VDD),.Y(I11701),.A(g7065));
  NOT NOT1_4996(.VSS(VSS),.VDD(VDD),.Y(I11534),.A(g6917));
  NOT NOT1_4997(.VSS(VSS),.VDD(VDD),.Y(g10787),.A(I16487));
  NOT NOT1_4998(.VSS(VSS),.VDD(VDD),.Y(g5291),.A(g4384));
  NOT NOT1_4999(.VSS(VSS),.VDD(VDD),.Y(g3392),.A(g3121));
  NOT NOT1_5000(.VSS(VSS),.VDD(VDD),.Y(I11272),.A(g6546));
  NOT NOT1_5001(.VSS(VSS),.VDD(VDD),.Y(g10282),.A(g10164));
  NOT NOT1_5002(.VSS(VSS),.VDD(VDD),.Y(g7750),.A(I12415));
  NOT NOT1_5003(.VSS(VSS),.VDD(VDD),.Y(g3485),.A(g2662));
  NOT NOT1_5004(.VSS(VSS),.VDD(VDD),.Y(g2562),.A(g1383));
  NOT NOT1_5005(.VSS(VSS),.VDD(VDD),.Y(g6697),.A(g5949));
  NOT NOT1_5006(.VSS(VSS),.VDD(VDD),.Y(g5144),.A(g4682));
  NOT NOT1_5007(.VSS(VSS),.VDD(VDD),.Y(g4592),.A(g3829));
  NOT NOT1_5008(.VSS(VSS),.VDD(VDD),.Y(g6914),.A(I11024));
  NOT NOT1_5009(.VSS(VSS),.VDD(VDD),.Y(I17444),.A(g11446));
  NOT NOT1_5010(.VSS(VSS),.VDD(VDD),.Y(g5344),.A(I8811));
  NOT NOT1_5011(.VSS(VSS),.VDD(VDD),.Y(g6210),.A(g5205));
  NOT NOT1_5012(.VSS(VSS),.VDD(VDD),.Y(I12150),.A(g7074));
  NOT NOT1_5013(.VSS(VSS),.VDD(VDD),.Y(g4746),.A(I8098));
  NOT NOT1_5014(.VSS(VSS),.VDD(VDD),.Y(g8181),.A(I13096));
  NOT NOT1_5015(.VSS(VSS),.VDD(VDD),.Y(g10827),.A(I16543));
  NOT NOT1_5016(.VSS(VSS),.VDD(VDD),.Y(g6596),.A(I10566));
  NOT NOT1_5017(.VSS(VSS),.VDD(VDD),.Y(I6738),.A(g3113));
  NOT NOT1_5018(.VSS(VSS),.VDD(VDD),.Y(g4221),.A(g3914));
  NOT NOT1_5019(.VSS(VSS),.VDD(VDD),.Y(g8381),.A(I13489));
  NOT NOT1_5020(.VSS(VSS),.VDD(VDD),.Y(g2101),.A(I4951));
  NOT NOT1_5021(.VSS(VSS),.VDD(VDD),.Y(g2817),.A(I5919));
  NOT NOT1_5022(.VSS(VSS),.VDD(VDD),.Y(g3941),.A(g3015));
  NOT NOT1_5023(.VSS(VSS),.VDD(VDD),.Y(g7040),.A(I11207));
  NOT NOT1_5024(.VSS(VSS),.VDD(VDD),.Y(g6413),.A(I10325));
  NOT NOT1_5025(.VSS(VSS),.VDD(VDD),.Y(I10831),.A(g6710));
  NOT NOT1_5026(.VSS(VSS),.VDD(VDD),.Y(g7440),.A(I11836));
  NOT NOT1_5027(.VSS(VSS),.VDD(VDD),.Y(g8197),.A(I13128));
  NOT NOT1_5028(.VSS(VSS),.VDD(VDD),.Y(g8700),.A(g8574));
  NOT NOT1_5029(.VSS(VSS),.VDD(VDD),.Y(I10445),.A(g5770));
  NOT NOT1_5030(.VSS(VSS),.VDD(VDD),.Y(I7523),.A(g4095));
  NOT NOT1_5031(.VSS(VSS),.VDD(VDD),.Y(I11140),.A(g6448));
  NOT NOT1_5032(.VSS(VSS),.VDD(VDD),.Y(I12196),.A(g7272));
  NOT NOT1_5033(.VSS(VSS),.VDD(VDD),.Y(g2605),.A(I5716));
  NOT NOT1_5034(.VSS(VSS),.VDD(VDD),.Y(g11441),.A(I17374));
  NOT NOT1_5035(.VSS(VSS),.VDD(VDD),.Y(I9150),.A(g5012));
  NOT NOT1_5036(.VSS(VSS),.VDD(VDD),.Y(I10499),.A(g6149));
  NOT NOT1_5037(.VSS(VSS),.VDD(VDD),.Y(g8421),.A(I13577));
  NOT NOT1_5038(.VSS(VSS),.VDD(VDD),.Y(g7123),.A(I11360));
  NOT NOT1_5039(.VSS(VSS),.VDD(VDD),.Y(g5088),.A(I8456));
  NOT NOT1_5040(.VSS(VSS),.VDD(VDD),.Y(g11206),.A(I16979));
  NOT NOT1_5041(.VSS(VSS),.VDD(VDD),.Y(g7323),.A(I11617));
  NOT NOT1_5042(.VSS(VSS),.VDD(VDD),.Y(I14499),.A(g8889));
  NOT NOT1_5043(.VSS(VSS),.VDD(VDD),.Y(I6907),.A(g2994));
  NOT NOT1_5044(.VSS(VSS),.VDD(VDD),.Y(I12526),.A(g7648));
  NOT NOT1_5045(.VSS(VSS),.VDD(VDD),.Y(g10803),.A(g10708));
  NOT NOT1_5046(.VSS(VSS),.VDD(VDD),.Y(I7205),.A(g2632));
  NOT NOT1_5047(.VSS(VSS),.VDD(VDD),.Y(I9773),.A(g4934));
  NOT NOT1_5048(.VSS(VSS),.VDD(VDD),.Y(I15759),.A(g10267));
  NOT NOT1_5049(.VSS(VSS),.VDD(VDD),.Y(I11061),.A(g6641));
  NOT NOT1_5050(.VSS(VSS),.VDD(VDD),.Y(I15725),.A(g10251));
  NOT NOT1_5051(.VSS(VSS),.VDD(VDD),.Y(g5701),.A(I9240));
  NOT NOT1_5052(.VSS(VSS),.VDD(VDD),.Y(g3708),.A(I6867));
  NOT NOT1_5053(.VSS(VSS),.VDD(VDD),.Y(g4953),.A(I8324));
  NOT NOT1_5054(.VSS(VSS),.VDD(VDD),.Y(g2751),.A(I5821));
  NOT NOT1_5055(.VSS(VSS),.VDD(VDD),.Y(g3520),.A(g2779));
  NOT NOT1_5056(.VSS(VSS),.VDD(VDD),.Y(g8950),.A(I14303));
  NOT NOT1_5057(.VSS(VSS),.VDD(VDD),.Y(I16500),.A(g10711));
  NOT NOT1_5058(.VSS(VSS),.VDD(VDD),.Y(g3219),.A(I6395));
  NOT NOT1_5059(.VSS(VSS),.VDD(VDD),.Y(I6517),.A(g3271));
  NOT NOT1_5060(.VSS(VSS),.VDD(VDD),.Y(I6690),.A(g2743));
  NOT NOT1_5061(.VSS(VSS),.VDD(VDD),.Y(I9409),.A(g5013));
  NOT NOT1_5062(.VSS(VSS),.VDD(VDD),.Y(I15114),.A(g9875));
  NOT NOT1_5063(.VSS(VSS),.VDD(VDD),.Y(I5427),.A(g913));
  NOT NOT1_5064(.VSS(VSS),.VDD(VDD),.Y(g4468),.A(I7837));
  NOT NOT1_5065(.VSS(VSS),.VDD(VDD),.Y(I15082),.A(g9719));
  NOT NOT1_5066(.VSS(VSS),.VDD(VDD),.Y(g6117),.A(I9804));
  NOT NOT1_5067(.VSS(VSS),.VDD(VDD),.Y(I14989),.A(g9813));
  NOT NOT1_5068(.VSS(VSS),.VDD(VDD),.Y(I17158),.A(g11312));
  NOT NOT1_5069(.VSS(VSS),.VDD(VDD),.Y(g3252),.A(I6414));
  NOT NOT1_5070(.VSS(VSS),.VDD(VDD),.Y(g10881),.A(I16613));
  NOT NOT1_5071(.VSS(VSS),.VDD(VDD),.Y(I7104),.A(g3186));
  NOT NOT1_5072(.VSS(VSS),.VDD(VDD),.Y(g11435),.A(I17356));
  NOT NOT1_5073(.VSS(VSS),.VDD(VDD),.Y(I6876),.A(g2956));
  NOT NOT1_5074(.VSS(VSS),.VDD(VDD),.Y(I9769),.A(g5287));
  NOT NOT1_5075(.VSS(VSS),.VDD(VDD),.Y(g11082),.A(I16859));
  NOT NOT1_5076(.VSS(VSS),.VDD(VDD),.Y(g3812),.A(g3228));
  NOT NOT1_5077(.VSS(VSS),.VDD(VDD),.Y(I7099),.A(g3228));
  NOT NOT1_5078(.VSS(VSS),.VDD(VDD),.Y(I12457),.A(g7559));
  NOT NOT1_5079(.VSS(VSS),.VDD(VDD),.Y(I10924),.A(g6736));
  NOT NOT1_5080(.VSS(VSS),.VDD(VDD),.Y(g5886),.A(g5361));
  NOT NOT1_5081(.VSS(VSS),.VDD(VDD),.Y(g11107),.A(g10974));
  NOT NOT1_5082(.VSS(VSS),.VDD(VDD),.Y(I9836),.A(g5405));
  NOT NOT1_5083(.VSS(VSS),.VDD(VDD),.Y(I14080),.A(g8714));
  NOT NOT1_5084(.VSS(VSS),.VDD(VDD),.Y(g7351),.A(I11701));
  NOT NOT1_5085(.VSS(VSS),.VDD(VDD),.Y(g2041),.A(g1791));
  NOT NOT1_5086(.VSS(VSS),.VDD(VDD),.Y(g7648),.A(I12255));
  NOT NOT1_5087(.VSS(VSS),.VDD(VDD),.Y(g7530),.A(I11926));
  NOT NOT1_5088(.VSS(VSS),.VDD(VDD),.Y(I11360),.A(g6351));
  NOT NOT1_5089(.VSS(VSS),.VDD(VDD),.Y(g8562),.A(I13779));
  NOT NOT1_5090(.VSS(VSS),.VDD(VDD),.Y(I15744),.A(g10261));
  NOT NOT1_5091(.VSS(VSS),.VDD(VDD),.Y(I13360),.A(g8126));
  NOT NOT1_5092(.VSS(VSS),.VDD(VDD),.Y(I17353),.A(g11381));
  NOT NOT1_5093(.VSS(VSS),.VDD(VDD),.Y(g3405),.A(g3144));
  NOT NOT1_5094(.VSS(VSS),.VDD(VDD),.Y(g5114),.A(I8506));
  NOT NOT1_5095(.VSS(VSS),.VDD(VDD),.Y(I5403),.A(g636));
  NOT NOT1_5096(.VSS(VSS),.VDD(VDD),.Y(g9778),.A(g9474));
  NOT NOT1_5097(.VSS(VSS),.VDD(VDD),.Y(g5314),.A(g4387));
  NOT NOT1_5098(.VSS(VSS),.VDD(VDD),.Y(I11447),.A(g6431));
  NOT NOT1_5099(.VSS(VSS),.VDD(VDD),.Y(g11345),.A(I17158));
  NOT NOT1_5100(.VSS(VSS),.VDD(VDD),.Y(g9894),.A(I15085));
  NOT NOT1_5101(.VSS(VSS),.VDD(VDD),.Y(g8723),.A(g8585));
  NOT NOT1_5102(.VSS(VSS),.VDD(VDD),.Y(g4716),.A(g3546));
  NOT NOT1_5103(.VSS(VSS),.VDD(VDD),.Y(I11162),.A(g6479));
  NOT NOT1_5104(.VSS(VSS),.VDD(VDD),.Y(I16613),.A(g10794));
  NOT NOT1_5105(.VSS(VSS),.VDD(VDD),.Y(g11399),.A(I17240));
  NOT NOT1_5106(.VSS(VSS),.VDD(VDD),.Y(g3765),.A(g3120));
  NOT NOT1_5107(.VSS(VSS),.VDD(VDD),.Y(I10753),.A(g5814));
  NOT NOT1_5108(.VSS(VSS),.VDD(VDD),.Y(I10461),.A(g5849));
  NOT NOT1_5109(.VSS(VSS),.VDD(VDD),.Y(I5391),.A(g1101));
  NOT NOT1_5110(.VSS(VSS),.VDD(VDD),.Y(g3911),.A(g3015));
  NOT NOT1_5111(.VSS(VSS),.VDD(VDD),.Y(I9229),.A(g4954));
  NOT NOT1_5112(.VSS(VSS),.VDD(VDD),.Y(g7010),.A(I11155));
  NOT NOT1_5113(.VSS(VSS),.VDD(VDD),.Y(g6581),.A(I10531));
  NOT NOT1_5114(.VSS(VSS),.VDD(VDD),.Y(g10890),.A(I16632));
  NOT NOT1_5115(.VSS(VSS),.VDD(VDD),.Y(g5650),.A(I9111));
  NOT NOT1_5116(.VSS(VSS),.VDD(VDD),.Y(g7410),.A(I11790));
  NOT NOT1_5117(.VSS(VSS),.VDD(VDD),.Y(g9782),.A(I14933));
  NOT NOT1_5118(.VSS(VSS),.VDD(VDD),.Y(g11398),.A(I17237));
  NOT NOT1_5119(.VSS(VSS),.VDD(VDD),.Y(I15804),.A(g10283));
  NOT NOT1_5120(.VSS(VSS),.VDD(VDD),.Y(I16947),.A(g11080));
  NOT NOT1_5121(.VSS(VSS),.VDD(VDD),.Y(I5695),.A(g575));
  NOT NOT1_5122(.VSS(VSS),.VDD(VDD),.Y(g10249),.A(g10135));
  NOT NOT1_5123(.VSS(VSS),.VDD(VDD),.Y(g2168),.A(I5111));
  NOT NOT1_5124(.VSS(VSS),.VDD(VDD),.Y(g2669),.A(g2015));
  NOT NOT1_5125(.VSS(VSS),.VDD(VDD),.Y(g6060),.A(I9695));
  NOT NOT1_5126(.VSS(VSS),.VDD(VDD),.Y(I16273),.A(g10559));
  NOT NOT1_5127(.VSS(VSS),.VDD(VDD),.Y(g2368),.A(I5445));
  NOT NOT1_5128(.VSS(VSS),.VDD(VDD),.Y(I11629),.A(g6914));
  NOT NOT1_5129(.VSS(VSS),.VDD(VDD),.Y(g11652),.A(I17758));
  NOT NOT1_5130(.VSS(VSS),.VDD(VDD),.Y(I9822),.A(g5219));
  NOT NOT1_5131(.VSS(VSS),.VDD(VDD),.Y(g9661),.A(I14786));
  NOT NOT1_5132(.VSS(VSS),.VDD(VDD),.Y(g4198),.A(I7411));
  NOT NOT1_5133(.VSS(VSS),.VDD(VDD),.Y(g4747),.A(g3586));
  NOT NOT1_5134(.VSS(VSS),.VDD(VDD),.Y(I11472),.A(g6488));
  NOT NOT1_5135(.VSS(VSS),.VDD(VDD),.Y(I10736),.A(g6104));
  NOT NOT1_5136(.VSS(VSS),.VDD(VDD),.Y(g4398),.A(g3914));
  NOT NOT1_5137(.VSS(VSS),.VDD(VDD),.Y(I13451),.A(g8152));
  NOT NOT1_5138(.VSS(VSS),.VDD(VDD),.Y(g3733),.A(I6917));
  NOT NOT1_5139(.VSS(VSS),.VDD(VDD),.Y(I7444),.A(g3683));
  NOT NOT1_5140(.VSS(VSS),.VDD(VDD),.Y(g10248),.A(g10134));
  NOT NOT1_5141(.VSS(VSS),.VDD(VDD),.Y(g2772),.A(g2508));
  NOT NOT1_5142(.VSS(VSS),.VDD(VDD),.Y(I7269),.A(g2851));
  NOT NOT1_5143(.VSS(VSS),.VDD(VDD),.Y(I15263),.A(g9995));
  NOT NOT1_5144(.VSS(VSS),.VDD(VDD),.Y(I10198),.A(g6118));
  NOT NOT1_5145(.VSS(VSS),.VDD(VDD),.Y(I12300),.A(g7240));
  NOT NOT1_5146(.VSS(VSS),.VDD(VDD),.Y(g10552),.A(I16217));
  NOT NOT1_5147(.VSS(VSS),.VDD(VDD),.Y(g8751),.A(g8632));
  NOT NOT1_5148(.VSS(VSS),.VDD(VDD),.Y(I15332),.A(g10001));
  NOT NOT1_5149(.VSS(VSS),.VDD(VDD),.Y(g10204),.A(g10174));
  NOT NOT1_5150(.VSS(VSS),.VDD(VDD),.Y(g2743),.A(I5801));
  NOT NOT1_5151(.VSS(VSS),.VDD(VDD),.Y(g4241),.A(g3664));
  NOT NOT1_5152(.VSS(VSS),.VDD(VDD),.Y(g2890),.A(I6052));
  NOT NOT1_5153(.VSS(VSS),.VDD(VDD),.Y(g5768),.A(I9352));
  NOT NOT1_5154(.VSS(VSS),.VDD(VDD),.Y(I10843),.A(g6723));
  NOT NOT1_5155(.VSS(VSS),.VDD(VDD),.Y(g8585),.A(I13828));
  NOT NOT1_5156(.VSS(VSS),.VDD(VDD),.Y(I5858),.A(g2529));
  NOT NOT1_5157(.VSS(VSS),.VDD(VDD),.Y(g5594),.A(I9016));
  NOT NOT1_5158(.VSS(VSS),.VDD(VDD),.Y(I14528),.A(g9270));
  NOT NOT1_5159(.VSS(VSS),.VDD(VDD),.Y(g3473),.A(I6676));
  NOT NOT1_5160(.VSS(VSS),.VDD(VDD),.Y(g7278),.A(I11524));
  NOT NOT1_5161(.VSS(VSS),.VDD(VDD),.Y(I14330),.A(g8819));
  NOT NOT1_5162(.VSS(VSS),.VDD(VDD),.Y(g9526),.A(g9256));
  NOT NOT1_5163(.VSS(VSS),.VDD(VDD),.Y(I4938),.A(g261));
  NOT NOT1_5164(.VSS(VSS),.VDD(VDD),.Y(I8250),.A(g4589));
  NOT NOT1_5165(.VSS(VSS),.VDD(VDD),.Y(I11071),.A(g6656));
  NOT NOT1_5166(.VSS(VSS),.VDD(VDD),.Y(I15406),.A(g10065));
  NOT NOT1_5167(.VSS(VSS),.VDD(VDD),.Y(I15962),.A(g10405));
  NOT NOT1_5168(.VSS(VSS),.VDD(VDD),.Y(g2011),.A(g976));
  NOT NOT1_5169(.VSS(VSS),.VDD(VDD),.Y(g6995),.A(g6482));
  NOT NOT1_5170(.VSS(VSS),.VDD(VDD),.Y(g7618),.A(I12202));
  NOT NOT1_5171(.VSS(VSS),.VDD(VDD),.Y(g3980),.A(g3121));
  NOT NOT1_5172(.VSS(VSS),.VDD(VDD),.Y(g8441),.A(I13621));
  NOT NOT1_5173(.VSS(VSS),.VDD(VDD),.Y(g11406),.A(I17261));
  NOT NOT1_5174(.VSS(VSS),.VDD(VDD),.Y(g5943),.A(I9581));
  NOT NOT1_5175(.VSS(VSS),.VDD(VDD),.Y(g7343),.A(I11677));
  NOT NOT1_5176(.VSS(VSS),.VDD(VDD),.Y(g2411),.A(I5494));
  NOT NOT1_5177(.VSS(VSS),.VDD(VDD),.Y(I10132),.A(g5696));
  NOT NOT1_5178(.VSS(VSS),.VDD(VDD),.Y(g10786),.A(I16484));
  NOT NOT1_5179(.VSS(VSS),.VDD(VDD),.Y(g3069),.A(I6277));
  NOT NOT1_5180(.VSS(VSS),.VDD(VDD),.Y(I13776),.A(g8513));
  NOT NOT1_5181(.VSS(VSS),.VDD(VDD),.Y(I13785),.A(g8516));
  NOT NOT1_5182(.VSS(VSS),.VDD(VDD),.Y(g1982),.A(g736));
  NOT NOT1_5183(.VSS(VSS),.VDD(VDD),.Y(g4524),.A(g3946));
  NOT NOT1_5184(.VSS(VSS),.VDD(VDD),.Y(g6294),.A(I10141));
  NOT NOT1_5185(.VSS(VSS),.VDD(VDD),.Y(I15500),.A(g10051));
  NOT NOT1_5186(.VSS(VSS),.VDD(VDD),.Y(I5251),.A(g1424));
  NOT NOT1_5187(.VSS(VSS),.VDD(VDD),.Y(I6590),.A(g3186));
  NOT NOT1_5188(.VSS(VSS),.VDD(VDD),.Y(g3540),.A(g3307));
  NOT NOT1_5189(.VSS(VSS),.VDD(VDD),.Y(I7729),.A(g3757));
  NOT NOT1_5190(.VSS(VSS),.VDD(VDD),.Y(g5887),.A(I9510));
  NOT NOT1_5191(.VSS(VSS),.VDD(VDD),.Y(g10356),.A(I15832));
  NOT NOT1_5192(.VSS(VSS),.VDD(VDD),.Y(I5047),.A(g1185));
  NOT NOT1_5193(.VSS(VSS),.VDD(VDD),.Y(g5122),.A(g4682));
  NOT NOT1_5194(.VSS(VSS),.VDD(VDD),.Y(g11500),.A(I17519));
  NOT NOT1_5195(.VSS(VSS),.VDD(VDD),.Y(g6190),.A(g5426));
  NOT NOT1_5196(.VSS(VSS),.VDD(VDD),.Y(g2074),.A(g1377));
  NOT NOT1_5197(.VSS(VSS),.VDD(VDD),.Y(g4319),.A(g4144));
  NOT NOT1_5198(.VSS(VSS),.VDD(VDD),.Y(g7693),.A(I12326));
  NOT NOT1_5199(.VSS(VSS),.VDD(VDD),.Y(g11049),.A(I16808));
  NOT NOT1_5200(.VSS(VSS),.VDD(VDD),.Y(I11950),.A(g6906));
  NOT NOT1_5201(.VSS(VSS),.VDD(VDD),.Y(I16514),.A(g10717));
  NOT NOT1_5202(.VSS(VSS),.VDD(VDD),.Y(g10826),.A(I16540));
  NOT NOT1_5203(.VSS(VSS),.VDD(VDD),.Y(I9062),.A(g4759));
  NOT NOT1_5204(.VSS(VSS),.VDD(VDD),.Y(g7334),.A(I11650));
  NOT NOT1_5205(.VSS(VSS),.VDD(VDD),.Y(g10380),.A(I15864));
  NOT NOT1_5206(.VSS(VSS),.VDD(VDD),.Y(g3206),.A(g2055));
  NOT NOT1_5207(.VSS(VSS),.VDD(VDD),.Y(I13825),.A(g8488));
  NOT NOT1_5208(.VSS(VSS),.VDD(VDD),.Y(I13370),.A(g8128));
  NOT NOT1_5209(.VSS(VSS),.VDD(VDD),.Y(I9620),.A(g5189));
  NOT NOT1_5210(.VSS(VSS),.VDD(VDD),.Y(g4258),.A(I7509));
  NOT NOT1_5211(.VSS(VSS),.VDD(VDD),.Y(I16507),.A(g10712));
  NOT NOT1_5212(.VSS(VSS),.VDD(VDD),.Y(g4352),.A(I7633));
  NOT NOT1_5213(.VSS(VSS),.VDD(VDD),.Y(I11858),.A(g6888));
  NOT NOT1_5214(.VSS(VSS),.VDD(VDD),.Y(g11048),.A(I16805));
  NOT NOT1_5215(.VSS(VSS),.VDD(VDD),.Y(g4577),.A(I7984));
  NOT NOT1_5216(.VSS(VSS),.VDD(VDD),.Y(g4867),.A(I8204));
  NOT NOT1_5217(.VSS(VSS),.VDD(VDD),.Y(I14709),.A(g9267));
  NOT NOT1_5218(.VSS(VSS),.VDD(VDD),.Y(g5033),.A(I8406));
  NOT NOT1_5219(.VSS(VSS),.VDD(VDD),.Y(g10233),.A(g10187));
  NOT NOT1_5220(.VSS(VSS),.VDD(VDD),.Y(g6156),.A(g5426));
  NOT NOT1_5221(.VSS(VSS),.VDD(VDD),.Y(g4717),.A(g3829));
  NOT NOT1_5222(.VSS(VSS),.VDD(VDD),.Y(I7014),.A(g2919));
  NOT NOT1_5223(.VSS(VSS),.VDD(VDD),.Y(I12511),.A(g7733));
  NOT NOT1_5224(.VSS(VSS),.VDD(VDD),.Y(g10182),.A(I15530));
  NOT NOT1_5225(.VSS(VSS),.VDD(VDD),.Y(g7555),.A(I11989));
  NOT NOT1_5226(.VSS(VSS),.VDD(VDD),.Y(g7804),.A(I12577));
  NOT NOT1_5227(.VSS(VSS),.VDD(VDD),.Y(I7414),.A(g4156));
  NOT NOT1_5228(.VSS(VSS),.VDD(VDD),.Y(I10087),.A(g5753));
  NOT NOT1_5229(.VSS(VSS),.VDD(VDD),.Y(g9919),.A(I15114));
  NOT NOT1_5230(.VSS(VSS),.VDD(VDD),.Y(g2080),.A(I4894));
  NOT NOT1_5231(.VSS(VSS),.VDD(VDD),.Y(I7946),.A(g3417));
  NOT NOT1_5232(.VSS(VSS),.VDD(VDD),.Y(I10258),.A(g6134));
  NOT NOT1_5233(.VSS(VSS),.VDD(VDD),.Y(I14087),.A(g8770));
  NOT NOT1_5234(.VSS(VSS),.VDD(VDD),.Y(g7792),.A(I12541));
  NOT NOT1_5235(.VSS(VSS),.VDD(VDD),.Y(g2480),.A(I5561));
  NOT NOT1_5236(.VSS(VSS),.VDD(VDD),.Y(I11367),.A(g6392));
  NOT NOT1_5237(.VSS(VSS),.VDD(VDD),.Y(I11394),.A(g6621));
  NOT NOT1_5238(.VSS(VSS),.VDD(VDD),.Y(g5096),.A(g4840));
  NOT NOT1_5239(.VSS(VSS),.VDD(VDD),.Y(g6942),.A(I11076));
  NOT NOT1_5240(.VSS(VSS),.VDD(VDD),.Y(g8890),.A(I14236));
  NOT NOT1_5241(.VSS(VSS),.VDD(VDD),.Y(g2713),.A(g2042));
  NOT NOT1_5242(.VSS(VSS),.VDD(VDD),.Y(I13367),.A(g8221));
  NOT NOT1_5243(.VSS(VSS),.VDD(VDD),.Y(I13394),.A(g8137));
  NOT NOT1_5244(.VSS(VSS),.VDD(VDD),.Y(g4211),.A(I7450));
  NOT NOT1_5245(.VSS(VSS),.VDD(VDD),.Y(g4186),.A(I7375));
  NOT NOT1_5246(.VSS(VSS),.VDD(VDD),.Y(g6704),.A(g5949));
  NOT NOT1_5247(.VSS(VSS),.VDD(VDD),.Y(I17687),.A(g11610));
  NOT NOT1_5248(.VSS(VSS),.VDD(VDD),.Y(g4386),.A(I7713));
  NOT NOT1_5249(.VSS(VSS),.VDD(VDD),.Y(g10932),.A(g10827));
  NOT NOT1_5250(.VSS(VSS),.VDD(VDD),.Y(I8929),.A(g4582));
  NOT NOT1_5251(.VSS(VSS),.VDD(VDD),.Y(g5845),.A(g5320));
  NOT NOT1_5252(.VSS(VSS),.VDD(VDD),.Y(g4975),.A(I8351));
  NOT NOT1_5253(.VSS(VSS),.VDD(VDD),.Y(g2569),.A(I5695));
  NOT NOT1_5254(.VSS(VSS),.VDD(VDD),.Y(I7513),.A(g4144));
  NOT NOT1_5255(.VSS(VSS),.VDD(VDD),.Y(g8011),.A(I12853));
  NOT NOT1_5256(.VSS(VSS),.VDD(VDD),.Y(I17752),.A(g11645));
  NOT NOT1_5257(.VSS(VSS),.VDD(VDD),.Y(g5195),.A(g4453));
  NOT NOT1_5258(.VSS(VSS),.VDD(VDD),.Y(g5395),.A(I8831));
  NOT NOT1_5259(.VSS(VSS),.VDD(VDD),.Y(g5891),.A(g5361));
  NOT NOT1_5260(.VSS(VSS),.VDD(VDD),.Y(I9842),.A(g5405));
  NOT NOT1_5261(.VSS(VSS),.VDD(VDD),.Y(I17374),.A(g11411));
  NOT NOT1_5262(.VSS(VSS),.VDD(VDD),.Y(g7113),.A(I11348));
  NOT NOT1_5263(.VSS(VSS),.VDD(VDD),.Y(g11106),.A(g10974));
  NOT NOT1_5264(.VSS(VSS),.VDD(VDD),.Y(g7313),.A(I11587));
  NOT NOT1_5265(.VSS(VSS),.VDD(VDD),.Y(I11420),.A(g6417));
  NOT NOT1_5266(.VSS(VSS),.VDD(VDD),.Y(g4426),.A(g3914));
  NOT NOT1_5267(.VSS(VSS),.VDD(VDD),.Y(g10897),.A(g10827));
  NOT NOT1_5268(.VSS(VSS),.VDD(VDD),.Y(I12916),.A(g7849));
  NOT NOT1_5269(.VSS(VSS),.VDD(VDD),.Y(I10069),.A(g5787));
  NOT NOT1_5270(.VSS(VSS),.VDD(VDD),.Y(g6954),.A(I11100));
  NOT NOT1_5271(.VSS(VSS),.VDD(VDD),.Y(g6250),.A(I10009));
  NOT NOT1_5272(.VSS(VSS),.VDD(VDD),.Y(g4170),.A(g3328));
  NOT NOT1_5273(.VSS(VSS),.VDD(VDD),.Y(g6810),.A(I10840));
  NOT NOT1_5274(.VSS(VSS),.VDD(VDD),.Y(g4614),.A(g3829));
  NOT NOT1_5275(.VSS(VSS),.VDD(VDD),.Y(g9527),.A(I14668));
  NOT NOT1_5276(.VSS(VSS),.VDD(VDD),.Y(g4370),.A(I7671));
  NOT NOT1_5277(.VSS(VSS),.VDD(VDD),.Y(I12550),.A(g7675));
  NOT NOT1_5278(.VSS(VSS),.VDD(VDD),.Y(I7378),.A(g4067));
  NOT NOT1_5279(.VSS(VSS),.VDD(VDD),.Y(I10810),.A(g6539));
  NOT NOT1_5280(.VSS(VSS),.VDD(VDD),.Y(I11318),.A(g6488));
  NOT NOT1_5281(.VSS(VSS),.VDD(VDD),.Y(g4125),.A(I7272));
  NOT NOT1_5282(.VSS(VSS),.VDD(VDD),.Y(I15371),.A(g9990));
  NOT NOT1_5283(.VSS(VSS),.VDD(VDD),.Y(g6432),.A(g6146));
  NOT NOT1_5284(.VSS(VSS),.VDD(VDD),.Y(g7908),.A(g7454));
  NOT NOT1_5285(.VSS(VSS),.VDD(VDD),.Y(I13227),.A(g8264));
  NOT NOT1_5286(.VSS(VSS),.VDD(VDD),.Y(g6053),.A(I9684));
  NOT NOT1_5287(.VSS(VSS),.VDD(VDD),.Y(I14955),.A(g9765));
  NOT NOT1_5288(.VSS(VSS),.VDD(VDD),.Y(I17669),.A(g11604));
  NOT NOT1_5289(.VSS(VSS),.VDD(VDD),.Y(g8992),.A(I14397));
  NOT NOT1_5290(.VSS(VSS),.VDD(VDD),.Y(g9764),.A(g9432));
  NOT NOT1_5291(.VSS(VSS),.VDD(VDD),.Y(I16920),.A(g11084));
  NOT NOT1_5292(.VSS(VSS),.VDD(VDD),.Y(g11033),.A(I16760));
  NOT NOT1_5293(.VSS(VSS),.VDD(VDD),.Y(g3291),.A(g2161));
  NOT NOT1_5294(.VSS(VSS),.VDD(VDD),.Y(I12307),.A(g7245));
  NOT NOT1_5295(.VSS(VSS),.VDD(VDD),.Y(I5935),.A(g2174));
  NOT NOT1_5296(.VSS(VSS),.VDD(VDD),.Y(I6844),.A(g2915));
  NOT NOT1_5297(.VSS(VSS),.VDD(VDD),.Y(g6453),.A(g5817));
  NOT NOT1_5298(.VSS(VSS),.VDD(VDD),.Y(I9854),.A(g5557));
  NOT NOT1_5299(.VSS(VSS),.VDD(VDD),.Y(I14970),.A(g9732));
  NOT NOT1_5300(.VSS(VSS),.VDD(VDD),.Y(g4280),.A(g4013));
  NOT NOT1_5301(.VSS(VSS),.VDD(VDD),.Y(I7182),.A(g2645));
  NOT NOT1_5302(.VSS(VSS),.VDD(VDD),.Y(I7288),.A(g2873));
  NOT NOT1_5303(.VSS(VSS),.VDD(VDD),.Y(g4939),.A(I8303));
  NOT NOT1_5304(.VSS(VSS),.VDD(VDD),.Y(I11540),.A(g6877));
  NOT NOT1_5305(.VSS(VSS),.VDD(VDD),.Y(I5982),.A(g2510));
  NOT NOT1_5306(.VSS(VSS),.VDD(VDD),.Y(g3144),.A(g2462));
  NOT NOT1_5307(.VSS(VSS),.VDD(VDD),.Y(I11058),.A(g6641));
  NOT NOT1_5308(.VSS(VSS),.VDD(VDD),.Y(I15795),.A(g10280));
  NOT NOT1_5309(.VSS(VSS),.VDD(VDD),.Y(g3344),.A(I6528));
  NOT NOT1_5310(.VSS(VSS),.VDD(VDD),.Y(I16121),.A(g10396));
  NOT NOT1_5311(.VSS(VSS),.VDD(VDD),.Y(g6568),.A(g5797));
  NOT NOT1_5312(.VSS(VSS),.VDD(VDD),.Y(I10171),.A(g5992));
  NOT NOT1_5313(.VSS(VSS),.VDD(VDD),.Y(g4083),.A(I7216));
  NOT NOT1_5314(.VSS(VSS),.VDD(VDD),.Y(g8080),.A(I12942));
  NOT NOT1_5315(.VSS(VSS),.VDD(VDD),.Y(I4879),.A(g256));
  NOT NOT1_5316(.VSS(VSS),.VDD(VDD),.Y(g4544),.A(g3880));
  NOT NOT1_5317(.VSS(VSS),.VDD(VDD),.Y(g3207),.A(g2439));
  NOT NOT1_5318(.VSS(VSS),.VDD(VDD),.Y(g8573),.A(I13812));
  NOT NOT1_5319(.VSS(VSS),.VDD(VDD),.Y(I7916),.A(g3664));
  NOT NOT1_5320(.VSS(VSS),.VDD(VDD),.Y(I7022),.A(g2941));
  NOT NOT1_5321(.VSS(VSS),.VDD(VDD),.Y(I13203),.A(g8196));
  NOT NOT1_5322(.VSS(VSS),.VDD(VDD),.Y(g8480),.A(I13682));
  NOT NOT1_5323(.VSS(VSS),.VDD(VDD),.Y(g7776),.A(I12493));
  NOT NOT1_5324(.VSS(VSS),.VDD(VDD),.Y(g2000),.A(g810));
  NOT NOT1_5325(.VSS(VSS),.VDD(VDD),.Y(I7749),.A(g3764));
  NOT NOT1_5326(.VSS(VSS),.VDD(VDD),.Y(I6557),.A(g3086));
  NOT NOT1_5327(.VSS(VSS),.VDD(VDD),.Y(g8713),.A(g8684));
  NOT NOT1_5328(.VSS(VSS),.VDD(VDD),.Y(I17525),.A(g11486));
  NOT NOT1_5329(.VSS(VSS),.VDD(VDD),.Y(g2126),.A(g12));
  NOT NOT1_5330(.VSS(VSS),.VDD(VDD),.Y(g4636),.A(I8036));
  NOT NOT1_5331(.VSS(VSS),.VDD(VDD),.Y(I15514),.A(g10122));
  NOT NOT1_5332(.VSS(VSS),.VDD(VDD),.Y(I17424),.A(g11424));
  NOT NOT1_5333(.VSS(VSS),.VDD(VDD),.Y(g3694),.A(I6851));
  NOT NOT1_5334(.VSS(VSS),.VDD(VDD),.Y(g6157),.A(I9880));
  NOT NOT1_5335(.VSS(VSS),.VDD(VDD),.Y(I6071),.A(g2269));
  NOT NOT1_5336(.VSS(VSS),.VDD(VDD),.Y(I14967),.A(g9763));
  NOT NOT1_5337(.VSS(VSS),.VDD(VDD),.Y(I12773),.A(g7581));
  NOT NOT1_5338(.VSS(VSS),.VDD(VDD),.Y(I16682),.A(g10799));
  NOT NOT1_5339(.VSS(VSS),.VDD(VDD),.Y(I17558),.A(g11504));
  NOT NOT1_5340(.VSS(VSS),.VDD(VDD),.Y(I15507),.A(g10047));
  NOT NOT1_5341(.VSS(VSS),.VDD(VDD),.Y(g5081),.A(I8449));
  NOT NOT1_5342(.VSS(VSS),.VDD(VDD),.Y(I12942),.A(g7982));
  NOT NOT1_5343(.VSS(VSS),.VDD(VDD),.Y(g3088),.A(I6294));
  NOT NOT1_5344(.VSS(VSS),.VDD(VDD),.Y(g5815),.A(I9421));
  NOT NOT1_5345(.VSS(VSS),.VDD(VDD),.Y(g8569),.A(I13800));
  NOT NOT1_5346(.VSS(VSS),.VDD(VDD),.Y(g4306),.A(g3586));
  NOT NOT1_5347(.VSS(VSS),.VDD(VDD),.Y(g7965),.A(I12759));
  NOT NOT1_5348(.VSS(VSS),.VDD(VDD),.Y(I12268),.A(g7107));
  NOT NOT1_5349(.VSS(VSS),.VDD(VDD),.Y(g5481),.A(I8900));
  NOT NOT1_5350(.VSS(VSS),.VDD(VDD),.Y(g11507),.A(I17540));
  NOT NOT1_5351(.VSS(VSS),.VDD(VDD),.Y(I12156),.A(g6878));
  NOT NOT1_5352(.VSS(VSS),.VDD(VDD),.Y(g4790),.A(g3337));
  NOT NOT1_5353(.VSS(VSS),.VDD(VDD),.Y(I12655),.A(g7402));
  NOT NOT1_5354(.VSS(VSS),.VDD(VDD),.Y(g5692),.A(I9221));
  NOT NOT1_5355(.VSS(VSS),.VDD(VDD),.Y(I15421),.A(g10083));
  NOT NOT1_5356(.VSS(VSS),.VDD(VDD),.Y(g1964),.A(g114));
  NOT NOT1_5357(.VSS(VSS),.VDD(VDD),.Y(g10387),.A(g10357));
  NOT NOT1_5358(.VSS(VSS),.VDD(VDD),.Y(g97),.A(I4780));
  NOT NOT1_5359(.VSS(VSS),.VDD(VDD),.Y(g7264),.A(I11501));
  NOT NOT1_5360(.VSS(VSS),.VDD(VDD),.Y(I12180),.A(g7263));
  NOT NOT1_5361(.VSS(VSS),.VDD(VDD),.Y(g10620),.A(I16295));
  NOT NOT1_5362(.VSS(VSS),.VDD(VDD),.Y(g4187),.A(I7378));
  NOT NOT1_5363(.VSS(VSS),.VDD(VDD),.Y(g4061),.A(I7182));
  NOT NOT1_5364(.VSS(VSS),.VDD(VDD),.Y(g10148),.A(g10121));
  NOT NOT1_5365(.VSS(VSS),.VDD(VDD),.Y(g11421),.A(I17318));
  NOT NOT1_5366(.VSS(VSS),.VDD(VDD),.Y(g4387),.A(I7716));
  NOT NOT1_5367(.VSS(VSS),.VDD(VDD),.Y(g4461),.A(g3829));
  NOT NOT1_5368(.VSS(VSS),.VDD(VDD),.Y(I6955),.A(g2871));
  NOT NOT1_5369(.VSS(VSS),.VDD(VDD),.Y(g7360),.A(I11728));
  NOT NOT1_5370(.VSS(VSS),.VDD(VDD),.Y(g11163),.A(I16920));
  NOT NOT1_5371(.VSS(VSS),.VDD(VDD),.Y(g10104),.A(I15338));
  NOT NOT1_5372(.VSS(VSS),.VDD(VDD),.Y(I11146),.A(g6439));
  NOT NOT1_5373(.VSS(VSS),.VDD(VDD),.Y(g4756),.A(g3440));
  NOT NOT1_5374(.VSS(VSS),.VDD(VDD),.Y(I17713),.A(g11621));
  NOT NOT1_5375(.VSS(VSS),.VDD(VDD),.Y(I13738),.A(g8295));
  NOT NOT1_5376(.VSS(VSS),.VDD(VDD),.Y(I13645),.A(g8379));
  NOT NOT1_5377(.VSS(VSS),.VDD(VDD),.Y(g8688),.A(g8507));
  NOT NOT1_5378(.VSS(VSS),.VDD(VDD),.Y(I12335),.A(g7133));
  NOT NOT1_5379(.VSS(VSS),.VDD(VDD),.Y(g7521),.A(I11901));
  NOT NOT1_5380(.VSS(VSS),.VDD(VDD),.Y(g10343),.A(I15795));
  NOT NOT1_5381(.VSS(VSS),.VDD(VDD),.Y(I14010),.A(g8642));
  NOT NOT1_5382(.VSS(VSS),.VDD(VDD),.Y(I14918),.A(g9535));
  NOT NOT1_5383(.VSS(VSS),.VDD(VDD),.Y(g8976),.A(I14349));
  NOT NOT1_5384(.VSS(VSS),.VDD(VDD),.Y(g2608),.A(I5725));
  NOT NOT1_5385(.VSS(VSS),.VDD(VDD),.Y(I9829),.A(g5013));
  NOT NOT1_5386(.VSS(VSS),.VDD(VDD),.Y(I16760),.A(g10888));
  NOT NOT1_5387(.VSS(VSS),.VDD(VDD),.Y(g2220),.A(g104));
  NOT NOT1_5388(.VSS(VSS),.VDD(VDD),.Y(g4427),.A(g3638));
  NOT NOT1_5389(.VSS(VSS),.VDD(VDD),.Y(I12930),.A(g7896));
  NOT NOT1_5390(.VSS(VSS),.VDD(VDD),.Y(g7450),.A(g7148));
  NOT NOT1_5391(.VSS(VSS),.VDD(VDD),.Y(I12993),.A(g8044));
  NOT NOT1_5392(.VSS(VSS),.VDD(VDD),.Y(I15473),.A(g10087));
  NOT NOT1_5393(.VSS(VSS),.VDD(VDD),.Y(I13290),.A(g8254));
  NOT NOT1_5394(.VSS(VSS),.VDD(VDD),.Y(g2779),.A(g1974));
  NOT NOT1_5395(.VSS(VSS),.VDD(VDD),.Y(I6150),.A(g2122));
  NOT NOT1_5396(.VSS(VSS),.VDD(VDD),.Y(g9987),.A(I15187));
  NOT NOT1_5397(.VSS(VSS),.VDD(VDD),.Y(g11541),.A(g11519));
  NOT NOT1_5398(.VSS(VSS),.VDD(VDD),.Y(I17610),.A(g11549));
  NOT NOT1_5399(.VSS(VSS),.VDD(VDD),.Y(I11698),.A(g7057));
  NOT NOT1_5400(.VSS(VSS),.VDD(VDD),.Y(g4200),.A(I7417));
  NOT NOT1_5401(.VSS(VSS),.VDD(VDD),.Y(g9771),.A(g9432));
  NOT NOT1_5402(.VSS(VSS),.VDD(VDD),.Y(I12694),.A(g7374));
  NOT NOT1_5403(.VSS(VSS),.VDD(VDD),.Y(I12838),.A(g7682));
  NOT NOT1_5404(.VSS(VSS),.VDD(VDD),.Y(g11473),.A(I17456));
  NOT NOT1_5405(.VSS(VSS),.VDD(VDD),.Y(g2023),.A(g1357));
  NOT NOT1_5406(.VSS(VSS),.VDD(VDD),.Y(I10078),.A(g5729));
  NOT NOT1_5407(.VSS(VSS),.VDD(VDD),.Y(I17255),.A(g11344));
  NOT NOT1_5408(.VSS(VSS),.VDD(VDD),.Y(g4514),.A(g3946));
  NOT NOT1_5409(.VSS(VSS),.VDD(VDD),.Y(I10598),.A(g5874));
  NOT NOT1_5410(.VSS(VSS),.VDD(VDD),.Y(g5783),.A(I9377));
  NOT NOT1_5411(.VSS(VSS),.VDD(VDD),.Y(g4003),.A(g3144));
  NOT NOT1_5412(.VSS(VSS),.VDD(VDD),.Y(g7724),.A(I12357));
  NOT NOT1_5413(.VSS(VSS),.VDD(VDD),.Y(I15359),.A(g10019));
  NOT NOT1_5414(.VSS(VSS),.VDD(VDD),.Y(I6409),.A(g2356));
  NOT NOT1_5415(.VSS(VSS),.VDD(VDD),.Y(g8126),.A(I12989));
  NOT NOT1_5416(.VSS(VSS),.VDD(VDD),.Y(I7719),.A(g3752));
  NOT NOT1_5417(.VSS(VSS),.VDD(VDD),.Y(g5112),.A(g4682));
  NOT NOT1_5418(.VSS(VSS),.VDD(VDD),.Y(g7379),.A(g6863));
  NOT NOT1_5419(.VSS(VSS),.VDD(VDD),.Y(g5218),.A(I8647));
  NOT NOT1_5420(.VSS(VSS),.VDD(VDD),.Y(g8326),.A(I13360));
  NOT NOT1_5421(.VSS(VSS),.VDD(VDD),.Y(I17188),.A(g11313));
  NOT NOT1_5422(.VSS(VSS),.VDD(VDD),.Y(I17124),.A(g11232));
  NOT NOT1_5423(.VSS(VSS),.VDD(VDD),.Y(g5267),.A(I8711));
  NOT NOT1_5424(.VSS(VSS),.VDD(VDD),.Y(I17678),.A(g11607));
  NOT NOT1_5425(.VSS(VSS),.VDD(VDD),.Y(I11427),.A(g6573));
  NOT NOT1_5426(.VSS(VSS),.VDD(VDD),.Y(I12487),.A(g7723));
  NOT NOT1_5427(.VSS(VSS),.VDD(VDD),.Y(I15829),.A(g10203));
  NOT NOT1_5428(.VSS(VSS),.VDD(VDD),.Y(I13427),.A(g8241));
  NOT NOT1_5429(.VSS(VSS),.VDD(VDD),.Y(g9892),.A(I15079));
  NOT NOT1_5430(.VSS(VSS),.VDD(VDD),.Y(I8039),.A(g3506));
  NOT NOT1_5431(.VSS(VSS),.VDD(VDD),.Y(I7752),.A(g3407));
  NOT NOT1_5432(.VSS(VSS),.VDD(VDD),.Y(g4763),.A(g3586));
  NOT NOT1_5433(.VSS(VSS),.VDD(VDD),.Y(I12502),.A(g7726));
  NOT NOT1_5434(.VSS(VSS),.VDD(VDD),.Y(g4191),.A(I7390));
  NOT NOT1_5435(.VSS(VSS),.VDD(VDD),.Y(I11632),.A(g6931));
  NOT NOT1_5436(.VSS(VSS),.VDD(VDD),.Y(g7878),.A(g7479));
  NOT NOT1_5437(.VSS(VSS),.VDD(VDD),.Y(g10850),.A(I16550));
  NOT NOT1_5438(.VSS(VSS),.VDD(VDD),.Y(g8760),.A(g8670));
  NOT NOT1_5439(.VSS(VSS),.VDD(VDD),.Y(g11434),.A(I17353));
  NOT NOT1_5440(.VSS(VSS),.VDD(VDD),.Y(g4391),.A(g3638));
  NOT NOT1_5441(.VSS(VSS),.VDD(VDD),.Y(g1989),.A(g770));
  NOT NOT1_5442(.VSS(VSS),.VDD(VDD),.Y(I10322),.A(g6193));
  NOT NOT1_5443(.VSS(VSS),.VDD(VDD),.Y(g7289),.A(I11543));
  NOT NOT1_5444(.VSS(VSS),.VDD(VDD),.Y(g7777),.A(I12496));
  NOT NOT1_5445(.VSS(VSS),.VDD(VDD),.Y(g7658),.A(I12271));
  NOT NOT1_5446(.VSS(VSS),.VDD(VDD),.Y(g5401),.A(I8839));
  NOT NOT1_5447(.VSS(VSS),.VDD(VDD),.Y(g3408),.A(g3108));
  NOT NOT1_5448(.VSS(VSS),.VDD(VDD),.Y(I10159),.A(g5936));
  NOT NOT1_5449(.VSS(VSS),.VDD(VDD),.Y(g10133),.A(g10064));
  NOT NOT1_5450(.VSS(VSS),.VDD(VDD),.Y(g5676),.A(I9185));
  NOT NOT1_5451(.VSS(VSS),.VDD(VDD),.Y(g2451),.A(g248));
  NOT NOT1_5452(.VSS(VSS),.VDD(VDD),.Y(I10901),.A(g6620));
  NOT NOT1_5453(.VSS(VSS),.VDD(VDD),.Y(g4637),.A(I8039));
  NOT NOT1_5454(.VSS(VSS),.VDD(VDD),.Y(I12279),.A(g7225));
  NOT NOT1_5455(.VSS(VSS),.VDD(VDD),.Y(I5348),.A(g746));
  NOT NOT1_5456(.VSS(VSS),.VDD(VDD),.Y(g3336),.A(I6523));
  NOT NOT1_5457(.VSS(VSS),.VDD(VDD),.Y(I15344),.A(g10025));
  NOT NOT1_5458(.VSS(VSS),.VDD(VDD),.Y(g6778),.A(g5987));
  NOT NOT1_5459(.VSS(VSS),.VDD(VDD),.Y(g7882),.A(g7479));
  NOT NOT1_5460(.VSS(VSS),.VDD(VDD),.Y(g3768),.A(I6979));
  NOT NOT1_5461(.VSS(VSS),.VDD(VDD),.Y(g10896),.A(I16650));
  NOT NOT1_5462(.VSS(VSS),.VDD(VDD),.Y(I13403),.A(g8236));
  NOT NOT1_5463(.VSS(VSS),.VDD(VDD),.Y(g11344),.A(I17155));
  NOT NOT1_5464(.VSS(VSS),.VDD(VDD),.Y(g4307),.A(g4013));
  NOT NOT1_5465(.VSS(VSS),.VDD(VDD),.Y(g4536),.A(g3880));
  NOT NOT1_5466(.VSS(VSS),.VDD(VDD),.Y(g10228),.A(I15604));
  NOT NOT1_5467(.VSS(VSS),.VDD(VDD),.Y(g4159),.A(I7300));
  NOT NOT1_5468(.VSS(VSS),.VDD(VDD),.Y(g2346),.A(I5414));
  NOT NOT1_5469(.VSS(VSS),.VDD(VDD),.Y(g4359),.A(g3880));
  NOT NOT1_5470(.VSS(VSS),.VDD(VDD),.Y(I12469),.A(g7531));
  NOT NOT1_5471(.VSS(VSS),.VDD(VDD),.Y(g6735),.A(I10736));
  NOT NOT1_5472(.VSS(VSS),.VDD(VDD),.Y(g8183),.A(I13102));
  NOT NOT1_5473(.VSS(VSS),.VDD(VDD),.Y(g8608),.A(g8482));
  NOT NOT1_5474(.VSS(VSS),.VDD(VDD),.Y(g8924),.A(I14249));
  NOT NOT1_5475(.VSS(VSS),.VDD(VDD),.Y(g5830),.A(I9446));
  NOT NOT1_5476(.VSS(VSS),.VDD(VDD),.Y(g7611),.A(I12183));
  NOT NOT1_5477(.VSS(VSS),.VDD(VDD),.Y(g8220),.A(g7826));
  NOT NOT1_5478(.VSS(VSS),.VDD(VDD),.Y(I12286),.A(g7231));
  NOT NOT1_5479(.VSS(VSS),.VDD(VDD),.Y(I14561),.A(g9025));
  NOT NOT1_5480(.VSS(VSS),.VDD(VDD),.Y(g5727),.A(I9273));
  NOT NOT1_5481(.VSS(VSS),.VDD(VDD),.Y(g2103),.A(I4961));
  NOT NOT1_5482(.VSS(VSS),.VDD(VDD),.Y(I8919),.A(g4576));
  NOT NOT1_5483(.VSS(VSS),.VDD(VDD),.Y(g3943),.A(g2779));
  NOT NOT1_5484(.VSS(VSS),.VDD(VDD),.Y(I9177),.A(g4904));
  NOT NOT1_5485(.VSS(VSS),.VDD(VDD),.Y(I7233),.A(g2817));
  NOT NOT1_5486(.VSS(VSS),.VDD(VDD),.Y(I10144),.A(g5689));
  NOT NOT1_5487(.VSS(VSS),.VDD(VDD),.Y(g9340),.A(I14525));
  NOT NOT1_5488(.VSS(VSS),.VDD(VDD),.Y(I14295),.A(g8806));
  NOT NOT1_5489(.VSS(VSS),.VDD(VDD),.Y(I9377),.A(g5576));
  NOT NOT1_5490(.VSS(VSS),.VDD(VDD),.Y(I17219),.A(g11292));
  NOT NOT1_5491(.VSS(VSS),.VDD(VDD),.Y(g7799),.A(I12562));
  NOT NOT1_5492(.VSS(VSS),.VDD(VDD),.Y(g4757),.A(I8109));
  NOT NOT1_5493(.VSS(VSS),.VDD(VDD),.Y(I16604),.A(g10786));
  NOT NOT1_5494(.VSS(VSS),.VDD(VDD),.Y(I7054),.A(g3093));
  NOT NOT1_5495(.VSS(VSS),.VDD(VDD),.Y(I11572),.A(g6822));
  NOT NOT1_5496(.VSS(VSS),.VDD(VDD),.Y(g8423),.A(I13583));
  NOT NOT1_5497(.VSS(VSS),.VDD(VDD),.Y(g6475),.A(g5987));
  NOT NOT1_5498(.VSS(VSS),.VDD(VDD),.Y(g4416),.A(g3638));
  NOT NOT1_5499(.VSS(VSS),.VDD(VDD),.Y(g7981),.A(g7624));
  NOT NOT1_5500(.VSS(VSS),.VDD(VDD),.Y(g6949),.A(I11091));
  NOT NOT1_5501(.VSS(VSS),.VDD(VDD),.Y(g3228),.A(I6409));
  NOT NOT1_5502(.VSS(VSS),.VDD(VDD),.Y(g8977),.A(I14352));
  NOT NOT1_5503(.VSS(VSS),.VDD(VDD),.Y(g2732),.A(I5792));
  NOT NOT1_5504(.VSS(VSS),.VDD(VDD),.Y(I9287),.A(g5576));
  NOT NOT1_5505(.VSS(VSS),.VDD(VDD),.Y(g9082),.A(g8892));
  NOT NOT1_5506(.VSS(VSS),.VDD(VDD),.Y(g10310),.A(I15736));
  NOT NOT1_5507(.VSS(VSS),.VDD(VDD),.Y(g8588),.A(I13831));
  NOT NOT1_5508(.VSS(VSS),.VDD(VDD),.Y(g7997),.A(g7697));
  NOT NOT1_5509(.VSS(VSS),.VDD(VDD),.Y(g2753),.A(I5827));
  NOT NOT1_5510(.VSS(VSS),.VDD(VDD),.Y(I12601),.A(g7629));
  NOT NOT1_5511(.VSS(VSS),.VDD(VDD),.Y(g6292),.A(I10135));
  NOT NOT1_5512(.VSS(VSS),.VDD(VDD),.Y(I11127),.A(g6452));
  NOT NOT1_5513(.VSS(VSS),.VDD(VDD),.Y(g4315),.A(g3863));
  NOT NOT1_5514(.VSS(VSS),.VDD(VDD),.Y(g4811),.A(g3661));
  NOT NOT1_5515(.VSS(VSS),.VDD(VDD),.Y(g2508),.A(g940));
  NOT NOT1_5516(.VSS(VSS),.VDD(VDD),.Y(g8361),.A(I13463));
  NOT NOT1_5517(.VSS(VSS),.VDD(VDD),.Y(g10379),.A(I15861));
  NOT NOT1_5518(.VSS(VSS),.VDD(VDD),.Y(I10966),.A(g6561));
  NOT NOT1_5519(.VSS(VSS),.VDD(VDD),.Y(g2240),.A(g88));
  NOT NOT1_5520(.VSS(VSS),.VDD(VDD),.Y(I8004),.A(g3967));
  NOT NOT1_5521(.VSS(VSS),.VDD(VDD),.Y(g2072),.A(I4876));
  NOT NOT1_5522(.VSS(VSS),.VDD(VDD),.Y(g3433),.A(I6648));
  NOT NOT1_5523(.VSS(VSS),.VDD(VDD),.Y(I6921),.A(g2839));
  NOT NOT1_5524(.VSS(VSS),.VDD(VDD),.Y(I5279),.A(g73));
  NOT NOT1_5525(.VSS(VSS),.VDD(VDD),.Y(g7332),.A(I11644));
  NOT NOT1_5526(.VSS(VSS),.VDD(VDD),.Y(g10050),.A(I15269));
  NOT NOT1_5527(.VSS(VSS),.VDD(VDD),.Y(I9199),.A(g4935));
  NOT NOT1_5528(.VSS(VSS),.VDD(VDD),.Y(g10378),.A(I15858));
  NOT NOT1_5529(.VSS(VSS),.VDD(VDD),.Y(I8647),.A(g4219));
  NOT NOT1_5530(.VSS(VSS),.VDD(VDD),.Y(I9399),.A(g5013));
  NOT NOT1_5531(.VSS(VSS),.VDD(VDD),.Y(g5624),.A(I9056));
  NOT NOT1_5532(.VSS(VSS),.VDD(VDD),.Y(g7680),.A(g7148));
  NOT NOT1_5533(.VSS(VSS),.VDD(VDD),.Y(g11506),.A(I17537));
  NOT NOT1_5534(.VSS(VSS),.VDD(VDD),.Y(g7353),.A(I11707));
  NOT NOT1_5535(.VSS(VSS),.VDD(VDD),.Y(g2043),.A(g1801));
  NOT NOT1_5536(.VSS(VSS),.VDD(VDD),.Y(g6084),.A(I9731));
  NOT NOT1_5537(.VSS(VSS),.VDD(VDD),.Y(g8327),.A(g8164));
  NOT NOT1_5538(.VSS(VSS),.VDD(VDD),.Y(I14364),.A(g8952));
  NOT NOT1_5539(.VSS(VSS),.VDD(VDD),.Y(g4874),.A(I8215));
  NOT NOT1_5540(.VSS(VSS),.VDD(VDD),.Y(g6039),.A(I9652));
  NOT NOT1_5541(.VSS(VSS),.VDD(VDD),.Y(g5068),.A(g4840));
  NOT NOT1_5542(.VSS(VSS),.VDD(VDD),.Y(I11956),.A(g6912));
  NOT NOT1_5543(.VSS(VSS),.VDD(VDD),.Y(g3096),.A(g2482));
  NOT NOT1_5544(.VSS(VSS),.VDD(VDD),.Y(I13956),.A(g8451));
  NOT NOT1_5545(.VSS(VSS),.VDD(VDD),.Y(I13376),.A(g8226));
  NOT NOT1_5546(.VSS(VSS),.VDD(VDD),.Y(I13385),.A(g8230));
  NOT NOT1_5547(.VSS(VSS),.VDD(VDD),.Y(I11103),.A(g6667));
  NOT NOT1_5548(.VSS(VSS),.VDD(VDD),.Y(g3496),.A(I6686));
  NOT NOT1_5549(.VSS(VSS),.VDD(VDD),.Y(g7744),.A(I12397));
  NOT NOT1_5550(.VSS(VSS),.VDD(VDD),.Y(I11889),.A(g6898));
  NOT NOT1_5551(.VSS(VSS),.VDD(VDD),.Y(I17470),.A(g11452));
  NOT NOT1_5552(.VSS(VSS),.VDD(VDD),.Y(g7802),.A(I12571));
  NOT NOT1_5553(.VSS(VSS),.VDD(VDD),.Y(I5652),.A(g554));
  NOT NOT1_5554(.VSS(VSS),.VDD(VDD),.Y(g8146),.A(g8033));
  NOT NOT1_5555(.VSS(VSS),.VDD(VDD),.Y(I5057),.A(g1961));
  NOT NOT1_5556(.VSS(VSS),.VDD(VDD),.Y(I11354),.A(g6553));
  NOT NOT1_5557(.VSS(VSS),.VDD(VDD),.Y(g2116),.A(I5020));
  NOT NOT1_5558(.VSS(VSS),.VDD(VDD),.Y(g8346),.A(I13418));
  NOT NOT1_5559(.VSS(VSS),.VDD(VDD),.Y(I5843),.A(g2509));
  NOT NOT1_5560(.VSS(VSS),.VDD(VDD),.Y(I13354),.A(g8214));
  NOT NOT1_5561(.VSS(VSS),.VDD(VDD),.Y(I8503),.A(g4445));
  NOT NOT1_5562(.VSS(VSS),.VDD(VDD),.Y(I5989),.A(g2252));
  NOT NOT1_5563(.VSS(VSS),.VDD(VDD),.Y(I9510),.A(g5421));
  NOT NOT1_5564(.VSS(VSS),.VDD(VDD),.Y(I11824),.A(g7246));
  NOT NOT1_5565(.VSS(VSS),.VDD(VDD),.Y(g2034),.A(g1766));
  NOT NOT1_5566(.VSS(VSS),.VDD(VDD),.Y(g5677),.A(I9188));
  NOT NOT1_5567(.VSS(VSS),.VDD(VDD),.Y(g8103),.A(g7994));
  NOT NOT1_5568(.VSS(VSS),.VDD(VDD),.Y(g3395),.A(I6601));
  NOT NOT1_5569(.VSS(VSS),.VDD(VDD),.Y(g2434),.A(g1362));
  NOT NOT1_5570(.VSS(VSS),.VDD(VDD),.Y(g3337),.A(g2745));
  NOT NOT1_5571(.VSS(VSS),.VDD(VDD),.Y(g3913),.A(g2920));
  NOT NOT1_5572(.VSS(VSS),.VDD(VDD),.Y(I10289),.A(g6003));
  NOT NOT1_5573(.VSS(VSS),.VDD(VDD),.Y(I17277),.A(g11390));
  NOT NOT1_5574(.VSS(VSS),.VDD(VDD),.Y(I12168),.A(g7256));
  NOT NOT1_5575(.VSS(VSS),.VDD(VDD),.Y(I11671),.A(g7047));
  NOT NOT1_5576(.VSS(VSS),.VDD(VDD),.Y(g9310),.A(I14503));
  NOT NOT1_5577(.VSS(VSS),.VDD(VDD),.Y(g6583),.A(I10535));
  NOT NOT1_5578(.VSS(VSS),.VDD(VDD),.Y(g6702),.A(g5949));
  NOT NOT1_5579(.VSS(VSS),.VDD(VDD),.Y(g4880),.A(g3638));
  NOT NOT1_5580(.VSS(VSS),.VDD(VDD),.Y(g5866),.A(g5361));
  NOT NOT1_5581(.VSS(VSS),.VDD(VDD),.Y(g8696),.A(g8656));
  NOT NOT1_5582(.VSS(VSS),.VDD(VDD),.Y(I5549),.A(g868));
  NOT NOT1_5583(.VSS(VSS),.VDD(VDD),.Y(I7029),.A(g2946));
  NOT NOT1_5584(.VSS(VSS),.VDD(VDD),.Y(I14309),.A(g8813));
  NOT NOT1_5585(.VSS(VSS),.VDD(VDD),.Y(g2347),.A(g1945));
  NOT NOT1_5586(.VSS(VSS),.VDD(VDD),.Y(I7429),.A(g3344));
  NOT NOT1_5587(.VSS(VSS),.VDD(VDD),.Y(g10802),.A(I16510));
  NOT NOT1_5588(.VSS(VSS),.VDD(VDD),.Y(g5149),.A(I8551));
  NOT NOT1_5589(.VSS(VSS),.VDD(VDD),.Y(I9144),.A(g5007));
  NOT NOT1_5590(.VSS(VSS),.VDD(VDD),.Y(I14224),.A(g8794));
  NOT NOT1_5591(.VSS(VSS),.VDD(VDD),.Y(g6919),.A(g6453));
  NOT NOT1_5592(.VSS(VSS),.VDD(VDD),.Y(I10308),.A(g6003));
  NOT NOT1_5593(.VSS(VSS),.VDD(VDD),.Y(I12363),.A(g7187));
  NOT NOT1_5594(.VSS(VSS),.VDD(VDD),.Y(I7956),.A(g3428));
  NOT NOT1_5595(.VSS(VSS),.VDD(VDD),.Y(g7901),.A(g7712));
  NOT NOT1_5596(.VSS(VSS),.VDD(VDD),.Y(g4272),.A(g3586));
  NOT NOT1_5597(.VSS(VSS),.VDD(VDD),.Y(I8320),.A(g4452));
  NOT NOT1_5598(.VSS(VSS),.VDD(VDD),.Y(g10730),.A(I16407));
  NOT NOT1_5599(.VSS(VSS),.VDD(VDD),.Y(I12478),.A(g7560));
  NOT NOT1_5600(.VSS(VSS),.VDD(VDD),.Y(I12015),.A(g6924));
  NOT NOT1_5601(.VSS(VSS),.VDD(VDD),.Y(g6276),.A(I10087));
  NOT NOT1_5602(.VSS(VSS),.VDD(VDD),.Y(g11649),.A(I17749));
  NOT NOT1_5603(.VSS(VSS),.VDD(VDD),.Y(g9824),.A(I14973));
  NOT NOT1_5604(.VSS(VSS),.VDD(VDD),.Y(g4243),.A(g3524));
  NOT NOT1_5605(.VSS(VSS),.VDD(VDD),.Y(g3266),.A(I6436));
  NOT NOT1_5606(.VSS(VSS),.VDD(VDD),.Y(I9259),.A(g5301));
  NOT NOT1_5607(.VSS(VSS),.VDD(VDD),.Y(g8240),.A(g7972));
  NOT NOT1_5608(.VSS(VSS),.VDD(VDD),.Y(g2914),.A(I6091));
  NOT NOT1_5609(.VSS(VSS),.VDD(VDD),.Y(g5198),.A(I8614));
  NOT NOT1_5610(.VSS(VSS),.VDD(VDD),.Y(g5747),.A(I9317));
  NOT NOT1_5611(.VSS(VSS),.VDD(VDD),.Y(I15491),.A(g10093));
  NOT NOT1_5612(.VSS(VSS),.VDD(VDD),.Y(g2210),.A(g103));
  NOT NOT1_5613(.VSS(VSS),.VDD(VDD),.Y(g4417),.A(I7757));
  NOT NOT1_5614(.VSS(VSS),.VDD(VDD),.Y(I10495),.A(g6144));
  NOT NOT1_5615(.VSS(VSS),.VDD(VDD),.Y(g8472),.A(I13666));
  NOT NOT1_5616(.VSS(VSS),.VDD(VDD),.Y(g6561),.A(g5773));
  NOT NOT1_5617(.VSS(VSS),.VDD(VDD),.Y(g11648),.A(I17746));
  NOT NOT1_5618(.VSS(VSS),.VDD(VDD),.Y(g4935),.A(g4420));
  NOT NOT1_5619(.VSS(VSS),.VDD(VDD),.Y(g9762),.A(I14903));
  NOT NOT1_5620(.VSS(VSS),.VDD(VDD),.Y(I17419),.A(g11421));
  NOT NOT1_5621(.VSS(VSS),.VDD(VDD),.Y(I12556),.A(g7678));
  NOT NOT1_5622(.VSS(VSS),.VDD(VDD),.Y(I15604),.A(g10148));
  NOT NOT1_5623(.VSS(VSS),.VDD(VDD),.Y(I10816),.A(g6406));
  NOT NOT1_5624(.VSS(VSS),.VDD(VDD),.Y(I9923),.A(g5308));
  NOT NOT1_5625(.VSS(VSS),.VDD(VDD),.Y(g2013),.A(g1101));
  NOT NOT1_5626(.VSS(VSS),.VDD(VDD),.Y(g8443),.A(I13627));
  NOT NOT1_5627(.VSS(VSS),.VDD(VDD),.Y(g7600),.A(I12150));
  NOT NOT1_5628(.VSS(VSS),.VDD(VDD),.Y(I12580),.A(g7540));
  NOT NOT1_5629(.VSS(VSS),.VDD(VDD),.Y(g7574),.A(g6995));
  NOT NOT1_5630(.VSS(VSS),.VDD(VDD),.Y(I6085),.A(g2234));
  NOT NOT1_5631(.VSS(VSS),.VDD(VDD),.Y(g10548),.A(I16209));
  NOT NOT1_5632(.VSS(VSS),.VDD(VDD),.Y(I17155),.A(g11310));
  NOT NOT1_5633(.VSS(VSS),.VDD(VDD),.Y(g3142),.A(I6360));
  NOT NOT1_5634(.VSS(VSS),.VDD(VDD),.Y(g5241),.A(g4386));
  NOT NOT1_5635(.VSS(VSS),.VDD(VDD),.Y(g6527),.A(I10445));
  NOT NOT1_5636(.VSS(VSS),.VDD(VDD),.Y(I12223),.A(g7049));
  NOT NOT1_5637(.VSS(VSS),.VDD(VDD),.Y(g4328),.A(g4130));
  NOT NOT1_5638(.VSS(VSS),.VDD(VDD),.Y(I14687),.A(g9258));
  NOT NOT1_5639(.VSS(VSS),.VDD(VDD),.Y(I17170),.A(g11294));
  NOT NOT1_5640(.VSS(VSS),.VDD(VDD),.Y(I14976),.A(g9670));
  NOT NOT1_5641(.VSS(VSS),.VDD(VDD),.Y(g8116),.A(I12971));
  NOT NOT1_5642(.VSS(VSS),.VDD(VDD),.Y(g3255),.A(I6421));
  NOT NOT1_5643(.VSS(VSS),.VDD(VDD),.Y(I7639),.A(g3722));
  NOT NOT1_5644(.VSS(VSS),.VDD(VDD),.Y(g8316),.A(I13332));
  NOT NOT1_5645(.VSS(VSS),.VDD(VDD),.Y(g3815),.A(g3228));
  NOT NOT1_5646(.VSS(VSS),.VDD(VDD),.Y(I11211),.A(g6527));
  NOT NOT1_5647(.VSS(VSS),.VDD(VDD),.Y(I10374),.A(g5852));
  NOT NOT1_5648(.VSS(VSS),.VDD(VDD),.Y(g6764),.A(g5987));
  NOT NOT1_5649(.VSS(VSS),.VDD(VDD),.Y(I7109),.A(g2970));
  NOT NOT1_5650(.VSS(VSS),.VDD(VDD),.Y(I5909),.A(g2207));
  NOT NOT1_5651(.VSS(VSS),.VDD(VDD),.Y(I16534),.A(g10747));
  NOT NOT1_5652(.VSS(VSS),.VDD(VDD),.Y(I10643),.A(g6026));
  NOT NOT1_5653(.VSS(VSS),.VDD(VDD),.Y(I11088),.A(g6434));
  NOT NOT1_5654(.VSS(VSS),.VDD(VDD),.Y(I11024),.A(g6399));
  NOT NOT1_5655(.VSS(VSS),.VDD(VDD),.Y(g9556),.A(I14701));
  NOT NOT1_5656(.VSS(VSS),.VDD(VDD),.Y(I16098),.A(g10369));
  NOT NOT1_5657(.VSS(VSS),.VDD(VDD),.Y(g10317),.A(I15749));
  NOT NOT1_5658(.VSS(VSS),.VDD(VDD),.Y(g8565),.A(I13788));
  NOT NOT1_5659(.VSS(VSS),.VDD(VDD),.Y(g2820),.A(I5926));
  NOT NOT1_5660(.VSS(VSS),.VDD(VDD),.Y(g3097),.A(g2482));
  NOT NOT1_5661(.VSS(VSS),.VDD(VDD),.Y(I9886),.A(g5286));
  NOT NOT1_5662(.VSS(VSS),.VDD(VDD),.Y(I6941),.A(g2858));
  NOT NOT1_5663(.VSS(VSS),.VDD(VDD),.Y(g3726),.A(I6898));
  NOT NOT1_5664(.VSS(VSS),.VDD(VDD),.Y(g7580),.A(I12056));
  NOT NOT1_5665(.VSS(VSS),.VDD(VDD),.Y(g6503),.A(I10421));
  NOT NOT1_5666(.VSS(VSS),.VDD(VDD),.Y(g5644),.A(I9093));
  NOT NOT1_5667(.VSS(VSS),.VDD(VDD),.Y(I5740),.A(g2341));
  NOT NOT1_5668(.VSS(VSS),.VDD(VDD),.Y(g6970),.A(I11122));
  NOT NOT1_5669(.VSS(VSS),.VDD(VDD),.Y(g8347),.A(I13421));
  NOT NOT1_5670(.VSS(VSS),.VDD(VDD),.Y(I15395),.A(g10058));
  NOT NOT1_5671(.VSS(VSS),.VDD(VDD),.Y(g2317),.A(g622));
  NOT NOT1_5672(.VSS(VSS),.VDD(VDD),.Y(I8892),.A(g4554));
  NOT NOT1_5673(.VSS(VSS),.VDD(VDD),.Y(g10129),.A(I15389));
  NOT NOT1_5674(.VSS(VSS),.VDD(VDD),.Y(g9930),.A(I15127));
  NOT NOT1_5675(.VSS(VSS),.VDD(VDD),.Y(I9114),.A(g5603));
  NOT NOT1_5676(.VSS(VSS),.VDD(VDD),.Y(g6925),.A(I11043));
  NOT NOT1_5677(.VSS(VSS),.VDD(VDD),.Y(I17194),.A(g11317));
  NOT NOT1_5678(.VSS(VSS),.VDD(VDD),.Y(I7707),.A(g3370));
  NOT NOT1_5679(.VSS(VSS),.VDD(VDD),.Y(g11395),.A(I17228));
  NOT NOT1_5680(.VSS(VSS),.VDD(VDD),.Y(g1962),.A(g27));
  NOT NOT1_5681(.VSS(VSS),.VDD(VDD),.Y(g10057),.A(I15278));
  NOT NOT1_5682(.VSS(VSS),.VDD(VDD),.Y(g2601),.A(I5704));
  NOT NOT1_5683(.VSS(VSS),.VDD(VDD),.Y(g10128),.A(I15386));
  NOT NOT1_5684(.VSS(VSS),.VDD(VDD),.Y(g5818),.A(g5320));
  NOT NOT1_5685(.VSS(VSS),.VDD(VDD),.Y(g8697),.A(g8660));
  NOT NOT1_5686(.VSS(VSS),.VDD(VDD),.Y(I6520),.A(g3186));
  NOT NOT1_5687(.VSS(VSS),.VDD(VDD),.Y(I14668),.A(g9309));
  NOT NOT1_5688(.VSS(VSS),.VDD(VDD),.Y(g4213),.A(I7456));
  NOT NOT1_5689(.VSS(VSS),.VDD(VDD),.Y(g11633),.A(I17713));
  NOT NOT1_5690(.VSS(VSS),.VDD(VDD),.Y(I11659),.A(g7097));
  NOT NOT1_5691(.VSS(VSS),.VDD(VDD),.Y(I12186),.A(g7264));
  NOT NOT1_5692(.VSS(VSS),.VDD(VDD),.Y(g6120),.A(I9813));
  NOT NOT1_5693(.VSS(VSS),.VDD(VDD),.Y(I10195),.A(g6116));
  NOT NOT1_5694(.VSS(VSS),.VDD(VDD),.Y(I6031),.A(g2209));
  NOT NOT1_5695(.VSS(VSS),.VDD(VDD),.Y(I12953),.A(g8024));
  NOT NOT1_5696(.VSS(VSS),.VDD(VDD),.Y(g10323),.A(I15763));
  NOT NOT1_5697(.VSS(VSS),.VDD(VDD),.Y(g11191),.A(g11112));
  NOT NOT1_5698(.VSS(VSS),.VDD(VDD),.Y(g2775),.A(I5862));
  NOT NOT1_5699(.VSS(VSS),.VDD(VDD),.Y(g7076),.A(I11303));
  NOT NOT1_5700(.VSS(VSS),.VDD(VDD),.Y(I6812),.A(g3290));
  NOT NOT1_5701(.VSS(VSS),.VDD(VDD),.Y(g3783),.A(I7009));
  NOT NOT1_5702(.VSS(VSS),.VDD(VDD),.Y(g7476),.A(g6933));
  NOT NOT1_5703(.VSS(VSS),.VDD(VDD),.Y(I6958),.A(g2872));
  NOT NOT1_5704(.VSS(VSS),.VDD(VDD),.Y(g5893),.A(g5106));
  NOT NOT1_5705(.VSS(VSS),.VDD(VDD),.Y(g6277),.A(I10090));
  NOT NOT1_5706(.VSS(VSS),.VDD(VDD),.Y(I14525),.A(g9109));
  NOT NOT1_5707(.VSS(VSS),.VDD(VDD),.Y(I14424),.A(g8945));
  NOT NOT1_5708(.VSS(VSS),.VDD(VDD),.Y(g3112),.A(g2482));
  NOT NOT1_5709(.VSS(VSS),.VDD(VDD),.Y(g3267),.A(I6439));
  NOT NOT1_5710(.VSS(VSS),.VDD(VDD),.Y(g10775),.A(I16461));
  NOT NOT1_5711(.VSS(VSS),.VDD(VDD),.Y(I16766),.A(g10892));
  NOT NOT1_5712(.VSS(VSS),.VDD(VDD),.Y(I12936),.A(g7983));
  NOT NOT1_5713(.VSS(VSS),.VDD(VDD),.Y(I15832),.A(g10206));
  NOT NOT1_5714(.VSS(VSS),.VDD(VDD),.Y(I8340),.A(g4804));
  NOT NOT1_5715(.VSS(VSS),.VDD(VDD),.Y(I11296),.A(g6525));
  NOT NOT1_5716(.VSS(VSS),.VDD(VDD),.Y(g2060),.A(g1380));
  NOT NOT1_5717(.VSS(VSS),.VDD(VDD),.Y(g6617),.A(g6019));
  NOT NOT1_5718(.VSS(VSS),.VDD(VDD),.Y(I14558),.A(g9024));
  NOT NOT1_5719(.VSS(VSS),.VDD(VDD),.Y(g6789),.A(I10789));
  NOT NOT1_5720(.VSS(VSS),.VDD(VDD),.Y(I17749),.A(g11644));
  NOT NOT1_5721(.VSS(VSS),.VDD(VDD),.Y(I11644),.A(g6970));
  NOT NOT1_5722(.VSS(VSS),.VDD(VDD),.Y(I17616),.A(g11561));
  NOT NOT1_5723(.VSS(VSS),.VDD(VDD),.Y(I16871),.A(g10973));
  NOT NOT1_5724(.VSS(VSS),.VDD(VDD),.Y(I11338),.A(g6680));
  NOT NOT1_5725(.VSS(VSS),.VDD(VDD),.Y(I13338),.A(g8210));
  NOT NOT1_5726(.VSS(VSS),.VDD(VDD),.Y(I9594),.A(g5083));
  NOT NOT1_5727(.VSS(VSS),.VDD(VDD),.Y(g4166),.A(I7315));
  NOT NOT1_5728(.VSS(VSS),.VDD(VDD),.Y(g11440),.A(I17371));
  NOT NOT1_5729(.VSS(VSS),.VDD(VDD),.Y(g4366),.A(I7659));
  NOT NOT1_5730(.VSS(VSS),.VDD(VDD),.Y(g5426),.A(I8869));
  NOT NOT1_5731(.VSS(VSS),.VDD(VDD),.Y(I15861),.A(g10339));
  NOT NOT1_5732(.VSS(VSS),.VDD(VDD),.Y(I16360),.A(g10590));
  NOT NOT1_5733(.VSS(VSS),.VDD(VDD),.Y(I6911),.A(g2825));
  NOT NOT1_5734(.VSS(VSS),.VDD(VDD),.Y(I13969),.A(g8451));
  NOT NOT1_5735(.VSS(VSS),.VDD(VDD),.Y(I7833),.A(g3585));
  NOT NOT1_5736(.VSS(VSS),.VDD(VDD),.Y(g7285),.A(I11531));
  NOT NOT1_5737(.VSS(VSS),.VDD(VDD),.Y(g3329),.A(I6504));
  NOT NOT1_5738(.VSS(VSS),.VDD(VDD),.Y(I15247),.A(g10032));
  NOT NOT1_5739(.VSS(VSS),.VDD(VDD),.Y(g11573),.A(g11561));
  NOT NOT1_5740(.VSS(VSS),.VDD(VDD),.Y(I5525),.A(g589));
  NOT NOT1_5741(.VSS(VSS),.VDD(VDD),.Y(I5710),.A(g2431));
  NOT NOT1_5742(.VSS(VSS),.VDD(VDD),.Y(g3761),.A(I6962));
  NOT NOT1_5743(.VSS(VSS),.VDD(VDD),.Y(g5614),.A(I9040));
  NOT NOT1_5744(.VSS(VSS),.VDD(VDD),.Y(I12762),.A(g7541));
  NOT NOT1_5745(.VSS(VSS),.VDD(VDD),.Y(I17704),.A(g11618));
  NOT NOT1_5746(.VSS(VSS),.VDD(VDD),.Y(g4056),.A(I7173));
  NOT NOT1_5747(.VSS(VSS),.VDD(VDD),.Y(g7500),.A(g6943));
  NOT NOT1_5748(.VSS(VSS),.VDD(VDD),.Y(I10713),.A(g6003));
  NOT NOT1_5749(.VSS(VSS),.VDD(VDD),.Y(g8317),.A(I13335));
  NOT NOT1_5750(.VSS(VSS),.VDD(VDD),.Y(I15389),.A(g10110));
  NOT NOT1_5751(.VSS(VSS),.VDD(VDD),.Y(g4456),.A(g3375));
  NOT NOT1_5752(.VSS(VSS),.VDD(VDD),.Y(I14713),.A(g9052));
  NOT NOT1_5753(.VSS(VSS),.VDD(VDD),.Y(g6299),.A(I10156));
  NOT NOT1_5754(.VSS(VSS),.VDD(VDD),.Y(g5821),.A(I9433));
  NOT NOT1_5755(.VSS(VSS),.VDD(VDD),.Y(g3828),.A(g2920));
  NOT NOT1_5756(.VSS(VSS),.VDD(VDD),.Y(g10697),.A(I16370));
  NOT NOT1_5757(.VSS(VSS),.VDD(VDD),.Y(g6547),.A(g5893));
  NOT NOT1_5758(.VSS(VSS),.VDD(VDD),.Y(I13197),.A(g8186));
  NOT NOT1_5759(.VSS(VSS),.VDD(VDD),.Y(g11389),.A(I17216));
  NOT NOT1_5760(.VSS(VSS),.VDD(VDD),.Y(g11045),.A(I16796));
  NOT NOT1_5761(.VSS(VSS),.VDD(VDD),.Y(I6733),.A(g3321));
  NOT NOT1_5762(.VSS(VSS),.VDD(VDD),.Y(I9065),.A(g4760));
  NOT NOT1_5763(.VSS(VSS),.VDD(VDD),.Y(I17466),.A(g11447));
  NOT NOT1_5764(.VSS(VSS),.VDD(VDD),.Y(g8601),.A(g8477));
  NOT NOT1_5765(.VSS(VSS),.VDD(VDD),.Y(g10261),.A(g10126));
  NOT NOT1_5766(.VSS(VSS),.VDD(VDD),.Y(g2937),.A(I6106));
  NOT NOT1_5767(.VSS(VSS),.VDD(VDD),.Y(g3727),.A(I6901));
  NOT NOT1_5768(.VSS(VSS),.VDD(VDD),.Y(g2079),.A(I4891));
  NOT NOT1_5769(.VSS(VSS),.VDD(VDD),.Y(g5984),.A(I9602));
  NOT NOT1_5770(.VSS(VSS),.VDD(VDD),.Y(I10610),.A(g5879));
  NOT NOT1_5771(.VSS(VSS),.VDD(VDD),.Y(g10880),.A(I16610));
  NOT NOT1_5772(.VSS(VSS),.VDD(VDD),.Y(I15701),.A(g10236));
  NOT NOT1_5773(.VSS(VSS),.VDD(VDD),.Y(g4355),.A(I7642));
  NOT NOT1_5774(.VSS(VSS),.VDD(VDD),.Y(g11388),.A(I17213));
  NOT NOT1_5775(.VSS(VSS),.VDD(VDD),.Y(g7339),.A(I11665));
  NOT NOT1_5776(.VSS(VSS),.VDD(VDD),.Y(g2479),.A(g26));
  NOT NOT1_5777(.VSS(VSS),.VDD(VDD),.Y(I10042),.A(g5723));
  NOT NOT1_5778(.VSS(VSS),.VDD(VDD),.Y(I15272),.A(g10019));
  NOT NOT1_5779(.VSS(VSS),.VDD(VDD),.Y(I16629),.A(g10860));
  NOT NOT1_5780(.VSS(VSS),.VDD(VDD),.Y(g2840),.A(I5960));
  NOT NOT1_5781(.VSS(VSS),.VDD(VDD),.Y(I10189),.A(g6112));
  NOT NOT1_5782(.VSS(VSS),.VDD(VDD),.Y(g7024),.A(I11169));
  NOT NOT1_5783(.VSS(VSS),.VDD(VDD),.Y(I16220),.A(g10502));
  NOT NOT1_5784(.VSS(VSS),.VDD(VDD),.Y(g2190),.A(I5149));
  NOT NOT1_5785(.VSS(VSS),.VDD(VDD),.Y(g4260),.A(I7513));
  NOT NOT1_5786(.VSS(VSS),.VDD(VDD),.Y(g2390),.A(I5475));
  NOT NOT1_5787(.VSS(VSS),.VDD(VDD),.Y(g7795),.A(I12550));
  NOT NOT1_5788(.VSS(VSS),.VDD(VDD),.Y(I9433),.A(g5069));
  NOT NOT1_5789(.VSS(VSS),.VDD(VDD),.Y(I17642),.A(g11579));
  NOT NOT1_5790(.VSS(VSS),.VDD(VDD),.Y(I10678),.A(g5777));
  NOT NOT1_5791(.VSS(VSS),.VDD(VDD),.Y(g7737),.A(I12388));
  NOT NOT1_5792(.VSS(VSS),.VDD(VDD),.Y(g7809),.A(I12592));
  NOT NOT1_5793(.VSS(VSS),.VDD(VDD),.Y(g3703),.A(g2920));
  NOT NOT1_5794(.VSS(VSS),.VDD(VDD),.Y(I14188),.A(g8792));
  NOT NOT1_5795(.VSS(VSS),.VDD(VDD),.Y(I14678),.A(g9265));
  NOT NOT1_5796(.VSS(VSS),.VDD(VDD),.Y(g5106),.A(I8490));
  NOT NOT1_5797(.VSS(VSS),.VDD(VDD),.Y(g4463),.A(g3829));
  NOT NOT1_5798(.VSS(VSS),.VDD(VDD),.Y(I9096),.A(g5568));
  NOT NOT1_5799(.VSS(VSS),.VDD(VDD),.Y(g2156),.A(I5073));
  NOT NOT1_5800(.VSS(VSS),.VDD(VDD),.Y(g7672),.A(I12293));
  NOT NOT1_5801(.VSS(VSS),.VDD(VDD),.Y(I14939),.A(g9454));
  NOT NOT1_5802(.VSS(VSS),.VDD(VDD),.Y(g2356),.A(I5438));
  NOT NOT1_5803(.VSS(VSS),.VDD(VDD),.Y(g7077),.A(I11306));
  NOT NOT1_5804(.VSS(VSS),.VDD(VDD),.Y(g6709),.A(g5949));
  NOT NOT1_5805(.VSS(VSS),.VDD(VDD),.Y(I17733),.A(g11639));
  NOT NOT1_5806(.VSS(VSS),.VDD(VDD),.Y(g9814),.A(g9490));
  NOT NOT1_5807(.VSS(VSS),.VDD(VDD),.Y(g5790),.A(I9388));
  NOT NOT1_5808(.VSS(VSS),.VDD(VDD),.Y(I9550),.A(g5030));
  NOT NOT1_5809(.VSS(VSS),.VDD(VDD),.Y(I10030),.A(g5685));
  NOT NOT1_5810(.VSS(VSS),.VDD(VDD),.Y(g7477),.A(I11869));
  NOT NOT1_5811(.VSS(VSS),.VDD(VDD),.Y(I10093),.A(g5779));
  NOT NOT1_5812(.VSS(VSS),.VDD(VDD),.Y(I9845),.A(g5405));
  NOT NOT1_5813(.VSS(VSS),.VDD(VDD),.Y(g3624),.A(I6767));
  NOT NOT1_5814(.VSS(VSS),.VDD(VDD),.Y(g6140),.A(I9851));
  NOT NOT1_5815(.VSS(VSS),.VDD(VDD),.Y(g6340),.A(I10243));
  NOT NOT1_5816(.VSS(VSS),.VDD(VDD),.Y(I5111),.A(g39));
  NOT NOT1_5817(.VSS(VSS),.VDD(VDD),.Y(I11581),.A(g6826));
  NOT NOT1_5818(.VSS(VSS),.VDD(VDD),.Y(I11450),.A(g6488));
  NOT NOT1_5819(.VSS(VSS),.VDD(VDD),.Y(I12568),.A(g7502));
  NOT NOT1_5820(.VSS(VSS),.VDD(VDD),.Y(g9350),.A(I14555));
  NOT NOT1_5821(.VSS(VSS),.VDD(VDD),.Y(g10499),.A(I16124));
  NOT NOT1_5822(.VSS(VSS),.VDD(VDD),.Y(I5311),.A(g98));
  NOT NOT1_5823(.VSS(VSS),.VDD(VDD),.Y(g3068),.A(g2303));
  NOT NOT1_5824(.VSS(VSS),.VDD(VDD),.Y(I13714),.A(g8351));
  NOT NOT1_5825(.VSS(VSS),.VDD(VDD),.Y(I11315),.A(g6644));
  NOT NOT1_5826(.VSS(VSS),.VDD(VDD),.Y(g8784),.A(I14087));
  NOT NOT1_5827(.VSS(VSS),.VDD(VDD),.Y(g2942),.A(I6121));
  NOT NOT1_5828(.VSS(VSS),.VDD(VDD),.Y(g8739),.A(g8640));
  NOT NOT1_5829(.VSS(VSS),.VDD(VDD),.Y(I12242),.A(g7089));
  NOT NOT1_5830(.VSS(VSS),.VDD(VDD),.Y(g4279),.A(I7536));
  NOT NOT1_5831(.VSS(VSS),.VDD(VDD),.Y(I11707),.A(g7009));
  NOT NOT1_5832(.VSS(VSS),.VDD(VDD),.Y(g7205),.A(I11433));
  NOT NOT1_5833(.VSS(VSS),.VDD(VDD),.Y(g9773),.A(g9474));
  NOT NOT1_5834(.VSS(VSS),.VDD(VDD),.Y(I7086),.A(g3142));
  NOT NOT1_5835(.VSS(VSS),.VDD(VDD),.Y(I13819),.A(g8488));
  NOT NOT1_5836(.VSS(VSS),.VDD(VDD),.Y(g11061),.A(g10974));
  NOT NOT1_5837(.VSS(VSS),.VDD(VDD),.Y(g10498),.A(I16121));
  NOT NOT1_5838(.VSS(VSS),.VDD(VDD),.Y(g9009),.A(I14405));
  NOT NOT1_5839(.VSS(VSS),.VDD(VDD),.Y(g6435),.A(I10355));
  NOT NOT1_5840(.VSS(VSS),.VDD(VDD),.Y(g4167),.A(I7318));
  NOT NOT1_5841(.VSS(VSS),.VDD(VDD),.Y(g5027),.A(I8396));
  NOT NOT1_5842(.VSS(VSS),.VDD(VDD),.Y(g6517),.A(I10434));
  NOT NOT1_5843(.VSS(VSS),.VDD(VDD),.Y(g6082),.A(I9727));
  NOT NOT1_5844(.VSS(VSS),.VDD(VDD),.Y(I12123),.A(g6861));
  NOT NOT1_5845(.VSS(VSS),.VDD(VDD),.Y(g4318),.A(g4130));
  NOT NOT1_5846(.VSS(VSS),.VDD(VDD),.Y(g4367),.A(I7662));
  NOT NOT1_5847(.VSS(VSS),.VDD(VDD),.Y(I16859),.A(g10911));
  NOT NOT1_5848(.VSS(VSS),.VDD(VDD),.Y(g4872),.A(I8211));
  NOT NOT1_5849(.VSS(VSS),.VDD(VDD),.Y(g7634),.A(I12242));
  NOT NOT1_5850(.VSS(VSS),.VDD(VDD),.Y(I5174),.A(g52));
  NOT NOT1_5851(.VSS(VSS),.VDD(VDD),.Y(I16950),.A(g11081));
  NOT NOT1_5852(.VSS(VSS),.VDD(VDD),.Y(g8079),.A(I12939));
  NOT NOT1_5853(.VSS(VSS),.VDD(VDD),.Y(I16370),.A(g10592));
  NOT NOT1_5854(.VSS(VSS),.VDD(VDD),.Y(g6482),.A(I10412));
  NOT NOT1_5855(.VSS(VSS),.VDD(VDD),.Y(I11055),.A(g6419));
  NOT NOT1_5856(.VSS(VSS),.VDD(VDD),.Y(g10056),.A(I15275));
  NOT NOT1_5857(.VSS(VSS),.VDD(VDD),.Y(I9807),.A(g5419));
  NOT NOT1_5858(.VSS(VSS),.VDD(VDD),.Y(g8479),.A(g8319));
  NOT NOT1_5859(.VSS(VSS),.VDD(VDD),.Y(I7185),.A(g2626));
  NOT NOT1_5860(.VSS(VSS),.VDD(VDD),.Y(I12751),.A(g7626));
  NOT NOT1_5861(.VSS(VSS),.VDD(VDD),.Y(g9769),.A(I14918));
  NOT NOT1_5862(.VSS(VSS),.VDD(VDD),.Y(g4057),.A(I7176));
  NOT NOT1_5863(.VSS(VSS),.VDD(VDD),.Y(g5904),.A(I9539));
  NOT NOT1_5864(.VSS(VSS),.VDD(VDD),.Y(g7304),.A(I11560));
  NOT NOT1_5865(.VSS(VSS),.VDD(VDD),.Y(g5200),.A(g4567));
  NOT NOT1_5866(.VSS(VSS),.VDD(VDD),.Y(g10080),.A(I15308));
  NOT NOT1_5867(.VSS(VSS),.VDD(VDD),.Y(g8294),.A(I13236));
  NOT NOT1_5868(.VSS(VSS),.VDD(VDD),.Y(I13978),.A(g8575));
  NOT NOT1_5869(.VSS(VSS),.VDD(VDD),.Y(g4457),.A(g3829));
  NOT NOT1_5870(.VSS(VSS),.VDD(VDD),.Y(g2163),.A(I5092));
  NOT NOT1_5871(.VSS(VSS),.VDD(VDD),.Y(I8877),.A(g4421));
  NOT NOT1_5872(.VSS(VSS),.VDD(VDD),.Y(g2363),.A(I5441));
  NOT NOT1_5873(.VSS(VSS),.VDD(VDD),.Y(I7070),.A(g3138));
  NOT NOT1_5874(.VSS(VSS),.VDD(VDD),.Y(g5446),.A(I8877));
  NOT NOT1_5875(.VSS(VSS),.VDD(VDD),.Y(I11590),.A(g6829));
  NOT NOT1_5876(.VSS(VSS),.VDD(VDD),.Y(I16172),.A(g10498));
  NOT NOT1_5877(.VSS(VSS),.VDD(VDD),.Y(g4193),.A(I7396));
  NOT NOT1_5878(.VSS(VSS),.VDD(VDD),.Y(g3716),.A(I6876));
  NOT NOT1_5879(.VSS(VSS),.VDD(VDD),.Y(g11360),.A(I17185));
  NOT NOT1_5880(.VSS(VSS),.VDD(VDD),.Y(g4393),.A(I7726));
  NOT NOT1_5881(.VSS(VSS),.VDD(VDD),.Y(I10837),.A(g6717));
  NOT NOT1_5882(.VSS(VSS),.VDD(VDD),.Y(g2432),.A(I5513));
  NOT NOT1_5883(.VSS(VSS),.VDD(VDD),.Y(I12293),.A(g7116));
  NOT NOT1_5884(.VSS(VSS),.VDD(VDD),.Y(g10271),.A(I15665));
  NOT NOT1_5885(.VSS(VSS),.VDD(VDD),.Y(I12638),.A(g7708));
  NOT NOT1_5886(.VSS(VSS),.VDD(VDD),.Y(g11447),.A(I17390));
  NOT NOT1_5887(.VSS(VSS),.VDD(VDD),.Y(I13741),.A(g8296));
  NOT NOT1_5888(.VSS(VSS),.VDD(VDD),.Y(I15162),.A(g9958));
  NOT NOT1_5889(.VSS(VSS),.VDD(VDD),.Y(g4549),.A(I7956));
  NOT NOT1_5890(.VSS(VSS),.VDD(VDD),.Y(I17555),.A(g11503));
  NOT NOT1_5891(.VSS(VSS),.VDD(VDD),.Y(I6898),.A(g2964));
  NOT NOT1_5892(.VSS(VSS),.VDD(VDD),.Y(I12265),.A(g7211));
  NOT NOT1_5893(.VSS(VSS),.VDD(VDD),.Y(g11162),.A(g10950));
  NOT NOT1_5894(.VSS(VSS),.VDD(VDD),.Y(g7754),.A(I12427));
  NOT NOT1_5895(.VSS(VSS),.VDD(VDD),.Y(g10461),.A(I15974));
  NOT NOT1_5896(.VSS(VSS),.VDD(VDD),.Y(g5191),.A(g4640));
  NOT NOT1_5897(.VSS(VSS),.VDD(VDD),.Y(g8156),.A(I13051));
  NOT NOT1_5898(.VSS(VSS),.VDD(VDD),.Y(I9248),.A(g4954));
  NOT NOT1_5899(.VSS(VSS),.VDD(VDD),.Y(g3747),.A(g3015));
  NOT NOT1_5900(.VSS(VSS),.VDD(VDD),.Y(I11094),.A(g6657));
  NOT NOT1_5901(.VSS(VSS),.VDD(VDD),.Y(g1973),.A(g466));
  NOT NOT1_5902(.VSS(VSS),.VDD(VDD),.Y(g5391),.A(I8827));
  NOT NOT1_5903(.VSS(VSS),.VDD(VDD),.Y(g8356),.A(I13448));
  NOT NOT1_5904(.VSS(VSS),.VDD(VDD),.Y(g10342),.A(I15792));
  NOT NOT1_5905(.VSS(VSS),.VDD(VDD),.Y(g3398),.A(g2896));
  NOT NOT1_5906(.VSS(VSS),.VDD(VDD),.Y(g6214),.A(g5446));
  NOT NOT1_5907(.VSS(VSS),.VDD(VDD),.Y(g7273),.A(g6365));
  NOT NOT1_5908(.VSS(VSS),.VDD(VDD),.Y(I5020),.A(g1176));
  NOT NOT1_5909(.VSS(VSS),.VDD(VDD),.Y(I6510),.A(g3267));
  NOT NOT1_5910(.VSS(VSS),.VDD(VDD),.Y(g9993),.A(I15193));
  NOT NOT1_5911(.VSS(VSS),.VDD(VDD),.Y(g10145),.A(I15437));
  NOT NOT1_5912(.VSS(VSS),.VDD(VDD),.Y(g10031),.A(I15229));
  NOT NOT1_5913(.VSS(VSS),.VDD(VDD),.Y(g6110),.A(I9783));
  NOT NOT1_5914(.VSS(VSS),.VDD(VDD),.Y(g5637),.A(I9074));
  NOT NOT1_5915(.VSS(VSS),.VDD(VDD),.Y(g6310),.A(I10189));
  NOT NOT1_5916(.VSS(VSS),.VDD(VDD),.Y(g11629),.A(I17701));
  NOT NOT1_5917(.VSS(VSS),.VDD(VDD),.Y(g9822),.A(I14967));
  NOT NOT1_5918(.VSS(VSS),.VDD(VDD),.Y(g10199),.A(g10172));
  NOT NOT1_5919(.VSS(VSS),.VDD(VDD),.Y(g11451),.A(I17410));
  NOT NOT1_5920(.VSS(VSS),.VDD(VDD),.Y(g11472),.A(I17453));
  NOT NOT1_5921(.VSS(VSS),.VDD(VDD),.Y(g7044),.A(I11217));
  NOT NOT1_5922(.VSS(VSS),.VDD(VDD),.Y(g10887),.A(I16623));
  NOT NOT1_5923(.VSS(VSS),.VDD(VDD),.Y(g2912),.A(I6085));
  NOT NOT1_5924(.VSS(VSS),.VDD(VDD),.Y(I13735),.A(g8293));
  NOT NOT1_5925(.VSS(VSS),.VDD(VDD),.Y(g1969),.A(g456));
  NOT NOT1_5926(.VSS(VSS),.VDD(VDD),.Y(g4121),.A(I7264));
  NOT NOT1_5927(.VSS(VSS),.VDD(VDD),.Y(g5107),.A(g4459));
  NOT NOT1_5928(.VSS(VSS),.VDD(VDD),.Y(g8704),.A(g8667));
  NOT NOT1_5929(.VSS(VSS),.VDD(VDD),.Y(g4321),.A(g3863));
  NOT NOT1_5930(.VSS(VSS),.VDD(VDD),.Y(g2157),.A(g1703));
  NOT NOT1_5931(.VSS(VSS),.VDD(VDD),.Y(g11628),.A(I17698));
  NOT NOT1_5932(.VSS(VSS),.VDD(VDD),.Y(g10198),.A(I15568));
  NOT NOT1_5933(.VSS(VSS),.VDD(VDD),.Y(I7131),.A(g2640));
  NOT NOT1_5934(.VSS(VSS),.VDD(VDD),.Y(I7006),.A(g2912));
  NOT NOT1_5935(.VSS(VSS),.VDD(VDD),.Y(g7983),.A(I12793));
  NOT NOT1_5936(.VSS(VSS),.VDD(VDD),.Y(I10201),.A(g5998));
  NOT NOT1_5937(.VSS(VSS),.VDD(VDD),.Y(g5223),.A(g4640));
  NOT NOT1_5938(.VSS(VSS),.VDD(VDD),.Y(I11695),.A(g7052));
  NOT NOT1_5939(.VSS(VSS),.VDD(VDD),.Y(g10528),.A(g10464));
  NOT NOT1_5940(.VSS(VSS),.VDD(VDD),.Y(g10696),.A(g10621));
  NOT NOT1_5941(.VSS(VSS),.VDD(VDD),.Y(g4232),.A(I7487));
  NOT NOT1_5942(.VSS(VSS),.VDD(VDD),.Y(I12835),.A(g7660));
  NOT NOT1_5943(.VSS(VSS),.VDD(VDD),.Y(I13695),.A(g8363));
  NOT NOT1_5944(.VSS(VSS),.VDD(VDD),.Y(g10330),.A(I15778));
  NOT NOT1_5945(.VSS(VSS),.VDD(VDD),.Y(g5858),.A(I9475));
  NOT NOT1_5946(.VSS(VSS),.VDD(VDD),.Y(g10393),.A(g10317));
  NOT NOT1_5947(.VSS(VSS),.VDD(VDD),.Y(I10075),.A(g5724));
  NOT NOT1_5948(.VSS(VSS),.VDD(VDD),.Y(I7766),.A(g3770));
  NOT NOT1_5949(.VSS(VSS),.VDD(VDD),.Y(g8954),.A(I14315));
  NOT NOT1_5950(.VSS(VSS),.VDD(VDD),.Y(I16540),.A(g10722));
  NOT NOT1_5951(.VSS(VSS),.VDD(VDD),.Y(g6236),.A(I9981));
  NOT NOT1_5952(.VSS(VSS),.VDD(VDD),.Y(I6694),.A(g2749));
  NOT NOT1_5953(.VSS(VSS),.VDD(VDD),.Y(g7543),.A(I11961));
  NOT NOT1_5954(.VSS(VSS),.VDD(VDD),.Y(I12586),.A(g7561));
  NOT NOT1_5955(.VSS(VSS),.VDD(VDD),.Y(g11071),.A(g10913));
  NOT NOT1_5956(.VSS(VSS),.VDD(VDD),.Y(g8363),.A(I13469));
  NOT NOT1_5957(.VSS(VSS),.VDD(VDD),.Y(I7487),.A(g3371));
  NOT NOT1_5958(.VSS(VSS),.VDD(VDD),.Y(I8237),.A(g4295));
  NOT NOT1_5959(.VSS(VSS),.VDD(VDD),.Y(g5416),.A(I8851));
  NOT NOT1_5960(.VSS(VSS),.VDD(VDD),.Y(I14494),.A(g8887));
  NOT NOT1_5961(.VSS(VSS),.VDD(VDD),.Y(g3119),.A(I6347));
  NOT NOT1_5962(.VSS(VSS),.VDD(VDD),.Y(g10132),.A(g10063));
  NOT NOT1_5963(.VSS(VSS),.VDD(VDD),.Y(I17519),.A(g11484));
  NOT NOT1_5964(.VSS(VSS),.VDD(VDD),.Y(g10869),.A(I16577));
  NOT NOT1_5965(.VSS(VSS),.VDD(VDD),.Y(I6088),.A(g2235));
  NOT NOT1_5966(.VSS(VSS),.VDD(VDD),.Y(I17176),.A(g11286));
  NOT NOT1_5967(.VSS(VSS),.VDD(VDD),.Y(I17185),.A(g11311));
  NOT NOT1_5968(.VSS(VSS),.VDD(VDD),.Y(I10623),.A(g6002));
  NOT NOT1_5969(.VSS(VSS),.VDD(VDD),.Y(I12442),.A(g7672));
  NOT NOT1_5970(.VSS(VSS),.VDD(VDD),.Y(I17675),.A(g11606));
  NOT NOT1_5971(.VSS(VSS),.VDD(VDD),.Y(I17092),.A(g11217));
  NOT NOT1_5972(.VSS(VSS),.VDD(VDD),.Y(I16203),.A(g10454));
  NOT NOT1_5973(.VSS(VSS),.VDD(VDD),.Y(g4519),.A(I7920));
  NOT NOT1_5974(.VSS(VSS),.VDD(VDD),.Y(g5251),.A(g4640));
  NOT NOT1_5975(.VSS(VSS),.VDD(VDD),.Y(g6590),.A(g5949));
  NOT NOT1_5976(.VSS(VSS),.VDD(VDD),.Y(g6877),.A(I10963));
  NOT NOT1_5977(.VSS(VSS),.VDD(VDD),.Y(I4777),.A(g18));
  NOT NOT1_5978(.VSS(VSS),.VDD(VDD),.Y(g10868),.A(I16574));
  NOT NOT1_5979(.VSS(VSS),.VDD(VDD),.Y(g5811),.A(I9415));
  NOT NOT1_5980(.VSS(VSS),.VDD(VDD),.Y(g5642),.A(I9087));
  NOT NOT1_5981(.VSS(VSS),.VDD(VDD),.Y(g3352),.A(I6538));
  NOT NOT1_5982(.VSS(VSS),.VDD(VDD),.Y(I9783),.A(g5395));
  NOT NOT1_5983(.VSS(VSS),.VDD(VDD),.Y(g2626),.A(g2000));
  NOT NOT1_5984(.VSS(VSS),.VDD(VDD),.Y(g7534),.A(I11942));
  NOT NOT1_5985(.VSS(VSS),.VDD(VDD),.Y(g7729),.A(I12372));
  NOT NOT1_5986(.VSS(VSS),.VDD(VDD),.Y(g7961),.A(g7664));
  NOT NOT1_5987(.VSS(VSS),.VDD(VDD),.Y(g5047),.A(g4354));
  NOT NOT1_5988(.VSS(VSS),.VDD(VDD),.Y(I13457),.A(g8184));
  NOT NOT1_5989(.VSS(VSS),.VDD(VDD),.Y(I10984),.A(g6757));
  NOT NOT1_5990(.VSS(VSS),.VDD(VDD),.Y(g9895),.A(I15088));
  NOT NOT1_5991(.VSS(VSS),.VDD(VDD),.Y(g6657),.A(I10620));
  NOT NOT1_5992(.VSS(VSS),.VDD(VDD),.Y(g10161),.A(I15479));
  NOT NOT1_5993(.VSS(VSS),.VDD(VDD),.Y(g4552),.A(g3880));
  NOT NOT1_5994(.VSS(VSS),.VDD(VDD),.Y(g4606),.A(g3829));
  NOT NOT1_5995(.VSS(VSS),.VDD(VDD),.Y(I15858),.A(g10336));
  NOT NOT1_5996(.VSS(VSS),.VDD(VDD),.Y(g8568),.A(I13797));
  NOT NOT1_5997(.VSS(VSS),.VDD(VDD),.Y(I8089),.A(g3545));
  NOT NOT1_5998(.VSS(VSS),.VDD(VDD),.Y(I10352),.A(g6216));
  NOT NOT1_5999(.VSS(VSS),.VDD(VDD),.Y(g6556),.A(g5747));
  NOT NOT1_6000(.VSS(VSS),.VDD(VDD),.Y(I14352),.A(g8946));
  NOT NOT1_6001(.VSS(VSS),.VDD(VDD),.Y(g7927),.A(g7500));
  NOT NOT1_6002(.VSS(VSS),.VDD(VDD),.Y(I10822),.A(g6584));
  NOT NOT1_6003(.VSS(VSS),.VDD(VDD),.Y(g5874),.A(I9491));
  NOT NOT1_6004(.VSS(VSS),.VDD(VDD),.Y(I9001),.A(g4762));
  NOT NOT1_6005(.VSS(VSS),.VDD(VDD),.Y(g10259),.A(g10141));
  NOT NOT1_6006(.VSS(VSS),.VDD(VDD),.Y(I14418),.A(g8941));
  NOT NOT1_6007(.VSS(VSS),.VDD(VDD),.Y(g10708),.A(I16387));
  NOT NOT1_6008(.VSS(VSS),.VDD(VDD),.Y(I16739),.A(g10856));
  NOT NOT1_6009(.VSS(VSS),.VDD(VDD),.Y(I12430),.A(g7649));
  NOT NOT1_6010(.VSS(VSS),.VDD(VDD),.Y(g3186),.A(I6373));
  NOT NOT1_6011(.VSS(VSS),.VDD(VDD),.Y(g5654),.A(I9123));
  NOT NOT1_6012(.VSS(VSS),.VDD(VDD),.Y(I12493),.A(g7650));
  NOT NOT1_6013(.VSS(VSS),.VDD(VDD),.Y(g10471),.A(g10378));
  NOT NOT1_6014(.VSS(VSS),.VDD(VDD),.Y(g7414),.A(I11794));
  NOT NOT1_6015(.VSS(VSS),.VDD(VDD),.Y(I9293),.A(g5486));
  NOT NOT1_6016(.VSS(VSS),.VDD(VDD),.Y(g3386),.A(g3144));
  NOT NOT1_6017(.VSS(VSS),.VDD(VDD),.Y(g10087),.A(I15314));
  NOT NOT1_6018(.VSS(VSS),.VDD(VDD),.Y(g8357),.A(I13451));
  NOT NOT1_6019(.VSS(VSS),.VDD(VDD),.Y(I9129),.A(g4892));
  NOT NOT1_6020(.VSS(VSS),.VDD(VDD),.Y(g7946),.A(g7416));
  NOT NOT1_6021(.VSS(VSS),.VDD(VDD),.Y(g10258),.A(g10198));
  NOT NOT1_6022(.VSS(VSS),.VDD(VDD),.Y(g3975),.A(g3121));
  NOT NOT1_6023(.VSS(VSS),.VDD(VDD),.Y(I7173),.A(g2644));
  NOT NOT1_6024(.VSS(VSS),.VDD(VDD),.Y(I9329),.A(g5504));
  NOT NOT1_6025(.VSS(VSS),.VDD(VDD),.Y(I5973),.A(g2247));
  NOT NOT1_6026(.VSS(VSS),.VDD(VDD),.Y(g4586),.A(g4089));
  NOT NOT1_6027(.VSS(VSS),.VDD(VDD),.Y(g11394),.A(I17225));
  NOT NOT1_6028(.VSS(VSS),.VDD(VDD),.Y(g6464),.A(I10398));
  NOT NOT1_6029(.VSS(VSS),.VDD(VDD),.Y(g7903),.A(g7446));
  NOT NOT1_6030(.VSS(VSS),.VDD(VDD),.Y(g2683),.A(g2037));
  NOT NOT1_6031(.VSS(VSS),.VDD(VDD),.Y(I11689),.A(g7044));
  NOT NOT1_6032(.VSS(VSS),.VDD(VDD),.Y(I6870),.A(g2852));
  NOT NOT1_6033(.VSS(VSS),.VDD(VDD),.Y(g3274),.A(I6454));
  NOT NOT1_6034(.VSS(VSS),.VDD(VDD),.Y(g3426),.A(g3121));
  NOT NOT1_6035(.VSS(VSS),.VDD(VDD),.Y(g5880),.A(g5361));
  NOT NOT1_6036(.VSS(VSS),.VDD(VDD),.Y(I12035),.A(g6930));
  NOT NOT1_6037(.VSS(VSS),.VDD(VDD),.Y(I13280),.A(g8250));
  NOT NOT1_6038(.VSS(VSS),.VDD(VDD),.Y(g2778),.A(g2276));
  NOT NOT1_6039(.VSS(VSS),.VDD(VDD),.Y(g10244),.A(g10131));
  NOT NOT1_6040(.VSS(VSS),.VDD(VDD),.Y(I9727),.A(g5250));
  NOT NOT1_6041(.VSS(VSS),.VDD(VDD),.Y(I7369),.A(g4051));
  NOT NOT1_6042(.VSS(VSS),.VDD(VDD),.Y(g3370),.A(I6560));
  NOT NOT1_6043(.VSS(VSS),.VDD(VDD),.Y(I10589),.A(g5763));
  NOT NOT1_6044(.VSS(VSS),.VDD(VDD),.Y(I13624),.A(g8320));
  NOT NOT1_6045(.VSS(VSS),.VDD(VDD),.Y(I14194),.A(g8798));
  NOT NOT1_6046(.VSS(VSS),.VDD(VDD),.Y(g11420),.A(I17315));
  NOT NOT1_6047(.VSS(VSS),.VDD(VDD),.Y(g6563),.A(g5783));
  NOT NOT1_6048(.VSS(VSS),.VDD(VDD),.Y(I7920),.A(g3440));
  NOT NOT1_6049(.VSS(VSS),.VDD(VDD),.Y(g5272),.A(I8724));
  NOT NOT1_6050(.VSS(VSS),.VDD(VDD),.Y(g11319),.A(I17116));
  NOT NOT1_6051(.VSS(VSS),.VDD(VDD),.Y(g7036),.A(g6420));
  NOT NOT1_6052(.VSS(VSS),.VDD(VDD),.Y(g9085),.A(g8892));
  NOT NOT1_6053(.VSS(VSS),.VDD(VDD),.Y(g10069),.A(I15296));
  NOT NOT1_6054(.VSS(VSS),.VDD(VDD),.Y(I7459),.A(g3720));
  NOT NOT1_6055(.VSS(VSS),.VDD(VDD),.Y(I9221),.A(g5236));
  NOT NOT1_6056(.VSS(VSS),.VDD(VDD),.Y(g4525),.A(g3880));
  NOT NOT1_6057(.VSS(VSS),.VDD(VDD),.Y(g7436),.A(g7227));
  NOT NOT1_6058(.VSS(VSS),.VDD(VDD),.Y(g8626),.A(g8498));
  NOT NOT1_6059(.VSS(VSS),.VDD(VDD),.Y(g6295),.A(I10144));
  NOT NOT1_6060(.VSS(VSS),.VDD(VDD),.Y(I12517),.A(g7737));
  NOT NOT1_6061(.VSS(VSS),.VDD(VDD),.Y(I13102),.A(g7928));
  NOT NOT1_6062(.VSS(VSS),.VDD(VDD),.Y(g6237),.A(I9984));
  NOT NOT1_6063(.VSS(VSS),.VDD(VDD),.Y(g11446),.A(I17387));
  NOT NOT1_6064(.VSS(VSS),.VDD(VDD),.Y(g10774),.A(I16458));
  NOT NOT1_6065(.VSS(VSS),.VDD(VDD),.Y(I17438),.A(g11444));
  NOT NOT1_6066(.VSS(VSS),.VDD(VDD),.Y(I10477),.A(g6049));
  NOT NOT1_6067(.VSS(VSS),.VDD(VDD),.Y(I16366),.A(g10591));
  NOT NOT1_6068(.VSS(VSS),.VDD(VDD),.Y(g5417),.A(I8854));
  NOT NOT1_6069(.VSS(VSS),.VDD(VDD),.Y(g2075),.A(I4883));
  NOT NOT1_6070(.VSS(VSS),.VDD(VDD),.Y(I14477),.A(g8943));
  NOT NOT1_6071(.VSS(VSS),.VDD(VDD),.Y(g10879),.A(I16607));
  NOT NOT1_6072(.VSS(VSS),.VDD(VDD),.Y(I16632),.A(g10861));
  NOT NOT1_6073(.VSS(VSS),.VDD(VDD),.Y(g11059),.A(g10974));
  NOT NOT1_6074(.VSS(VSS),.VDD(VDD),.Y(g6844),.A(I10904));
  NOT NOT1_6075(.VSS(VSS),.VDD(VDD),.Y(g7335),.A(I11653));
  NOT NOT1_6076(.VSS(VSS),.VDD(VDD),.Y(g2475),.A(g192));
  NOT NOT1_6077(.VSS(VSS),.VDD(VDD),.Y(I14119),.A(g8779));
  NOT NOT1_6078(.VSS(VSS),.VDD(VDD),.Y(g1988),.A(g766));
  NOT NOT1_6079(.VSS(VSS),.VDD(VDD),.Y(g3544),.A(g3164));
  NOT NOT1_6080(.VSS(VSS),.VDD(VDD),.Y(g2949),.A(I6150));
  NOT NOT1_6081(.VSS(VSS),.VDD(VDD),.Y(g7288),.A(I11540));
  NOT NOT1_6082(.VSS(VSS),.VDD(VDD),.Y(g11540),.A(g11519));
  NOT NOT1_6083(.VSS(VSS),.VDD(VDD),.Y(g5982),.A(I9598));
  NOT NOT1_6084(.VSS(VSS),.VDD(VDD),.Y(g10878),.A(I16604));
  NOT NOT1_6085(.VSS(VSS),.VDD(VDD),.Y(I7793),.A(g3783));
  NOT NOT1_6086(.VSS(VSS),.VDD(VDD),.Y(I10864),.A(g6634));
  NOT NOT1_6087(.VSS(VSS),.VDD(VDD),.Y(g3636),.A(I6815));
  NOT NOT1_6088(.VSS(VSS),.VDD(VDD),.Y(g5629),.A(I9065));
  NOT NOT1_6089(.VSS(VSS),.VDD(VDD),.Y(I9953),.A(g5484));
  NOT NOT1_6090(.VSS(VSS),.VDD(VDD),.Y(g6089),.A(g4977));
  NOT NOT1_6091(.VSS(VSS),.VDD(VDD),.Y(I12193),.A(g7270));
  NOT NOT1_6092(.VSS(VSS),.VDD(VDD),.Y(g10171),.A(I15507));
  NOT NOT1_6093(.VSS(VSS),.VDD(VDD),.Y(g6731),.A(g6001));
  NOT NOT1_6094(.VSS(VSS),.VDD(VDD),.Y(I9068),.A(g4768));
  NOT NOT1_6095(.VSS(VSS),.VDD(VDD),.Y(g7805),.A(I12580));
  NOT NOT1_6096(.VSS(VSS),.VDD(VDD),.Y(I5655),.A(g557));
  NOT NOT1_6097(.VSS(VSS),.VDD(VDD),.Y(g7916),.A(g7651));
  NOT NOT1_6098(.VSS(VSS),.VDD(VDD),.Y(g11203),.A(g11112));
  NOT NOT1_6099(.VSS(VSS),.VDD(VDD),.Y(g5542),.A(I8967));
  NOT NOT1_6100(.VSS(VSS),.VDD(VDD),.Y(g7022),.A(g6389));
  NOT NOT1_6101(.VSS(VSS),.VDD(VDD),.Y(g3306),.A(I6477));
  NOT NOT1_6102(.VSS(VSS),.VDD(VDD),.Y(g2998),.A(g2462));
  NOT NOT1_6103(.VSS(VSS),.VDD(VDD),.Y(g2646),.A(g1992));
  NOT NOT1_6104(.VSS(VSS),.VDD(VDD),.Y(g4158),.A(g3304));
  NOT NOT1_6105(.VSS(VSS),.VDD(VDD),.Y(g7422),.A(I11810));
  NOT NOT1_6106(.VSS(VSS),.VDD(VDD),.Y(g7749),.A(I12412));
  NOT NOT1_6107(.VSS(VSS),.VDD(VDD),.Y(I6065),.A(g2226));
  NOT NOT1_6108(.VSS(VSS),.VDD(VDD),.Y(g6557),.A(g5748));
  NOT NOT1_6109(.VSS(VSS),.VDD(VDD),.Y(I12165),.A(g6882));
  NOT NOT1_6110(.VSS(VSS),.VDD(VDD),.Y(I12523),.A(g7421));
  NOT NOT1_6111(.VSS(VSS),.VDD(VDD),.Y(g10792),.A(I16492));
  NOT NOT1_6112(.VSS(VSS),.VDD(VDD),.Y(g11044),.A(I16793));
  NOT NOT1_6113(.VSS(VSS),.VDD(VDD),.Y(g3790),.A(g3228));
  NOT NOT1_6114(.VSS(VSS),.VDD(VDD),.Y(I15281),.A(g10025));
  NOT NOT1_6115(.VSS(VSS),.VDD(VDD),.Y(g2084),.A(I4900));
  NOT NOT1_6116(.VSS(VSS),.VDD(VDD),.Y(g2603),.A(I5710));
  NOT NOT1_6117(.VSS(VSS),.VDD(VDD),.Y(I8967),.A(g4482));
  NOT NOT1_6118(.VSS(VSS),.VDD(VDD),.Y(g6705),.A(I10682));
  NOT NOT1_6119(.VSS(VSS),.VDD(VDD),.Y(g2039),.A(g1781));
  NOT NOT1_6120(.VSS(VSS),.VDD(VDD),.Y(I9677),.A(g5190));
  NOT NOT1_6121(.VSS(VSS),.VDD(VDD),.Y(g3387),.A(I6587));
  NOT NOT1_6122(.VSS(VSS),.VDD(VDD),.Y(I10305),.A(g6180));
  NOT NOT1_6123(.VSS(VSS),.VDD(VDD),.Y(g5800),.A(I9402));
  NOT NOT1_6124(.VSS(VSS),.VDD(VDD),.Y(I5410),.A(g901));
  NOT NOT1_6125(.VSS(VSS),.VDD(VDD),.Y(g3461),.A(I6671));
  NOT NOT1_6126(.VSS(VSS),.VDD(VDD),.Y(I15377),.A(g10104));
  NOT NOT1_6127(.VSS(VSS),.VDD(VDD),.Y(g6242),.A(I9995));
  NOT NOT1_6128(.VSS(VSS),.VDD(VDD),.Y(g2850),.A(I5976));
  NOT NOT1_6129(.VSS(VSS),.VDD(VDD),.Y(g9431),.A(g9085));
  NOT NOT1_6130(.VSS(VSS),.VDD(VDD),.Y(g7798),.A(I12559));
  NOT NOT1_6131(.VSS(VSS),.VDD(VDD),.Y(g11301),.A(I17084));
  NOT NOT1_6132(.VSS(VSS),.VDD(VDD),.Y(g10459),.A(I15968));
  NOT NOT1_6133(.VSS(VSS),.VDD(VDD),.Y(g9812),.A(g9490));
  NOT NOT1_6134(.VSS(VSS),.VDD(VDD),.Y(g3756),.A(g3015));
  NOT NOT1_6135(.VSS(VSS),.VDD(VDD),.Y(g4587),.A(g3829));
  NOT NOT1_6136(.VSS(VSS),.VDD(VDD),.Y(I12475),.A(g7545));
  NOT NOT1_6137(.VSS(VSS),.VDD(VDD),.Y(g11377),.A(I17202));
  NOT NOT1_6138(.VSS(VSS),.VDD(VDD),.Y(I9866),.A(g5274));
  NOT NOT1_6139(.VSS(VSS),.VDD(VDD),.Y(g6948),.A(I11088));
  NOT NOT1_6140(.VSS(VSS),.VDD(VDD),.Y(g3622),.A(I6757));
  NOT NOT1_6141(.VSS(VSS),.VDD(VDD),.Y(g9958),.A(I15157));
  NOT NOT1_6142(.VSS(VSS),.VDD(VDD),.Y(g7560),.A(I12012));
  NOT NOT1_6143(.VSS(VSS),.VDD(VDD),.Y(g4275),.A(g3664));
  NOT NOT1_6144(.VSS(VSS),.VDD(VDD),.Y(g4311),.A(g4130));
  NOT NOT1_6145(.VSS(VSS),.VDD(VDD),.Y(g10458),.A(I15965));
  NOT NOT1_6146(.VSS(VSS),.VDD(VDD),.Y(g8782),.A(I14083));
  NOT NOT1_6147(.VSS(VSS),.VDD(VDD),.Y(g3427),.A(g3144));
  NOT NOT1_6148(.VSS(VSS),.VDD(VDD),.Y(I15562),.A(g10098));
  NOT NOT1_6149(.VSS(VSS),.VDD(VDD),.Y(I9349),.A(g5515));
  NOT NOT1_6150(.VSS(VSS),.VDD(VDD),.Y(g6955),.A(I11103));
  NOT NOT1_6151(.VSS(VSS),.VDD(VDD),.Y(I10036),.A(g5701));
  NOT NOT1_6152(.VSS(VSS),.VDD(VDD),.Y(g4615),.A(I8024));
  NOT NOT1_6153(.VSS(VSS),.VDD(VDD),.Y(g5213),.A(g4640));
  NOT NOT1_6154(.VSS(VSS),.VDD(VDD),.Y(g11645),.A(I17739));
  NOT NOT1_6155(.VSS(VSS),.VDD(VDD),.Y(I10177),.A(g6103));
  NOT NOT1_6156(.VSS(VSS),.VDD(VDD),.Y(I10560),.A(g5887));
  NOT NOT1_6157(.VSS(VSS),.VDD(VDD),.Y(I11456),.A(g6440));
  NOT NOT1_6158(.VSS(VSS),.VDD(VDD),.Y(I14101),.A(g8774));
  NOT NOT1_6159(.VSS(VSS),.VDD(VDD),.Y(I9848),.A(g5557));
  NOT NOT1_6160(.VSS(VSS),.VDD(VDD),.Y(I15290),.A(g9984));
  NOT NOT1_6161(.VSS(VSS),.VDD(VDD),.Y(g6254),.A(I10021));
  NOT NOT1_6162(.VSS(VSS),.VDD(VDD),.Y(g8475),.A(g8314));
  NOT NOT1_6163(.VSS(VSS),.VDD(VDD),.Y(g4174),.A(I7339));
  NOT NOT1_6164(.VSS(VSS),.VDD(VDD),.Y(g6814),.A(I10852));
  NOT NOT1_6165(.VSS(VSS),.VDD(VDD),.Y(g9765),.A(I14910));
  NOT NOT1_6166(.VSS(VSS),.VDD(VDD),.Y(I17636),.A(g11577));
  NOT NOT1_6167(.VSS(VSS),.VDD(VDD),.Y(I15698),.A(g10235));
  NOT NOT1_6168(.VSS(VSS),.VDD(VDD),.Y(g10545),.A(I16200));
  NOT NOT1_6169(.VSS(VSS),.VDD(VDD),.Y(g2919),.A(I6102));
  NOT NOT1_6170(.VSS(VSS),.VDD(VDD),.Y(g7037),.A(I11198));
  NOT NOT1_6171(.VSS(VSS),.VDD(VDD),.Y(g10079),.A(I15305));
  NOT NOT1_6172(.VSS(VSS),.VDD(VDD),.Y(g10444),.A(g10325));
  NOT NOT1_6173(.VSS(VSS),.VDD(VDD),.Y(I9699),.A(g5426));
  NOT NOT1_6174(.VSS(VSS),.VDD(VDD),.Y(g6150),.A(I9869));
  NOT NOT1_6175(.VSS(VSS),.VDD(VDD),.Y(I14642),.A(g9088));
  NOT NOT1_6176(.VSS(VSS),.VDD(VDD),.Y(g7437),.A(I11829));
  NOT NOT1_6177(.VSS(VSS),.VDD(VDD),.Y(I16784),.A(g10895));
  NOT NOT1_6178(.VSS(VSS),.VDD(VDD),.Y(I5667),.A(g566));
  NOT NOT1_6179(.VSS(VSS),.VDD(VDD),.Y(I6395),.A(g2334));
  NOT NOT1_6180(.VSS(VSS),.VDD(VDD),.Y(I6891),.A(g2962));
  NOT NOT1_6181(.VSS(VSS),.VDD(VDD),.Y(g8292),.A(I13230));
  NOT NOT1_6182(.VSS(VSS),.VDD(VDD),.Y(g2952),.A(g2455));
  NOT NOT1_6183(.VSS(VSS),.VDD(VDD),.Y(I16956),.A(g11096));
  NOT NOT1_6184(.VSS(VSS),.VDD(VDD),.Y(g3345),.A(I6531));
  NOT NOT1_6185(.VSS(VSS),.VDD(VDD),.Y(I16376),.A(g10596));
  NOT NOT1_6186(.VSS(VSS),.VDD(VDD),.Y(I13314),.A(g8260));
  NOT NOT1_6187(.VSS(VSS),.VDD(VDD),.Y(g4284),.A(g3664));
  NOT NOT1_6188(.VSS(VSS),.VDD(VDD),.Y(g7579),.A(I12053));
  NOT NOT1_6189(.VSS(VSS),.VDD(VDD),.Y(g8526),.A(I13735));
  NOT NOT1_6190(.VSS(VSS),.VDD(VDD),.Y(g10598),.A(I16273));
  NOT NOT1_6191(.VSS(VSS),.VDD(VDD),.Y(g3763),.A(I6968));
  NOT NOT1_6192(.VSS(VSS),.VDD(VDD),.Y(I10733),.A(g6099));
  NOT NOT1_6193(.VSS(VSS),.VDD(VDD),.Y(g4545),.A(I7952));
  NOT NOT1_6194(.VSS(VSS),.VDD(VDD),.Y(I11076),.A(g6649));
  NOT NOT1_6195(.VSS(VSS),.VDD(VDD),.Y(I11085),.A(g6433));
  NOT NOT1_6196(.VSS(VSS),.VDD(VDD),.Y(g3391),.A(g2896));
  NOT NOT1_6197(.VSS(VSS),.VDD(VDD),.Y(g9733),.A(I14876));
  NOT NOT1_6198(.VSS(VSS),.VDD(VDD),.Y(I15427),.A(g10088));
  NOT NOT1_6199(.VSS(VSS),.VDD(VDD),.Y(I16095),.A(g10401));
  NOT NOT1_6200(.VSS(VSS),.VDD(VDD),.Y(g4180),.A(I7357));
  NOT NOT1_6201(.VSS(VSS),.VDD(VDD),.Y(g5490),.A(I8911));
  NOT NOT1_6202(.VSS(VSS),.VDD(VDD),.Y(g9270),.A(I14485));
  NOT NOT1_6203(.VSS(VSS),.VDD(VDD),.Y(g4380),.A(I7701));
  NOT NOT1_6204(.VSS(VSS),.VDD(VDD),.Y(g11427),.A(I17334));
  NOT NOT1_6205(.VSS(VSS),.VDD(VDD),.Y(g5166),.A(g4682));
  NOT NOT1_6206(.VSS(VSS),.VDD(VDD),.Y(I11596),.A(g6831));
  NOT NOT1_6207(.VSS(VSS),.VDD(VDD),.Y(g4591),.A(g3829));
  NOT NOT1_6208(.VSS(VSS),.VDD(VDD),.Y(I15632),.A(g10184));
  NOT NOT1_6209(.VSS(VSS),.VDD(VDD),.Y(g11366),.A(I17191));
  NOT NOT1_6210(.VSS(VSS),.VDD(VDD),.Y(g3637),.A(I6818));
  NOT NOT1_6211(.VSS(VSS),.VDD(VDD),.Y(I7216),.A(g2952));
  NOT NOT1_6212(.VSS(VSS),.VDD(VDD),.Y(g7752),.A(I12421));
  NOT NOT1_6213(.VSS(VSS),.VDD(VDD),.Y(g11632),.A(I17710));
  NOT NOT1_6214(.VSS(VSS),.VDD(VDD),.Y(g8484),.A(g8336));
  NOT NOT1_6215(.VSS(VSS),.VDD(VDD),.Y(I16181),.A(g10491));
  NOT NOT1_6216(.VSS(VSS),.VDD(VDD),.Y(I10630),.A(g5889));
  NOT NOT1_6217(.VSS(VSS),.VDD(VDD),.Y(g8439),.A(I13615));
  NOT NOT1_6218(.VSS(VSS),.VDD(VDD),.Y(g2004),.A(I4820));
  NOT NOT1_6219(.VSS(VSS),.VDD(VDD),.Y(I10693),.A(g6068));
  NOT NOT1_6220(.VSS(VSS),.VDD(VDD),.Y(g6836),.A(I10888));
  NOT NOT1_6221(.VSS(VSS),.VDD(VDD),.Y(I12372),.A(g7137));
  NOT NOT1_6222(.VSS(VSS),.VDD(VDD),.Y(g7917),.A(g7497));
  NOT NOT1_6223(.VSS(VSS),.VDD(VDD),.Y(g2986),.A(I6220));
  NOT NOT1_6224(.VSS(VSS),.VDD(VDD),.Y(g3307),.A(I6480));
  NOT NOT1_6225(.VSS(VSS),.VDD(VDD),.Y(g9473),.A(g9103));
  NOT NOT1_6226(.VSS(VSS),.VDD(VDD),.Y(I7671),.A(g3351));
  NOT NOT1_6227(.VSS(VSS),.VDD(VDD),.Y(g2647),.A(g1993));
  NOT NOT1_6228(.VSS(VSS),.VDD(VDD),.Y(g10159),.A(I15473));
  NOT NOT1_6229(.VSS(VSS),.VDD(VDD),.Y(g4420),.A(I7766));
  NOT NOT1_6230(.VSS(VSS),.VDD(VDD),.Y(g10125),.A(I15377));
  NOT NOT1_6231(.VSS(VSS),.VDD(VDD),.Y(g10532),.A(g10473));
  NOT NOT1_6232(.VSS(VSS),.VDD(VDD),.Y(g10901),.A(g10802));
  NOT NOT1_6233(.VSS(VSS),.VDD(VDD),.Y(I10009),.A(g5542));
  NOT NOT1_6234(.VSS(VSS),.VDD(VDD),.Y(g5649),.A(I9108));
  NOT NOT1_6235(.VSS(VSS),.VDD(VDD),.Y(g3359),.A(I6543));
  NOT NOT1_6236(.VSS(VSS),.VDD(VDD),.Y(I15403),.A(g10069));
  NOT NOT1_6237(.VSS(VSS),.VDD(VDD),.Y(g1965),.A(g119));
  NOT NOT1_6238(.VSS(VSS),.VDD(VDD),.Y(g4507),.A(g3546));
  NOT NOT1_6239(.VSS(VSS),.VDD(VDD),.Y(g5348),.A(I8815));
  NOT NOT1_6240(.VSS(VSS),.VDD(VDD),.Y(g6967),.A(I11119));
  NOT NOT1_6241(.VSS(VSS),.VDD(VDD),.Y(I5555),.A(g110));
  NOT NOT1_6242(.VSS(VSS),.VDD(VDD),.Y(I11269),.A(g6545));
  NOT NOT1_6243(.VSS(VSS),.VDD(VDD),.Y(g9980),.A(I15181));
  NOT NOT1_6244(.VSS(VSS),.VDD(VDD),.Y(g2764),.A(I5850));
  NOT NOT1_6245(.VSS(VSS),.VDD(VDD),.Y(I8462),.A(g4475));
  NOT NOT1_6246(.VSS(VSS),.VDD(VDD),.Y(g11403),.A(I17252));
  NOT NOT1_6247(.VSS(VSS),.VDD(VDD),.Y(g10158),.A(I15470));
  NOT NOT1_6248(.VSS(VSS),.VDD(VDD),.Y(g11547),.A(g11519));
  NOT NOT1_6249(.VSS(VSS),.VDD(VDD),.Y(g7042),.A(I11211));
  NOT NOT1_6250(.VSS(VSS),.VDD(VDD),.Y(I11773),.A(g7257));
  NOT NOT1_6251(.VSS(VSS),.VDD(VDD),.Y(g10783),.A(I16479));
  NOT NOT1_6252(.VSS(VSS),.VDD(VDD),.Y(g4794),.A(I8164));
  NOT NOT1_6253(.VSS(VSS),.VDD(VDD),.Y(I11942),.A(g6909));
  NOT NOT1_6254(.VSS(VSS),.VDD(VDD),.Y(I13773),.A(g8384));
  NOT NOT1_6255(.VSS(VSS),.VDD(VDD),.Y(I5792),.A(g2080));
  NOT NOT1_6256(.VSS(VSS),.VDD(VDD),.Y(g7442),.A(g7237));
  NOT NOT1_6257(.VSS(VSS),.VDD(VDD),.Y(g8702),.A(g8664));
  NOT NOT1_6258(.VSS(VSS),.VDD(VDD),.Y(I13341),.A(g8210));
  NOT NOT1_6259(.VSS(VSS),.VDD(VDD),.Y(I12790),.A(g7618));
  NOT NOT1_6260(.VSS(VSS),.VDD(VDD),.Y(g7786),.A(I12523));
  NOT NOT1_6261(.VSS(VSS),.VDD(VDD),.Y(g2503),.A(g1872));
  NOT NOT1_6262(.VSS(VSS),.VDD(VDD),.Y(g3757),.A(I6952));
  NOT NOT1_6263(.VSS(VSS),.VDD(VDD),.Y(I9352),.A(g4944));
  NOT NOT1_6264(.VSS(VSS),.VDD(VDD),.Y(I17312),.A(g11392));
  NOT NOT1_6265(.VSS(VSS),.VDD(VDD),.Y(g10353),.A(I15823));
  NOT NOT1_6266(.VSS(VSS),.VDD(VDD),.Y(g3416),.A(g3144));
  NOT NOT1_6267(.VSS(VSS),.VDD(VDD),.Y(g6993),.A(I11135));
  NOT NOT1_6268(.VSS(VSS),.VDD(VDD),.Y(I11180),.A(g6506));
  NOT NOT1_6269(.VSS(VSS),.VDD(VDD),.Y(I16190),.A(g10493));
  NOT NOT1_6270(.VSS(VSS),.VDD(VDD),.Y(I14485),.A(g8883));
  NOT NOT1_6271(.VSS(VSS),.VDD(VDD),.Y(g7364),.A(I11740));
  NOT NOT1_6272(.VSS(VSS),.VDD(VDD),.Y(I6815),.A(g2755));
  NOT NOT1_6273(.VSS(VSS),.VDD(VDD),.Y(I9717),.A(g5426));
  NOT NOT1_6274(.VSS(VSS),.VDD(VDD),.Y(I15551),.A(g10080));
  NOT NOT1_6275(.VSS(VSS),.VDD(VDD),.Y(I14555),.A(g9009));
  NOT NOT1_6276(.VSS(VSS),.VDD(VDD),.Y(g3522),.A(g3164));
  NOT NOT1_6277(.VSS(VSS),.VDD(VDD),.Y(g8952),.A(I14309));
  NOT NOT1_6278(.VSS(VSS),.VDD(VDD),.Y(g11572),.A(g11561));
  NOT NOT1_6279(.VSS(VSS),.VDD(VDD),.Y(I11734),.A(g7024));
  NOT NOT1_6280(.VSS(VSS),.VDD(VDD),.Y(g8276),.A(I13200));
  NOT NOT1_6281(.VSS(VSS),.VDD(VDD),.Y(g3811),.A(I7029));
  NOT NOT1_6282(.VSS(VSS),.VDD(VDD),.Y(g2224),.A(g695));
  NOT NOT1_6283(.VSS(VSS),.VDD(VDD),.Y(I6097),.A(g2391));
  NOT NOT1_6284(.VSS(VSS),.VDD(VDD),.Y(g5063),.A(g4363));
  NOT NOT1_6285(.VSS(VSS),.VDD(VDD),.Y(I10914),.A(g6728));
  NOT NOT1_6286(.VSS(VSS),.VDD(VDD),.Y(g7454),.A(g7148));
  NOT NOT1_6287(.VSS(VSS),.VDD(VDD),.Y(I6726),.A(g3306));
  NOT NOT1_6288(.VSS(VSS),.VDD(VDD),.Y(I14570),.A(g9028));
  NOT NOT1_6289(.VSS(VSS),.VDD(VDD),.Y(I9893),.A(g5557));
  NOT NOT1_6290(.VSS(VSS),.VDD(VDD),.Y(I13335),.A(g8206));
  NOT NOT1_6291(.VSS(VSS),.VDD(VDD),.Y(g7770),.A(I12475));
  NOT NOT1_6292(.VSS(VSS),.VDD(VDD),.Y(I14914),.A(g9533));
  NOT NOT1_6293(.VSS(VSS),.VDD(VDD),.Y(g4515),.A(I7916));
  NOT NOT1_6294(.VSS(VSS),.VDD(VDD),.Y(g4204),.A(I7429));
  NOT NOT1_6295(.VSS(VSS),.VDD(VDD),.Y(I15127),.A(g9919));
  NOT NOT1_6296(.VSS(VSS),.VDD(VDD),.Y(I16546),.A(g10724));
  NOT NOT1_6297(.VSS(VSS),.VDD(VDD),.Y(g8561),.A(I13776));
  NOT NOT1_6298(.VSS(VSS),.VDD(VDD),.Y(g2320),.A(g18));
  NOT NOT1_6299(.VSS(VSS),.VDD(VDD),.Y(I10907),.A(g6705));
  NOT NOT1_6300(.VSS(VSS),.VDD(VDD),.Y(g7725),.A(I12360));
  NOT NOT1_6301(.VSS(VSS),.VDD(VDD),.Y(I8842),.A(g4556));
  NOT NOT1_6302(.VSS(VSS),.VDD(VDD),.Y(g7532),.A(I11932));
  NOT NOT1_6303(.VSS(VSS),.VDD(VDD),.Y(I7308),.A(g3070));
  NOT NOT1_6304(.VSS(VSS),.VDD(VDD),.Y(g3874),.A(g2920));
  NOT NOT1_6305(.VSS(VSS),.VDD(VDD),.Y(I8192),.A(g3566));
  NOT NOT1_6306(.VSS(VSS),.VDD(VDD),.Y(I12208),.A(g7124));
  NOT NOT1_6307(.VSS(VSS),.VDD(VDD),.Y(I8298),.A(g4437));
  NOT NOT1_6308(.VSS(VSS),.VDD(VDD),.Y(I8085),.A(g3664));
  NOT NOT1_6309(.VSS(VSS),.VDD(VDD),.Y(I13965),.A(g8451));
  NOT NOT1_6310(.VSS(VSS),.VDD(VDD),.Y(g8004),.A(I12838));
  NOT NOT1_6311(.VSS(VSS),.VDD(VDD),.Y(g6921),.A(I11037));
  NOT NOT1_6312(.VSS(VSS),.VDD(VDD),.Y(g8986),.A(I14379));
  NOT NOT1_6313(.VSS(VSS),.VDD(VDD),.Y(I5494),.A(g1690));
  NOT NOT1_6314(.VSS(VSS),.VDD(VDD),.Y(I13131),.A(g7979));
  NOT NOT1_6315(.VSS(VSS),.VDD(VDD),.Y(I14239),.A(g8803));
  NOT NOT1_6316(.VSS(VSS),.VDD(VDD),.Y(I15956),.A(g10402));
  NOT NOT1_6317(.VSS(VSS),.VDD(VDD),.Y(g2617),.A(g1997));
  NOT NOT1_6318(.VSS(VSS),.VDD(VDD),.Y(g2906),.A(I6071));
  NOT NOT1_6319(.VSS(VSS),.VDD(VDD),.Y(I14567),.A(g9027));
  NOT NOT1_6320(.VSS(VSS),.VDD(VDD),.Y(g2789),.A(g2276));
  NOT NOT1_6321(.VSS(VSS),.VDD(VDD),.Y(g5619),.A(g4840));
  NOT NOT1_6322(.VSS(VSS),.VDD(VDD),.Y(g5167),.A(g4682));
  NOT NOT1_6323(.VSS(VSS),.VDD(VDD),.Y(I15980),.A(g10414));
//
  AND2 AND2_0(.VSS(VSS),.VDD(VDD),.Y(g11103),.A(g2250),.B(g10937));
  AND2 AND2_1(.VSS(VSS),.VDD(VDD),.Y(g9900),.A(g9845),.B(g8327));
  AND2 AND2_2(.VSS(VSS),.VDD(VDD),.Y(g11095),.A(g845),.B(g10950));
  AND2 AND2_3(.VSS(VSS),.VDD(VDD),.Y(g3880),.A(g3186),.B(g2023));
  AND2 AND2_4(.VSS(VSS),.VDD(VDD),.Y(g4973),.A(g1645),.B(g4467));
  AND2 AND2_5(.VSS(VSS),.VDD(VDD),.Y(g7389),.A(g7001),.B(g3880));
  AND2 AND2_6(.VSS(VSS),.VDD(VDD),.Y(g7888),.A(g7465),.B(g7025));
  AND2 AND2_7(.VSS(VSS),.VDD(VDD),.Y(g4969),.A(g1642),.B(g4463));
  AND2 AND2_8(.VSS(VSS),.VDD(VDD),.Y(g8224),.A(g1882),.B(g7887));
  AND2 AND2_9(.VSS(VSS),.VDD(VDD),.Y(g2892),.A(g1980),.B(g1976));
  AND2 AND2_10(.VSS(VSS),.VDD(VDD),.Y(g5686),.A(g158),.B(g5361));
  AND2 AND2_11(.VSS(VSS),.VDD(VDD),.Y(g10308),.A(g10217),.B(g9085));
  AND2 AND2_12(.VSS(VSS),.VDD(VDD),.Y(g4123),.A(g2695),.B(g3037));
  AND2 AND2_13(.VSS(VSS),.VDD(VDD),.Y(g8120),.A(g1909),.B(g7944));
  AND2 AND2_14(.VSS(VSS),.VDD(VDD),.Y(g6788),.A(g287),.B(g5876));
  AND2 AND2_15(.VSS(VSS),.VDD(VDD),.Y(g5598),.A(g778),.B(g4824));
  AND2 AND2_16(.VSS(VSS),.VDD(VDD),.Y(g9694),.A(g278),.B(g9432));
  AND2 AND2_17(.VSS(VSS),.VDD(VDD),.Y(g10495),.A(g10431),.B(g3971));
  AND2 AND2_18(.VSS(VSS),.VDD(VDD),.Y(g2945),.A(g2411),.B(g1684));
  AND2 AND2_19(.VSS(VSS),.VDD(VDD),.Y(g11190),.A(g5623),.B(g11065));
  AND2 AND2_20(.VSS(VSS),.VDD(VDD),.Y(g8789),.A(g8639),.B(g8719));
  AND2 AND2_21(.VSS(VSS),.VDD(VDD),.Y(g9852),.A(g9728),.B(g9563));
  AND2 AND2_22(.VSS(VSS),.VDD(VDD),.Y(g5625),.A(g1053),.B(g4399));
  AND2 AND2_23(.VSS(VSS),.VDD(VDD),.Y(g4875),.A(g995),.B(g3914));
  AND2 AND2_24(.VSS(VSS),.VDD(VDD),.Y(g9701),.A(g1574),.B(g9474));
  AND2 AND2_25(.VSS(VSS),.VDD(VDD),.Y(g7138),.A(g6055),.B(g6707));
  AND2 AND2_26(.VSS(VSS),.VDD(VDD),.Y(g10752),.A(g10692),.B(g3586));
  AND2 AND2_27(.VSS(VSS),.VDD(VDD),.Y(g11211),.A(g11058),.B(g5534));
  AND2 AND2_28(.VSS(VSS),.VDD(VDD),.Y(g11024),.A(g435),.B(g10974));
  AND2 AND2_29(.VSS(VSS),.VDD(VDD),.Y(g8547),.A(g8307),.B(g7693));
  AND2 AND2_30(.VSS(VSS),.VDD(VDD),.Y(g10669),.A(g10577),.B(g9429));
  AND2 AND2_31(.VSS(VSS),.VDD(VDD),.Y(g7707),.A(g691),.B(g7206));
  AND2 AND2_32(.VSS(VSS),.VDD(VDD),.Y(g4884),.A(g3813),.B(g2971));
  AND2 AND2_33(.VSS(VSS),.VDD(VDD),.Y(g4839),.A(g225),.B(g3946));
  AND2 AND2_34(.VSS(VSS),.VDD(VDD),.Y(g9870),.A(g1561),.B(g9816));
  AND2 AND2_35(.VSS(VSS),.VDD(VDD),.Y(g6640),.A(g5281),.B(g5801));
  AND2 AND2_36(.VSS(VSS),.VDD(VDD),.Y(g9650),.A(g2797),.B(g9240));
  AND2 AND2_37(.VSS(VSS),.VDD(VDD),.Y(g5687),.A(g139),.B(g5361));
  AND2 AND2_38(.VSS(VSS),.VDD(VDD),.Y(g7957),.A(g2885),.B(g7527));
  AND2 AND2_39(.VSS(VSS),.VDD(VDD),.Y(g3512),.A(g2050),.B(g2971));
  AND2 AND2_40(.VSS(VSS),.VDD(VDD),.Y(g8244),.A(g7847),.B(g4336));
  AND2 AND2_41(.VSS(VSS),.VDD(VDD),.Y(g7449),.A(g6868),.B(g4355));
  AND2 AND2_42(.VSS(VSS),.VDD(VDD),.Y(g4235),.A(g1011),.B(g3914));
  AND2 AND2_43(.VSS(VSS),.VDD(VDD),.Y(g4343),.A(g345),.B(g3586));
  AND2 AND2_44(.VSS(VSS),.VDD(VDD),.Y(g11296),.A(g5482),.B(g11241));
  AND2 AND2_45(.VSS(VSS),.VDD(VDD),.Y(g9594),.A(g1),.B(g9292));
  AND2 AND2_46(.VSS(VSS),.VDD(VDD),.Y(g6829),.A(g213),.B(g6596));
  AND2 AND2_47(.VSS(VSS),.VDD(VDD),.Y(g4334),.A(g1160),.B(g3703));
  AND2 AND2_48(.VSS(VSS),.VDD(VDD),.Y(g9943),.A(g9923),.B(g9367));
  AND2 AND2_49(.VSS(VSS),.VDD(VDD),.Y(g5525),.A(g1721),.B(g4292));
  AND2 AND2_50(.VSS(VSS),.VDD(VDD),.Y(g4548),.A(g440),.B(g3990));
  AND3 AND3_0(.VSS(VSS),.VDD(VDD),.Y(g8876),.A(g8105),.B(g6764),.C(g8858));
  AND2 AND2_51(.VSS(VSS),.VDD(VDD),.Y(g6733),.A(g5678),.B(g4324));
  AND2 AND2_52(.VSS(VSS),.VDD(VDD),.Y(g4804),.A(g476),.B(g3458));
  AND2 AND2_53(.VSS(VSS),.VDD(VDD),.Y(g10705),.A(g10564),.B(g4840));
  AND2 AND2_54(.VSS(VSS),.VDD(VDD),.Y(g9934),.A(g9913),.B(g9624));
  AND2 AND2_55(.VSS(VSS),.VDD(VDD),.Y(g6225),.A(g566),.B(g5082));
  AND2 AND2_56(.VSS(VSS),.VDD(VDD),.Y(g6324),.A(g1240),.B(g5949));
  AND2 AND2_57(.VSS(VSS),.VDD(VDD),.Y(g10686),.A(g10612),.B(g3863));
  AND2 AND2_58(.VSS(VSS),.VDD(VDD),.Y(g6540),.A(g1223),.B(g6072));
  AND2 AND2_59(.VSS(VSS),.VDD(VDD),.Y(g8663),.A(g8538),.B(g4013));
  AND2 AND2_60(.VSS(VSS),.VDD(VDD),.Y(g11581),.A(g1308),.B(g11539));
  AND2 AND2_61(.VSS(VSS),.VDD(VDD),.Y(g6206),.A(g560),.B(g5068));
  AND2 AND2_62(.VSS(VSS),.VDD(VDD),.Y(g4518),.A(g452),.B(g3975));
  AND2 AND2_63(.VSS(VSS),.VDD(VDD),.Y(g3989),.A(g248),.B(g3164));
  AND2 AND2_64(.VSS(VSS),.VDD(VDD),.Y(g7730),.A(g7260),.B(g2347));
  AND2 AND2_65(.VSS(VSS),.VDD(VDD),.Y(g5174),.A(g1235),.B(g4681));
  AND2 AND2_66(.VSS(VSS),.VDD(VDD),.Y(g7504),.A(g7148),.B(g2847));
  AND2 AND2_67(.VSS(VSS),.VDD(VDD),.Y(g7185),.A(g1887),.B(g6724));
  AND2 AND2_68(.VSS(VSS),.VDD(VDD),.Y(g2563),.A(I5689),.B(I5690));
  AND2 AND2_69(.VSS(VSS),.VDD(VDD),.Y(g7881),.A(g7612),.B(g3810));
  AND2 AND2_70(.VSS(VSS),.VDD(VDD),.Y(g11070),.A(g2008),.B(g10913));
  AND2 AND2_71(.VSS(VSS),.VDD(VDD),.Y(g9859),.A(g9736),.B(g9573));
  AND3 AND3_1(.VSS(VSS),.VDD(VDD),.Y(g8877),.A(g8103),.B(g6764),.C(g8858));
  AND2 AND2_72(.VSS(VSS),.VDD(VDD),.Y(g11590),.A(g2274),.B(g11561));
  AND2 AND2_73(.VSS(VSS),.VDD(VDD),.Y(g6199),.A(g557),.B(g5062));
  AND2 AND2_74(.VSS(VSS),.VDD(VDD),.Y(g9266),.A(g8932),.B(g3398));
  AND2 AND2_75(.VSS(VSS),.VDD(VDD),.Y(g5545),.A(g1730),.B(g4321));
  AND2 AND2_76(.VSS(VSS),.VDD(VDD),.Y(g5180),.A(g4541),.B(g4533));
  AND2 AND2_77(.VSS(VSS),.VDD(VDD),.Y(g5591),.A(g1615),.B(g4514));
  AND2 AND2_78(.VSS(VSS),.VDD(VDD),.Y(g8556),.A(g8412),.B(g8029));
  AND2 AND2_79(.VSS(VSS),.VDD(VDD),.Y(g11094),.A(g374),.B(g10883));
  AND2 AND2_80(.VSS(VSS),.VDD(VDD),.Y(g5853),.A(g5044),.B(g1927));
  AND2 AND2_81(.VSS(VSS),.VDD(VDD),.Y(g6245),.A(g575),.B(g5098));
  AND2 AND2_82(.VSS(VSS),.VDD(VDD),.Y(g4360),.A(g1861),.B(g3748));
  AND3 AND3_2(.VSS(VSS),.VDD(VDD),.Y(g8930),.A(g8100),.B(g6368),.C(g8828));
  AND2 AND2_83(.VSS(VSS),.VDD(VDD),.Y(g5507),.A(g4310),.B(g3528));
  AND2 AND2_84(.VSS(VSS),.VDD(VDD),.Y(g11150),.A(g3087),.B(g10913));
  AND2 AND2_85(.VSS(VSS),.VDD(VDD),.Y(g8464),.A(g8302),.B(g7416));
  AND2 AND2_86(.VSS(VSS),.VDD(VDD),.Y(g9692),.A(g272),.B(g9432));
  AND2 AND2_87(.VSS(VSS),.VDD(VDD),.Y(g4996),.A(g1428),.B(g4682));
  AND2 AND2_88(.VSS(VSS),.VDD(VDD),.Y(g7131),.A(g6044),.B(g6700));
  AND2 AND2_89(.VSS(VSS),.VDD(VDD),.Y(g11019),.A(g421),.B(g10974));
  AND2 AND2_90(.VSS(VSS),.VDD(VDD),.Y(g9960),.A(g9951),.B(g9536));
  AND2 AND2_91(.VSS(VSS),.VDD(VDD),.Y(g11196),.A(g4912),.B(g11068));
  AND2 AND2_92(.VSS(VSS),.VDD(VDD),.Y(g11018),.A(g7286),.B(g10974));
  AND2 AND2_93(.VSS(VSS),.VDD(VDD),.Y(g6819),.A(g243),.B(g6596));
  AND2 AND2_94(.VSS(VSS),.VDD(VDD),.Y(g10595),.A(g10550),.B(g4347));
  AND2 AND2_95(.VSS(VSS),.VDD(VDD),.Y(g10494),.A(g10433),.B(g3945));
  AND2 AND2_96(.VSS(VSS),.VDD(VDD),.Y(g10623),.A(g10544),.B(g4536));
  AND2 AND2_97(.VSS(VSS),.VDD(VDD),.Y(g4878),.A(g1868),.B(g3531));
  AND2 AND2_98(.VSS(VSS),.VDD(VDD),.Y(g5204),.A(g4838),.B(g2126));
  AND2 AND2_99(.VSS(VSS),.VDD(VDD),.Y(g8844),.A(g8609),.B(g8709));
  AND2 AND2_100(.VSS(VSS),.VDD(VDD),.Y(g6701),.A(g6185),.B(g4228));
  AND2 AND2_101(.VSS(VSS),.VDD(VDD),.Y(g10782),.A(g10725),.B(g5146));
  AND2 AND2_102(.VSS(VSS),.VDD(VDD),.Y(g5100),.A(g1791),.B(g4606));
  AND2 AND2_103(.VSS(VSS),.VDD(VDD),.Y(g4882),.A(g1089),.B(g3638));
  AND2 AND2_104(.VSS(VSS),.VDD(VDD),.Y(g8731),.A(g8622),.B(g7918));
  AND2 AND2_105(.VSS(VSS),.VDD(VDD),.Y(g6215),.A(g1504),.B(g5128));
  AND2 AND2_106(.VSS(VSS),.VDD(VDD),.Y(g6886),.A(g1932),.B(g6420));
  AND2 AND2_107(.VSS(VSS),.VDD(VDD),.Y(g3586),.A(g3323),.B(g2191));
  AND2 AND2_108(.VSS(VSS),.VDD(VDD),.Y(g8557),.A(g8415),.B(g8033));
  AND3 AND3_3(.VSS(VSS),.VDD(VDD),.Y(g8966),.A(g8081),.B(g6778),.C(g8849));
  AND2 AND2_109(.VSS(VSS),.VDD(VDD),.Y(g8071),.A(g691),.B(g7826));
  AND2 AND2_110(.VSS(VSS),.VDD(VDD),.Y(g11597),.A(g11576),.B(g5446));
  AND2 AND2_111(.VSS(VSS),.VDD(VDD),.Y(g9828),.A(g9722),.B(g9785));
  AND2 AND2_112(.VSS(VSS),.VDD(VDD),.Y(g2918),.A(g2411),.B(g1672));
  AND2 AND2_113(.VSS(VSS),.VDD(VDD),.Y(g9830),.A(g9725),.B(g9785));
  AND3 AND3_4(.VSS(VSS),.VDD(VDD),.Y(g8955),.A(g8110),.B(g6368),.C(g8828));
  AND2 AND2_114(.VSS(VSS),.VDD(VDD),.Y(g9592),.A(g4),.B(g9292));
  AND2 AND2_115(.VSS(VSS),.VDD(VDD),.Y(g5123),.A(g1618),.B(g4669));
  AND2 AND2_116(.VSS(VSS),.VDD(VDD),.Y(g7059),.A(g6078),.B(g6714));
  AND2 AND2_117(.VSS(VSS),.VDD(VDD),.Y(g8254),.A(g2773),.B(g7909));
  AND2 AND2_118(.VSS(VSS),.VDD(VDD),.Y(g7459),.A(g7148),.B(g2814));
  AND2 AND2_119(.VSS(VSS),.VDD(VDD),.Y(g11102),.A(g861),.B(g10950));
  AND2 AND2_120(.VSS(VSS),.VDD(VDD),.Y(g7718),.A(g709),.B(g7221));
  AND2 AND2_121(.VSS(VSS),.VDD(VDD),.Y(g7535),.A(g7148),.B(g2874));
  AND2 AND2_122(.VSS(VSS),.VDD(VDD),.Y(g9703),.A(g1577),.B(g9474));
  AND2 AND2_123(.VSS(VSS),.VDD(VDD),.Y(g5528),.A(g4322),.B(g3537));
  AND2 AND2_124(.VSS(VSS),.VDD(VDD),.Y(g5151),.A(g4478),.B(g2733));
  AND2 AND2_125(.VSS(VSS),.VDD(VDD),.Y(g9932),.A(g9911),.B(g9624));
  AND2 AND2_126(.VSS(VSS),.VDD(VDD),.Y(g5530),.A(g1636),.B(g4305));
  AND2 AND2_127(.VSS(VSS),.VDD(VDD),.Y(g3506),.A(g986),.B(g2760));
  AND2 AND2_128(.VSS(VSS),.VDD(VDD),.Y(g8769),.A(g8629),.B(g5151));
  AND2 AND2_129(.VSS(VSS),.VDD(VDD),.Y(g6887),.A(g6187),.B(g6566));
  AND2 AND2_130(.VSS(VSS),.VDD(VDD),.Y(g6228),.A(g5605),.B(g713));
  AND2 AND2_131(.VSS(VSS),.VDD(VDD),.Y(g6322),.A(g1275),.B(g5949));
  AND2 AND2_132(.VSS(VSS),.VDD(VDD),.Y(g3111),.A(I6337),.B(I6338));
  AND3 AND3_5(.VSS(VSS),.VDD(VDD),.Y(g8967),.A(g8085),.B(g6778),.C(g8849));
  AND2 AND2_133(.VSS(VSS),.VDD(VDD),.Y(g5010),.A(g1458),.B(g4640));
  AND2 AND2_134(.VSS(VSS),.VDD(VDD),.Y(g3275),.A(g115),.B(g2356));
  AND2 AND2_135(.VSS(VSS),.VDD(VDD),.Y(g10809),.A(g4811),.B(g10754));
  AND2 AND2_136(.VSS(VSS),.VDD(VDD),.Y(g2895),.A(g2411),.B(g1678));
  AND2 AND2_137(.VSS(VSS),.VDD(VDD),.Y(g7721),.A(g736),.B(g7237));
  AND2 AND2_138(.VSS(VSS),.VDD(VDD),.Y(g9866),.A(g1549),.B(g9802));
  AND2 AND2_139(.VSS(VSS),.VDD(VDD),.Y(g9716),.A(g1534),.B(g9490));
  AND2 AND2_140(.VSS(VSS),.VDD(VDD),.Y(g10808),.A(g10744),.B(g3829));
  AND2 AND2_141(.VSS(VSS),.VDD(VDD),.Y(g3374),.A(g1231),.B(g3047));
  AND2 AND2_142(.VSS(VSS),.VDD(VDD),.Y(g4492),.A(g1786),.B(g3685));
  AND2 AND2_143(.VSS(VSS),.VDD(VDD),.Y(g8822),.A(g8614),.B(g8752));
  AND2 AND2_144(.VSS(VSS),.VDD(VDD),.Y(g10560),.A(g10487),.B(g4575));
  AND3 AND3_6(.VSS(VSS),.VDD(VDD),.Y(g11456),.A(g3765),.B(g3517),.C(g11422));
  AND2 AND2_145(.VSS(VSS),.VDD(VDD),.Y(g9848),.A(g9724),.B(g9557));
  AND2 AND2_146(.VSS(VSS),.VDD(VDD),.Y(g4714),.A(g646),.B(g3333));
  AND2 AND2_147(.VSS(VSS),.VDD(VDD),.Y(g6550),.A(g1231),.B(g6089));
  AND2 AND2_148(.VSS(VSS),.VDD(VDD),.Y(g5172),.A(g4555),.B(g4549));
  AND2 AND2_149(.VSS(VSS),.VDD(VDD),.Y(g10642),.A(g10612),.B(g3829));
  AND2 AND2_150(.VSS(VSS),.VDD(VDD),.Y(g3284),.A(g2531),.B(g677));
  AND2 AND2_151(.VSS(VSS),.VDD(VDD),.Y(g9699),.A(g284),.B(g9432));
  AND2 AND2_152(.VSS(VSS),.VDD(VDD),.Y(g9855),.A(g302),.B(g9772));
  AND2 AND2_153(.VSS(VSS),.VDD(VDD),.Y(g5618),.A(g1630),.B(g4551));
  AND2 AND2_154(.VSS(VSS),.VDD(VDD),.Y(g6891),.A(g1950),.B(g6435));
  AND2 AND2_155(.VSS(VSS),.VDD(VDD),.Y(g7940),.A(g7620),.B(g4013));
  AND2 AND2_156(.VSS(VSS),.VDD(VDD),.Y(g11085),.A(g312),.B(g10897));
  AND2 AND2_157(.VSS(VSS),.VDD(VDD),.Y(g4736),.A(g396),.B(g3379));
  AND2 AND2_158(.VSS(VSS),.VDD(VDD),.Y(g4968),.A(g1432),.B(g4682));
  AND2 AND2_159(.VSS(VSS),.VDD(VDD),.Y(g8837),.A(g8646),.B(g8697));
  AND2 AND2_160(.VSS(VSS),.VDD(VDD),.Y(g9644),.A(g1182),.B(g9125));
  AND2 AND2_161(.VSS(VSS),.VDD(VDD),.Y(g5804),.A(g1546),.B(g5261));
  AND2 AND2_162(.VSS(VSS),.VDD(VDD),.Y(g8462),.A(g8300),.B(g7406));
  AND4 AND4_0(.VSS(VSS),.VDD(VDD),.Y(I6330),.A(g2549),.B(g2556),.C(g2562),.D(g2570));
  AND2 AND2_163(.VSS(VSS),.VDD(VDD),.Y(g11156),.A(g333),.B(g10934));
  AND2 AND2_164(.VSS(VSS),.VDD(VDD),.Y(g6342),.A(g293),.B(g5886));
  AND2 AND2_165(.VSS(VSS),.VDD(VDD),.Y(g9867),.A(g1552),.B(g9807));
  AND2 AND2_166(.VSS(VSS),.VDD(VDD),.Y(g9717),.A(g1537),.B(g9490));
  AND2 AND2_167(.VSS(VSS),.VDD(VDD),.Y(g4871),.A(g1864),.B(g3523));
  AND2 AND2_168(.VSS(VSS),.VDD(VDD),.Y(g10454),.A(g10435),.B(g3411));
  AND2 AND2_169(.VSS(VSS),.VDD(VDD),.Y(g4722),.A(g426),.B(g3353));
  AND2 AND2_170(.VSS(VSS),.VDD(VDD),.Y(g7741),.A(g6961),.B(g3880));
  AND2 AND2_171(.VSS(VSS),.VDD(VDD),.Y(g4500),.A(g1357),.B(g3941));
  AND2 AND2_172(.VSS(VSS),.VDD(VDD),.Y(g9386),.A(g1327),.B(g9151));
  AND2 AND2_173(.VSS(VSS),.VDD(VDD),.Y(g8842),.A(g8607),.B(g8707));
  AND2 AND2_174(.VSS(VSS),.VDD(VDD),.Y(g9599),.A(g8),.B(g9292));
  AND2 AND2_175(.VSS(VSS),.VDD(VDD),.Y(g9274),.A(g8974),.B(g5708));
  AND2 AND2_176(.VSS(VSS),.VDD(VDD),.Y(g5518),.A(g4317),.B(g3532));
  AND2 AND2_177(.VSS(VSS),.VDD(VDD),.Y(g9614),.A(g1197),.B(g9111));
  AND2 AND2_178(.VSS(VSS),.VDD(VDD),.Y(g4838),.A(g3275),.B(g4122));
  AND2 AND2_179(.VSS(VSS),.VDD(VDD),.Y(g9125),.A(g8966),.B(g6674));
  AND2 AND2_180(.VSS(VSS),.VDD(VDD),.Y(g7217),.A(g4610),.B(g6432));
  AND2 AND2_181(.VSS(VSS),.VDD(VDD),.Y(g11557),.A(g2707),.B(g11519));
  AND2 AND2_182(.VSS(VSS),.VDD(VDD),.Y(g2911),.A(g2411),.B(g1675));
  AND2 AND2_183(.VSS(VSS),.VDD(VDD),.Y(g11210),.A(g11078),.B(g4515));
  AND2 AND2_184(.VSS(VSS),.VDD(VDD),.Y(g7466),.A(g7148),.B(g2821));
  AND2 AND2_185(.VSS(VSS),.VDD(VDD),.Y(g9939),.A(g9918),.B(g9367));
  AND2 AND2_186(.VSS(VSS),.VDD(VDD),.Y(g11279),.A(g4939),.B(g11200));
  AND3 AND3_7(.VSS(VSS),.VDD(VDD),.Y(g10518),.A(g10513),.B(g10440),.C(I16145));
  AND2 AND2_187(.VSS(VSS),.VDD(VDD),.Y(g4477),.A(g1129),.B(g3878));
  AND2 AND2_188(.VSS(VSS),.VDD(VDD),.Y(g8708),.A(g7605),.B(g8592));
  AND2 AND2_189(.VSS(VSS),.VDD(VDD),.Y(g7055),.A(g5900),.B(g6579));
  AND2 AND2_190(.VSS(VSS),.VDD(VDD),.Y(g5264),.A(g1095),.B(g4763));
  AND2 AND2_191(.VSS(VSS),.VDD(VDD),.Y(g6329),.A(g1265),.B(g5949));
  AND2 AND2_192(.VSS(VSS),.VDD(VDD),.Y(g6828),.A(g1377),.B(g6596));
  AND2 AND2_193(.VSS(VSS),.VDD(VDD),.Y(g8176),.A(g5299),.B(g7853));
  AND2 AND2_194(.VSS(VSS),.VDD(VDD),.Y(g6830),.A(g1380),.B(g6596));
  AND2 AND2_195(.VSS(VSS),.VDD(VDD),.Y(g8005),.A(g7510),.B(g6871));
  AND2 AND2_196(.VSS(VSS),.VDD(VDD),.Y(g4099),.A(g770),.B(g3281));
  AND2 AND2_197(.VSS(VSS),.VDD(VDD),.Y(g11601),.A(g1351),.B(g11574));
  AND2 AND2_198(.VSS(VSS),.VDD(VDD),.Y(g11187),.A(g5597),.B(g11061));
  AND2 AND2_199(.VSS(VSS),.VDD(VDD),.Y(g6746),.A(g6228),.B(g6166));
  AND2 AND2_200(.VSS(VSS),.VDD(VDD),.Y(g6221),.A(g782),.B(g5598));
  AND2 AND2_201(.VSS(VSS),.VDD(VDD),.Y(g8765),.A(g8630),.B(g5151));
  AND2 AND2_202(.VSS(VSS),.VDD(VDD),.Y(g9622),.A(g1200),.B(g9111));
  AND2 AND2_203(.VSS(VSS),.VDD(VDD),.Y(g11143),.A(g10923),.B(g4567));
  AND2 AND2_204(.VSS(VSS),.VDD(VDD),.Y(g9904),.A(g9886),.B(g9676));
  AND2 AND2_205(.VSS(VSS),.VDD(VDD),.Y(g8733),.A(g8625),.B(g7920));
  AND3 AND3_8(.VSS(VSS),.VDD(VDD),.Y(g8974),.A(g8094),.B(g6368),.C(g8858));
  AND2 AND2_206(.VSS(VSS),.VDD(VDD),.Y(g6624),.A(g348),.B(g6171));
  AND2 AND2_207(.VSS(VSS),.VDD(VDD),.Y(g11169),.A(g530),.B(g11112));
  AND2 AND2_208(.VSS(VSS),.VDD(VDD),.Y(g8073),.A(g709),.B(g7826));
  AND2 AND2_209(.VSS(VSS),.VDD(VDD),.Y(g9841),.A(g9706),.B(g9512));
  AND2 AND2_210(.VSS(VSS),.VDD(VDD),.Y(g5882),.A(g5592),.B(g3829));
  AND2 AND2_211(.VSS(VSS),.VDD(VDD),.Y(g8796),.A(g8645),.B(g8725));
  AND2 AND2_212(.VSS(VSS),.VDD(VDD),.Y(g11168),.A(g534),.B(g11112));
  AND2 AND2_213(.VSS(VSS),.VDD(VDD),.Y(g4269),.A(g1015),.B(g3914));
  AND2 AND2_214(.VSS(VSS),.VDD(VDD),.Y(g5271),.A(g727),.B(g4772));
  AND2 AND2_215(.VSS(VSS),.VDD(VDD),.Y(g10348),.A(g10272),.B(g3705));
  AND2 AND2_216(.VSS(VSS),.VDD(VDD),.Y(g5611),.A(g1047),.B(g4382));
  AND2 AND2_217(.VSS(VSS),.VDD(VDD),.Y(g8069),.A(g673),.B(g7826));
  AND2 AND2_218(.VSS(VSS),.VDD(VDD),.Y(g9695),.A(g1567),.B(g9474));
  AND2 AND2_219(.VSS(VSS),.VDD(VDD),.Y(g10304),.A(g10211),.B(g9079));
  AND2 AND2_220(.VSS(VSS),.VDD(VDD),.Y(g8469),.A(g8305),.B(g7422));
  AND2 AND2_221(.VSS(VSS),.VDD(VDD),.Y(g4712),.A(g1071),.B(g3638));
  AND2 AND2_222(.VSS(VSS),.VDD(VDD),.Y(g6576),.A(g5762),.B(g5503));
  AND2 AND2_223(.VSS(VSS),.VDD(VDD),.Y(g10622),.A(g10543),.B(g4525));
  AND2 AND2_224(.VSS(VSS),.VDD(VDD),.Y(g11015),.A(g5217),.B(g10827));
  AND2 AND2_225(.VSS(VSS),.VDD(VDD),.Y(g5674),.A(g148),.B(g5361));
  AND2 AND2_226(.VSS(VSS),.VDD(VDD),.Y(g9359),.A(g1308),.B(g9173));
  AND2 AND2_227(.VSS(VSS),.VDD(VDD),.Y(g9223),.A(g6454),.B(g8960));
  AND2 AND2_228(.VSS(VSS),.VDD(VDD),.Y(g11556),.A(g2701),.B(g11519));
  AND2 AND2_229(.VSS(VSS),.VDD(VDD),.Y(g9858),.A(g1595),.B(g9774));
  AND2 AND2_230(.VSS(VSS),.VDD(VDD),.Y(g5541),.A(g4331),.B(g3582));
  AND2 AND2_231(.VSS(VSS),.VDD(VDD),.Y(g4534),.A(g363),.B(g3586));
  AND2 AND2_232(.VSS(VSS),.VDD(VDD),.Y(g6198),.A(g1499),.B(g5128));
  AND2 AND2_233(.VSS(VSS),.VDD(VDD),.Y(g6747),.A(g2214),.B(g5897));
  AND2 AND2_234(.VSS(VSS),.VDD(VDD),.Y(g6699),.A(g6177),.B(g4221));
  AND2 AND2_235(.VSS(VSS),.VDD(VDD),.Y(g6855),.A(g1964),.B(g6392));
  AND2 AND2_236(.VSS(VSS),.VDD(VDD),.Y(g3804),.A(g3098),.B(g2203));
  AND2 AND2_237(.VSS(VSS),.VDD(VDD),.Y(g5680),.A(g153),.B(g5361));
  AND2 AND2_238(.VSS(VSS),.VDD(VDD),.Y(g9642),.A(g2654),.B(g9240));
  AND2 AND2_239(.VSS(VSS),.VDD(VDD),.Y(g5744),.A(g1528),.B(g5191));
  AND2 AND2_240(.VSS(VSS),.VDD(VDD),.Y(g10333),.A(g10262),.B(g3307));
  AND2 AND2_241(.VSS(VSS),.VDD(VDD),.Y(g8399),.A(g6094),.B(g8229));
  AND2 AND2_242(.VSS(VSS),.VDD(VDD),.Y(g9447),.A(g1762),.B(g9030));
  AND2 AND2_243(.VSS(VSS),.VDD(VDD),.Y(g4903),.A(g1849),.B(g4243));
  AND2 AND2_244(.VSS(VSS),.VDD(VDD),.Y(g11178),.A(g516),.B(g11112));
  AND2 AND2_245(.VSS(VSS),.VDD(VDD),.Y(g8510),.A(g8414),.B(g7972));
  AND2 AND2_246(.VSS(VSS),.VDD(VDD),.Y(g8245),.A(g7850),.B(g4339));
  AND2 AND2_247(.VSS(VSS),.VDD(VDD),.Y(g6319),.A(g1296),.B(g5949));
  AND2 AND2_248(.VSS(VSS),.VDD(VDD),.Y(g11186),.A(g5594),.B(g11059));
  AND2 AND2_249(.VSS(VSS),.VDD(VDD),.Y(g3908),.A(g186),.B(g3164));
  AND2 AND2_250(.VSS(VSS),.VDD(VDD),.Y(g2951),.A(g2411),.B(g1681));
  AND2 AND2_251(.VSS(VSS),.VDD(VDD),.Y(g6352),.A(g278),.B(g5894));
  AND2 AND2_252(.VSS(VSS),.VDD(VDD),.Y(g9595),.A(g901),.B(g9205));
  AND2 AND2_253(.VSS(VSS),.VDD(VDD),.Y(g4831),.A(g810),.B(g4109));
  AND2 AND2_254(.VSS(VSS),.VDD(VDD),.Y(g5492),.A(g1654),.B(g4263));
  AND2 AND2_255(.VSS(VSS),.VDD(VDD),.Y(g9272),.A(g8934),.B(g3424));
  AND2 AND2_256(.VSS(VSS),.VDD(VDD),.Y(g10312),.A(g10220),.B(g9094));
  AND2 AND2_257(.VSS(VSS),.VDD(VDD),.Y(g6186),.A(g546),.B(g5042));
  AND2 AND2_258(.VSS(VSS),.VDD(VDD),.Y(g9612),.A(g2652),.B(g9240));
  AND2 AND2_259(.VSS(VSS),.VDD(VDD),.Y(g9417),.A(g1738),.B(g9052));
  AND2 AND2_260(.VSS(VSS),.VDD(VDD),.Y(g9935),.A(g9914),.B(g9624));
  AND2 AND2_261(.VSS(VSS),.VDD(VDD),.Y(g8701),.A(g7597),.B(g8582));
  AND2 AND2_262(.VSS(VSS),.VDD(VDD),.Y(g10745),.A(g10658),.B(g3586));
  AND2 AND2_263(.VSS(VSS),.VDD(VDD),.Y(g11216),.A(g956),.B(g11162));
  AND2 AND2_264(.VSS(VSS),.VDD(VDD),.Y(g9328),.A(g8971),.B(g5708));
  AND2 AND2_265(.VSS(VSS),.VDD(VDD),.Y(g11587),.A(g1327),.B(g11546));
  AND2 AND2_266(.VSS(VSS),.VDD(VDD),.Y(g6821),.A(g237),.B(g6596));
  AND2 AND2_267(.VSS(VSS),.VDD(VDD),.Y(g6325),.A(g1245),.B(g5949));
  AND2 AND2_268(.VSS(VSS),.VDD(VDD),.Y(g4560),.A(g431),.B(g4002));
  AND2 AND2_269(.VSS(VSS),.VDD(VDD),.Y(g7368),.A(g6980),.B(g3880));
  AND2 AND2_270(.VSS(VSS),.VDD(VDD),.Y(g6083),.A(g552),.B(g5619));
  AND2 AND2_271(.VSS(VSS),.VDD(VDD),.Y(g6544),.A(g1227),.B(g6081));
  AND2 AND2_272(.VSS(VSS),.VDD(VDD),.Y(g5476),.A(g1615),.B(g4237));
  AND2 AND2_273(.VSS(VSS),.VDD(VDD),.Y(g7743),.A(g6967),.B(g3880));
  AND2 AND2_274(.VSS(VSS),.VDD(VDD),.Y(g4869),.A(g1083),.B(g3638));
  AND2 AND2_275(.VSS(VSS),.VDD(VDD),.Y(g5722),.A(g1598),.B(g5144));
  AND2 AND2_276(.VSS(VSS),.VDD(VDD),.Y(g6790),.A(g5813),.B(g4398));
  AND2 AND2_277(.VSS(VSS),.VDD(VDD),.Y(g8408),.A(g704),.B(g8139));
  AND2 AND2_278(.VSS(VSS),.VDD(VDD),.Y(g10761),.A(g10700),.B(g10699));
  AND2 AND2_279(.VSS(VSS),.VDD(VDD),.Y(g7734),.A(g6944),.B(g3880));
  AND2 AND2_280(.VSS(VSS),.VDD(VDD),.Y(g8136),.A(g7926),.B(g7045));
  AND2 AND2_281(.VSS(VSS),.VDD(VDD),.Y(g6187),.A(g5569),.B(g2340));
  AND2 AND2_282(.VSS(VSS),.VDD(VDD),.Y(g4752),.A(g401),.B(g3385));
  AND2 AND2_283(.VSS(VSS),.VDD(VDD),.Y(g9902),.A(g9894),.B(g9392));
  AND2 AND2_284(.VSS(VSS),.VDD(VDD),.Y(g8768),.A(g8623),.B(g5151));
  AND2 AND2_285(.VSS(VSS),.VDD(VDD),.Y(g5500),.A(g1657),.B(g4272));
  AND2 AND2_286(.VSS(VSS),.VDD(VDD),.Y(g2496),.A(g374),.B(g369));
  AND2 AND2_287(.VSS(VSS),.VDD(VDD),.Y(g6756),.A(g3010),.B(g5877));
  AND3 AND3_9(.VSS(VSS),.VDD(VDD),.Y(g8972),.A(g8085),.B(g6764),.C(g8858));
  AND2 AND2_288(.VSS(VSS),.VDD(VDD),.Y(g6622),.A(g336),.B(g6165));
  AND2 AND2_289(.VSS(VSS),.VDD(VDD),.Y(g11639),.A(g11612),.B(g7897));
  AND2 AND2_290(.VSS(VSS),.VDD(VDD),.Y(g9366),.A(g1311),.B(g9173));
  AND2 AND2_291(.VSS(VSS),.VDD(VDD),.Y(g11230),.A(g471),.B(g11062));
  AND2 AND2_292(.VSS(VSS),.VDD(VDD),.Y(g10328),.A(g10252),.B(g3307));
  AND2 AND2_293(.VSS(VSS),.VDD(VDD),.Y(g5024),.A(g1284),.B(g4513));
  AND2 AND2_294(.VSS(VSS),.VDD(VDD),.Y(g4364),.A(g1215),.B(g3756));
  AND2 AND2_295(.VSS(VSS),.VDD(VDD),.Y(g9649),.A(g916),.B(g9205));
  AND2 AND2_296(.VSS(VSS),.VDD(VDD),.Y(g5795),.A(g1543),.B(g5251));
  AND2 AND2_297(.VSS(VSS),.VDD(VDD),.Y(g5737),.A(g1524),.B(g5183));
  AND2 AND2_298(.VSS(VSS),.VDD(VDD),.Y(g6841),.A(g1400),.B(g6596));
  AND2 AND2_299(.VSS(VSS),.VDD(VDD),.Y(g4054),.A(g1753),.B(g2793));
  AND2 AND2_300(.VSS(VSS),.VDD(VDD),.Y(g6345),.A(g5823),.B(g4426));
  AND2 AND2_301(.VSS(VSS),.VDD(VDD),.Y(g11391),.A(g11275),.B(g7912));
  AND2 AND2_302(.VSS(VSS),.VDD(VDD),.Y(g9851),.A(g296),.B(g9770));
  AND2 AND2_303(.VSS(VSS),.VDD(VDD),.Y(g6763),.A(g5802),.B(g4381));
  AND2 AND2_304(.VSS(VSS),.VDD(VDD),.Y(g4770),.A(g416),.B(g3415));
  AND3 AND3_10(.VSS(VSS),.VDD(VDD),.Y(I16142),.A(g10511),.B(g10509),.C(g10507));
  AND2 AND2_305(.VSS(VSS),.VDD(VDD),.Y(g9698),.A(g1571),.B(g9474));
  AND2 AND2_306(.VSS(VSS),.VDD(VDD),.Y(g4725),.A(g1032),.B(g3914));
  AND2 AND2_307(.VSS(VSS),.VDD(VDD),.Y(g5477),.A(g1887),.B(g4241));
  AND2 AND2_308(.VSS(VSS),.VDD(VDD),.Y(g9964),.A(g9954),.B(g9536));
  AND2 AND2_309(.VSS(VSS),.VDD(VDD),.Y(g5523),.A(g1663),.B(g4290));
  AND2 AND2_310(.VSS(VSS),.VDD(VDD),.Y(g4553),.A(g435),.B(g3995));
  AND2 AND2_311(.VSS(VSS),.VDD(VDD),.Y(g8550),.A(g8402),.B(g8011));
  AND2 AND2_312(.VSS(VSS),.VDD(VDD),.Y(g8845),.A(g8611),.B(g8711));
  AND2 AND2_313(.VSS(VSS),.VDD(VDD),.Y(g2081),.A(g932),.B(g928));
  AND2 AND2_314(.VSS(VSS),.VDD(VDD),.Y(g6359),.A(g281),.B(g5898));
  AND2 AND2_315(.VSS(VSS),.VDD(VDD),.Y(g11586),.A(g1324),.B(g11545));
  AND2 AND2_316(.VSS(VSS),.VDD(VDD),.Y(g11007),.A(g5147),.B(g10827));
  AND2 AND2_317(.VSS(VSS),.VDD(VDD),.Y(g5104),.A(g1796),.B(g4608));
  AND2 AND2_318(.VSS(VSS),.VDD(VDD),.Y(g5099),.A(g4821),.B(g3829));
  AND2 AND2_319(.VSS(VSS),.VDD(VDD),.Y(g6757),.A(g2221),.B(g5919));
  AND2 AND2_320(.VSS(VSS),.VDD(VDD),.Y(g5499),.A(g1627),.B(g4270));
  AND2 AND2_321(.VSS(VSS),.VDD(VDD),.Y(g4389),.A(g3529),.B(g3092));
  AND2 AND2_322(.VSS(VSS),.VDD(VDD),.Y(g6416),.A(g3497),.B(g5774));
  AND2 AND2_323(.VSS(VSS),.VDD(VDD),.Y(g9720),.A(g1546),.B(g9490));
  AND2 AND2_324(.VSS(VSS),.VDD(VDD),.Y(g4990),.A(g1444),.B(g4682));
  AND2 AND2_325(.VSS(VSS),.VDD(VDD),.Y(g9619),.A(g2772),.B(g9010));
  AND4 AND4_1(.VSS(VSS),.VDD(VDD),.Y(I6630),.A(g2677),.B(g2683),.C(g2689),.D(g2701));
  AND2 AND2_326(.VSS(VSS),.VDD(VDD),.Y(g6047),.A(g2017),.B(g4977));
  AND2 AND2_327(.VSS(VSS),.VDD(VDD),.Y(g9652),.A(g953),.B(g9223));
  AND3 AND3_11(.VSS(VSS),.VDD(VDD),.Y(g10515),.A(g10505),.B(g10469),.C(I16142));
  AND2 AND2_328(.VSS(VSS),.VDD(VDD),.Y(g9843),.A(g9711),.B(g9519));
  AND2 AND2_329(.VSS(VSS),.VDD(VDD),.Y(g5273),.A(g1074),.B(g4776));
  AND2 AND2_330(.VSS(VSS),.VDD(VDD),.Y(g11465),.A(g11434),.B(g5446));
  AND2 AND2_331(.VSS(VSS),.VDD(VDD),.Y(g5044),.A(g4348),.B(g1918));
  AND2 AND2_332(.VSS(VSS),.VDD(VDD),.Y(g11237),.A(g5472),.B(g11109));
  AND2 AND2_333(.VSS(VSS),.VDD(VDD),.Y(g9834),.A(g9731),.B(g9785));
  AND2 AND2_334(.VSS(VSS),.VDD(VDD),.Y(g6654),.A(g363),.B(g6214));
  AND2 AND2_335(.VSS(VSS),.VDD(VDD),.Y(g5444),.A(g1041),.B(g4880));
  AND2 AND2_336(.VSS(VSS),.VDD(VDD),.Y(g3714),.A(g1690),.B(g2991));
  AND2 AND2_337(.VSS(VSS),.VDD(VDD),.Y(g11340),.A(g11285),.B(g4424));
  AND2 AND2_338(.VSS(VSS),.VDD(VDD),.Y(g9598),.A(g2086),.B(g9274));
  AND2 AND2_339(.VSS(VSS),.VDD(VDD),.Y(g8097),.A(g6200),.B(g7851));
  AND2 AND2_340(.VSS(VSS),.VDD(VDD),.Y(g8726),.A(g8608),.B(g7913));
  AND2 AND2_341(.VSS(VSS),.VDD(VDD),.Y(g6880),.A(g4816),.B(g6562));
  AND2 AND2_342(.VSS(VSS),.VDD(VDD),.Y(g4338),.A(g1157),.B(g3707));
  AND2 AND2_343(.VSS(VSS),.VDD(VDD),.Y(g5543),.A(g4874),.B(g4312));
  AND3 AND3_12(.VSS(VSS),.VDD(VDD),.Y(g8960),.A(g8085),.B(g6368),.C(g8828));
  AND2 AND2_344(.VSS(VSS),.VDD(VDD),.Y(g4109),.A(g806),.B(g3287));
  AND2 AND2_345(.VSS(VSS),.VDD(VDD),.Y(g10759),.A(g10698),.B(g10697));
  AND2 AND2_346(.VSS(VSS),.VDD(VDD),.Y(g9938),.A(g9917),.B(g9367));
  AND2 AND2_347(.VSS(VSS),.VDD(VDD),.Y(g10758),.A(g10652),.B(g4013));
  AND2 AND2_348(.VSS(VSS),.VDD(VDD),.Y(g4759),.A(g406),.B(g3392));
  AND2 AND2_349(.VSS(VSS),.VDD(VDD),.Y(g9909),.A(g9891),.B(g9804));
  AND2 AND2_350(.VSS(VSS),.VDD(VDD),.Y(g7127),.A(g6663),.B(g2241));
  AND2 AND2_351(.VSS(VSS),.VDD(VDD),.Y(g11165),.A(g476),.B(g11112));
  AND2 AND2_352(.VSS(VSS),.VDD(VDD),.Y(g6234),.A(g2244),.B(g5151));
  AND2 AND2_353(.VSS(VSS),.VDD(VDD),.Y(g6328),.A(g1260),.B(g5949));
  AND2 AND2_354(.VSS(VSS),.VDD(VDD),.Y(g8401),.A(g677),.B(g8124));
  AND2 AND2_355(.VSS(VSS),.VDD(VDD),.Y(g11006),.A(g5125),.B(g10827));
  AND2 AND2_356(.VSS(VSS),.VDD(VDD),.Y(g4865),.A(g1080),.B(g3638));
  AND2 AND2_357(.VSS(VSS),.VDD(VDD),.Y(g4715),.A(g1077),.B(g3638));
  AND3 AND3_13(.VSS(VSS),.VDD(VDD),.Y(g4604),.A(g3056),.B(g3753),.C(g2325));
  AND2 AND2_358(.VSS(VSS),.VDD(VDD),.Y(g5513),.A(g1675),.B(g4282));
  AND2 AND2_359(.VSS(VSS),.VDD(VDD),.Y(g11222),.A(g965),.B(g11055));
  AND2 AND2_360(.VSS(VSS),.VDD(VDD),.Y(g4498),.A(g1145),.B(g3940));
  AND2 AND2_361(.VSS(VSS),.VDD(VDD),.Y(g6554),.A(g5075),.B(g6183));
  AND2 AND2_362(.VSS(VSS),.VDD(VDD),.Y(g7732),.A(g6935),.B(g3880));
  AND2 AND2_363(.VSS(VSS),.VDD(VDD),.Y(g9586),.A(g2727),.B(g9173));
  AND3 AND3_14(.VSS(VSS),.VDD(VDD),.Y(g5178),.A(g2047),.B(g4401),.C(g4104));
  AND2 AND2_364(.VSS(VSS),.VDD(VDD),.Y(g4584),.A(g3710),.B(g2322));
  AND2 AND2_365(.VSS(VSS),.VDD(VDD),.Y(g7472),.A(g7148),.B(g2829));
  AND2 AND2_366(.VSS(VSS),.VDD(VDD),.Y(g11253),.A(g981),.B(g11072));
  AND2 AND2_367(.VSS(VSS),.VDD(VDD),.Y(g5182),.A(g1240),.B(g4713));
  AND2 AND2_368(.VSS(VSS),.VDD(VDD),.Y(g9860),.A(g1598),.B(g9775));
  AND2 AND2_369(.VSS(VSS),.VDD(VDD),.Y(g8703),.A(g7601),.B(g8585));
  AND2 AND2_370(.VSS(VSS),.VDD(VDD),.Y(g11600),.A(g1346),.B(g11573));
  AND2 AND2_371(.VSS(VSS),.VDD(VDD),.Y(g9710),.A(g1586),.B(g9474));
  AND2 AND2_372(.VSS(VSS),.VDD(VDD),.Y(g9645),.A(g1203),.B(g9111));
  AND2 AND2_373(.VSS(VSS),.VDD(VDD),.Y(g11236),.A(g5469),.B(g11108));
  AND2 AND2_374(.VSS(VSS),.VDD(VDD),.Y(g4162),.A(g3106),.B(g2971));
  AND2 AND2_375(.VSS(VSS),.VDD(VDD),.Y(g6090),.A(g553),.B(g5627));
  AND2 AND2_376(.VSS(VSS),.VDD(VDD),.Y(g9691),.A(g269),.B(g9432));
  AND2 AND2_377(.VSS(VSS),.VDD(VDD),.Y(g11372),.A(g11316),.B(g4266));
  AND2 AND2_378(.VSS(VSS),.VDD(VDD),.Y(g6823),.A(g1368),.B(g6596));
  AND2 AND2_379(.VSS(VSS),.VDD(VDD),.Y(g11175),.A(g501),.B(g11112));
  AND2 AND2_380(.VSS(VSS),.VDD(VDD),.Y(g8068),.A(g664),.B(g7826));
  AND2 AND2_381(.VSS(VSS),.VDD(VDD),.Y(g9607),.A(g12),.B(g9274));
  AND2 AND2_382(.VSS(VSS),.VDD(VDD),.Y(g9962),.A(g9952),.B(g9536));
  AND2 AND2_383(.VSS(VSS),.VDD(VDD),.Y(g6348),.A(g296),.B(g5891));
  AND2 AND2_384(.VSS(VSS),.VDD(VDD),.Y(g9659),.A(g956),.B(g9223));
  AND2 AND2_385(.VSS(VSS),.VDD(VDD),.Y(g9358),.A(g1318),.B(g9151));
  AND2 AND2_386(.VSS(VSS),.VDD(VDD),.Y(g3104),.A(I6316),.B(I6317));
  AND2 AND2_387(.VSS(VSS),.VDD(VDD),.Y(g4486),.A(g1711),.B(g3910));
  AND2 AND2_388(.VSS(VSS),.VDD(VDD),.Y(g9587),.A(g892),.B(g8995));
  AND2 AND2_389(.VSS(VSS),.VDD(VDD),.Y(g5632),.A(g1636),.B(g4563));
  AND2 AND2_390(.VSS(VSS),.VDD(VDD),.Y(g9111),.A(g8965),.B(g6674));
  AND2 AND2_391(.VSS(VSS),.VDD(VDD),.Y(g4881),.A(g991),.B(g3914));
  AND2 AND2_392(.VSS(VSS),.VDD(VDD),.Y(g11209),.A(g11074),.B(g9448));
  AND2 AND2_393(.VSS(VSS),.VDD(VDD),.Y(g8848),.A(g8715),.B(g8713));
  AND2 AND2_394(.VSS(VSS),.VDD(VDD),.Y(g4070),.A(g3263),.B(g2330));
  AND2 AND2_395(.VSS(VSS),.VDD(VDD),.Y(g6463),.A(g5052),.B(g6210));
  AND2 AND2_396(.VSS(VSS),.VDD(VDD),.Y(g8699),.A(g7595),.B(g8579));
  AND4 AND4_2(.VSS(VSS),.VDD(VDD),.Y(I5689),.A(g1419),.B(g1424),.C(g1428),.D(g1432));
  AND2 AND2_397(.VSS(VSS),.VDD(VDD),.Y(g7820),.A(g1896),.B(g7479));
  AND2 AND2_398(.VSS(VSS),.VDD(VDD),.Y(g11021),.A(g448),.B(g10974));
  AND2 AND2_399(.VSS(VSS),.VDD(VDD),.Y(g5917),.A(g1044),.B(g5320));
  AND2 AND2_400(.VSS(VSS),.VDD(VDD),.Y(g6619),.A(g49),.B(g6156));
  AND2 AND2_401(.VSS(VSS),.VDD(VDD),.Y(g6318),.A(g1300),.B(g5949));
  AND2 AND2_402(.VSS(VSS),.VDD(VDD),.Y(g6872),.A(g1896),.B(g6389));
  AND2 AND2_403(.VSS(VSS),.VDD(VDD),.Y(g11320),.A(g11201),.B(g4379));
  AND2 AND2_404(.VSS(VSS),.VDD(VDD),.Y(g10514),.A(g10489),.B(g4580));
  AND2 AND2_405(.VSS(VSS),.VDD(VDD),.Y(g4006),.A(g201),.B(g3228));
  AND2 AND2_406(.VSS(VSS),.VDD(VDD),.Y(g9853),.A(g299),.B(g9771));
  AND2 AND2_407(.VSS(VSS),.VDD(VDD),.Y(g11274),.A(g4913),.B(g11197));
  AND2 AND2_408(.VSS(VSS),.VDD(VDD),.Y(g6193),.A(g2206),.B(g5151));
  AND2 AND2_409(.VSS(VSS),.VDD(VDD),.Y(g8119),.A(g6239),.B(g7890));
  AND2 AND2_410(.VSS(VSS),.VDD(VDD),.Y(g9420),.A(g1747),.B(g9030));
  AND2 AND2_411(.VSS(VSS),.VDD(VDD),.Y(g5233),.A(g1791),.B(g4492));
  AND2 AND2_412(.VSS(VSS),.VDD(VDD),.Y(g7581),.A(g7092),.B(g5420));
  AND2 AND2_413(.VSS(VSS),.VDD(VDD),.Y(g6549),.A(g5515),.B(g6175));
  AND2 AND2_414(.VSS(VSS),.VDD(VDD),.Y(g11464),.A(g11433),.B(g5446));
  AND2 AND2_415(.VSS(VSS),.VDD(VDD),.Y(g4801),.A(g516),.B(g3439));
  AND2 AND2_416(.VSS(VSS),.VDD(VDD),.Y(g6834),.A(g1365),.B(g6596));
  AND2 AND2_417(.VSS(VSS),.VDD(VDD),.Y(g4487),.A(g1718),.B(g3911));
  AND2 AND2_418(.VSS(VSS),.VDD(VDD),.Y(g2939),.A(g2411),.B(g1687));
  AND2 AND2_419(.VSS(VSS),.VDD(VDD),.Y(g7060),.A(g6739),.B(g5521));
  AND2 AND2_420(.VSS(VSS),.VDD(VDD),.Y(g5770),.A(g4466),.B(g5128));
  AND2 AND2_421(.VSS(VSS),.VDD(VDD),.Y(g5725),.A(g1580),.B(g5166));
  AND2 AND2_422(.VSS(VSS),.VDD(VDD),.Y(g11641),.A(g11615),.B(g7901));
  AND2 AND2_423(.VSS(VSS),.VDD(VDD),.Y(g2544),.A(g1341),.B(g1336));
  AND2 AND2_424(.VSS(VSS),.VDD(VDD),.Y(g11292),.A(g11252),.B(g4250));
  AND2 AND2_425(.VSS(VSS),.VDD(VDD),.Y(g5532),.A(g1681),.B(g4307));
  AND2 AND2_426(.VSS(VSS),.VDD(VDD),.Y(g11153),.A(g3771),.B(g10913));
  AND2 AND2_427(.VSS(VSS),.VDD(VDD),.Y(g9905),.A(g9872),.B(g9680));
  AND2 AND2_428(.VSS(VSS),.VDD(VDD),.Y(g7739),.A(g6957),.B(g3880));
  AND2 AND2_429(.VSS(VSS),.VDD(VDD),.Y(g6321),.A(g1284),.B(g5949));
  AND2 AND2_430(.VSS(VSS),.VDD(VDD),.Y(g8386),.A(g6085),.B(g8219));
  AND3 AND3_15(.VSS(VSS),.VDD(VDD),.Y(g8975),.A(g8089),.B(g6764),.C(g8858));
  AND2 AND2_431(.VSS(VSS),.VDD(VDD),.Y(g2306),.A(g1223),.B(g1218));
  AND2 AND2_432(.VSS(VSS),.VDD(VDD),.Y(g6625),.A(g1218),.B(g6178));
  AND2 AND2_433(.VSS(VSS),.VDD(VDD),.Y(g7937),.A(g7606),.B(g4013));
  AND2 AND2_434(.VSS(VSS),.VDD(VDD),.Y(g10788),.A(g8303),.B(g10754));
  AND2 AND2_435(.VSS(VSS),.VDD(VDD),.Y(g10325),.A(g10248),.B(g3307));
  AND2 AND2_436(.VSS(VSS),.VDD(VDD),.Y(g8170),.A(g5270),.B(g7853));
  AND2 AND2_437(.VSS(VSS),.VDD(VDD),.Y(g5706),.A(g1574),.B(g5121));
  AND2 AND2_438(.VSS(VSS),.VDD(VDD),.Y(g2756),.A(g936),.B(g2081));
  AND2 AND2_439(.VSS(VSS),.VDD(VDD),.Y(g8821),.A(g8643),.B(g8751));
  AND2 AND2_440(.VSS(VSS),.VDD(VDD),.Y(g10946),.A(g5225),.B(g10827));
  AND2 AND2_441(.VSS(VSS),.VDD(VDD),.Y(g4169),.A(g2765),.B(g3066));
  AND2 AND2_442(.VSS(VSS),.VDD(VDD),.Y(g5029),.A(g1077),.B(g4521));
  AND2 AND2_443(.VSS(VSS),.VDD(VDD),.Y(g11164),.A(g4889),.B(g11112));
  AND2 AND2_444(.VSS(VSS),.VDD(VDD),.Y(g4007),.A(g2683),.B(g2276));
  AND2 AND2_445(.VSS(VSS),.VDD(VDD),.Y(g4059),.A(g1756),.B(g2796));
  AND2 AND2_446(.VSS(VSS),.VDD(VDD),.Y(g4868),.A(g1027),.B(g3914));
  AND2 AND2_447(.VSS(VSS),.VDD(VDD),.Y(g5675),.A(g131),.B(g5361));
  AND2 AND2_448(.VSS(VSS),.VDD(VDD),.Y(g4718),.A(g650),.B(g3343));
  AND2 AND2_449(.VSS(VSS),.VDD(VDD),.Y(g10682),.A(g10600),.B(g3863));
  AND2 AND2_450(.VSS(VSS),.VDD(VDD),.Y(g6687),.A(g5486),.B(g5840));
  AND2 AND2_451(.VSS(VSS),.VDD(VDD),.Y(g7704),.A(g682),.B(g7197));
  AND2 AND2_452(.VSS(VSS),.VDD(VDD),.Y(g4582),.A(g525),.B(g4055));
  AND2 AND2_453(.VSS(VSS),.VDD(VDD),.Y(g4261),.A(g1019),.B(g3914));
  AND2 AND2_454(.VSS(VSS),.VDD(VDD),.Y(g3422),.A(g225),.B(g3228));
  AND2 AND2_455(.VSS(VSS),.VDD(VDD),.Y(g5745),.A(g1549),.B(g5192));
  AND2 AND2_456(.VSS(VSS),.VDD(VDD),.Y(g8387),.A(g6086),.B(g8220));
  AND2 AND2_457(.VSS(VSS),.VDD(VDD),.Y(g7954),.A(g2874),.B(g7512));
  AND2 AND2_458(.VSS(VSS),.VDD(VDD),.Y(g11283),.A(g4966),.B(g11205));
  AND2 AND2_459(.VSS(VSS),.VDD(VDD),.Y(g8461),.A(g8298),.B(g7403));
  AND2 AND2_460(.VSS(VSS),.VDD(VDD),.Y(g10760),.A(g10695),.B(g10691));
  AND2 AND2_461(.VSS(VSS),.VDD(VDD),.Y(g11492),.A(g11480),.B(g4807));
  AND3 AND3_16(.VSS(VSS),.VDD(VDD),.Y(g7032),.A(g2965),.B(g6626),.C(g5292));
  AND2 AND2_462(.VSS(VSS),.VDD(VDD),.Y(g8756),.A(g7431),.B(g8674));
  AND2 AND2_463(.VSS(VSS),.VDD(VDD),.Y(g9151),.A(g8967),.B(g6674));
  AND2 AND2_464(.VSS(VSS),.VDD(VDD),.Y(g6341),.A(g272),.B(g5885));
  AND2 AND2_465(.VSS(VSS),.VDD(VDD),.Y(g10506),.A(g10390),.B(g2135));
  AND2 AND2_466(.VSS(VSS),.VDD(VDD),.Y(g9648),.A(g16),.B(g9274));
  AND2 AND2_467(.VSS(VSS),.VDD(VDD),.Y(g7453),.A(g7148),.B(g2809));
  AND2 AND2_468(.VSS(VSS),.VDD(VDD),.Y(g6525),.A(g5995),.B(g3102));
  AND2 AND2_469(.VSS(VSS),.VDD(VDD),.Y(g6645),.A(g67),.B(g6202));
  AND2 AND2_470(.VSS(VSS),.VDD(VDD),.Y(g5707),.A(g1595),.B(g5122));
  AND2 AND2_471(.VSS(VSS),.VDD(VDD),.Y(g8046),.A(g7548),.B(g5128));
  AND2 AND2_472(.VSS(VSS),.VDD(VDD),.Y(g11091),.A(g833),.B(g10950));
  AND2 AND2_473(.VSS(VSS),.VDD(VDD),.Y(g11174),.A(g496),.B(g11112));
  AND2 AND2_474(.VSS(VSS),.VDD(VDD),.Y(g9010),.A(g6454),.B(g8930));
  AND2 AND2_475(.VSS(VSS),.VDD(VDD),.Y(g8403),.A(g6101),.B(g8239));
  AND2 AND2_476(.VSS(VSS),.VDD(VDD),.Y(g5201),.A(g1250),.B(g4721));
  AND2 AND2_477(.VSS(VSS),.VDD(VDD),.Y(g8841),.A(g8605),.B(g8704));
  AND2 AND2_478(.VSS(VSS),.VDD(VDD),.Y(g6879),.A(g1914),.B(g6407));
  AND2 AND2_479(.VSS(VSS),.VDD(VDD),.Y(g8763),.A(g7440),.B(g8680));
  AND2 AND2_480(.VSS(VSS),.VDD(VDD),.Y(g4502),.A(g2031),.B(g3938));
  AND2 AND2_481(.VSS(VSS),.VDD(VDD),.Y(g9839),.A(g9702),.B(g9742));
  AND2 AND2_482(.VSS(VSS),.VDD(VDD),.Y(g6358),.A(g5841),.B(g4441));
  AND2 AND2_483(.VSS(VSS),.VDD(VDD),.Y(g5575),.A(g1618),.B(g4501));
  AND2 AND2_484(.VSS(VSS),.VDD(VDD),.Y(g4940),.A(g3500),.B(g4440));
  AND2 AND2_485(.VSS(VSS),.VDD(VDD),.Y(g8107),.A(g6226),.B(g7882));
  AND2 AND2_486(.VSS(VSS),.VDD(VDD),.Y(g10240),.A(g10150),.B(g9103));
  AND2 AND2_487(.VSS(VSS),.VDD(VDD),.Y(g11192),.A(g5628),.B(g11066));
  AND2 AND2_488(.VSS(VSS),.VDD(VDD),.Y(g9618),.A(g910),.B(g9205));
  AND2 AND2_489(.VSS(VSS),.VDD(VDD),.Y(g5539),.A(g1684),.B(g4314));
  AND2 AND2_490(.VSS(VSS),.VDD(VDD),.Y(g8416),.A(g731),.B(g8151));
  AND2 AND2_491(.VSS(VSS),.VDD(VDD),.Y(g9693),.A(g275),.B(g9432));
  AND2 AND2_492(.VSS(VSS),.VDD(VDD),.Y(g11553),.A(g2683),.B(g11519));
  AND2 AND2_493(.VSS(VSS),.VDD(VDD),.Y(g8047),.A(g7557),.B(g5919));
  AND2 AND2_494(.VSS(VSS),.VDD(VDD),.Y(g5268),.A(g1098),.B(g4769));
  AND2 AND2_495(.VSS(VSS),.VDD(VDD),.Y(g9555),.A(g9107),.B(g3391));
  AND2 AND2_496(.VSS(VSS),.VDD(VDD),.Y(g6180),.A(g2190),.B(g5128));
  AND2 AND2_497(.VSS(VSS),.VDD(VDD),.Y(g6832),.A(g1383),.B(g6596));
  AND2 AND2_498(.VSS(VSS),.VDD(VDD),.Y(g10633),.A(g10600),.B(g3829));
  AND2 AND2_499(.VSS(VSS),.VDD(VDD),.Y(g7894),.A(g7617),.B(g3816));
  AND2 AND2_500(.VSS(VSS),.VDD(VDD),.Y(g8654),.A(g8529),.B(g4013));
  AND2 AND2_501(.VSS(VSS),.VDD(VDD),.Y(g9621),.A(g1179),.B(g9125));
  AND2 AND2_502(.VSS(VSS),.VDD(VDD),.Y(g6794),.A(g5819),.B(g4415));
  AND2 AND2_503(.VSS(VSS),.VDD(VDD),.Y(g9313),.A(g8876),.B(g5708));
  AND2 AND2_504(.VSS(VSS),.VDD(VDD),.Y(g4883),.A(g248),.B(g3946));
  AND2 AND2_505(.VSS(VSS),.VDD(VDD),.Y(g3412),.A(g219),.B(g3228));
  AND2 AND2_506(.VSS(VSS),.VDD(VDD),.Y(g7661),.A(g7127),.B(g2251));
  AND3 AND3_17(.VSS(VSS),.VDD(VDD),.Y(g2800),.A(g2399),.B(g2369),.C(g591));
  AND2 AND2_507(.VSS(VSS),.VDD(VDD),.Y(g3389),.A(g207),.B(g3228));
  AND2 AND2_508(.VSS(VSS),.VDD(VDD),.Y(g3706),.A(g471),.B(g3268));
  AND2 AND2_509(.VSS(VSS),.VDD(VDD),.Y(g9908),.A(g9890),.B(g9782));
  AND2 AND2_510(.VSS(VSS),.VDD(VDD),.Y(g3429),.A(g231),.B(g3228));
  AND2 AND2_511(.VSS(VSS),.VDD(VDD),.Y(g6628),.A(g351),.B(g6182));
  AND2 AND2_512(.VSS(VSS),.VDD(VDD),.Y(g5470),.A(g1044),.B(g4222));
  AND2 AND2_513(.VSS(VSS),.VDD(VDD),.Y(g7526),.A(g7148),.B(g2868));
  AND2 AND2_514(.VSS(VSS),.VDD(VDD),.Y(g5897),.A(g2204),.B(g5354));
  AND2 AND2_515(.VSS(VSS),.VDD(VDD),.Y(g5025),.A(g1482),.B(g4640));
  AND2 AND2_516(.VSS(VSS),.VDD(VDD),.Y(g6204),.A(g3738),.B(g4921));
  AND2 AND2_517(.VSS(VSS),.VDD(VDD),.Y(g4048),.A(g1750),.B(g2790));
  AND3 AND3_18(.VSS(VSS),.VDD(VDD),.Y(g8935),.A(g8106),.B(g6778),.C(g8849));
  AND2 AND2_518(.VSS(VSS),.VDD(VDD),.Y(g3281),.A(g766),.B(g2525));
  AND2 AND2_519(.VSS(VSS),.VDD(VDD),.Y(g9593),.A(g898),.B(g9205));
  AND2 AND2_520(.VSS(VSS),.VDD(VDD),.Y(g4827),.A(g213),.B(g3946));
  AND2 AND2_521(.VSS(VSS),.VDD(VDD),.Y(g10701),.A(g10620),.B(g10619));
  AND2 AND2_522(.VSS(VSS),.VDD(VDD),.Y(g10777),.A(g10733),.B(g3015));
  AND2 AND2_523(.VSS(VSS),.VDD(VDD),.Y(g8130),.A(g1936),.B(g7952));
  AND2 AND2_524(.VSS(VSS),.VDD(VDD),.Y(g9965),.A(g9955),.B(g9536));
  AND2 AND2_525(.VSS(VSS),.VDD(VDD),.Y(g3684),.A(g1710),.B(g3015));
  AND2 AND2_526(.VSS(VSS),.VDD(VDD),.Y(g11213),.A(g947),.B(g11157));
  AND2 AND2_527(.VSS(VSS),.VDD(VDD),.Y(g5006),.A(g1462),.B(g4640));
  AND2 AND2_528(.VSS(VSS),.VDD(VDD),.Y(g9933),.A(g9912),.B(g9624));
  AND2 AND2_529(.VSS(VSS),.VDD(VDD),.Y(g8554),.A(g8407),.B(g8020));
  AND2 AND2_530(.VSS(VSS),.VDD(VDD),.Y(g9641),.A(g913),.B(g9205));
  AND2 AND2_531(.VSS(VSS),.VDD(VDD),.Y(g6123),.A(g5630),.B(g4311));
  AND2 AND2_532(.VSS(VSS),.VDD(VDD),.Y(g6323),.A(g1235),.B(g5949));
  AND2 AND2_533(.VSS(VSS),.VDD(VDD),.Y(g10766),.A(g10646),.B(g4840));
  AND2 AND2_534(.VSS(VSS),.VDD(VDD),.Y(g6666),.A(g5301),.B(g5818));
  AND2 AND2_535(.VSS(VSS),.VDD(VDD),.Y(g4994),.A(g1504),.B(g4640));
  AND2 AND2_536(.VSS(VSS),.VDD(VDD),.Y(g5755),.A(g5103),.B(g5354));
  AND2 AND2_537(.VSS(VSS),.VDD(VDD),.Y(g11592),.A(g3717),.B(g11561));
  AND2 AND2_538(.VSS(VSS),.VDD(VDD),.Y(g6351),.A(g6210),.B(g5052));
  AND2 AND2_539(.VSS(VSS),.VDD(VDD),.Y(g6875),.A(g1905),.B(g6400));
  AND2 AND2_540(.VSS(VSS),.VDD(VDD),.Y(g4816),.A(g4070),.B(g2336));
  AND2 AND2_541(.VSS(VSS),.VDD(VDD),.Y(g9658),.A(g947),.B(g9240));
  AND2 AND2_542(.VSS(VSS),.VDD(VDD),.Y(g6530),.A(g6207),.B(g3829));
  AND2 AND2_543(.VSS(VSS),.VDD(VDD),.Y(g8366),.A(g8199),.B(g7265));
  AND2 AND2_544(.VSS(VSS),.VDD(VDD),.Y(g9835),.A(g9735),.B(g9785));
  AND2 AND2_545(.VSS(VSS),.VDD(VDD),.Y(g6655),.A(g5296),.B(g5812));
  AND3 AND3_19(.VSS(VSS),.VDD(VDD),.Y(g5445),.A(g4631),.B(g3875),.C(g2733));
  AND2 AND2_546(.VSS(VSS),.VDD(VDD),.Y(g5173),.A(g3094),.B(g4676));
  AND2 AND2_547(.VSS(VSS),.VDD(VDD),.Y(g7970),.A(g7384),.B(g7703));
  AND2 AND2_548(.VSS(VSS),.VDD(VDD),.Y(g3098),.A(g2331),.B(g2198));
  AND2 AND2_549(.VSS(VSS),.VDD(VDD),.Y(g5491),.A(g1624),.B(g4262));
  AND2 AND2_550(.VSS(VSS),.VDD(VDD),.Y(g9271),.A(g6681),.B(g8949));
  AND2 AND2_551(.VSS(VSS),.VDD(VDD),.Y(g11152),.A(g369),.B(g10903));
  AND2 AND2_552(.VSS(VSS),.VDD(VDD),.Y(g9611),.A(g2651),.B(g9010));
  AND2 AND2_553(.VSS(VSS),.VDD(VDD),.Y(g6410),.A(g2804),.B(g5759));
  AND2 AND2_554(.VSS(VSS),.VDD(VDD),.Y(g10451),.A(g10444),.B(g3365));
  AND2 AND2_555(.VSS(VSS),.VDD(VDD),.Y(g4397),.A(g3475),.B(g2181));
  AND2 AND2_556(.VSS(VSS),.VDD(VDD),.Y(g7224),.A(g5398),.B(g6441));
  AND2 AND2_557(.VSS(VSS),.VDD(VDD),.Y(g5602),.A(g1624),.B(g4535));
  AND2 AND2_558(.VSS(VSS),.VDD(VDD),.Y(g4421),.A(g4112),.B(g2980));
  AND2 AND2_559(.VSS(VSS),.VDD(VDD),.Y(g6884),.A(g5569),.B(g6564));
  AND2 AND2_560(.VSS(VSS),.VDD(VDD),.Y(g6839),.A(g1397),.B(g6596));
  AND2 AND2_561(.VSS(VSS),.VDD(VDD),.Y(g8698),.A(g7591),.B(g8576));
  AND3 AND3_20(.VSS(VSS),.VDD(VDD),.Y(g8964),.A(g8255),.B(g6368),.C(g8849));
  AND2 AND2_562(.VSS(VSS),.VDD(VDD),.Y(g8260),.A(g2775),.B(g7911));
  AND2 AND2_563(.VSS(VSS),.VDD(VDD),.Y(g11413),.A(g11354),.B(g10679));
  AND2 AND2_564(.VSS(VSS),.VDD(VDD),.Y(g4950),.A(g1415),.B(g4682));
  AND2 AND2_565(.VSS(VSS),.VDD(VDD),.Y(g5535),.A(g4327),.B(g3544));
  AND2 AND2_566(.VSS(VSS),.VDD(VDD),.Y(g7277),.A(g6772),.B(g731));
  AND2 AND2_567(.VSS(VSS),.VDD(VDD),.Y(g8463),.A(g8301),.B(g7410));
  AND2 AND2_568(.VSS(VSS),.VDD(VDD),.Y(g3268),.A(g466),.B(g2511));
  AND2 AND2_569(.VSS(VSS),.VDD(VDD),.Y(g10785),.A(g10728),.B(g5177));
  AND2 AND2_570(.VSS(VSS),.VDD(VDD),.Y(g6618),.A(g658),.B(g6016));
  AND2 AND2_571(.VSS(VSS),.VDD(VDD),.Y(g6235),.A(g569),.B(g5089));
  AND2 AND2_572(.VSS(VSS),.VDD(VDD),.Y(g10950),.A(g10788),.B(g6355));
  AND2 AND2_573(.VSS(VSS),.VDD(VDD),.Y(g4723),.A(g3626),.B(g2779));
  AND2 AND2_574(.VSS(VSS),.VDD(VDD),.Y(g8720),.A(g8601),.B(g7905));
  AND2 AND2_575(.VSS(VSS),.VDD(VDD),.Y(g6693),.A(g5494),.B(g5845));
  AND2 AND2_576(.VSS(VSS),.VDD(VDD),.Y(g11020),.A(g452),.B(g10974));
  AND2 AND2_577(.VSS(VSS),.VDD(VDD),.Y(g11583),.A(g1314),.B(g11541));
  AND2 AND2_578(.VSS(VSS),.VDD(VDD),.Y(g8118),.A(g1900),.B(g7941));
  AND2 AND2_579(.VSS(VSS),.VDD(VDD),.Y(g8167),.A(g5253),.B(g7853));
  AND2 AND2_580(.VSS(VSS),.VDD(VDD),.Y(g6334),.A(g1389),.B(g5904));
  AND2 AND2_581(.VSS(VSS),.VDD(VDD),.Y(g7892),.A(g7616),.B(g3815));
  AND2 AND2_582(.VSS(VSS),.VDD(VDD),.Y(g8652),.A(g8523),.B(g4013));
  AND2 AND2_583(.VSS(VSS),.VDD(VDD),.Y(g5721),.A(g1577),.B(g5143));
  AND2 AND2_584(.VSS(VSS),.VDD(VDD),.Y(g10367),.A(g10362),.B(g3375));
  AND2 AND2_585(.VSS(VSS),.VDD(VDD),.Y(g9901),.A(g9893),.B(g9392));
  AND2 AND2_586(.VSS(VSS),.VDD(VDD),.Y(g6792),.A(g290),.B(g5881));
  AND2 AND2_587(.VSS(VSS),.VDD(VDD),.Y(g11282),.A(g4958),.B(g11203));
  AND2 AND2_588(.VSS(VSS),.VDD(VDD),.Y(g7945),.A(g2847),.B(g7473));
  AND3 AND3_21(.VSS(VSS),.VDD(VDD),.Y(g8971),.A(g8081),.B(g6764),.C(g8858));
  AND2 AND2_589(.VSS(VSS),.VDD(VDD),.Y(g11302),.A(g5508),.B(g11244));
  AND2 AND2_590(.VSS(VSS),.VDD(VDD),.Y(g4585),.A(g521),.B(g4060));
  AND2 AND2_591(.VSS(VSS),.VDD(VDD),.Y(g6621),.A(g52),.B(g6164));
  AND2 AND2_592(.VSS(VSS),.VDD(VDD),.Y(g5502),.A(g1932),.B(g4275));
  AND2 AND2_593(.VSS(VSS),.VDD(VDD),.Y(g11105),.A(g3634),.B(g10937));
  AND2 AND2_594(.VSS(VSS),.VDD(VDD),.Y(g7709),.A(g6856),.B(g4333));
  AND2 AND2_595(.VSS(VSS),.VDD(VDD),.Y(g8598),.A(g8471),.B(g7432));
  AND2 AND2_596(.VSS(VSS),.VDD(VDD),.Y(g7140),.A(g6069),.B(g6711));
  AND2 AND2_597(.VSS(VSS),.VDD(VDD),.Y(g9600),.A(g904),.B(g9205));
  AND2 AND2_598(.VSS(VSS),.VDD(VDD),.Y(g9864),.A(g1604),.B(g9778));
  AND2 AND2_599(.VSS(VSS),.VDD(VDD),.Y(g11640),.A(g11613),.B(g7900));
  AND2 AND2_600(.VSS(VSS),.VDD(VDD),.Y(g5188),.A(g4504),.B(g4496));
  AND2 AND2_601(.VSS(VSS),.VDD(VDD),.Y(g7435),.A(g7260),.B(g6572));
  AND2 AND2_602(.VSS(VSS),.VDD(VDD),.Y(g7876),.A(g7609),.B(g3790));
  AND2 AND2_603(.VSS(VSS),.VDD(VDD),.Y(g5030),.A(g1280),.B(g4523));
  AND2 AND2_604(.VSS(VSS),.VDD(VDD),.Y(g4058),.A(g2707),.B(g2276));
  AND2 AND2_605(.VSS(VSS),.VDD(VDD),.Y(g6776),.A(g5809),.B(g4390));
  AND2 AND2_606(.VSS(VSS),.VDD(VDD),.Y(g4890),.A(g630),.B(g4739));
  AND2 AND2_607(.VSS(VSS),.VDD(VDD),.Y(g2525),.A(g762),.B(g758));
  AND2 AND2_608(.VSS(VSS),.VDD(VDD),.Y(g10301),.A(g8892),.B(g10223));
  AND2 AND2_609(.VSS(VSS),.VDD(VDD),.Y(g4505),.A(g354),.B(g3586));
  AND2 AND2_610(.VSS(VSS),.VDD(VDD),.Y(g9623),.A(g17),.B(g9274));
  AND2 AND2_611(.VSS(VSS),.VDD(VDD),.Y(g10739),.A(g10676),.B(g3368));
  AND2 AND2_612(.VSS(VSS),.VDD(VDD),.Y(g11027),.A(g391),.B(g10974));
  AND2 AND2_613(.VSS(VSS),.VDD(VDD),.Y(g10738),.A(g10692),.B(g4840));
  AND2 AND2_614(.VSS(VSS),.VDD(VDD),.Y(g8687),.A(g8558),.B(g8036));
  AND2 AND2_615(.VSS(VSS),.VDD(VDD),.Y(g6360),.A(g302),.B(g5899));
  AND2 AND2_616(.VSS(VSS),.VDD(VDD),.Y(g9871),.A(g1564),.B(g9668));
  AND2 AND2_617(.VSS(VSS),.VDD(VDD),.Y(g5108),.A(g1801),.B(g4614));
  AND2 AND2_618(.VSS(VSS),.VDD(VDD),.Y(g11248),.A(g976),.B(g11071));
  AND2 AND2_619(.VSS(VSS),.VDD(VDD),.Y(g4992),.A(g1407),.B(g4682));
  AND2 AND2_620(.VSS(VSS),.VDD(VDD),.Y(g11552),.A(g2677),.B(g11519));
  AND2 AND2_621(.VSS(VSS),.VDD(VDD),.Y(g9651),.A(g944),.B(g9240));
  AND2 AND2_622(.VSS(VSS),.VDD(VDD),.Y(g11204),.A(g971),.B(g11083));
  AND2 AND2_623(.VSS(VSS),.VDD(VDD),.Y(g7824),.A(g1932),.B(g7479));
  AND2 AND2_624(.VSS(VSS),.VDD(VDD),.Y(g4480),.A(g1133),.B(g3905));
  AND2 AND2_625(.VSS(VSS),.VDD(VDD),.Y(g6179),.A(g5115),.B(g5354));
  AND2 AND2_626(.VSS(VSS),.VDD(VDD),.Y(g8710),.A(g7607),.B(g8595));
  AND2 AND2_627(.VSS(VSS),.VDD(VDD),.Y(g7590),.A(g7102),.B(g5425));
  AND2 AND2_628(.VSS(VSS),.VDD(VDD),.Y(g9384),.A(g968),.B(g9223));
  AND2 AND2_629(.VSS(VSS),.VDD(VDD),.Y(g3407),.A(g2561),.B(g3012));
  AND2 AND2_630(.VSS(VSS),.VDD(VDD),.Y(g9838),.A(g9700),.B(g9754));
  AND2 AND2_631(.VSS(VSS),.VDD(VDD),.Y(g3718),.A(g192),.B(g3164));
  AND2 AND2_632(.VSS(VSS),.VDD(VDD),.Y(g10661),.A(g10594),.B(g3015));
  AND2 AND2_633(.VSS(VSS),.VDD(VDD),.Y(g11380),.A(g11321),.B(g4285));
  AND3 AND3_22(.VSS(VSS),.VDD(VDD),.Y(g8879),.A(g8110),.B(g6764),.C(g8858));
  AND2 AND2_634(.VSS(VSS),.VDD(VDD),.Y(g7930),.A(g7621),.B(g3110));
  AND3 AND3_23(.VSS(VSS),.VDD(VDD),.Y(g8962),.A(g8089),.B(g6368),.C(g8828));
  AND2 AND2_635(.VSS(VSS),.VDD(VDD),.Y(g10715),.A(g2272),.B(g10630));
  AND2 AND2_636(.VSS(VSS),.VDD(VDD),.Y(g8659),.A(g8535),.B(g4013));
  AND2 AND2_637(.VSS(VSS),.VDD(VDD),.Y(g3015),.A(g2028),.B(g2191));
  AND2 AND2_638(.VSS(VSS),.VDD(VDD),.Y(g9643),.A(g950),.B(g9223));
  AND2 AND2_639(.VSS(VSS),.VDD(VDD),.Y(g9205),.A(g6454),.B(g8957));
  AND2 AND2_640(.VSS(VSS),.VDD(VDD),.Y(g5538),.A(g1669),.B(g4313));
  AND2 AND2_641(.VSS(VSS),.VDD(VDD),.Y(g4000),.A(g1744),.B(g2778));
  AND2 AND2_642(.VSS(VSS),.VDD(VDD),.Y(g4126),.A(g2701),.B(g3040));
  AND2 AND2_643(.VSS(VSS),.VDD(VDD),.Y(g4400),.A(g4088),.B(g3829));
  AND2 AND2_644(.VSS(VSS),.VDD(VDD),.Y(g2794),.A(I5886),.B(I5887));
  AND2 AND2_645(.VSS(VSS),.VDD(VDD),.Y(g4760),.A(g486),.B(g3393));
  AND2 AND2_646(.VSS(VSS),.VDD(VDD),.Y(g6238),.A(g572),.B(g5096));
  AND2 AND2_647(.VSS(VSS),.VDD(VDD),.Y(g10784),.A(g10727),.B(g5169));
  AND2 AND2_648(.VSS(VSS),.VDD(VDD),.Y(g8174),.A(g5284),.B(g7853));
  AND2 AND2_649(.VSS(VSS),.VDD(VDD),.Y(g6332),.A(g1374),.B(g5904));
  AND2 AND2_650(.VSS(VSS),.VDD(VDD),.Y(g5067),.A(g305),.B(g4811));
  AND2 AND2_651(.VSS(VSS),.VDD(VDD),.Y(g5418),.A(g1512),.B(g4344));
  AND2 AND2_652(.VSS(VSS),.VDD(VDD),.Y(g10297),.A(g8892),.B(g10211));
  AND2 AND2_653(.VSS(VSS),.VDD(VDD),.Y(g6353),.A(g299),.B(g5895));
  AND2 AND2_654(.VSS(VSS),.VDD(VDD),.Y(g11026),.A(g386),.B(g10974));
  AND2 AND2_655(.VSS(VSS),.VDD(VDD),.Y(g11212),.A(g944),.B(g11155));
  AND2 AND2_656(.VSS(VSS),.VDD(VDD),.Y(g6744),.A(g4828),.B(g6151));
  AND2 AND2_657(.VSS(VSS),.VDD(VDD),.Y(g5493),.A(g1923),.B(g4265));
  AND2 AND2_658(.VSS(VSS),.VDD(VDD),.Y(g10671),.A(g10578),.B(g9431));
  AND2 AND2_659(.VSS(VSS),.VDD(VDD),.Y(g4383),.A(g2517),.B(g3829));
  AND2 AND2_660(.VSS(VSS),.VDD(VDD),.Y(g5256),.A(g4297),.B(g2779));
  AND2 AND2_661(.VSS(VSS),.VDD(VDD),.Y(g4220),.A(g105),.B(g3539));
  AND2 AND2_662(.VSS(VSS),.VDD(VDD),.Y(g8380),.A(g8252),.B(g4240));
  AND2 AND2_663(.VSS(VSS),.VDD(VDD),.Y(g7071),.A(g5916),.B(g6590));
  AND2 AND2_664(.VSS(VSS),.VDD(VDD),.Y(g4779),.A(g501),.B(g3427));
  AND2 AND2_665(.VSS(VSS),.VDD(VDD),.Y(g9613),.A(g1176),.B(g9125));
  AND2 AND2_666(.VSS(VSS),.VDD(VDD),.Y(g7705),.A(g6853),.B(g4328));
  AND2 AND2_667(.VSS(VSS),.VDD(VDD),.Y(g9269),.A(g8933),.B(g3413));
  AND2 AND2_668(.VSS(VSS),.VDD(VDD),.Y(g5181),.A(g4520),.B(g4510));
  AND2 AND2_669(.VSS(VSS),.VDD(VDD),.Y(g4977),.A(g4567),.B(g4807));
  AND2 AND2_670(.VSS(VSS),.VDD(VDD),.Y(g7948),.A(g2855),.B(g7497));
  AND2 AND2_671(.VSS(VSS),.VDD(VDD),.Y(g11149),.A(g324),.B(g10930));
  AND2 AND2_672(.VSS(VSS),.VDD(VDD),.Y(g9862),.A(g1601),.B(g9777));
  AND2 AND2_673(.VSS(VSS),.VDD(VDD),.Y(g11387),.A(g11284),.B(g3629));
  AND2 AND2_674(.VSS(VSS),.VDD(VDD),.Y(g7955),.A(g2877),.B(g7516));
  AND2 AND2_675(.VSS(VSS),.VDD(VDD),.Y(g4161),.A(g2719),.B(g3060));
  AND2 AND2_676(.VSS(VSS),.VDD(VDD),.Y(g11148),.A(g2321),.B(g10913));
  AND2 AND2_677(.VSS(VSS),.VDD(VDD),.Y(g9712),.A(g1528),.B(g9490));
  AND2 AND2_678(.VSS(VSS),.VDD(VDD),.Y(g8931),.A(g8807),.B(g8164));
  AND2 AND2_679(.VSS(VSS),.VDD(VDD),.Y(g11097),.A(g378),.B(g10884));
  AND3 AND3_24(.VSS(VSS),.VDD(VDD),.Y(g5421),.A(g4631),.B(g2733),.C(g3819));
  AND2 AND2_680(.VSS(VSS),.VDD(VDD),.Y(g11104),.A(g2963),.B(g10937));
  AND2 AND2_681(.VSS(VSS),.VDD(VDD),.Y(g5263),.A(g709),.B(g4761));
  AND2 AND2_682(.VSS(VSS),.VDD(VDD),.Y(g6092),.A(g1059),.B(g5320));
  AND2 AND2_683(.VSS(VSS),.VDD(VDD),.Y(g4999),.A(g1499),.B(g4640));
  AND4 AND4_3(.VSS(VSS),.VDD(VDD),.Y(I6338),.A(g2475),.B(g2456),.C(g2451),.D(g2446));
  AND3 AND3_25(.VSS(VSS),.VDD(VDD),.Y(g7409),.A(g4976),.B(g632),.C(g6858));
  AND2 AND2_684(.VSS(VSS),.VDD(VDD),.Y(g4103),.A(g2683),.B(g2997));
  AND4 AND4_4(.VSS(VSS),.VDD(VDD),.Y(I6309),.A(g2446),.B(g2451),.C(g2456),.D(g2475));
  AND2 AND2_685(.VSS(VSS),.VDD(VDD),.Y(g6580),.A(g1801),.B(g5944));
  AND2 AND2_686(.VSS(VSS),.VDD(VDD),.Y(g5631),.A(g1056),.B(g4416));
  AND2 AND2_687(.VSS(VSS),.VDD(VDD),.Y(g9414),.A(g1730),.B(g9052));
  AND2 AND2_688(.VSS(VSS),.VDD(VDD),.Y(g9660),.A(g1188),.B(g9125));
  AND2 AND2_689(.VSS(VSS),.VDD(VDD),.Y(g9946),.A(g9926),.B(g9392));
  AND2 AND2_690(.VSS(VSS),.VDD(VDD),.Y(g5257),.A(g691),.B(g4755));
  AND2 AND2_691(.VSS(VSS),.VDD(VDD),.Y(g4732),.A(g391),.B(g3372));
  AND2 AND2_692(.VSS(VSS),.VDD(VDD),.Y(g3108),.A(I6330),.B(I6331));
  AND2 AND2_693(.VSS(VSS),.VDD(VDD),.Y(g4753),.A(g481),.B(g3386));
  AND2 AND2_694(.VSS(VSS),.VDD(VDD),.Y(g9903),.A(g9885),.B(g9673));
  AND2 AND2_695(.VSS(VSS),.VDD(VDD),.Y(g10625),.A(g10546),.B(g4552));
  AND2 AND2_696(.VSS(VSS),.VDD(VDD),.Y(g5605),.A(g4828),.B(g704));
  AND2 AND2_697(.VSS(VSS),.VDD(VDD),.Y(g6623),.A(g55),.B(g6170));
  AND2 AND2_698(.VSS(VSS),.VDD(VDD),.Y(g11228),.A(g466),.B(g11060));
  AND2 AND2_699(.VSS(VSS),.VDD(VDD),.Y(g11011),.A(g1968),.B(g10809));
  AND2 AND2_700(.VSS(VSS),.VDD(VDD),.Y(g6889),.A(g1941),.B(g6427));
  AND2 AND2_701(.VSS(VSS),.VDD(VDD),.Y(g8040),.A(g7523),.B(g5128));
  AND2 AND2_702(.VSS(VSS),.VDD(VDD),.Y(g7822),.A(g1914),.B(g7479));
  AND2 AND2_703(.VSS(VSS),.VDD(VDD),.Y(g8123),.A(g1918),.B(g7946));
  AND2 AND2_704(.VSS(VSS),.VDD(VDD),.Y(g11582),.A(g1311),.B(g11540));
  AND2 AND2_705(.VSS(VSS),.VDD(VDD),.Y(g4316),.A(g1965),.B(g3400));
  AND2 AND2_706(.VSS(VSS),.VDD(VDD),.Y(g10969),.A(g3625),.B(g10809));
  AND2 AND2_707(.VSS(VSS),.VDD(VDD),.Y(g5041),.A(g3983),.B(g4401));
  AND2 AND2_708(.VSS(VSS),.VDD(VDD),.Y(g9335),.A(g8975),.B(g5708));
  AND2 AND2_709(.VSS(VSS),.VDD(VDD),.Y(g9831),.A(g9727),.B(g9785));
  AND2 AND2_710(.VSS(VSS),.VDD(VDD),.Y(g4565),.A(g534),.B(g4010));
  AND2 AND2_711(.VSS(VSS),.VDD(VDD),.Y(g9422),.A(g1750),.B(g9030));
  AND2 AND2_712(.VSS(VSS),.VDD(VDD),.Y(g8648),.A(g4588),.B(g8511));
  AND3 AND3_26(.VSS(VSS),.VDD(VDD),.Y(g8875),.A(g8255),.B(g6368),.C(g8858));
  AND2 AND2_713(.VSS(VSS),.VDD(VDD),.Y(g5168),.A(g1512),.B(g4679));
  AND2 AND2_714(.VSS(VSS),.VDD(VDD),.Y(g7895),.A(g7503),.B(g7036));
  AND2 AND2_715(.VSS(VSS),.VDD(VDD),.Y(g8655),.A(g8532),.B(g4013));
  AND2 AND2_716(.VSS(VSS),.VDD(VDD),.Y(g3396),.A(g213),.B(g3228));
  AND2 AND2_717(.VSS(VSS),.VDD(VDD),.Y(g4914),.A(g1062),.B(g4436));
  AND2 AND2_718(.VSS(VSS),.VDD(VDD),.Y(g9947),.A(g9927),.B(g9392));
  AND2 AND2_719(.VSS(VSS),.VDD(VDD),.Y(g5772),.A(g1555),.B(g5214));
  AND2 AND2_720(.VSS(VSS),.VDD(VDD),.Y(g6838),.A(g192),.B(g6596));
  AND2 AND2_721(.VSS(VSS),.VDD(VDD),.Y(g5531),.A(g1666),.B(g4306));
  AND2 AND2_722(.VSS(VSS),.VDD(VDD),.Y(g6795),.A(g5036),.B(g5878));
  AND2 AND2_723(.VSS(VSS),.VDD(VDD),.Y(g10503),.A(g10388),.B(g2135));
  AND2 AND2_724(.VSS(VSS),.VDD(VDD),.Y(g8010),.A(g7738),.B(g7413));
  AND2 AND2_725(.VSS(VSS),.VDD(VDD),.Y(g8410),.A(g713),.B(g8143));
  AND2 AND2_726(.VSS(VSS),.VDD(VDD),.Y(g6231),.A(g818),.B(g5608));
  AND2 AND2_727(.VSS(VSS),.VDD(VDD),.Y(g10581),.A(g10531),.B(g9453));
  AND2 AND2_728(.VSS(VSS),.VDD(VDD),.Y(g10450),.A(g10364),.B(g3359));
  AND2 AND2_729(.VSS(VSS),.VDD(VDD),.Y(g2804),.A(g2132),.B(g1891));
  AND2 AND2_730(.VSS(VSS),.VDD(VDD),.Y(g3418),.A(g2379),.B(g3012));
  AND2 AND2_731(.VSS(VSS),.VDD(VDD),.Y(g4820),.A(g186),.B(g3946));
  AND2 AND2_732(.VSS(VSS),.VDD(VDD),.Y(g9653),.A(g1185),.B(g9125));
  AND2 AND2_733(.VSS(VSS),.VDD(VDD),.Y(g6205),.A(g1515),.B(g5151));
  AND2 AND2_734(.VSS(VSS),.VDD(VDD),.Y(g10818),.A(g10730),.B(g4545));
  AND2 AND2_735(.VSS(VSS),.VDD(VDD),.Y(g8172),.A(g5275),.B(g7853));
  AND2 AND2_736(.VSS(VSS),.VDD(VDD),.Y(g10496),.A(g10429),.B(g3977));
  AND2 AND2_737(.VSS(VSS),.VDD(VDD),.Y(g5074),.A(g1771),.B(g4587));
  AND2 AND2_738(.VSS(VSS),.VDD(VDD),.Y(g9869),.A(g1558),.B(g9814));
  AND2 AND2_739(.VSS(VSS),.VDD(VDD),.Y(g9719),.A(g1543),.B(g9490));
  AND2 AND2_740(.VSS(VSS),.VDD(VDD),.Y(g10741),.A(g10635),.B(g4013));
  AND2 AND2_741(.VSS(VSS),.VDD(VDD),.Y(g3381),.A(g940),.B(g2756));
  AND2 AND2_742(.VSS(VSS),.VDD(VDD),.Y(g5863),.A(g5272),.B(g2173));
  AND2 AND2_743(.VSS(VSS),.VDD(VDD),.Y(g8693),.A(g3738),.B(g8509));
  AND2 AND2_744(.VSS(VSS),.VDD(VDD),.Y(g5480),.A(g4279),.B(g3519));
  AND2 AND2_745(.VSS(VSS),.VDD(VDD),.Y(g4581),.A(g3766),.B(g3254));
  AND2 AND2_746(.VSS(VSS),.VDD(VDD),.Y(g3685),.A(g1781),.B(g2981));
  AND2 AND2_747(.VSS(VSS),.VDD(VDD),.Y(g5569),.A(g4816),.B(g2338));
  AND2 AND2_748(.VSS(VSS),.VDD(VDD),.Y(g8555),.A(g8409),.B(g8025));
  AND2 AND2_749(.VSS(VSS),.VDD(VDD),.Y(g3263),.A(g2503),.B(g2328));
  AND2 AND2_750(.VSS(VSS),.VDD(VDD),.Y(g9364),.A(g965),.B(g9223));
  AND2 AND2_751(.VSS(VSS),.VDD(VDD),.Y(g4784),.A(g506),.B(g3432));
  AND2 AND2_752(.VSS(VSS),.VDD(VDD),.Y(g9454),.A(g8994),.B(g5708));
  AND4 AND4_5(.VSS(VSS),.VDD(VDD),.Y(I6331),.A(g2060),.B(g2070),.C(g2074),.D(g2077));
  AND2 AND2_753(.VSS(VSS),.VDD(VDD),.Y(g11299),.A(g5498),.B(g11243));
  AND2 AND2_754(.VSS(VSS),.VDD(VDD),.Y(g6983),.A(g6592),.B(g3105));
  AND2 AND2_755(.VSS(VSS),.VDD(VDD),.Y(g7958),.A(g736),.B(g7697));
  AND2 AND2_756(.VSS(VSS),.VDD(VDD),.Y(g4995),.A(g1474),.B(g4640));
  AND2 AND2_757(.VSS(VSS),.VDD(VDD),.Y(g4079),.A(g2765),.B(g2276));
  AND2 AND2_758(.VSS(VSS),.VDD(VDD),.Y(g2264),.A(g1771),.B(g1766));
  AND2 AND2_759(.VSS(VSS),.VDD(VDD),.Y(g2160),.A(g745),.B(g746));
  AND2 AND2_760(.VSS(VSS),.VDD(VDD),.Y(g3257),.A(g378),.B(g2496));
  AND2 AND2_761(.VSS(VSS),.VDD(VDD),.Y(g3101),.A(I6309),.B(I6310));
  AND2 AND2_762(.VSS(VSS),.VDD(VDD),.Y(g5000),.A(g1470),.B(g4640));
  AND2 AND2_763(.VSS(VSS),.VDD(VDD),.Y(g3301),.A(g1346),.B(g2544));
  AND2 AND2_764(.VSS(VSS),.VDD(VDD),.Y(g5126),.A(g3076),.B(g4638));
  AND4 AND4_6(.VSS(VSS),.VDD(VDD),.Y(I5084),.A(g1462),.B(g1470),.C(g1474),.D(g1478));
  AND2 AND2_765(.VSS(VSS),.VDD(VDD),.Y(g9412),.A(g1727),.B(g9052));
  AND2 AND2_766(.VSS(VSS),.VDD(VDD),.Y(g9389),.A(g1330),.B(g9151));
  AND2 AND2_767(.VSS(VSS),.VDD(VDD),.Y(g2379),.A(g744),.B(g743));
  AND2 AND2_768(.VSS(VSS),.VDD(VDD),.Y(g10706),.A(g10567),.B(g4840));
  AND3 AND3_27(.VSS(VSS),.VDD(VDD),.Y(I16145),.A(g10366),.B(g10447),.C(g10446));
  AND2 AND2_769(.VSS(VSS),.VDD(VDD),.Y(g10597),.A(g10533),.B(g4359));
  AND3 AND3_28(.VSS(VSS),.VDD(VDD),.Y(g8965),.A(g8110),.B(g6778),.C(g8849));
  AND2 AND2_770(.VSS(VSS),.VDD(VDD),.Y(g5608),.A(g814),.B(g4831));
  AND2 AND2_771(.VSS(VSS),.VDD(VDD),.Y(g5220),.A(g1083),.B(g4729));
  AND2 AND2_772(.VSS(VSS),.VDD(VDD),.Y(g10624),.A(g10545),.B(g4544));
  AND2 AND2_773(.VSS(VSS),.VDD(VDD),.Y(g10300),.A(g8892),.B(g10220));
  AND2 AND2_774(.VSS(VSS),.VDD(VDD),.Y(g5023),.A(g1071),.B(g4511));
  AND2 AND2_775(.VSS(VSS),.VDD(VDD),.Y(g4432),.A(g3723),.B(g1975));
  AND2 AND2_776(.VSS(VSS),.VDD(VDD),.Y(g4053),.A(g2701),.B(g2276));
  AND2 AND2_777(.VSS(VSS),.VDD(VDD),.Y(g8050),.A(g7596),.B(g5919));
  AND2 AND2_778(.VSS(VSS),.VDD(VDD),.Y(g5588),.A(g1639),.B(g4508));
  AND3 AND3_29(.VSS(VSS),.VDD(VDD),.Y(g6679),.A(g4631),.B(g6074),.C(g2733));
  AND2 AND2_779(.VSS(VSS),.VDD(VDD),.Y(g9963),.A(g9953),.B(g9536));
  AND2 AND2_780(.VSS(VSS),.VDD(VDD),.Y(g3772),.A(g2542),.B(g3089));
  AND2 AND2_781(.VSS(VSS),.VDD(VDD),.Y(g5051),.A(g4432),.B(g2834));
  AND2 AND2_782(.VSS(VSS),.VDD(VDD),.Y(g6831),.A(g207),.B(g6596));
  AND2 AND2_783(.VSS(VSS),.VDD(VDD),.Y(g2981),.A(g1776),.B(g2264));
  AND2 AND2_784(.VSS(VSS),.VDD(VDD),.Y(g8724),.A(g8606),.B(g7910));
  AND2 AND2_785(.VSS(VSS),.VDD(VDD),.Y(g4157),.A(g2713),.B(g3055));
  AND2 AND2_786(.VSS(VSS),.VDD(VDD),.Y(g9707),.A(g1583),.B(g9474));
  AND3 AND3_30(.VSS(VSS),.VDD(VDD),.Y(g8878),.A(g8099),.B(g6368),.C(g8858));
  AND2 AND2_787(.VSS(VSS),.VDD(VDD),.Y(g2132),.A(g1872),.B(g1882));
  AND2 AND2_788(.VSS(VSS),.VDD(VDD),.Y(g10763),.A(g10639),.B(g4840));
  AND3 AND3_31(.VSS(VSS),.VDD(VDD),.Y(g8289),.A(g6777),.B(g8109),.C(g6475));
  AND2 AND2_789(.VSS(VSS),.VDD(VDD),.Y(g7898),.A(g7511),.B(g7041));
  AND2 AND2_790(.VSS(VSS),.VDD(VDD),.Y(g11271),.A(g5624),.B(g11191));
  AND2 AND2_791(.VSS(VSS),.VDD(VDD),.Y(g11461),.A(g11429),.B(g5446));
  AND2 AND2_792(.VSS(VSS),.VDD(VDD),.Y(g5732),.A(g1604),.B(g5176));
  AND2 AND2_793(.VSS(VSS),.VDD(VDD),.Y(g11145),.A(g315),.B(g10927));
  AND2 AND2_794(.VSS(VSS),.VDD(VDD),.Y(g11031),.A(g411),.B(g10974));
  AND2 AND2_795(.VSS(VSS),.VDD(VDD),.Y(g9865),.A(g1607),.B(g9780));
  AND2 AND2_796(.VSS(VSS),.VDD(VDD),.Y(g5944),.A(g1796),.B(g5233));
  AND2 AND2_797(.VSS(VSS),.VDD(VDD),.Y(g9715),.A(g1531),.B(g9490));
  AND2 AND2_798(.VSS(VSS),.VDD(VDD),.Y(g9604),.A(g1194),.B(g9111));
  AND2 AND2_799(.VSS(VSS),.VDD(VDD),.Y(g8799),.A(g8647),.B(g8727));
  AND2 AND2_800(.VSS(VSS),.VDD(VDD),.Y(g11198),.A(g4919),.B(g11069));
  AND2 AND2_801(.VSS(VSS),.VDD(VDD),.Y(g6873),.A(g3263),.B(g6557));
  AND2 AND2_802(.VSS(VSS),.VDD(VDD),.Y(g6632),.A(g61),.B(g6190));
  AND2 AND2_803(.VSS(VSS),.VDD(VDD),.Y(g6095),.A(g1062),.B(g5320));
  AND2 AND2_804(.VSS(VSS),.VDD(VDD),.Y(g3863),.A(g3323),.B(g2728));
  AND2 AND2_805(.VSS(VSS),.VDD(VDD),.Y(g9833),.A(g9729),.B(g9785));
  AND2 AND2_806(.VSS(VSS),.VDD(VDD),.Y(g6653),.A(g70),.B(g6213));
  AND2 AND2_807(.VSS(VSS),.VDD(VDD),.Y(g6102),.A(g1038),.B(g5320));
  AND2 AND2_808(.VSS(VSS),.VDD(VDD),.Y(g7819),.A(g1887),.B(g7479));
  AND2 AND2_809(.VSS(VSS),.VDD(VDD),.Y(g11393),.A(g11280),.B(g7916));
  AND2 AND2_810(.VSS(VSS),.VDD(VDD),.Y(g2511),.A(g461),.B(g456));
  AND2 AND2_811(.VSS(VSS),.VDD(VDD),.Y(g7088),.A(g2331),.B(g6737));
  AND2 AND2_812(.VSS(VSS),.VDD(VDD),.Y(g9584),.A(g2726),.B(g9173));
  AND2 AND2_813(.VSS(VSS),.VDD(VDD),.Y(g9896),.A(g9883),.B(g9624));
  AND3 AND3_32(.VSS(VSS),.VDD(VDD),.Y(g8209),.A(g4094),.B(g3792),.C(g7980));
  AND2 AND2_814(.VSS(VSS),.VDD(VDD),.Y(g6752),.A(g6187),.B(g2343));
  AND2 AND2_815(.VSS(VSS),.VDD(VDD),.Y(g4778),.A(g421),.B(g3426));
  AND2 AND2_816(.VSS(VSS),.VDD(VDD),.Y(g11161),.A(g1969),.B(g10937));
  AND2 AND2_817(.VSS(VSS),.VDD(VDD),.Y(g9268),.A(g6681),.B(g8947));
  AND2 AND2_818(.VSS(VSS),.VDD(VDD),.Y(g5681),.A(g135),.B(g5361));
  AND2 AND2_819(.VSS(VSS),.VDD(VDD),.Y(g7951),.A(g2868),.B(g7505));
  AND2 AND2_820(.VSS(VSS),.VDD(VDD),.Y(g9419),.A(g1744),.B(g9030));
  AND2 AND2_821(.VSS(VSS),.VDD(VDD),.Y(g10268),.A(g10183),.B(g3307));
  AND2 AND2_822(.VSS(VSS),.VDD(VDD),.Y(g5533),.A(g1724),.B(g4308));
  AND2 AND2_823(.VSS(VSS),.VDD(VDD),.Y(g9052),.A(g8936),.B(g7192));
  AND2 AND2_824(.VSS(VSS),.VDD(VDD),.Y(g6786),.A(g178),.B(g5919));
  AND2 AND2_825(.VSS(VSS),.VDD(VDD),.Y(g10670),.A(g10571),.B(g9091));
  AND2 AND2_826(.VSS(VSS),.VDD(VDD),.Y(g11087),.A(g829),.B(g10950));
  AND2 AND2_827(.VSS(VSS),.VDD(VDD),.Y(g4949),.A(g3505),.B(g4449));
  AND2 AND2_828(.VSS(VSS),.VDD(VDD),.Y(g6364),.A(g5851),.B(g4454));
  AND2 AND2_829(.VSS(VSS),.VDD(VDD),.Y(g7825),.A(g1941),.B(g7479));
  AND2 AND2_830(.VSS(VSS),.VDD(VDD),.Y(g3400),.A(g115),.B(g3164));
  AND2 AND2_831(.VSS(VSS),.VDD(VDD),.Y(g4998),.A(g1304),.B(g4485));
  AND2 AND2_832(.VSS(VSS),.VDD(VDD),.Y(g10667),.A(g10576),.B(g9427));
  AND2 AND2_833(.VSS(VSS),.VDD(VDD),.Y(g7136),.A(g6050),.B(g6704));
  AND2 AND2_834(.VSS(VSS),.VDD(VDD),.Y(g6532),.A(g339),.B(g6057));
  AND2 AND2_835(.VSS(VSS),.VDD(VDD),.Y(g9385),.A(g1324),.B(g9151));
  AND4 AND4_7(.VSS(VSS),.VDD(VDD),.Y(I5690),.A(g1436),.B(g1440),.C(g1444),.D(g1448));
  AND2 AND2_836(.VSS(VSS),.VDD(VDD),.Y(g4484),.A(g1137),.B(g3909));
  AND2 AND2_837(.VSS(VSS),.VDD(VDD),.Y(g9897),.A(g9884),.B(g9624));
  AND2 AND2_838(.VSS(VSS),.VDD(VDD),.Y(g9425),.A(g1753),.B(g9030));
  AND2 AND2_839(.VSS(VSS),.VDD(VDD),.Y(g3383),.A(g186),.B(g3228));
  AND2 AND2_840(.VSS(VSS),.VDD(VDD),.Y(g5601),.A(g1035),.B(g4375));
  AND2 AND2_841(.VSS(VSS),.VDD(VDD),.Y(g7943),.A(g2840),.B(g7467));
  AND2 AND2_842(.VSS(VSS),.VDD(VDD),.Y(g11171),.A(g481),.B(g11112));
  AND2 AND2_843(.VSS(VSS),.VDD(VDD),.Y(g3423),.A(I6630),.B(I6631));
  AND2 AND2_844(.VSS(VSS),.VDD(VDD),.Y(g7230),.A(g6064),.B(g6444));
  AND2 AND2_845(.VSS(VSS),.VDD(VDD),.Y(g4952),.A(g1648),.B(g4457));
  AND2 AND2_846(.VSS(VSS),.VDD(VDD),.Y(g8736),.A(g7439),.B(g8635));
  AND2 AND2_847(.VSS(VSS),.VDD(VDD),.Y(g6787),.A(g266),.B(g5875));
  AND3 AND3_33(.VSS(VSS),.VDD(VDD),.Y(g8968),.A(g8089),.B(g6778),.C(g8849));
  AND2 AND2_848(.VSS(VSS),.VDD(VDD),.Y(g10306),.A(g10214),.B(g9082));
  AND2 AND2_849(.VSS(VSS),.VDD(VDD),.Y(g9331),.A(g8972),.B(g5708));
  AND2 AND2_850(.VSS(VSS),.VDD(VDD),.Y(g11459),.A(g11427),.B(g5446));
  AND2 AND2_851(.VSS(VSS),.VDD(VDD),.Y(g4561),.A(g538),.B(g4003));
  AND2 AND2_852(.VSS(VSS),.VDD(VDD),.Y(g11425),.A(g11350),.B(g10899));
  AND2 AND2_853(.VSS(VSS),.VDD(VDD),.Y(g11458),.A(g11426),.B(g5446));
  AND2 AND2_854(.VSS(VSS),.VDD(VDD),.Y(g5739),.A(g1607),.B(g5185));
  AND2 AND2_855(.VSS(VSS),.VDD(VDD),.Y(g7496),.A(g7148),.B(g2840));
  AND2 AND2_856(.VSS(VSS),.VDD(VDD),.Y(g4986),.A(g1411),.B(g4682));
  AND2 AND2_857(.VSS(VSS),.VDD(VDD),.Y(g11010),.A(g5187),.B(g10827));
  AND2 AND2_858(.VSS(VSS),.VDD(VDD),.Y(g3999),.A(g1741),.B(g2777));
  AND2 AND2_859(.VSS(VSS),.VDD(VDD),.Y(g8175),.A(g5291),.B(g7853));
  AND2 AND2_860(.VSS(VSS),.VDD(VDD),.Y(g8722),.A(g8604),.B(g7908));
  AND2 AND2_861(.VSS(VSS),.VDD(VDD),.Y(g4764),.A(g411),.B(g3404));
  AND2 AND2_862(.VSS(VSS),.VDD(VDD),.Y(g7137),.A(g5590),.B(g6361));
  AND2 AND2_863(.VSS(VSS),.VDD(VDD),.Y(g7891),.A(g7471),.B(g7028));
  AND2 AND2_864(.VSS(VSS),.VDD(VDD),.Y(g8651),.A(g8520),.B(g4013));
  AND2 AND2_865(.VSS(VSS),.VDD(VDD),.Y(g5479),.A(g1845),.B(g4243));
  AND2 AND2_866(.VSS(VSS),.VDD(VDD),.Y(g11599),.A(g1341),.B(g11572));
  AND2 AND2_867(.VSS(VSS),.VDD(VDD),.Y(g6684),.A(g5314),.B(g5836));
  AND2 AND2_868(.VSS(VSS),.VDD(VDD),.Y(g6745),.A(g5605),.B(g6158));
  AND2 AND2_869(.VSS(VSS),.VDD(VDD),.Y(g6639),.A(g357),.B(g6196));
  AND2 AND2_870(.VSS(VSS),.VDD(VDD),.Y(g10937),.A(g4822),.B(g10822));
  AND2 AND2_871(.VSS(VSS),.VDD(VDD),.Y(g3696),.A(g1713),.B(g3015));
  AND2 AND2_872(.VSS(VSS),.VDD(VDD),.Y(g4503),.A(g654),.B(g3943));
  AND2 AND2_873(.VSS(VSS),.VDD(VDD),.Y(g6791),.A(g269),.B(g5880));
  AND2 AND2_874(.VSS(VSS),.VDD(VDD),.Y(g5190),.A(g1245),.B(g4716));
  AND2 AND2_875(.VSS(VSS),.VDD(VDD),.Y(g5390),.A(g3220),.B(g4819));
  AND2 AND2_876(.VSS(VSS),.VDD(VDD),.Y(g8384),.A(g8180),.B(g3397));
  AND2 AND2_877(.VSS(VSS),.VDD(VDD),.Y(g4224),.A(g1092),.B(g3638));
  AND2 AND2_878(.VSS(VSS),.VDD(VDD),.Y(g5501),.A(g1672),.B(g4273));
  AND2 AND2_879(.VSS(VSS),.VDD(VDD),.Y(g9173),.A(g8968),.B(g6674));
  AND2 AND2_880(.VSS(VSS),.VDD(VDD),.Y(g6759),.A(g148),.B(g5919));
  AND2 AND2_881(.VSS(VSS),.VDD(VDD),.Y(g8838),.A(g8602),.B(g8702));
  AND2 AND2_882(.VSS(VSS),.VDD(VDD),.Y(g8024),.A(g7394),.B(g4337));
  AND2 AND2_883(.VSS(VSS),.VDD(VDD),.Y(g10666),.A(g10575),.B(g9424));
  AND2 AND2_884(.VSS(VSS),.VDD(VDD),.Y(g11158),.A(g309),.B(g10935));
  AND2 AND2_885(.VSS(VSS),.VDD(VDD),.Y(g9602),.A(g2650),.B(g9010));
  AND2 AND2_886(.VSS(VSS),.VDD(VDD),.Y(g5704),.A(g143),.B(g5361));
  AND2 AND2_887(.VSS(VSS),.VDD(VDD),.Y(g4617),.A(g3275),.B(g3879));
  AND2 AND2_888(.VSS(VSS),.VDD(VDD),.Y(g11561),.A(g11518),.B(g3015));
  AND2 AND2_889(.VSS(VSS),.VDD(VDD),.Y(g9868),.A(g1555),.B(g9812));
  AND2 AND2_890(.VSS(VSS),.VDD(VDD),.Y(g11295),.A(g5475),.B(g11239));
  AND2 AND2_891(.VSS(VSS),.VDD(VDD),.Y(g11144),.A(g305),.B(g10926));
  AND2 AND2_892(.VSS(VSS),.VDD(VDD),.Y(g9718),.A(g1540),.B(g9490));
  AND2 AND2_893(.VSS(VSS),.VDD(VDD),.Y(g3434),.A(g237),.B(g3228));
  AND2 AND2_894(.VSS(VSS),.VDD(VDD),.Y(g4987),.A(g1440),.B(g4682));
  AND2 AND2_895(.VSS(VSS),.VDD(VDD),.Y(g4771),.A(g496),.B(g3416));
  AND2 AND2_896(.VSS(VSS),.VDD(VDD),.Y(g5250),.A(g1270),.B(g4748));
  AND2 AND2_897(.VSS(VSS),.VDD(VDD),.Y(g6098),.A(g1065),.B(g5320));
  AND2 AND2_898(.VSS(VSS),.VDD(VDD),.Y(g9582),.A(g2725),.B(g9173));
  AND2 AND2_899(.VSS(VSS),.VDD(VDD),.Y(g6833),.A(g186),.B(g6596));
  AND2 AND2_900(.VSS(VSS),.VDD(VDD),.Y(g3533),.A(g1981),.B(g2892));
  AND2 AND2_901(.VSS(VSS),.VDD(VDD),.Y(g4892),.A(g632),.B(g4739));
  AND2 AND2_902(.VSS(VSS),.VDD(VDD),.Y(g8104),.A(g6218),.B(g7880));
  AND2 AND2_903(.VSS(VSS),.VDD(VDD),.Y(g9415),.A(g1733),.B(g9052));
  AND2 AND2_904(.VSS(VSS),.VDD(VDD),.Y(g8499),.A(g8377),.B(g4737));
  AND2 AND2_905(.VSS(VSS),.VDD(VDD),.Y(g9664),.A(g1191),.B(g9125));
  AND2 AND2_906(.VSS(VSS),.VDD(VDD),.Y(g10740),.A(g10676),.B(g3384));
  AND2 AND2_907(.VSS(VSS),.VDD(VDD),.Y(g2534),.A(g798),.B(g794));
  AND2 AND2_908(.VSS(VSS),.VDD(VDD),.Y(g8754),.A(g7420),.B(g8667));
  AND2 AND2_909(.VSS(VSS),.VDD(VDD),.Y(g9721),.A(g9413),.B(g4785));
  AND2 AND2_910(.VSS(VSS),.VDD(VDD),.Y(g6162),.A(g3584),.B(g5200));
  AND2 AND2_911(.VSS(VSS),.VDD(VDD),.Y(g4991),.A(g1508),.B(g4640));
  AND2 AND2_912(.VSS(VSS),.VDD(VDD),.Y(g6362),.A(g5846),.B(g4450));
  AND4 AND4_8(.VSS(VSS),.VDD(VDD),.Y(I6631),.A(g2707),.B(g2713),.C(g2719),.D(g2765));
  AND2 AND2_913(.VSS(VSS),.VDD(VDD),.Y(g10685),.A(g10608),.B(g3863));
  AND2 AND2_914(.VSS(VSS),.VDD(VDD),.Y(g4340),.A(g1153),.B(g3715));
  AND2 AND2_915(.VSS(VSS),.VDD(VDD),.Y(g11023),.A(g440),.B(g10974));
  AND2 AND2_916(.VSS(VSS),.VDD(VDD),.Y(g8044),.A(g7598),.B(g5919));
  AND2 AND2_917(.VSS(VSS),.VDD(VDD),.Y(g11224),.A(g968),.B(g11056));
  AND2 AND2_918(.VSS(VSS),.VDD(VDD),.Y(g11571),.A(g2018),.B(g11561));
  AND2 AND2_919(.VSS(VSS),.VDD(VDD),.Y(g4959),.A(g1520),.B(g4682));
  AND2 AND2_920(.VSS(VSS),.VDD(VDD),.Y(g10334),.A(g10265),.B(g3307));
  AND2 AND2_921(.VSS(VSS),.VDD(VDD),.Y(g5626),.A(g1633),.B(g4557));
  AND2 AND2_922(.VSS(VSS),.VDD(VDD),.Y(g9940),.A(g9920),.B(g9367));
  AND2 AND2_923(.VSS(VSS),.VDD(VDD),.Y(g4876),.A(g1086),.B(g3638));
  AND2 AND2_924(.VSS(VSS),.VDD(VDD),.Y(g6728),.A(g6250),.B(g4318));
  AND2 AND2_925(.VSS(VSS),.VDD(VDD),.Y(g6730),.A(g1872),.B(g6128));
  AND2 AND2_926(.VSS(VSS),.VDD(VDD),.Y(g9689),.A(g263),.B(g9432));
  AND2 AND2_927(.VSS(VSS),.VDD(VDD),.Y(g10762),.A(g10635),.B(g4840));
  AND2 AND2_928(.VSS(VSS),.VDD(VDD),.Y(g6070),.A(g1050),.B(g5320));
  AND2 AND2_929(.VSS(VSS),.VDD(VDD),.Y(g9428),.A(g1756),.B(g9030));
  AND2 AND2_930(.VSS(VSS),.VDD(VDD),.Y(g9030),.A(g8935),.B(g7192));
  AND2 AND2_931(.VSS(VSS),.VDD(VDD),.Y(g9430),.A(g1759),.B(g9030));
  AND2 AND2_932(.VSS(VSS),.VDD(VDD),.Y(g8927),.A(g7872),.B(g8807));
  AND2 AND2_933(.VSS(VSS),.VDD(VDD),.Y(g7068),.A(g5912),.B(g6586));
  AND2 AND2_934(.VSS(VSS),.VDD(VDD),.Y(g8014),.A(g7740),.B(g7419));
  AND2 AND2_935(.VSS(VSS),.VDD(VDD),.Y(g11392),.A(g11278),.B(g7914));
  AND2 AND2_936(.VSS(VSS),.VDD(VDD),.Y(g5782),.A(g1558),.B(g5223));
  AND2 AND2_937(.VSS(VSS),.VDD(VDD),.Y(g9910),.A(g9892),.B(g9809));
  AND2 AND2_938(.VSS(VSS),.VDD(VDD),.Y(g4824),.A(g774),.B(g4099));
  AND2 AND2_939(.VSS(VSS),.VDD(VDD),.Y(g6331),.A(g201),.B(g5904));
  AND2 AND2_940(.VSS(VSS),.VDD(VDD),.Y(g4236),.A(g1098),.B(g3638));
  AND2 AND2_941(.VSS(VSS),.VDD(VDD),.Y(g11559),.A(g2719),.B(g11519));
  AND2 AND2_942(.VSS(VSS),.VDD(VDD),.Y(g9609),.A(g907),.B(g9205));
  AND2 AND2_943(.VSS(VSS),.VDD(VDD),.Y(g11558),.A(g2713),.B(g11519));
  AND2 AND2_944(.VSS(VSS),.VDD(VDD),.Y(g6087),.A(g1056),.B(g5320));
  AND2 AND2_945(.VSS(VSS),.VDD(VDD),.Y(g4877),.A(g243),.B(g3946));
  AND2 AND2_946(.VSS(VSS),.VDD(VDD),.Y(g5526),.A(g1950),.B(g4294));
  AND2 AND2_947(.VSS(VSS),.VDD(VDD),.Y(g10751),.A(g10646),.B(g4013));
  AND2 AND2_948(.VSS(VSS),.VDD(VDD),.Y(g10772),.A(g10655),.B(g4840));
  AND2 AND2_949(.VSS(VSS),.VDD(VDD),.Y(g8135),.A(g1945),.B(g7956));
  AND2 AND2_950(.VSS(VSS),.VDD(VDD),.Y(g11544),.A(g11515),.B(g10584));
  AND2 AND2_951(.VSS(VSS),.VDD(VDD),.Y(g5084),.A(g1776),.B(g4591));
  AND2 AND2_952(.VSS(VSS),.VDD(VDD),.Y(g8382),.A(g6077),.B(g8213));
  AND2 AND2_953(.VSS(VSS),.VDD(VDD),.Y(g10230),.A(g8892),.B(g10145));
  AND2 AND2_954(.VSS(VSS),.VDD(VDD),.Y(g5484),.A(g1896),.B(g4256));
  AND2 AND2_955(.VSS(VSS),.VDD(VDD),.Y(g7241),.A(g6772),.B(g6172));
  AND2 AND2_956(.VSS(VSS),.VDD(VDD),.Y(g3942),.A(g219),.B(g3164));
  AND2 AND2_957(.VSS(VSS),.VDD(VDD),.Y(g10638),.A(g10608),.B(g3829));
  AND2 AND2_958(.VSS(VSS),.VDD(VDD),.Y(g4064),.A(g1759),.B(g2799));
  AND2 AND2_959(.VSS(VSS),.VDD(VDD),.Y(g9365),.A(g1321),.B(g9151));
  AND2 AND2_960(.VSS(VSS),.VDD(VDD),.Y(g9861),.A(g9738),.B(g9579));
  AND2 AND2_961(.VSS(VSS),.VDD(VDD),.Y(g8749),.A(g7604),.B(g8660));
  AND2 AND2_962(.VSS(VSS),.VDD(VDD),.Y(g11255),.A(g456),.B(g11075));
  AND2 AND2_963(.VSS(VSS),.VDD(VDD),.Y(g11189),.A(g5616),.B(g11064));
  AND2 AND2_964(.VSS(VSS),.VDD(VDD),.Y(g10510),.A(g10393),.B(g2135));
  AND3 AND3_34(.VSS(VSS),.VDD(VDD),.Y(g8947),.A(g8056),.B(g6368),.C(g8828));
  AND2 AND2_965(.VSS(VSS),.VDD(VDD),.Y(g2917),.A(g2424),.B(g1657));
  AND2 AND2_966(.VSS(VSS),.VDD(VDD),.Y(g5919),.A(g5216),.B(g2965));
  AND2 AND2_967(.VSS(VSS),.VDD(VDD),.Y(g11188),.A(g5604),.B(g11063));
  AND2 AND2_968(.VSS(VSS),.VDD(VDD),.Y(g9846),.A(g287),.B(g9764));
  AND2 AND2_969(.VSS(VSS),.VDD(VDD),.Y(g7818),.A(g1878),.B(g7479));
  AND2 AND2_970(.VSS(VSS),.VDD(VDD),.Y(g11460),.A(g11428),.B(g5446));
  AND2 AND2_971(.VSS(VSS),.VDD(VDD),.Y(g5276),.A(g736),.B(g4780));
  AND2 AND2_972(.VSS(VSS),.VDD(VDD),.Y(g11030),.A(g406),.B(g10974));
  AND2 AND2_973(.VSS(VSS),.VDD(VDD),.Y(g11093),.A(g841),.B(g10950));
  AND2 AND2_974(.VSS(VSS),.VDD(VDD),.Y(g7893),.A(g7478),.B(g7031));
  AND2 AND2_975(.VSS(VSS),.VDD(VDD),.Y(g8653),.A(g8526),.B(g4013));
  AND2 AND2_976(.VSS(VSS),.VDD(VDD),.Y(g10442),.A(g10311),.B(g2135));
  AND2 AND2_977(.VSS(VSS),.VDD(VDD),.Y(g6535),.A(g345),.B(g6063));
  AND2 AND2_978(.VSS(VSS),.VDD(VDD),.Y(g8102),.A(g6209),.B(g7878));
  AND4 AND4_9(.VSS(VSS),.VDD(VDD),.Y(I5085),.A(g1490),.B(g1494),.C(g1504),.D(g1508));
  AND2 AND2_979(.VSS(VSS),.VDD(VDD),.Y(g5004),.A(g1296),.B(g4499));
  AND2 AND2_980(.VSS(VSS),.VDD(VDD),.Y(g3912),.A(g207),.B(g3164));
  AND2 AND2_981(.VSS(VSS),.VDD(VDD),.Y(g7186),.A(g2503),.B(g6403));
  AND2 AND2_982(.VSS(VSS),.VDD(VDD),.Y(g4489),.A(g348),.B(g3586));
  AND2 AND2_983(.VSS(VSS),.VDD(VDD),.Y(g9662),.A(g2094),.B(g9292));
  AND2 AND2_984(.VSS(VSS),.VDD(VDD),.Y(g9418),.A(g1741),.B(g9052));
  AND2 AND2_985(.VSS(VSS),.VDD(VDD),.Y(g11218),.A(g959),.B(g11053));
  AND2 AND2_986(.VSS(VSS),.VDD(VDD),.Y(g4471),.A(g1121),.B(g3862));
  AND2 AND2_987(.VSS(VSS),.VDD(VDD),.Y(g10746),.A(g10643),.B(g4013));
  AND2 AND2_988(.VSS(VSS),.VDD(VDD),.Y(g7125),.A(g1212),.B(g6648));
  AND2 AND2_989(.VSS(VSS),.VDD(VDD),.Y(g7821),.A(g1905),.B(g7479));
  AND2 AND2_990(.VSS(VSS),.VDD(VDD),.Y(g6246),.A(g178),.B(g5361));
  AND2 AND2_991(.VSS(VSS),.VDD(VDD),.Y(g9256),.A(g6689),.B(g8963));
  AND2 AND2_992(.VSS(VSS),.VDD(VDD),.Y(g8042),.A(g7533),.B(g5128));
  AND2 AND2_993(.VSS(VSS),.VDD(VDD),.Y(g10237),.A(g10145),.B(g9100));
  AND2 AND2_994(.VSS(VSS),.VDD(VDD),.Y(g7939),.A(g2829),.B(g7460));
  AND2 AND2_995(.VSS(VSS),.VDD(VDD),.Y(g8786),.A(g8638),.B(g8716));
  AND2 AND2_996(.VSS(VSS),.VDD(VDD),.Y(g10684),.A(g10604),.B(g3863));
  AND2 AND2_997(.VSS(VSS),.VDD(VDD),.Y(g11455),.A(g11435),.B(g5446));
  AND2 AND2_998(.VSS(VSS),.VDD(VDD),.Y(g8364),.A(g658),.B(g8235));
  AND3 AND3_35(.VSS(VSS),.VDD(VDD),.Y(g2990),.A(g2061),.B(g2557),.C(g1814));
  AND2 AND2_999(.VSS(VSS),.VDD(VDD),.Y(g9847),.A(g290),.B(g9766));
  AND2 AND2_1000(.VSS(VSS),.VDD(VDD),.Y(g8054),.A(g7584),.B(g5919));
  AND2 AND2_1001(.VSS(VSS),.VDD(VDD),.Y(g5617),.A(g1050),.B(g4391));
  AND2 AND2_1002(.VSS(VSS),.VDD(VDD),.Y(g6502),.A(g5981),.B(g3095));
  AND2 AND2_1003(.VSS(VSS),.VDD(VDD),.Y(g5789),.A(g1561),.B(g5232));
  AND2 AND2_1004(.VSS(VSS),.VDD(VDD),.Y(g4009),.A(g1747),.B(g2789));
  AND2 AND2_1005(.VSS(VSS),.VDD(VDD),.Y(g11277),.A(g4920),.B(g11199));
  AND2 AND2_1006(.VSS(VSS),.VDD(VDD),.Y(g6940),.A(g6472),.B(g1945));
  AND2 AND2_1007(.VSS(VSS),.VDD(VDD),.Y(g7061),.A(g790),.B(g6760));
  AND2 AND2_1008(.VSS(VSS),.VDD(VDD),.Y(g11595),.A(g1336),.B(g11575));
  AND2 AND2_1009(.VSS(VSS),.VDD(VDD),.Y(g5771),.A(g1534),.B(g5213));
  AND2 AND2_1010(.VSS(VSS),.VDD(VDD),.Y(g8553),.A(g8405),.B(g8015));
  AND2 AND2_1011(.VSS(VSS),.VDD(VDD),.Y(g4836),.A(g643),.B(g3520));
  AND2 AND2_1012(.VSS(VSS),.VDD(VDD),.Y(g5547),.A(g1733),.B(g4326));
  AND2 AND2_1013(.VSS(VSS),.VDD(VDD),.Y(g6216),.A(g2232),.B(g5151));
  AND2 AND2_1014(.VSS(VSS),.VDD(VDD),.Y(g4967),.A(g1515),.B(g4682));
  AND2 AND2_1015(.VSS(VSS),.VDD(VDD),.Y(g6671),.A(g342),.B(g6227));
  AND2 AND2_1016(.VSS(VSS),.VDD(VDD),.Y(g7200),.A(g3098),.B(g6418));
  AND2 AND2_1017(.VSS(VSS),.VDD(VDD),.Y(g3661),.A(g382),.B(g3257));
  AND2 AND2_1018(.VSS(VSS),.VDD(VDD),.Y(g7046),.A(g5892),.B(g6570));
  AND2 AND2_1019(.VSS(VSS),.VDD(VDD),.Y(g4229),.A(g999),.B(g3914));
  AND2 AND2_1020(.VSS(VSS),.VDD(VDD),.Y(g8389),.A(g6091),.B(g8225));
  AND2 AND2_1021(.VSS(VSS),.VDD(VDD),.Y(g6430),.A(g5044),.B(g5791));
  AND2 AND2_1022(.VSS(VSS),.VDD(VDD),.Y(g8706),.A(g7602),.B(g8589));
  AND2 AND2_1023(.VSS(VSS),.VDD(VDD),.Y(g4993),.A(g1448),.B(g4682));
  AND2 AND2_1024(.VSS(VSS),.VDD(VDD),.Y(g6247),.A(g127),.B(g5361));
  AND2 AND2_1025(.VSS(VSS),.VDD(VDD),.Y(g9257),.A(g6689),.B(g8964));
  AND2 AND2_1026(.VSS(VSS),.VDD(VDD),.Y(g11170),.A(g525),.B(g11112));
  AND2 AND2_1027(.VSS(VSS),.VDD(VDD),.Y(g7145),.A(g6082),.B(g6718));
  AND2 AND2_1028(.VSS(VSS),.VDD(VDD),.Y(g5738),.A(g1586),.B(g5184));
  AND2 AND2_1029(.VSS(VSS),.VDD(VDD),.Y(g6826),.A(g225),.B(g6596));
  AND2 AND2_1030(.VSS(VSS),.VDD(VDD),.Y(g7191),.A(g6343),.B(g4323));
  AND2 AND2_1031(.VSS(VSS),.VDD(VDD),.Y(g3998),.A(g2677),.B(g2276));
  AND2 AND2_1032(.VSS(VSS),.VDD(VDD),.Y(g6741),.A(g3284),.B(g6141));
  AND2 AND2_1033(.VSS(VSS),.VDD(VDD),.Y(g5478),.A(g1905),.B(g4242));
  AND2 AND2_1034(.VSS(VSS),.VDD(VDD),.Y(g11167),.A(g538),.B(g11112));
  AND2 AND2_1035(.VSS(VSS),.VDD(VDD),.Y(g11194),.A(g5637),.B(g11067));
  AND2 AND2_1036(.VSS(VSS),.VDD(VDD),.Y(g11589),.A(g1333),.B(g11548));
  AND2 AND2_1037(.VSS(VSS),.VDD(VDD),.Y(g6638),.A(g64),.B(g6195));
  AND2 AND2_1038(.VSS(VSS),.VDD(VDD),.Y(g4921),.A(g2779),.B(g4431));
  AND2 AND2_1039(.VSS(VSS),.VDD(VDD),.Y(g7536),.A(g7148),.B(g2877));
  AND2 AND2_1040(.VSS(VSS),.VDD(VDD),.Y(g9585),.A(g889),.B(g8995));
  AND2 AND2_1041(.VSS(VSS),.VDD(VDD),.Y(g2957),.A(g2424),.B(g1663));
  AND2 AND2_1042(.VSS(VSS),.VDD(VDD),.Y(g11588),.A(g1330),.B(g11547));
  AND2 AND2_1043(.VSS(VSS),.VDD(VDD),.Y(g5690),.A(g1567),.B(g5112));
  AND2 AND2_1044(.VSS(VSS),.VDD(VDD),.Y(g6883),.A(g1923),.B(g6413));
  AND2 AND2_1045(.VSS(VSS),.VDD(VDD),.Y(g4837),.A(g1068),.B(g3638));
  AND3 AND3_36(.VSS(VSS),.VDD(VDD),.Y(g8963),.A(g8056),.B(g6368),.C(g8849));
  AND2 AND2_1046(.VSS(VSS),.VDD(VDD),.Y(g8791),.A(g8641),.B(g8721));
  AND2 AND2_1047(.VSS(VSS),.VDD(VDD),.Y(g6217),.A(g563),.B(g5073));
  AND4 AND4_10(.VSS(VSS),.VDD(VDD),.Y(I6316),.A(g2082),.B(g2087),.C(g2381),.D(g2395));
  AND2 AND2_1048(.VSS(VSS),.VDD(VDD),.Y(g11022),.A(g444),.B(g10974));
  AND2 AND2_1049(.VSS(VSS),.VDD(VDD),.Y(g5915),.A(g4168),.B(g4977));
  AND2 AND2_1050(.VSS(VSS),.VDD(VDD),.Y(g4788),.A(g511),.B(g3436));
  AND2 AND2_1051(.VSS(VSS),.VDD(VDD),.Y(g8759),.A(g7437),.B(g8677));
  AND2 AND2_1052(.VSS(VSS),.VDD(VDD),.Y(g5110),.A(g1806),.B(g4618));
  AND2 AND2_1053(.VSS(VSS),.VDD(VDD),.Y(g11254),.A(g986),.B(g11073));
  AND2 AND2_1054(.VSS(VSS),.VDD(VDD),.Y(g6827),.A(g219),.B(g6596));
  AND3 AND3_37(.VSS(VSS),.VDD(VDD),.Y(g8957),.A(g8081),.B(g6368),.C(g8828));
  AND2 AND2_1055(.VSS(VSS),.VDD(VDD),.Y(g6333),.A(g197),.B(g5904));
  AND2 AND2_1056(.VSS(VSS),.VDD(VDD),.Y(g8049),.A(g7567),.B(g5919));
  AND2 AND2_1057(.VSS(VSS),.VDD(VDD),.Y(g4392),.A(g3273),.B(g3829));
  AND2 AND2_1058(.VSS(VSS),.VDD(VDD),.Y(g9856),.A(g1592),.B(g9773));
  AND2 AND2_1059(.VSS(VSS),.VDD(VDD),.Y(g9411),.A(g1724),.B(g9052));
  AND2 AND2_1060(.VSS(VSS),.VDD(VDD),.Y(g5002),.A(g1494),.B(g4640));
  AND2 AND2_1061(.VSS(VSS),.VDD(VDD),.Y(g11101),.A(g857),.B(g10950));
  AND2 AND2_1062(.VSS(VSS),.VDD(VDD),.Y(g11177),.A(g511),.B(g11112));
  AND2 AND2_1063(.VSS(VSS),.VDD(VDD),.Y(g11560),.A(g2765),.B(g11519));
  AND2 AND2_1064(.VSS(VSS),.VDD(VDD),.Y(g8098),.A(g6201),.B(g7852));
  AND2 AND2_1065(.VSS(VSS),.VDD(VDD),.Y(g3970),.A(g225),.B(g3164));
  AND2 AND2_1066(.VSS(VSS),.VDD(VDD),.Y(g4941),.A(g1038),.B(g4451));
  AND2 AND2_1067(.VSS(VSS),.VDD(VDD),.Y(g10453),.A(g10437),.B(g3395));
  AND2 AND2_1068(.VSS(VSS),.VDD(VDD),.Y(g5877),.A(g4921),.B(g639));
  AND2 AND2_1069(.VSS(VSS),.VDD(VDD),.Y(g6662),.A(g366),.B(g6220));
  AND2 AND2_1070(.VSS(VSS),.VDD(VDD),.Y(g7935),.A(g2821),.B(g7454));
  AND2 AND2_1071(.VSS(VSS),.VDD(VDD),.Y(g6067),.A(g1047),.B(g5320));
  AND4 AND4_11(.VSS(VSS),.VDD(VDD),.Y(I6317),.A(g2406),.B(g2420),.C(g2434),.D(g2438));
  AND2 AND2_1072(.VSS(VSS),.VDD(VDD),.Y(g9863),.A(g9740),.B(g9576));
  AND4 AND4_12(.VSS(VSS),.VDD(VDD),.Y(I5886),.A(g174),.B(g170),.C(g2249),.D(g2254));
  AND2 AND2_1073(.VSS(VSS),.VDD(VDD),.Y(g6994),.A(g6758),.B(g3829));
  AND2 AND2_1074(.VSS(VSS),.VDD(VDD),.Y(g9713),.A(g1589),.B(g9474));
  AND2 AND2_1075(.VSS(VSS),.VDD(VDD),.Y(g4431),.A(g2268),.B(g3533));
  AND2 AND2_1076(.VSS(VSS),.VDD(VDD),.Y(g4252),.A(g1007),.B(g3914));
  AND2 AND2_1077(.VSS(VSS),.VDD(VDD),.Y(g11166),.A(g542),.B(g11112));
  AND2 AND2_1078(.VSS(VSS),.VDD(VDD),.Y(g7130),.A(g6041),.B(g6697));
  AND2 AND2_1079(.VSS(VSS),.VDD(VDD),.Y(g11009),.A(g5179),.B(g10827));
  AND2 AND2_1080(.VSS(VSS),.VDD(VDD),.Y(g7542),.A(g7148),.B(g2885));
  AND2 AND2_1081(.VSS(VSS),.VDD(VDD),.Y(g8019),.A(g7386),.B(g4332));
  AND2 AND2_1082(.VSS(VSS),.VDD(VDD),.Y(g11008),.A(g5171),.B(g10827));
  AND2 AND2_1083(.VSS(VSS),.VDD(VDD),.Y(g3516),.A(g1209),.B(g3015));
  AND2 AND2_1084(.VSS(VSS),.VDD(VDD),.Y(g8052),.A(g7573),.B(g5128));
  AND2 AND2_1085(.VSS(VSS),.VDD(VDD),.Y(g3987),.A(g243),.B(g3164));
  AND2 AND2_1086(.VSS(VSS),.VDD(VDD),.Y(g4765),.A(g491),.B(g3405));
  AND2 AND2_1087(.VSS(VSS),.VDD(VDD),.Y(g11555),.A(g2695),.B(g11519));
  AND2 AND2_1088(.VSS(VSS),.VDD(VDD),.Y(g9857),.A(g9734),.B(g9569));
  AND2 AND2_1089(.VSS(VSS),.VDD(VDD),.Y(g8728),.A(g8610),.B(g7915));
  AND2 AND2_1090(.VSS(VSS),.VDD(VDD),.Y(g8730),.A(g8613),.B(g7917));
  AND2 AND2_1091(.VSS(VSS),.VDD(VDD),.Y(g8185),.A(g664),.B(g7997));
  AND2 AND2_1092(.VSS(VSS),.VDD(VDD),.Y(g5194),.A(g1610),.B(g4717));
  AND2 AND2_1093(.VSS(VSS),.VDD(VDD),.Y(g8385),.A(g6084),.B(g8218));
  AND2 AND2_1094(.VSS(VSS),.VDD(VDD),.Y(g4610),.A(g3804),.B(g2212));
  AND2 AND2_1095(.VSS(VSS),.VDD(VDD),.Y(g7902),.A(g7661),.B(g6587));
  AND2 AND2_1096(.VSS(VSS),.VDD(VDD),.Y(g4073),.A(g3200),.B(g3222));
  AND2 AND2_1097(.VSS(VSS),.VDD(VDD),.Y(g8070),.A(g682),.B(g7826));
  AND2 AND2_1098(.VSS(VSS),.VDD(VDD),.Y(g5731),.A(g1583),.B(g5175));
  AND2 AND2_1099(.VSS(VSS),.VDD(VDD),.Y(g11238),.A(g5474),.B(g11110));
  AND2 AND2_1100(.VSS(VSS),.VDD(VDD),.Y(g4473),.A(g1125),.B(g3874));
  AND2 AND2_1101(.VSS(VSS),.VDD(VDD),.Y(g8470),.A(g8308),.B(g7427));
  AND2 AND2_1102(.VSS(VSS),.VDD(VDD),.Y(g5489),.A(g4287),.B(g3521));
  AND2 AND2_1103(.VSS(VSS),.VDD(VDD),.Y(g3991),.A(g1738),.B(g2774));
  AND4 AND4_13(.VSS(VSS),.VDD(VDD),.Y(I5887),.A(g2078),.B(g2083),.C(g166),.D(g2095));
  AND2 AND2_1104(.VSS(VSS),.VDD(VDD),.Y(g7823),.A(g1923),.B(g7479));
  AND2 AND2_1105(.VSS(VSS),.VDD(VDD),.Y(g4069),.A(g1762),.B(g2802));
  AND3 AND3_38(.VSS(VSS),.VDD(VDD),.Y(g11519),.A(g1317),.B(g3015),.C(g11492));
  AND2 AND2_1106(.VSS(VSS),.VDD(VDD),.Y(g11176),.A(g506),.B(g11112));
  AND2 AND2_1107(.VSS(VSS),.VDD(VDD),.Y(g11092),.A(g837),.B(g10950));
  AND2 AND2_1108(.VSS(VSS),.VDD(VDD),.Y(g11154),.A(g330),.B(g10932));
  AND2 AND2_1109(.VSS(VSS),.VDD(VDD),.Y(g9608),.A(g7),.B(g9292));
  AND2 AND2_1110(.VSS(VSS),.VDD(VDD),.Y(g11637),.A(g11626),.B(g5446));
  AND2 AND2_1111(.VSS(VSS),.VDD(VDD),.Y(g2091),.A(g976),.B(g971));
  AND2 AND2_1112(.VSS(VSS),.VDD(VDD),.Y(g8406),.A(g695),.B(g8131));
  AND2 AND2_1113(.VSS(VSS),.VDD(VDD),.Y(g5254),.A(g4335),.B(g4165));
  AND2 AND2_1114(.VSS(VSS),.VDD(VDD),.Y(g7260),.A(g6752),.B(g2345));
  AND2 AND2_1115(.VSS(VSS),.VDD(VDD),.Y(g5150),.A(g1275),.B(g4678));
  AND2 AND2_1116(.VSS(VSS),.VDD(VDD),.Y(g8766),.A(g8612),.B(g5151));
  AND2 AND2_1117(.VSS(VSS),.VDD(VDD),.Y(g9588),.A(g3272),.B(g9173));
  AND2 AND2_1118(.VSS(VSS),.VDD(VDD),.Y(g8801),.A(g8742),.B(g8729));
  AND2 AND2_1119(.VSS(VSS),.VDD(VDD),.Y(g7063),.A(g5903),.B(g6582));
  AND2 AND2_1120(.VSS(VSS),.VDD(VDD),.Y(g10303),.A(g10208),.B(g9076));
  AND2 AND2_1121(.VSS(VSS),.VDD(VDD),.Y(g5009),.A(g1486),.B(g4640));
  AND2 AND2_1122(.VSS(VSS),.VDD(VDD),.Y(g9665),.A(g1314),.B(g9151));
  AND2 AND2_1123(.VSS(VSS),.VDD(VDD),.Y(g8748),.A(g7670),.B(g8656));
  AND2 AND2_1124(.VSS(VSS),.VDD(VDD),.Y(g11215),.A(g953),.B(g11160));
  AND2 AND2_1125(.VSS(VSS),.VDD(VDD),.Y(g10750),.A(g10687),.B(g3586));
  AND3 AND3_39(.VSS(VSS),.VDD(VDD),.Y(g5769),.A(g2112),.B(g4921),.C(g3818));
  AND2 AND2_1126(.VSS(VSS),.VDD(VDD),.Y(g8755),.A(g7426),.B(g8671));
  AND2 AND2_1127(.VSS(VSS),.VDD(VDD),.Y(g6673),.A(g5305),.B(g5822));
  AND2 AND2_1128(.VSS(VSS),.VDD(VDD),.Y(g5212),.A(g1255),.B(g4726));
  AND2 AND2_1129(.VSS(VSS),.VDD(VDD),.Y(g7720),.A(g727),.B(g7232));
  AND3 AND3_40(.VSS(VSS),.VDD(VDD),.Y(g5918),.A(g2965),.B(g5292),.C(g4609));
  AND2 AND2_1130(.VSS(VSS),.VDD(VDD),.Y(g8045),.A(g7547),.B(g5128));
  AND2 AND2_1131(.VSS(VSS),.VDD(VDD),.Y(g8173),.A(g7971),.B(g3112));
  AND2 AND2_1132(.VSS(VSS),.VDD(VDD),.Y(g11349),.A(g11288),.B(g7964));
  AND2 AND2_1133(.VSS(VSS),.VDD(VDD),.Y(g7843),.A(g7599),.B(g5919));
  AND2 AND2_1134(.VSS(VSS),.VDD(VDD),.Y(g9696),.A(g281),.B(g9432));
  AND2 AND2_1135(.VSS(VSS),.VDD(VDD),.Y(g6772),.A(g6228),.B(g722));
  AND2 AND2_1136(.VSS(VSS),.VDD(VDD),.Y(g6058),.A(g1035),.B(g5320));
  AND2 AND2_1137(.VSS(VSS),.VDD(VDD),.Y(g6531),.A(g79),.B(g6056));
  AND2 AND2_1138(.VSS(VSS),.VDD(VDD),.Y(g6743),.A(g4106),.B(g6146));
  AND2 AND2_1139(.VSS(VSS),.VDD(VDD),.Y(g6890),.A(g6752),.B(g6568));
  AND2 AND2_1140(.VSS(VSS),.VDD(VDD),.Y(g7549),.A(g7269),.B(g3829));
  AND2 AND2_1141(.VSS(VSS),.VDD(VDD),.Y(g8169),.A(g5265),.B(g7853));
  AND2 AND2_1142(.VSS(VSS),.VDD(VDD),.Y(g11304),.A(g5520),.B(g11245));
  AND2 AND2_1143(.VSS(VSS),.VDD(VDD),.Y(g9944),.A(g9924),.B(g9392));
  AND2 AND2_1144(.VSS(VSS),.VDD(VDD),.Y(g9240),.A(g6454),.B(g8962));
  AND2 AND2_1145(.VSS(VSS),.VDD(VDD),.Y(g8059),.A(g7592),.B(g5919));
  AND2 AND2_1146(.VSS(VSS),.VDD(VDD),.Y(g8718),.A(g8600),.B(g7903));
  AND2 AND2_1147(.VSS(VSS),.VDD(VDD),.Y(g8767),.A(g8616),.B(g5151));
  AND2 AND2_1148(.VSS(VSS),.VDD(VDD),.Y(g9316),.A(g8877),.B(g5708));
  AND2 AND2_1149(.VSS(VSS),.VDD(VDD),.Y(g7625),.A(g673),.B(g7085));
  AND2 AND2_1150(.VSS(VSS),.VDD(VDD),.Y(g8793),.A(g8644),.B(g8723));
  AND2 AND2_1151(.VSS(VSS),.VDD(VDD),.Y(g2940),.A(g2424),.B(g1654));
  AND2 AND2_1152(.VSS(VSS),.VDD(VDD),.Y(g4114),.A(g1351),.B(g3301));
  AND2 AND2_1153(.VSS(VSS),.VDD(VDD),.Y(g11636),.A(g11624),.B(g7936));
  AND2 AND2_1154(.VSS(VSS),.VDD(VDD),.Y(g10949),.A(g2947),.B(g10809));
  AND2 AND2_1155(.VSS(VSS),.VDD(VDD),.Y(g4870),.A(g237),.B(g3946));
  AND2 AND2_1156(.VSS(VSS),.VDD(VDD),.Y(g3563),.A(g3275),.B(g2126));
  AND2 AND2_1157(.VSS(VSS),.VDD(VDD),.Y(g10948),.A(g2223),.B(g10809));
  AND2 AND2_1158(.VSS(VSS),.VDD(VDD),.Y(g8246),.A(g7846),.B(g7442));
  AND2 AND2_1159(.VSS(VSS),.VDD(VDD),.Y(g5788),.A(g1540),.B(g5231));
  AND2 AND2_1160(.VSS(VSS),.VDD(VDD),.Y(g4008),.A(g2689),.B(g2276));
  AND2 AND2_1161(.VSS(VSS),.VDD(VDD),.Y(g9596),.A(g2649),.B(g9010));
  AND2 AND2_1162(.VSS(VSS),.VDD(VDD),.Y(g5249),.A(g1089),.B(g4747));
  AND2 AND2_1163(.VSS(VSS),.VDD(VDD),.Y(g11585),.A(g1321),.B(g11543));
  AND2 AND2_1164(.VSS(VSS),.VDD(VDD),.Y(g3089),.A(g2054),.B(g2050));
  AND2 AND2_1165(.VSS(VSS),.VDD(VDD),.Y(g4972),.A(g1436),.B(g4682));
  AND2 AND2_1166(.VSS(VSS),.VDD(VDD),.Y(g11554),.A(g2689),.B(g11519));
  AND2 AND2_1167(.VSS(VSS),.VDD(VDD),.Y(g7586),.A(g7096),.B(g5423));
  AND2 AND2_1168(.VSS(VSS),.VDD(VDD),.Y(g10673),.A(g10580),.B(g9450));
  AND3 AND3_41(.VSS(VSS),.VDD(VDD),.Y(g4806),.A(g3215),.B(g3992),.C(g2493));
  AND2 AND2_1169(.VSS(VSS),.VDD(VDD),.Y(g5485),.A(g1914),.B(g4257));
  AND2 AND2_1170(.VSS(VSS),.VDD(VDD),.Y(g9936),.A(g9915),.B(g9624));
  AND2 AND2_1171(.VSS(VSS),.VDD(VDD),.Y(g2910),.A(g2424),.B(g1660));
  AND2 AND2_1172(.VSS(VSS),.VDD(VDD),.Y(g9317),.A(g6109),.B(g8875));
  AND2 AND2_1173(.VSS(VSS),.VDD(VDD),.Y(g10933),.A(g10853),.B(g3982));
  AND2 AND2_1174(.VSS(VSS),.VDD(VDD),.Y(g8388),.A(g8177),.B(g7689));
  AND2 AND2_1175(.VSS(VSS),.VDD(VDD),.Y(g4465),.A(g1117),.B(g3828));
  AND2 AND2_1176(.VSS(VSS),.VDD(VDD),.Y(g7141),.A(g6073),.B(g6716));
  AND2 AND2_1177(.VSS(VSS),.VDD(VDD),.Y(g10508),.A(g10391),.B(g2135));
  AND2 AND2_1178(.VSS(VSS),.VDD(VDD),.Y(g4230),.A(g1095),.B(g3638));
  AND2 AND2_1179(.VSS(VSS),.VDD(VDD),.Y(g10634),.A(g10604),.B(g3829));
  AND2 AND2_1180(.VSS(VSS),.VDD(VDD),.Y(g9601),.A(g922),.B(g9192));
  AND2 AND2_1181(.VSS(VSS),.VDD(VDD),.Y(g6126),.A(g5639),.B(g4319));
  AND2 AND2_1182(.VSS(VSS),.VDD(VDD),.Y(g6326),.A(g1250),.B(g5949));
  AND2 AND2_1183(.VSS(VSS),.VDD(VDD),.Y(g7710),.A(g700),.B(g7214));
  AND2 AND2_1184(.VSS(VSS),.VDD(VDD),.Y(g8028),.A(g7375),.B(g7436));
  AND2 AND2_1185(.VSS(VSS),.VDD(VDD),.Y(g6760),.A(g786),.B(g6221));
  AND2 AND2_1186(.VSS(VSS),.VDD(VDD),.Y(g5640),.A(g1059),.B(g4427));
  AND2 AND2_1187(.VSS(VSS),.VDD(VDD),.Y(g5031),.A(g1478),.B(g4640));
  AND2 AND2_1188(.VSS(VSS),.VDD(VDD),.Y(g4550),.A(g342),.B(g3586));
  AND2 AND2_1189(.VSS(VSS),.VDD(VDD),.Y(g7879),.A(g7610),.B(g3798));
  AND2 AND2_1190(.VSS(VSS),.VDD(VDD),.Y(g7962),.A(g7730),.B(g6712));
  AND2 AND2_1191(.VSS(VSS),.VDD(VDD),.Y(g9597),.A(g1170),.B(g9125));
  AND2 AND2_1192(.VSS(VSS),.VDD(VDD),.Y(g10452),.A(g10439),.B(g3388));
  AND2 AND2_1193(.VSS(VSS),.VDD(VDD),.Y(g4891),.A(g631),.B(g4739));
  AND2 AND2_1194(.VSS(VSS),.VDD(VDD),.Y(g5005),.A(g1490),.B(g4640));
  AND2 AND2_1195(.VSS(VSS),.VDD(VDD),.Y(g6423),.A(g4348),.B(g5784));
  AND2 AND2_1196(.VSS(VSS),.VDD(VDD),.Y(g8108),.A(g1891),.B(g7938));
  AND3 AND3_42(.VSS(VSS),.VDD(VDD),.Y(g4807),.A(g3015),.B(g1289),.C(g3937));
  AND2 AND2_1197(.VSS(VSS),.VDD(VDD),.Y(g5911),.A(g3322),.B(g4977));
  AND2 AND2_1198(.VSS(VSS),.VDD(VDD),.Y(g9937),.A(g9916),.B(g9624));
  AND2 AND2_1199(.VSS(VSS),.VDD(VDD),.Y(g9840),.A(g9704),.B(g9747));
  AND2 AND2_1200(.VSS(VSS),.VDD(VDD),.Y(g10780),.A(g10723),.B(g5124));
  AND2 AND2_1201(.VSS(VSS),.VDD(VDD),.Y(g8217),.A(g1872),.B(g7883));
  AND2 AND2_1202(.VSS(VSS),.VDD(VDD),.Y(g11013),.A(g5209),.B(g10827));
  AND2 AND2_1203(.VSS(VSS),.VDD(VDD),.Y(g9390),.A(g1333),.B(g9151));
  AND2 AND2_1204(.VSS(VSS),.VDD(VDD),.Y(g11214),.A(g950),.B(g11159));
  AND2 AND2_1205(.VSS(VSS),.VDD(VDD),.Y(g6327),.A(g1255),.B(g5949));
  AND2 AND2_1206(.VSS(VSS),.VDD(VDD),.Y(g4342),.A(g1149),.B(g3719));
  AND2 AND2_1207(.VSS(VSS),.VDD(VDD),.Y(g5796),.A(g1564),.B(g5252));
  AND2 AND2_1208(.VSS(VSS),.VDD(VDD),.Y(g5473),.A(g4268),.B(g3518));
  AND2 AND2_1209(.VSS(VSS),.VDD(VDD),.Y(g6346),.A(g5038),.B(g5883));
  AND2 AND2_1210(.VSS(VSS),.VDD(VDD),.Y(g6633),.A(g354),.B(g6191));
  AND2 AND2_1211(.VSS(VSS),.VDD(VDD),.Y(g11005),.A(g5119),.B(g10827));
  AND2 AND2_1212(.VSS(VSS),.VDD(VDD),.Y(g8365),.A(g668),.B(g8240));
  AND2 AND2_1213(.VSS(VSS),.VDD(VDD),.Y(g8048),.A(g7558),.B(g5919));
  AND2 AND2_1214(.VSS(VSS),.VDD(VDD),.Y(g4481),.A(g1713),.B(g3906));
  AND2 AND2_1215(.VSS(VSS),.VDD(VDD),.Y(g4097),.A(g2677),.B(g2989));
  AND2 AND2_1216(.VSS(VSS),.VDD(VDD),.Y(g8055),.A(g7588),.B(g5128));
  AND2 AND2_1217(.VSS(VSS),.VDD(VDD),.Y(g4497),.A(g351),.B(g3586));
  AND2 AND2_1218(.VSS(VSS),.VDD(VDD),.Y(g9942),.A(g9922),.B(g9367));
  AND2 AND2_1219(.VSS(VSS),.VDD(VDD),.Y(g6696),.A(g5504),.B(g5850));
  AND3 AND3_43(.VSS(VSS),.VDD(VDD),.Y(g10731),.A(g5118),.B(g1850),.C(g10665));
  AND2 AND2_1220(.VSS(VSS),.VDD(VDD),.Y(g8827),.A(g8552),.B(g8696));
  AND2 AND2_1221(.VSS(VSS),.VDD(VDD),.Y(g5540),.A(g1727),.B(g4315));
  AND2 AND2_1222(.VSS(VSS),.VDD(VDD),.Y(g4960),.A(g1403),.B(g4682));
  AND2 AND2_1223(.VSS(VSS),.VDD(VDD),.Y(g8846),.A(g8615),.B(g8712));
  AND2 AND2_1224(.VSS(VSS),.VDD(VDD),.Y(g6508),.A(g5983),.B(g3096));
  AND2 AND2_1225(.VSS(VSS),.VDD(VDD),.Y(g6240),.A(g182),.B(g5361));
  AND2 AND2_1226(.VSS(VSS),.VDD(VDD),.Y(g7931),.A(g2809),.B(g7446));
  AND2 AND2_1227(.VSS(VSS),.VDD(VDD),.Y(g5287),.A(g3876),.B(g4782));
  AND2 AND2_1228(.VSS(VSS),.VDD(VDD),.Y(g6472),.A(g5853),.B(g1936));
  AND2 AND2_1229(.VSS(VSS),.VDD(VDD),.Y(g11100),.A(g853),.B(g10950));
  AND2 AND2_1230(.VSS(VSS),.VDD(VDD),.Y(g11235),.A(g5443),.B(g11107));
  AND2 AND2_1231(.VSS(VSS),.VDD(VDD),.Y(g5199),.A(g1068),.B(g4719));
  AND2 AND2_1232(.VSS(VSS),.VDD(VDD),.Y(g6316),.A(g1270),.B(g5949));
  AND2 AND2_1233(.VSS(VSS),.VDD(VDD),.Y(g7515),.A(g7148),.B(g2855));
  AND2 AND2_1234(.VSS(VSS),.VDD(VDD),.Y(g10583),.A(g10518),.B(g10515));
  AND2 AND2_1235(.VSS(VSS),.VDD(VDD),.Y(g5781),.A(g1537),.B(g5222));
  AND2 AND2_1236(.VSS(VSS),.VDD(VDD),.Y(g8018),.A(g7742),.B(g7425));
  AND2 AND2_1237(.VSS(VSS),.VDD(VDD),.Y(g4401),.A(g2971),.B(g3772));
  AND3 AND3_44(.VSS(VSS),.VDD(VDD),.Y(g8994),.A(g8110),.B(g6778),.C(g8925));
  AND2 AND2_1238(.VSS(VSS),.VDD(VDD),.Y(g2950),.A(g2424),.B(g1666));
  AND2 AND2_1239(.VSS(VSS),.VDD(VDD),.Y(g5510),.A(g1630),.B(g4280));
  AND2 AND2_1240(.VSS(VSS),.VDD(VDD),.Y(g6347),.A(g275),.B(g5890));
  AND2 AND2_1241(.VSS(VSS),.VDD(VDD),.Y(g9357),.A(g962),.B(g9223));
  AND2 AND2_1242(.VSS(VSS),.VDD(VDD),.Y(g4828),.A(g4106),.B(g695));
  AND2 AND2_1243(.VSS(VSS),.VDD(VDD),.Y(g11407),.A(g11339),.B(g5949));
  AND2 AND2_1244(.VSS(VSS),.VDD(VDD),.Y(g4727),.A(g386),.B(g3364));
  AND2 AND2_1245(.VSS(VSS),.VDD(VDD),.Y(g10357),.A(g10278),.B(g2462));
  AND2 AND2_1246(.VSS(VSS),.VDD(VDD),.Y(g10743),.A(g10639),.B(g4013));
  AND2 AND2_1247(.VSS(VSS),.VDD(VDD),.Y(g5259),.A(g627),.B(g4739));
  AND2 AND2_1248(.VSS(VSS),.VDD(VDD),.Y(g5694),.A(g162),.B(g5361));
  AND2 AND2_1249(.VSS(VSS),.VDD(VDD),.Y(g10769),.A(g10652),.B(g4840));
  AND2 AND2_1250(.VSS(VSS),.VDD(VDD),.Y(g11584),.A(g1318),.B(g11542));
  AND2 AND2_1251(.VSS(VSS),.VDD(VDD),.Y(g4932),.A(g1065),.B(g4442));
  AND2 AND2_1252(.VSS(VSS),.VDD(VDD),.Y(g10768),.A(g10649),.B(g4840));
  AND2 AND2_1253(.VSS(VSS),.VDD(VDD),.Y(g6820),.A(g1362),.B(g6596));
  AND2 AND2_1254(.VSS(VSS),.VDD(VDD),.Y(g4068),.A(g2719),.B(g2276));
  AND2 AND2_1255(.VSS(VSS),.VDD(VDD),.Y(g6317),.A(g1304),.B(g5949));
  AND2 AND2_1256(.VSS(VSS),.VDD(VDD),.Y(g5215),.A(g4276),.B(g3400));
  AND2 AND2_1257(.VSS(VSS),.VDD(VDD),.Y(g4576),.A(g530),.B(g4049));
  AND2 AND2_1258(.VSS(VSS),.VDD(VDD),.Y(g4866),.A(g231),.B(g3946));
  AND2 AND2_1259(.VSS(VSS),.VDD(VDD),.Y(g6775),.A(g822),.B(g6231));
  AND2 AND2_1260(.VSS(VSS),.VDD(VDD),.Y(g3829),.A(g2028),.B(g2728));
  AND2 AND2_1261(.VSS(VSS),.VDD(VDD),.Y(g10662),.A(g8892),.B(g10571));
  AND2 AND2_1262(.VSS(VSS),.VDD(VDD),.Y(g8101),.A(g6208),.B(g7877));
  AND2 AND2_1263(.VSS(VSS),.VDD(VDD),.Y(g5825),.A(g3204),.B(g5318));
  AND4 AND4_14(.VSS(VSS),.VDD(VDD),.Y(I6310),.A(g2396),.B(g2407),.C(g2421),.D(g2435));
  AND2 AND2_1264(.VSS(VSS),.VDD(VDD),.Y(g7884),.A(g7457),.B(g7022));
  AND2 AND2_1265(.VSS(VSS),.VDD(VDD),.Y(g5008),.A(g1292),.B(g4507));
  AND2 AND2_1266(.VSS(VSS),.VDD(VDD),.Y(g3974),.A(g231),.B(g3164));
  AND2 AND2_1267(.VSS(VSS),.VDD(VDD),.Y(g9949),.A(g9929),.B(g9392));
  AND2 AND2_1268(.VSS(VSS),.VDD(VDD),.Y(g2531),.A(g658),.B(g668));
  AND2 AND2_1269(.VSS(VSS),.VDD(VDD),.Y(g9292),.A(g8878),.B(g5708));
  AND2 AND2_1270(.VSS(VSS),.VDD(VDD),.Y(g10778),.A(g1027),.B(g10729));
  AND2 AND2_1271(.VSS(VSS),.VDD(VDD),.Y(g8041),.A(g7524),.B(g5128));
  AND2 AND2_1272(.VSS(VSS),.VDD(VDD),.Y(g6079),.A(g1053),.B(g5320));
  AND2 AND2_1273(.VSS(VSS),.VDD(VDD),.Y(g7235),.A(g6663),.B(g6447));
  AND2 AND2_1274(.VSS(VSS),.VDD(VDD),.Y(g9603),.A(g1173),.B(g9125));
  AND2 AND2_1275(.VSS(VSS),.VDD(VDD),.Y(g6840),.A(g248),.B(g6596));
  AND2 AND2_1276(.VSS(VSS),.VDD(VDD),.Y(g9850),.A(g9726),.B(g9560));
  AND2 AND2_1277(.VSS(VSS),.VDD(VDD),.Y(g7988),.A(g1878),.B(g7379));
  AND2 AND2_1278(.VSS(VSS),.VDD(VDD),.Y(g5228),.A(g1086),.B(g4734));
  AND2 AND2_1279(.VSS(VSS),.VDD(VDD),.Y(g7134),.A(g5587),.B(g6354));
  AND2 AND2_1280(.VSS(VSS),.VDD(VDD),.Y(g5934),.A(g5215),.B(g1965));
  AND2 AND2_1281(.VSS(VSS),.VDD(VDD),.Y(g5230),.A(g1265),.B(g4735));
  AND2 AND2_1282(.VSS(VSS),.VDD(VDD),.Y(g8168),.A(g5262),.B(g7853));
  AND2 AND2_1283(.VSS(VSS),.VDD(VDD),.Y(g9583),.A(g886),.B(g8995));
  AND2 AND2_1284(.VSS(VSS),.VDD(VDD),.Y(g10672),.A(g10579),.B(g9449));
  AND2 AND2_1285(.VSS(VSS),.VDD(VDD),.Y(g3287),.A(g802),.B(g2534));
  AND2 AND2_1286(.VSS(VSS),.VDD(VDD),.Y(g8772),.A(g8627),.B(g5151));
  AND2 AND2_1287(.VSS(VSS),.VDD(VDD),.Y(g4893),.A(g635),.B(g4739));
  AND2 AND2_1288(.VSS(VSS),.VDD(VDD),.Y(g10331),.A(g10256),.B(g3307));
  AND2 AND2_1289(.VSS(VSS),.VDD(VDD),.Y(g8505),.A(g8309),.B(g4789));
  AND2 AND2_1290(.VSS(VSS),.VDD(VDD),.Y(g10449),.A(g10420),.B(g3345));
  AND2 AND2_1291(.VSS(VSS),.VDD(VDD),.Y(g11273),.A(g5638),.B(g11195));
  AND2 AND2_1292(.VSS(VSS),.VDD(VDD),.Y(g8734),.A(g8626),.B(g7923));
  AND2 AND2_1293(.VSS(VSS),.VDD(VDD),.Y(g5913),.A(g1041),.B(g5320));
  AND2 AND2_1294(.VSS(VSS),.VDD(VDD),.Y(g10448),.A(g10421),.B(g3335));
  AND2 AND2_1295(.VSS(VSS),.VDD(VDD),.Y(g6163),.A(g4572),.B(g5354));
  AND2 AND2_1296(.VSS(VSS),.VDD(VDD),.Y(g6363),.A(g284),.B(g5901));
  AND2 AND2_1297(.VSS(VSS),.VDD(VDD),.Y(g7202),.A(g6349),.B(g4329));
  AND2 AND2_1298(.VSS(VSS),.VDD(VDD),.Y(g11463),.A(g11432),.B(g5446));
  AND2 AND2_1299(.VSS(VSS),.VDD(VDD),.Y(g8074),.A(g718),.B(g7826));
  AND2 AND2_1300(.VSS(VSS),.VDD(VDD),.Y(g4325),.A(g1166),.B(g3682));
  AND2 AND2_1301(.VSS(VSS),.VDD(VDD),.Y(g8474),.A(g8383),.B(g5285));
  AND2 AND2_1302(.VSS(VSS),.VDD(VDD),.Y(g11234),.A(g5424),.B(g11106));
  AND2 AND2_1303(.VSS(VSS),.VDD(VDD),.Y(g5266),.A(g718),.B(g4766));
  AND2 AND2_1304(.VSS(VSS),.VDD(VDD),.Y(g4483),.A(g336),.B(g3586));
  AND2 AND2_1305(.VSS(VSS),.VDD(VDD),.Y(g5248),.A(g673),.B(g4738));
  AND2 AND2_1306(.VSS(VSS),.VDD(VDD),.Y(g11514),.A(g11491),.B(g5151));
  AND2 AND2_1307(.VSS(VSS),.VDD(VDD),.Y(g5255),.A(g682),.B(g4754));
  AND2 AND2_1308(.VSS(VSS),.VDD(VDD),.Y(g4106),.A(g3284),.B(g686));
  AND2 AND2_1309(.VSS(VSS),.VDD(VDD),.Y(g2760),.A(g981),.B(g2091));
  AND2 AND2_1310(.VSS(VSS),.VDD(VDD),.Y(g5097),.A(g1786),.B(g4603));
  AND2 AND2_1311(.VSS(VSS),.VDD(VDD),.Y(g5726),.A(g1601),.B(g5167));
  AND2 AND2_1312(.VSS(VSS),.VDD(VDD),.Y(g5497),.A(g4296),.B(g3522));
  AND2 AND2_1313(.VSS(VSS),.VDD(VDD),.Y(g5354),.A(g2733),.B(g4460));
  AND2 AND2_1314(.VSS(VSS),.VDD(VDD),.Y(g7933),.A(g2814),.B(g7450));
  AND2 AND2_1315(.VSS(VSS),.VDD(VDD),.Y(g9617),.A(g9),.B(g9274));
  AND2 AND2_1316(.VSS(VSS),.VDD(VDD),.Y(g9906),.A(g9873),.B(g9683));
  AND2 AND2_1317(.VSS(VSS),.VDD(VDD),.Y(g11012),.A(g5196),.B(g10827));
  AND2 AND2_1318(.VSS(VSS),.VDD(VDD),.Y(g7050),.A(g5896),.B(g6575));
  AND2 AND2_1319(.VSS(VSS),.VDD(VDD),.Y(g10971),.A(g10849),.B(g3161));
  AND2 AND2_1320(.VSS(VSS),.VDD(VDD),.Y(g4904),.A(g1850),.B(g4243));
  AND2 AND2_1321(.VSS(VSS),.VDD(VDD),.Y(g10369),.A(g10361),.B(g3382));
  AND2 AND2_1322(.VSS(VSS),.VDD(VDD),.Y(g8400),.A(g6097),.B(g8234));
  AND2 AND2_1323(.VSS(VSS),.VDD(VDD),.Y(g4345),.A(g1169),.B(g3730));
  AND2 AND2_1324(.VSS(VSS),.VDD(VDD),.Y(g2161),.A(I5084),.B(I5085));
  AND2 AND2_1325(.VSS(VSS),.VDD(VDD),.Y(g5001),.A(g1300),.B(g4491));
  AND2 AND2_1326(.VSS(VSS),.VDD(VDD),.Y(g9945),.A(g9925),.B(g9392));
  AND2 AND2_1327(.VSS(VSS),.VDD(VDD),.Y(g7271),.A(g5028),.B(g6499));
  AND2 AND2_1328(.VSS(VSS),.VDD(VDD),.Y(g9709),.A(g1524),.B(g9490));
  AND2 AND2_1329(.VSS(VSS),.VDD(VDD),.Y(g4223),.A(g1003),.B(g3914));
  AND2 AND2_1330(.VSS(VSS),.VDD(VDD),.Y(g10716),.A(g10497),.B(g10675));
  AND2 AND2_1331(.VSS(VSS),.VDD(VDD),.Y(g11291),.A(g11247),.B(g4233));
  AND2 AND2_1332(.VSS(VSS),.VDD(VDD),.Y(g6661),.A(g73),.B(g6219));
  AND2 AND2_1333(.VSS(VSS),.VDD(VDD),.Y(g11173),.A(g491),.B(g11112));
  AND2 AND2_1334(.VSS(VSS),.VDD(VDD),.Y(g6075),.A(g549),.B(g5613));
  AND2 AND2_1335(.VSS(VSS),.VDD(VDD),.Y(g8023),.A(g7367),.B(g7430));
  AND2 AND2_1336(.VSS(VSS),.VDD(VDD),.Y(g9907),.A(g9888),.B(g9686));
  AND2 AND2_1337(.VSS(VSS),.VDD(VDD),.Y(g10582),.A(g10532),.B(g9473));
  AND2 AND2_1338(.VSS(VSS),.VDD(VDD),.Y(g5746),.A(g1589),.B(g5193));
  AND2 AND2_1339(.VSS(VSS),.VDD(VDD),.Y(g5221),.A(g1260),.B(g4730));
  AND2 AND2_1340(.VSS(VSS),.VDD(VDD),.Y(g9959),.A(g9950),.B(g9536));
  AND2 AND2_1341(.VSS(VSS),.VDD(VDD),.Y(g7674),.A(g7004),.B(g3880));
  AND2 AND2_1342(.VSS(VSS),.VDD(VDD),.Y(g9690),.A(g266),.B(g9432));
  AND2 AND2_1343(.VSS(VSS),.VDD(VDD),.Y(g6627),.A(g58),.B(g6181));
  AND2 AND2_1344(.VSS(VSS),.VDD(VDD),.Y(g5703),.A(g174),.B(g5361));
  AND2 AND2_1345(.VSS(VSS),.VDD(VDD),.Y(g4522),.A(g360),.B(g3586));
  AND2 AND2_1346(.VSS(VSS),.VDD(VDD),.Y(g4115),.A(g2689),.B(g3009));
  AND2 AND2_1347(.VSS(VSS),.VDD(VDD),.Y(g7541),.A(g7075),.B(g3109));
  AND2 AND2_1348(.VSS(VSS),.VDD(VDD),.Y(g10627),.A(g10548),.B(g4564));
  AND2 AND2_1349(.VSS(VSS),.VDD(VDD),.Y(g4047),.A(g2695),.B(g2276));
  AND2 AND2_1350(.VSS(VSS),.VDD(VDD),.Y(g6526),.A(g76),.B(g6052));
  AND2 AND2_1351(.VSS(VSS),.VDD(VDD),.Y(g2944),.A(g2424),.B(g1669));
  AND2 AND2_1352(.VSS(VSS),.VDD(VDD),.Y(g6646),.A(g360),.B(g6203));
  AND2 AND2_1353(.VSS(VSS),.VDD(VDD),.Y(g7132),.A(g6048),.B(g6702));
  AND2 AND2_1354(.VSS(VSS),.VDD(VDD),.Y(g11029),.A(g401),.B(g10974));
  AND2 AND2_1355(.VSS(VSS),.VDD(VDD),.Y(g8051),.A(g7572),.B(g5128));
  AND2 AND2_1356(.VSS(VSS),.VDD(VDD),.Y(g8127),.A(g1927),.B(g7949));
  AND2 AND2_1357(.VSS(VSS),.VDD(VDD),.Y(g7209),.A(g3804),.B(g6425));
  AND2 AND2_1358(.VSS(VSS),.VDD(VDD),.Y(g11028),.A(g396),.B(g10974));
  AND2 AND2_1359(.VSS(VSS),.VDD(VDD),.Y(g6439),.A(g4479),.B(g5919));
  AND2 AND2_1360(.VSS(VSS),.VDD(VDD),.Y(g10742),.A(g10655),.B(g3586));
  AND2 AND2_1361(.VSS(VSS),.VDD(VDD),.Y(g9110),.A(g8880),.B(g4790));
  AND2 AND2_1362(.VSS(VSS),.VDD(VDD),.Y(g10681),.A(g10567),.B(g3586));
  AND2 AND2_1363(.VSS(VSS),.VDD(VDD),.Y(g4537),.A(g444),.B(g3988));
  AND2 AND2_1364(.VSS(VSS),.VDD(VDD),.Y(g9663),.A(g959),.B(g9223));
  AND2 AND2_1365(.VSS(VSS),.VDD(VDD),.Y(g5349),.A(g2126),.B(g4617));
  AND2 AND2_1366(.VSS(VSS),.VDD(VDD),.Y(g8732),.A(g8624),.B(g7919));
  AND2 AND2_1367(.VSS(VSS),.VDD(VDD),.Y(g3807),.A(g3003),.B(g3062));
  AND2 AND2_1368(.VSS(VSS),.VDD(VDD),.Y(g8753),.A(g7414),.B(g8664));
  AND2 AND2_1369(.VSS(VSS),.VDD(VDD),.Y(g5848),.A(g3860),.B(g5519));
  AND2 AND2_1370(.VSS(VSS),.VDD(VDD),.Y(g8508),.A(g8411),.B(g7967));
  AND2 AND2_1371(.VSS(VSS),.VDD(VDD),.Y(g8072),.A(g700),.B(g7826));
  AND2 AND2_1372(.VSS(VSS),.VDD(VDD),.Y(g5699),.A(g1592),.B(g5117));
  AND2 AND2_1373(.VSS(VSS),.VDD(VDD),.Y(g11240),.A(g5481),.B(g11111));
  AND2 AND2_1374(.VSS(VSS),.VDD(VDD),.Y(g5398),.A(g4610),.B(g2224));
  AND2 AND2_1375(.VSS(VSS),.VDD(VDD),.Y(g6616),.A(g6105),.B(g3246));
  AND2 AND2_1376(.VSS(VSS),.VDD(VDD),.Y(g10690),.A(g10616),.B(g3863));
  AND2 AND2_1377(.VSS(VSS),.VDD(VDD),.Y(g8043),.A(g7582),.B(g5128));
  AND2 AND2_1378(.VSS(VSS),.VDD(VDD),.Y(g9590),.A(g895),.B(g8995));
  AND2 AND2_1379(.VSS(VSS),.VDD(VDD),.Y(g4128),.A(g1976),.B(g2779));
  AND2 AND2_1380(.VSS(VSS),.VDD(VDD),.Y(g6404),.A(g2132),.B(g5748));
  AND2 AND2_1381(.VSS(VSS),.VDD(VDD),.Y(g6647),.A(g5288),.B(g5808));
  AND2 AND2_1382(.VSS(VSS),.VDD(VDD),.Y(g10504),.A(g10389),.B(g2135));
  AND2 AND2_1383(.VSS(VSS),.VDD(VDD),.Y(g9657),.A(g919),.B(g9205));
  AND2 AND2_1384(.VSS(VSS),.VDD(VDD),.Y(g4542),.A(g366),.B(g3586));
  AND2 AND2_1385(.VSS(VSS),.VDD(VDD),.Y(g4330),.A(g1163),.B(g3693));
  AND2 AND2_1386(.VSS(VSS),.VDD(VDD),.Y(g3497),.A(g2804),.B(g1900));
  AND2 AND2_1387(.VSS(VSS),.VDD(VDD),.Y(g5524),.A(g1678),.B(g4291));
  AND2 AND2_1388(.VSS(VSS),.VDD(VDD),.Y(g8147),.A(g2955),.B(g7961));
  AND2 AND2_1389(.VSS(VSS),.VDD(VDD),.Y(g4554),.A(g542),.B(g3996));
  AND2 AND2_1390(.VSS(VSS),.VDD(VDD),.Y(g9899),.A(g9889),.B(g9367));
  AND2 AND2_1391(.VSS(VSS),.VDD(VDD),.Y(g5258),.A(g700),.B(g4756));
  AND2 AND2_1392(.VSS(VSS),.VDD(VDD),.Y(g7736),.A(g6951),.B(g3880));
  AND2 AND2_1393(.VSS(VSS),.VDD(VDD),.Y(g6224),.A(g1520),.B(g5151));
  AND2 AND2_1394(.VSS(VSS),.VDD(VDD),.Y(g10626),.A(g10547),.B(g4558));
  AND2 AND2_1395(.VSS(VSS),.VDD(VDD),.Y(g6320),.A(g1292),.B(g5949));
  AND2 AND2_1396(.VSS(VSS),.VDD(VDD),.Y(g7623),.A(g664),.B(g7079));
  AND2 AND2_1397(.VSS(VSS),.VDD(VDD),.Y(g10299),.A(g8892),.B(g10217));
  AND2 AND2_1398(.VSS(VSS),.VDD(VDD),.Y(g7889),.A(g7615),.B(g3814));
  AND2 AND2_1399(.VSS(VSS),.VDD(VDD),.Y(g10298),.A(g8892),.B(g10214));
  AND2 AND2_1400(.VSS(VSS),.VDD(VDD),.Y(g8413),.A(g722),.B(g8146));
  AND2 AND2_1401(.VSS(VSS),.VDD(VDD),.Y(g3979),.A(g237),.B(g3164));
  AND2 AND2_1402(.VSS(VSS),.VDD(VDD),.Y(g4902),.A(g1848),.B(g4243));
  AND2 AND2_1403(.VSS(VSS),.VDD(VDD),.Y(g5211),.A(g1080),.B(g4724));
  AND2 AND2_1404(.VSS(VSS),.VDD(VDD),.Y(g4512),.A(g357),.B(g3586));
  AND2 AND2_1405(.VSS(VSS),.VDD(VDD),.Y(g7722),.A(g7127),.B(g6449));
  AND2 AND2_1406(.VSS(VSS),.VDD(VDD),.Y(g9844),.A(g9714),.B(g9522));
  AND2 AND2_1407(.VSS(VSS),.VDD(VDD),.Y(g4490),.A(g1141),.B(g3913));
  AND2 AND2_1408(.VSS(VSS),.VDD(VDD),.Y(g4823),.A(g207),.B(g3946));
  AND2 AND2_1409(.VSS(VSS),.VDD(VDD),.Y(g6516),.A(g5993),.B(g3097));
  AND2 AND2_1410(.VSS(VSS),.VDD(VDD),.Y(g5026),.A(g1453),.B(g4640));
  AND2 AND2_1411(.VSS(VSS),.VDD(VDD),.Y(g8820),.A(g8705),.B(g5422));
  AND2 AND2_1412(.VSS(VSS),.VDD(VDD),.Y(g10737),.A(g10687),.B(g4840));
  AND3 AND3_45(.VSS(VSS),.VDD(VDD),.Y(g8936),.A(g8115),.B(g6778),.C(g8849));
  AND2 AND2_1413(.VSS(VSS),.VDD(VDD),.Y(g10232),.A(g8892),.B(g10150));
  AND2 AND2_1414(.VSS(VSS),.VDD(VDD),.Y(g6771),.A(g263),.B(g5866));
  AND2 AND2_1415(.VSS(VSS),.VDD(VDD),.Y(g5170),.A(g1811),.B(g4680));
  AND2 AND2_1416(.VSS(VSS),.VDD(VDD),.Y(g8117),.A(g6236),.B(g7886));
  AND2 AND2_1417(.VSS(VSS),.VDD(VDD),.Y(g4529),.A(g448),.B(g3980));
  AND2 AND2_1418(.VSS(VSS),.VDD(VDD),.Y(g4348),.A(g3497),.B(g1909));
  AND2 AND2_1419(.VSS(VSS),.VDD(VDD),.Y(g9966),.A(g9956),.B(g9536));
  AND2 AND2_1420(.VSS(VSS),.VDD(VDD),.Y(g5280),.A(g4593),.B(g3052));
  AND2 AND2_1421(.VSS(VSS),.VDD(VDD),.Y(g7139),.A(g6060),.B(g6709));
  AND2 AND2_1422(.VSS(VSS),.VDD(VDD),.Y(g11099),.A(g382),.B(g10885));
  AND2 AND2_1423(.VSS(VSS),.VDD(VDD),.Y(g6892),.A(g6472),.B(g5805));
  AND2 AND2_1424(.VSS(VSS),.VDD(VDD),.Y(g9705),.A(g1580),.B(g9474));
  AND2 AND2_1425(.VSS(VSS),.VDD(VDD),.Y(g10512),.A(g10395),.B(g2135));
  AND2 AND2_1426(.VSS(VSS),.VDD(VDD),.Y(g11098),.A(g849),.B(g10950));
  AND2 AND2_1427(.VSS(VSS),.VDD(VDD),.Y(g8775),.A(g8628),.B(g5151));
  AND2 AND2_1428(.VSS(VSS),.VDD(VDD),.Y(g5083),.A(g3709),.B(g4586));
  AND2 AND2_1429(.VSS(VSS),.VDD(VDD),.Y(g5544),.A(g1687),.B(g4320));
  AND2 AND2_1430(.VSS(VSS),.VDD(VDD),.Y(g11272),.A(g5629),.B(g11193));
  AND2 AND2_1431(.VSS(VSS),.VDD(VDD),.Y(g5483),.A(g1621),.B(g4254));
  AND2 AND2_1432(.VSS(VSS),.VDD(VDD),.Y(g9948),.A(g9928),.B(g9392));
  AND2 AND2_1433(.VSS(VSS),.VDD(VDD),.Y(g4063),.A(g2713),.B(g2276));
  AND2 AND2_1434(.VSS(VSS),.VDD(VDD),.Y(g11462),.A(g11431),.B(g5446));
  AND2 AND2_1435(.VSS(VSS),.VDD(VDD),.Y(g6738),.A(g2531),.B(g6137));
  AND2 AND2_1436(.VSS(VSS),.VDD(VDD),.Y(g8060),.A(g7593),.B(g5919));
  AND2 AND2_1437(.VSS(VSS),.VDD(VDD),.Y(g6244),.A(g2255),.B(g5151));
  AND2 AND2_1438(.VSS(VSS),.VDD(VDD),.Y(g11032),.A(g416),.B(g10974));
  AND2 AND2_1439(.VSS(VSS),.VDD(VDD),.Y(g10445),.A(g10315),.B(g2135));
  AND2 AND2_1440(.VSS(VSS),.VDD(VDD),.Y(g9150),.A(g8882),.B(g4805));
  AND2 AND2_1441(.VSS(VSS),.VDD(VDD),.Y(g10316),.A(g10223),.B(g9097));
  AND2 AND2_1442(.VSS(VSS),.VDD(VDD),.Y(g5756),.A(g1531),.B(g5202));
  AND2 AND2_1443(.VSS(VSS),.VDD(VDD),.Y(g4720),.A(g1023),.B(g3914));
  AND2 AND2_1444(.VSS(VSS),.VDD(VDD),.Y(g9409),.A(g1721),.B(g9052));
  AND2 AND2_1445(.VSS(VSS),.VDD(VDD),.Y(g8995),.A(g6454),.B(g8929));
  AND2 AND2_1446(.VSS(VSS),.VDD(VDD),.Y(g6876),.A(g4070),.B(g6560));
  AND2 AND2_1447(.VSS(VSS),.VDD(VDD),.Y(g4989),.A(g1424),.B(g4682));
  AND2 AND2_1448(.VSS(VSS),.VDD(VDD),.Y(g9836),.A(g9737),.B(g9785));
  AND3 AND3_46(.VSS(VSS),.VDD(VDD),.Y(g6656),.A(g2733),.B(g6061),.C(g4631));
  AND2 AND2_1449(.VSS(VSS),.VDD(VDD),.Y(g5514),.A(g1941),.B(g4284));
  AND2 AND2_1450(.VSS(VSS),.VDD(VDD),.Y(g8390),.A(g8268),.B(g6465));
  AND2 AND2_1451(.VSS(VSS),.VDD(VDD),.Y(g5003),.A(g1466),.B(g4640));
  AND2 AND2_1452(.VSS(VSS),.VDD(VDD),.Y(g9967),.A(g9957),.B(g9536));
  AND2 AND2_1453(.VSS(VSS),.VDD(VDD),.Y(g5145),.A(g1639),.B(g4673));
  AND2 AND2_1454(.VSS(VSS),.VDD(VDD),.Y(g4834),.A(g219),.B(g3946));
  AND2 AND2_1455(.VSS(VSS),.VDD(VDD),.Y(g4971),.A(g1419),.B(g4682));
  AND2 AND2_1456(.VSS(VSS),.VDD(VDD),.Y(g10753),.A(g10649),.B(g4013));
  AND2 AND2_1457(.VSS(VSS),.VDD(VDD),.Y(g5695),.A(g166),.B(g5361));
  AND2 AND2_1458(.VSS(VSS),.VDD(VDD),.Y(g7613),.A(g6940),.B(g5984));
  AND2 AND2_1459(.VSS(VSS),.VDD(VDD),.Y(g10736),.A(g10658),.B(g4840));
  AND2 AND2_1460(.VSS(VSS),.VDD(VDD),.Y(g11220),.A(g962),.B(g11054));
  AND2 AND2_1461(.VSS(VSS),.VDD(VDD),.Y(g7444),.A(g7277),.B(g5827));
  AND2 AND2_1462(.VSS(VSS),.VDD(VDD),.Y(g5536),.A(g4867),.B(g4298));
  AND2 AND2_1463(.VSS(VSS),.VDD(VDD),.Y(g6663),.A(g6064),.B(g2237));
  AND2 AND2_1464(.VSS(VSS),.VDD(VDD),.Y(g4670),.A(g192),.B(g3946));
  AND2 AND2_1465(.VSS(VSS),.VDD(VDD),.Y(g6824),.A(g1371),.B(g6596));
  AND2 AND2_1466(.VSS(VSS),.VDD(VDD),.Y(g4253),.A(g1074),.B(g3638));
  AND2 AND2_1467(.VSS(VSS),.VDD(VDD),.Y(g8250),.A(g2771),.B(g7907));
  AND2 AND2_1468(.VSS(VSS),.VDD(VDD),.Y(g8163),.A(g7960),.B(g3737));
  AND2 AND2_1469(.VSS(VSS),.VDD(VDD),.Y(g10764),.A(g10643),.B(g4840));
  AND2 AND2_1470(.VSS(VSS),.VDD(VDD),.Y(g5757),.A(g1552),.B(g5203));
  AND2 AND2_1471(.VSS(VSS),.VDD(VDD),.Y(g10365),.A(g10319),.B(g2135));
  AND2 AND2_1472(.VSS(VSS),.VDD(VDD),.Y(g8032),.A(g7385),.B(g7438));
  AND2 AND2_1473(.VSS(VSS),.VDD(VDD),.Y(g11591),.A(g2988),.B(g11561));
  AND2 AND2_1474(.VSS(VSS),.VDD(VDD),.Y(g8053),.A(g7583),.B(g5919));
  AND2 AND2_1475(.VSS(VSS),.VDD(VDD),.Y(g11147),.A(g321),.B(g10929));
  AND2 AND2_1476(.VSS(VSS),.VDD(VDD),.Y(g5522),.A(g1633),.B(g4289));
  AND2 AND2_1477(.VSS(VSS),.VDD(VDD),.Y(g5115),.A(g1394),.B(g4572));
  AND2 AND2_1478(.VSS(VSS),.VDD(VDD),.Y(g9837),.A(g9697),.B(g9751));
  AND2 AND2_1479(.VSS(VSS),.VDD(VDD),.Y(g9620),.A(g2653),.B(g9240));
  AND2 AND2_1480(.VSS(VSS),.VDD(VDD),.Y(g11151),.A(g327),.B(g10931));
  AND2 AND2_1481(.VSS(VSS),.VDD(VDD),.Y(g11172),.A(g486),.B(g11112));
  AND2 AND2_1482(.VSS(VSS),.VDD(VDD),.Y(g7885),.A(g7614),.B(g3812));
  AND2 AND2_1483(.VSS(VSS),.VDD(VDD),.Y(g6064),.A(g5398),.B(g2230));
  AND3 AND3_47(.VSS(VSS),.VDD(VDD),.Y(g8929),.A(g8095),.B(g6368),.C(g8828));
  AND2 AND2_1484(.VSS(VSS),.VDD(VDD),.Y(g5595),.A(g1621),.B(g4524));
  AND2 AND2_1485(.VSS(VSS),.VDD(VDD),.Y(g5537),.A(g4143),.B(g4299));
  AND2 AND2_1486(.VSS(VSS),.VDD(VDD),.Y(g9842),.A(g9708),.B(g9516));
  AND2 AND2_1487(.VSS(VSS),.VDD(VDD),.Y(g4141),.A(g2707),.B(g3051));
  AND2 AND2_1488(.VSS(VSS),.VDD(VDD),.Y(g4341),.A(g339),.B(g3586));
  AND2 AND2_1489(.VSS(VSS),.VDD(VDD),.Y(g9192),.A(g6454),.B(g8955));
  AND2 AND2_1490(.VSS(VSS),.VDD(VDD),.Y(g7679),.A(g1950),.B(g6863));
  AND2 AND2_1491(.VSS(VSS),.VDD(VDD),.Y(g7378),.A(g6990),.B(g3880));
  AND2 AND2_1492(.VSS(VSS),.VDD(VDD),.Y(g5612),.A(g1627),.B(g4543));
  AND2 AND2_1493(.VSS(VSS),.VDD(VDD),.Y(g3939),.A(g213),.B(g3164));
  AND2 AND2_1494(.VSS(VSS),.VDD(VDD),.Y(g7135),.A(g869),.B(g6355));
  AND2 AND2_1495(.VSS(VSS),.VDD(VDD),.Y(g10970),.A(g10852),.B(g3390));
  AND2 AND2_1496(.VSS(VSS),.VDD(VDD),.Y(g11025),.A(g426),.B(g10974));
  AND2 AND2_1497(.VSS(VSS),.VDD(VDD),.Y(g9854),.A(g9730),.B(g9566));
  AND2 AND2_1498(.VSS(VSS),.VDD(VDD),.Y(g7182),.A(g1878),.B(g6720));
  AND2 AND2_1499(.VSS(VSS),.VDD(VDD),.Y(g9941),.A(g9921),.B(g9367));
  AND2 AND2_1500(.VSS(VSS),.VDD(VDD),.Y(g6194),.A(g554),.B(g5043));
  AND2 AND2_1501(.VSS(VSS),.VDD(VDD),.Y(g5128),.A(g4474),.B(g2733));
  AND2 AND2_1502(.VSS(VSS),.VDD(VDD),.Y(g4962),.A(g1651),.B(g4461));
  AND2 AND2_1503(.VSS(VSS),.VDD(VDD),.Y(g4358),.A(g1209),.B(g3747));
  AND2 AND2_1504(.VSS(VSS),.VDD(VDD),.Y(g8683),.A(g4803),.B(g8549));
  AND2 AND2_1505(.VSS(VSS),.VDD(VDD),.Y(g4506),.A(g1113),.B(g3944));
  AND2 AND2_1506(.VSS(VSS),.VDD(VDD),.Y(g6471),.A(g5224),.B(g6014));
  AND2 AND2_1507(.VSS(VSS),.VDD(VDD),.Y(g8778),.A(g8688),.B(g2317));
  AND2 AND2_1508(.VSS(VSS),.VDD(VDD),.Y(g11281),.A(g4948),.B(g11202));
  AND2 AND2_1509(.VSS(VSS),.VDD(VDD),.Y(g8735),.A(g7600),.B(g8632));
  AND2 AND2_1510(.VSS(VSS),.VDD(VDD),.Y(g11146),.A(g318),.B(g10928));
  AND2 AND2_1511(.VSS(VSS),.VDD(VDD),.Y(g3904),.A(g2948),.B(g2779));
  AND2 AND2_1512(.VSS(VSS),.VDD(VDD),.Y(g8075),.A(g727),.B(g7826));
  AND2 AND2_1513(.VSS(VSS),.VDD(VDD),.Y(g9829),.A(g9723),.B(g9785));
  AND3 AND3_48(.VSS(VSS),.VDD(VDD),.Y(g8949),.A(g8255),.B(g6368),.C(g8828));
  AND2 AND2_1514(.VSS(VSS),.VDD(VDD),.Y(g7632),.A(g7184),.B(g5574));
  AND2 AND2_1515(.VSS(VSS),.VDD(VDD),.Y(g11290),.A(g11246),.B(g4226));
  AND2 AND2_1516(.VSS(VSS),.VDD(VDD),.Y(g6350),.A(g5837),.B(g4435));
  AND2 AND2_1517(.VSS(VSS),.VDD(VDD),.Y(g10599),.A(g10534),.B(g4365));
  AND2 AND2_1518(.VSS(VSS),.VDD(VDD),.Y(g5902),.A(g2555),.B(g4977));
  AND4 AND4_15(.VSS(VSS),.VDD(VDD),.Y(I6337),.A(g201),.B(g2421),.C(g2407),.D(g2396));
  AND2 AND2_1519(.VSS(VSS),.VDD(VDD),.Y(g2276),.A(g1765),.B(g1610));
  AND2 AND2_1520(.VSS(VSS),.VDD(VDD),.Y(g6438),.A(g5853),.B(g5797));
  AND2 AND2_1521(.VSS(VSS),.VDD(VDD),.Y(g5512),.A(g1660),.B(g4281));
  AND2 AND2_1522(.VSS(VSS),.VDD(VDD),.Y(g5090),.A(g1781),.B(g4592));
  AND2 AND2_1523(.VSS(VSS),.VDD(VDD),.Y(g7719),.A(g718),.B(g7227));
  AND2 AND2_1524(.VSS(VSS),.VDD(VDD),.Y(g2561),.A(g742),.B(g741));
  AND2 AND2_1525(.VSS(VSS),.VDD(VDD),.Y(g3695),.A(g1712),.B(g3015));
  AND2 AND2_1526(.VSS(VSS),.VDD(VDD),.Y(g8603),.A(g3983),.B(g8548));
  AND2 AND2_1527(.VSS(VSS),.VDD(VDD),.Y(g8039),.A(g7587),.B(g5128));
  AND2 AND2_1528(.VSS(VSS),.VDD(VDD),.Y(g9610),.A(g925),.B(g9192));
  AND2 AND2_1529(.VSS(VSS),.VDD(VDD),.Y(g3536),.A(g2390),.B(g3103));
  AND2 AND2_1530(.VSS(VSS),.VDD(VDD),.Y(g5529),.A(g4129),.B(g4288));
  AND2 AND2_1531(.VSS(VSS),.VDD(VDD),.Y(g5148),.A(g3088),.B(g4671));
  AND2 AND2_1532(.VSS(VSS),.VDD(VDD),.Y(g9124),.A(g8881),.B(g4802));
  AND2 AND2_1533(.VSS(VSS),.VDD(VDD),.Y(g9324),.A(g8879),.B(g5708));
  AND2 AND2_1534(.VSS(VSS),.VDD(VDD),.Y(g4559),.A(g2034),.B(g3829));
  AND2 AND2_1535(.VSS(VSS),.VDD(VDD),.Y(g10561),.A(g10549),.B(g4583));
  AND2 AND2_1536(.VSS(VSS),.VDD(VDD),.Y(g5698),.A(g1571),.B(g5116));
  AND2 AND2_1537(.VSS(VSS),.VDD(VDD),.Y(g11226),.A(g461),.B(g11057));
  AND2 AND2_1538(.VSS(VSS),.VDD(VDD),.Y(g10295),.A(g8892),.B(g10208));
  AND2 AND2_1539(.VSS(VSS),.VDD(VDD),.Y(g5260),.A(g1092),.B(g4758));
  AND2 AND2_1540(.VSS(VSS),.VDD(VDD),.Y(g10680),.A(g10564),.B(g3586));
  AND2 AND2_1541(.VSS(VSS),.VDD(VDD),.Y(g6822),.A(g231),.B(g6596));
  AND2 AND2_1542(.VSS(VSS),.VDD(VDD),.Y(g4905),.A(g1853),.B(g4243));
  AND2 AND2_1543(.VSS(VSS),.VDD(VDD),.Y(g11551),.A(g11538),.B(g4013));
  AND2 AND2_1544(.VSS(VSS),.VDD(VDD),.Y(g3047),.A(g1227),.B(g2306));
  AND2 AND2_1545(.VSS(VSS),.VDD(VDD),.Y(g9849),.A(g293),.B(g9768));
  AND2 AND2_1546(.VSS(VSS),.VDD(VDD),.Y(g5279),.A(g1766),.B(g4783));
  AND2 AND2_1547(.VSS(VSS),.VDD(VDD),.Y(g8404),.A(g686),.B(g8129));
  AND2 AND2_1548(.VSS(VSS),.VDD(VDD),.Y(g5720),.A(g170),.B(g5361));
  AND2 AND2_1549(.VSS(VSS),.VDD(VDD),.Y(g5318),.A(g4401),.B(g1857));
  AND2 AND2_1550(.VSS(VSS),.VDD(VDD),.Y(g8764),.A(g7443),.B(g8684));
  AND2 AND2_1551(.VSS(VSS),.VDD(VDD),.Y(g11376),.A(g11318),.B(g4277));
  AND2 AND2_1552(.VSS(VSS),.VDD(VDD),.Y(g11297),.A(g5490),.B(g11242));
  AND2 AND2_1553(.VSS(VSS),.VDD(VDD),.Y(g9898),.A(g9887),.B(g9367));
//
  OR2 OR2_0(.VSS(VSS),.VDD(VDD),.Y(g6895),.A(g6776),.B(g4875));
  OR2 OR2_1(.VSS(VSS),.VDD(VDD),.Y(g7189),.A(g6632),.B(g6053));
  OR2 OR2_2(.VSS(VSS),.VDD(VDD),.Y(g9510),.A(g9125),.B(g9111));
  OR2 OR2_3(.VSS(VSS),.VDD(VDD),.Y(g7297),.A(g7132),.B(g6323));
  OR2 OR2_4(.VSS(VSS),.VDD(VDD),.Y(g9088),.A(g8927),.B(g8381));
  OR2 OR2_5(.VSS(VSS),.VDD(VDD),.Y(g9923),.A(g9865),.B(g9707));
  OR2 OR2_6(.VSS(VSS),.VDD(VDD),.Y(g6485),.A(g5848),.B(g5067));
  OR2 OR2_7(.VSS(VSS),.VDD(VDD),.Y(g8771),.A(g5483),.B(g8652));
  OR2 OR2_8(.VSS(VSS),.VDD(VDD),.Y(g5813),.A(g5617),.B(g4869));
  OR2 OR2_9(.VSS(VSS),.VDD(VDD),.Y(g7963),.A(g7687),.B(g7182));
  OR2 OR2_10(.VSS(VSS),.VDD(VDD),.Y(g10643),.A(g10624),.B(g7736));
  OR3 OR3_0(.VSS(VSS),.VDD(VDD),.Y(g9886),.A(g9607),.B(g9592),.C(g9759));
  OR3 OR3_1(.VSS(VSS),.VDD(VDD),.Y(g9951),.A(g9902),.B(g9899),.C(g9803));
  OR2 OR2_11(.VSS(VSS),.VDD(VDD),.Y(g11625),.A(g6535),.B(g11597));
  OR2 OR2_12(.VSS(VSS),.VDD(VDD),.Y(g8945),.A(g8801),.B(g8710));
  OR2 OR2_13(.VSS(VSS),.VDD(VDD),.Y(g10489),.A(g4961),.B(g10367));
  OR2 OR2_14(.VSS(VSS),.VDD(VDD),.Y(g10559),.A(g4141),.B(g10512));
  OR2 OR2_15(.VSS(VSS),.VDD(VDD),.Y(g10558),.A(g4126),.B(g10510));
  OR2 OR2_16(.VSS(VSS),.VDD(VDD),.Y(g11338),.A(g11283),.B(g11178));
  OR2 OR2_17(.VSS(VSS),.VDD(VDD),.Y(g8435),.A(g8403),.B(g8075));
  OR2 OR2_18(.VSS(VSS),.VDD(VDD),.Y(g10544),.A(g5511),.B(g10495));
  OR2 OR2_19(.VSS(VSS),.VDD(VDD),.Y(g6911),.A(g6342),.B(g5681));
  OR2 OR2_20(.VSS(VSS),.VDD(VDD),.Y(g10865),.A(g5538),.B(g10752));
  OR2 OR2_21(.VSS(VSS),.VDD(VDD),.Y(g3698),.A(g3121),.B(g2480));
  OR2 OR2_22(.VSS(VSS),.VDD(VDD),.Y(g8214),.A(g7472),.B(g8004));
  OR2 OR2_23(.VSS(VSS),.VDD(VDD),.Y(g6124),.A(g5181),.B(g5188));
  OR2 OR2_24(.VSS(VSS),.VDD(VDD),.Y(g6469),.A(g5698),.B(g4959));
  OR2 OR2_25(.VSS(VSS),.VDD(VDD),.Y(g5587),.A(g4714),.B(g3904));
  OR2 OR2_26(.VSS(VSS),.VDD(VDD),.Y(g6177),.A(g5444),.B(g4712));
  OR3 OR3_2(.VSS(VSS),.VDD(VDD),.Y(I14585),.A(g8995),.B(g9205),.C(g9192));
  OR2 OR2_27(.VSS(VSS),.VDD(VDD),.Y(g9891),.A(g9741),.B(g9760));
  OR2 OR2_28(.VSS(VSS),.VDD(VDD),.Y(g9913),.A(g9849),.B(g9691));
  OR4 OR4_0(.VSS(VSS),.VDD(VDD),.Y(I5600),.A(g496),.B(g491),.C(g486),.D(g481));
  OR2 OR2_29(.VSS(VSS),.VDD(VDD),.Y(g11257),.A(g11234),.B(g11019));
  OR2 OR2_30(.VSS(VSS),.VDD(VDD),.Y(g8236),.A(g7526),.B(g8001));
  OR2 OR2_31(.VSS(VSS),.VDD(VDD),.Y(g7385),.A(g7235),.B(g6746));
  OR2 OR2_32(.VSS(VSS),.VDD(VDD),.Y(g6898),.A(g6790),.B(g4881));
  OR2 OR2_33(.VSS(VSS),.VDD(VDD),.Y(g6900),.A(g6787),.B(g6246));
  OR2 OR2_34(.VSS(VSS),.VDD(VDD),.Y(g4264),.A(g4048),.B(g4053));
  OR3 OR3_3(.VSS(VSS),.VDD(VDD),.Y(g9726),.A(g9411),.B(g9420),.C(g9489));
  OR2 OR2_35(.VSS(VSS),.VDD(VDD),.Y(g6088),.A(g5260),.B(g4522));
  OR2 OR2_36(.VSS(VSS),.VDD(VDD),.Y(g6923),.A(g6353),.B(g5695));
  OR2 OR2_37(.VSS(VSS),.VDD(VDD),.Y(g8194),.A(g5168),.B(g7940));
  OR3 OR3_4(.VSS(VSS),.VDD(VDD),.Y(g9676),.A(g9454),.B(g9292),.C(g9274));
  OR2 OR2_38(.VSS(VSS),.VDD(VDD),.Y(g11256),.A(g11186),.B(g11018));
  OR2 OR2_39(.VSS(VSS),.VDD(VDD),.Y(g3860),.A(g3107),.B(g2167));
  OR2 OR2_40(.VSS(VSS),.VDD(VDD),.Y(g11280),.A(g11254),.B(g11153));
  OR4 OR4_1(.VSS(VSS),.VDD(VDD),.Y(g9727),.A(g9650),.B(g9663),.C(g9362),.D(I14866));
  OR2 OR2_41(.VSS(VSS),.VDD(VDD),.Y(g4997),.A(g4581),.B(g4584));
  OR2 OR2_42(.VSS(VSS),.VDD(VDD),.Y(g11624),.A(g11595),.B(g11571));
  OR2 OR2_43(.VSS(VSS),.VDD(VDD),.Y(g11300),.A(g11213),.B(g11091));
  OR2 OR2_44(.VSS(VSS),.VDD(VDD),.Y(g4238),.A(g3999),.B(g4007));
  OR2 OR2_45(.VSS(VSS),.VDD(VDD),.Y(g8814),.A(g7945),.B(g8728));
  OR2 OR2_46(.VSS(VSS),.VDD(VDD),.Y(g10401),.A(g9317),.B(g10291));
  OR2 OR2_47(.VSS(VSS),.VDD(VDD),.Y(g8773),.A(g5491),.B(g8653));
  OR2 OR2_48(.VSS(VSS),.VDD(VDD),.Y(g11231),.A(g11156),.B(g11013));
  OR2 OR2_49(.VSS(VSS),.VDD(VDD),.Y(g10864),.A(g5532),.B(g10751));
  OR2 OR2_50(.VSS(VSS),.VDD(VDD),.Y(g9624),.A(g9316),.B(g9313));
  OR3 OR3_5(.VSS(VSS),.VDD(VDD),.Y(g9953),.A(g9945),.B(g9939),.C(g9669));
  OR2 OR2_51(.VSS(VSS),.VDD(VDD),.Y(g6122),.A(g5172),.B(g5180));
  OR2 OR2_52(.VSS(VSS),.VDD(VDD),.Y(g6465),.A(g5825),.B(g5041));
  OR2 OR2_53(.VSS(VSS),.VDD(VDD),.Y(g6934),.A(g6363),.B(g5720));
  OR2 OR2_54(.VSS(VSS),.VDD(VDD),.Y(g7664),.A(g6855),.B(g4084));
  OR2 OR2_55(.VSS(VSS),.VDD(VDD),.Y(g7246),.A(g6465),.B(g6003));
  OR2 OR2_56(.VSS(VSS),.VDD(VDD),.Y(g7203),.A(g6640),.B(g6058));
  OR2 OR2_57(.VSS(VSS),.VDD(VDD),.Y(g6096),.A(g5268),.B(g4542));
  OR2 OR2_58(.VSS(VSS),.VDD(VDD),.Y(g9747),.A(g9173),.B(g9509));
  OR2 OR2_59(.VSS(VSS),.VDD(VDD),.Y(g11314),.A(g11224),.B(g11102));
  OR2 OR2_60(.VSS(VSS),.VDD(VDD),.Y(g10733),.A(g5227),.B(g10674));
  OR2 OR2_61(.VSS(VSS),.VDD(VDD),.Y(g8921),.A(g8827),.B(g8748));
  OR4 OR4_2(.VSS(VSS),.VDD(VDD),.Y(I15054),.A(g7853),.B(g9782),.C(g9624),.D(g9785));
  OR2 OR2_62(.VSS(VSS),.VDD(VDD),.Y(g11269),.A(g11196),.B(g11031));
  OR2 OR2_63(.VSS(VSS),.VDD(VDD),.Y(g5555),.A(g4389),.B(g4397));
  OR2 OR2_64(.VSS(VSS),.VDD(VDD),.Y(g11268),.A(g11194),.B(g11030));
  OR2 OR2_65(.VSS(VSS),.VDD(VDD),.Y(g10485),.A(g9317),.B(g10376));
  OR2 OR2_66(.VSS(VSS),.VDD(VDD),.Y(g10555),.A(g4103),.B(g10504));
  OR2 OR2_67(.VSS(VSS),.VDD(VDD),.Y(g6481),.A(g5722),.B(g4972));
  OR2 OR2_68(.VSS(VSS),.VDD(VDD),.Y(g10712),.A(g10662),.B(g9531));
  OR2 OR2_69(.VSS(VSS),.VDD(VDD),.Y(g11335),.A(g11279),.B(g11175));
  OR2 OR2_70(.VSS(VSS),.VDD(VDD),.Y(g8249),.A(g8018),.B(g7710));
  OR2 OR2_71(.VSS(VSS),.VDD(VDD),.Y(g7638),.A(g7265),.B(g6488));
  OR2 OR2_72(.VSS(VSS),.VDD(VDD),.Y(g10567),.A(g10514),.B(g7378));
  OR2 OR2_73(.VSS(VSS),.VDD(VDD),.Y(g11487),.A(g6662),.B(g11464));
  OR4 OR4_3(.VSS(VSS),.VDD(VDD),.Y(I15210),.A(g9839),.B(g9964),.C(g9852),.D(g9882));
  OR4 OR4_4(.VSS(VSS),.VDD(VDD),.Y(I5805),.A(g2102),.B(g2099),.C(g2096),.D(g2088));
  OR2 OR2_74(.VSS(VSS),.VDD(VDD),.Y(g8941),.A(g8796),.B(g8706));
  OR2 OR2_75(.VSS(VSS),.VDD(VDD),.Y(g11443),.A(g7130),.B(g11407));
  OR2 OR2_76(.VSS(VSS),.VDD(VDD),.Y(g4231),.A(g3991),.B(g3998));
  OR2 OR2_77(.VSS(VSS),.VDD(VDD),.Y(g11278),.A(g11253),.B(g11150));
  OR4 OR4_5(.VSS(VSS),.VDD(VDD),.Y(I15039),.A(g7853),.B(g9809),.C(g9624),.D(g9785));
  OR2 OR2_78(.VSS(VSS),.VDD(VDD),.Y(g11286),.A(g10670),.B(g11209));
  OR2 OR2_79(.VSS(VSS),.VDD(VDD),.Y(g8431),.A(g8387),.B(g8071));
  OR2 OR2_80(.VSS(VSS),.VDD(VDD),.Y(g7133),.A(g6616),.B(g3067));
  OR2 OR2_81(.VSS(VSS),.VDD(VDD),.Y(g11306),.A(g11216),.B(g11095));
  OR2 OR2_82(.VSS(VSS),.VDD(VDD),.Y(g8252),.A(g7988),.B(g7679));
  OR2 OR2_83(.VSS(VSS),.VDD(VDD),.Y(g8812),.A(g7939),.B(g8724));
  OR2 OR2_84(.VSS(VSS),.VDD(VDD),.Y(g7846),.A(g7722),.B(g7241));
  OR2 OR2_85(.VSS(VSS),.VDD(VDD),.Y(g3875),.A(g3275),.B(g12));
  OR2 OR2_86(.VSS(VSS),.VDD(VDD),.Y(g5996),.A(g5473),.B(g3908));
  OR2 OR2_87(.VSS(VSS),.VDD(VDD),.Y(g6592),.A(g5100),.B(g5882));
  OR2 OR2_88(.VSS(VSS),.VDD(VDD),.Y(g8286),.A(g8107),.B(g7823));
  OR2 OR2_89(.VSS(VSS),.VDD(VDD),.Y(g10501),.A(g4161),.B(g10445));
  OR2 OR2_90(.VSS(VSS),.VDD(VDD),.Y(g10728),.A(g4973),.B(g10642));
  OR2 OR2_91(.VSS(VSS),.VDD(VDD),.Y(g8270),.A(g7894),.B(g3434));
  OR2 OR2_92(.VSS(VSS),.VDD(VDD),.Y(g7290),.A(g7046),.B(g6316));
  OR2 OR2_93(.VSS(VSS),.VDD(VDD),.Y(g6068),.A(g5220),.B(g4497));
  OR2 OR2_94(.VSS(VSS),.VDD(VDD),.Y(g6468),.A(g5690),.B(g4950));
  OR2 OR2_95(.VSS(VSS),.VDD(VDD),.Y(g11217),.A(g11144),.B(g11005));
  OR2 OR2_96(.VSS(VSS),.VDD(VDD),.Y(g11478),.A(g6532),.B(g11455));
  OR4 OR4_6(.VSS(VSS),.VDD(VDD),.Y(g9536),.A(g9335),.B(g9331),.C(g9328),.D(g9324));
  OR2 OR2_97(.VSS(VSS),.VDD(VDD),.Y(g5981),.A(g5074),.B(g4383));
  OR2 OR2_98(.VSS(VSS),.VDD(VDD),.Y(g11486),.A(g6654),.B(g11463));
  OR2 OR2_99(.VSS(VSS),.VDD(VDD),.Y(g8377),.A(g8185),.B(g7958));
  OR2 OR2_100(.VSS(VSS),.VDD(VDD),.Y(g8206),.A(g7459),.B(g8007));
  OR2 OR2_101(.VSS(VSS),.VDD(VDD),.Y(g11580),.A(g11413),.B(g11544));
  OR2 OR2_102(.VSS(VSS),.VDD(VDD),.Y(g8287),.A(g8117),.B(g7824));
  OR2 OR2_103(.VSS(VSS),.VDD(VDD),.Y(g11223),.A(g11147),.B(g11008));
  OR2 OR2_104(.VSS(VSS),.VDD(VDD),.Y(g9522),.A(g9173),.B(g9125));
  OR2 OR2_105(.VSS(VSS),.VDD(VDD),.Y(g8199),.A(g7902),.B(g7444));
  OR2 OR2_106(.VSS(VSS),.VDD(VDD),.Y(g5802),.A(g5601),.B(g4837));
  OR2 OR2_107(.VSS(VSS),.VDD(VDD),.Y(g11321),.A(g11230),.B(g11105));
  OR2 OR2_108(.VSS(VSS),.VDD(VDD),.Y(g6524),.A(g5746),.B(g4996));
  OR2 OR2_109(.VSS(VSS),.VDD(VDD),.Y(g10664),.A(g10240),.B(g10582));
  OR2 OR2_110(.VSS(VSS),.VDD(VDD),.Y(g7257),.A(g6701),.B(g4725));
  OR2 OR2_111(.VSS(VSS),.VDD(VDD),.Y(g7301),.A(g7140),.B(g6327));
  OR2 OR2_112(.VSS(VSS),.VDD(VDD),.Y(g10484),.A(g9317),.B(g10400));
  OR2 OR2_113(.VSS(VSS),.VDD(VDD),.Y(g10554),.A(g4097),.B(g10503));
  OR2 OR2_114(.VSS(VSS),.VDD(VDD),.Y(g8259),.A(g8028),.B(g7719));
  OR2 OR2_115(.VSS(VSS),.VDD(VDD),.Y(g11334),.A(g11277),.B(g11174));
  OR2 OR2_116(.VSS(VSS),.VDD(VDD),.Y(g8819),.A(g7957),.B(g8734));
  OR2 OR2_117(.VSS(VSS),.VDD(VDD),.Y(g8923),.A(g8846),.B(g8763));
  OR2 OR2_118(.VSS(VSS),.VDD(VDD),.Y(g8488),.A(g3664),.B(g8390));
  OR2 OR2_119(.VSS(VSS),.VDD(VDD),.Y(g7441),.A(g7271),.B(g6789));
  OR2 OR2_120(.VSS(VSS),.VDD(VDD),.Y(g6026),.A(g5507),.B(g3970));
  OR2 OR2_121(.VSS(VSS),.VDD(VDD),.Y(g10799),.A(g6225),.B(g10769));
  OR2 OR2_122(.VSS(VSS),.VDD(VDD),.Y(g10798),.A(g6217),.B(g10768));
  OR2 OR2_123(.VSS(VSS),.VDD(VDD),.Y(g10805),.A(g10759),.B(g10760));
  OR2 OR2_124(.VSS(VSS),.VDD(VDD),.Y(g10732),.A(g4358),.B(g10661));
  OR2 OR2_125(.VSS(VSS),.VDD(VDD),.Y(g6061),.A(g5204),.B(g4));
  OR2 OR2_126(.VSS(VSS),.VDD(VDD),.Y(g9512),.A(g9151),.B(g9125));
  OR2 OR2_127(.VSS(VSS),.VDD(VDD),.Y(g10013),.A(I15214),.B(I15215));
  OR2 OR2_128(.VSS(VSS),.VDD(VDD),.Y(g8806),.A(g7931),.B(g8718));
  OR2 OR2_129(.VSS(VSS),.VDD(VDD),.Y(g8943),.A(g8837),.B(g8749));
  OR2 OR2_130(.VSS(VSS),.VDD(VDD),.Y(g11293),.A(g11211),.B(g10818));
  OR2 OR2_131(.VSS(VSS),.VDD(VDD),.Y(g11265),.A(g11189),.B(g11027));
  OR2 OR2_132(.VSS(VSS),.VDD(VDD),.Y(g8887),.A(g8842),.B(g8755));
  OR2 OR2_133(.VSS(VSS),.VDD(VDD),.Y(g5838),.A(g5612),.B(g4866));
  OR2 OR2_134(.VSS(VSS),.VDD(VDD),.Y(g6514),.A(g5738),.B(g4992));
  OR2 OR2_135(.VSS(VSS),.VDD(VDD),.Y(g8322),.A(g8136),.B(g6891));
  OR2 OR2_136(.VSS(VSS),.VDD(VDD),.Y(g8230),.A(g7515),.B(g7991));
  OR2 OR2_137(.VSS(VSS),.VDD(VDD),.Y(g5809),.A(g5611),.B(g4865));
  OR2 OR2_138(.VSS(VSS),.VDD(VDD),.Y(g8433),.A(g8399),.B(g8073));
  OR2 OR2_139(.VSS(VSS),.VDD(VDD),.Y(g11579),.A(g5123),.B(g11551));
  OR2 OR2_140(.VSS(VSS),.VDD(VDD),.Y(g10771),.A(g5533),.B(g10684));
  OR2 OR2_141(.VSS(VSS),.VDD(VDD),.Y(g11615),.A(g11601),.B(g11592));
  OR2 OR2_142(.VSS(VSS),.VDD(VDD),.Y(g9367),.A(g9335),.B(g9331));
  OR3 OR3_6(.VSS(VSS),.VDD(VDD),.Y(g9872),.A(g9617),.B(g9594),.C(g9750));
  OR2 OR2_143(.VSS(VSS),.VDD(VDD),.Y(g6522),.A(g5744),.B(g4994));
  OR2 OR2_144(.VSS(VSS),.VDD(VDD),.Y(g8266),.A(g7885),.B(g3412));
  OR2 OR2_145(.VSS(VSS),.VDD(VDD),.Y(g10414),.A(g10300),.B(g9534));
  OR2 OR2_146(.VSS(VSS),.VDD(VDD),.Y(g11275),.A(g11248),.B(g11148));
  OR2 OR2_147(.VSS(VSS),.VDD(VDD),.Y(g11430),.A(g11387),.B(g4006));
  OR2 OR2_148(.VSS(VSS),.VDD(VDD),.Y(g8248),.A(g8014),.B(g7707));
  OR3 OR3_7(.VSS(VSS),.VDD(VDD),.Y(g9686),.A(g9454),.B(g9292),.C(g9274));
  OR2 OR2_149(.VSS(VSS),.VDD(VDD),.Y(g8815),.A(g7948),.B(g8730));
  OR2 OR2_150(.VSS(VSS),.VDD(VDD),.Y(g7183),.A(g6623),.B(g6046));
  OR2 OR2_151(.VSS(VSS),.VDD(VDD),.Y(g5983),.A(g5084),.B(g4392));
  OR2 OR2_152(.VSS(VSS),.VDD(VDD),.Y(g8154),.A(g7891),.B(g6879));
  OR2 OR2_153(.VSS(VSS),.VDD(VDD),.Y(g6537),.A(g5781),.B(g5005));
  OR2 OR2_154(.VSS(VSS),.VDD(VDD),.Y(g4309),.A(g4069),.B(g4079));
  OR2 OR2_155(.VSS(VSS),.VDD(VDD),.Y(g10725),.A(g4962),.B(g10634));
  OR2 OR2_156(.VSS(VSS),.VDD(VDD),.Y(g6243),.A(g5537),.B(g4774));
  OR4 OR4_7(.VSS(VSS),.VDD(VDD),.Y(I6351),.A(g2405),.B(g2389),.C(g2380),.D(g2372));
  OR3 OR3_8(.VSS(VSS),.VDD(VDD),.Y(g9519),.A(g9173),.B(g9151),.C(g9125));
  OR2 OR2_157(.VSS(VSS),.VDD(VDD),.Y(g9740),.A(g9418),.B(g9505));
  OR2 OR2_158(.VSS(VSS),.VDD(VDD),.Y(g8267),.A(g7889),.B(g3422));
  OR3 OR3_9(.VSS(VSS),.VDD(VDD),.Y(g10744),.A(g10600),.B(g10668),.C(I16427));
  OR2 OR2_159(.VSS(VSS),.VDD(VDD),.Y(g6542),.A(g5789),.B(g5010));
  OR2 OR2_160(.VSS(VSS),.VDD(VDD),.Y(g7303),.A(g7145),.B(g6329));
  OR2 OR2_161(.VSS(VSS),.VDD(VDD),.Y(g10652),.A(g10627),.B(g7743));
  OR2 OR2_162(.VSS(VSS),.VDD(VDD),.Y(g5036),.A(g4871),.B(g4162));
  OR2 OR2_163(.VSS(VSS),.VDD(VDD),.Y(g7240),.A(g6687),.B(g6095));
  OR2 OR2_164(.VSS(VSS),.VDD(VDD),.Y(g8221),.A(g7496),.B(g7993));
  OR2 OR2_165(.VSS(VSS),.VDD(VDD),.Y(g6902),.A(g6794),.B(g4223));
  OR3 OR3_10(.VSS(VSS),.VDD(VDD),.Y(I14776),.A(g8995),.B(g9205),.C(g9192));
  OR2 OR2_166(.VSS(VSS),.VDD(VDD),.Y(g10500),.A(g4157),.B(g10442));
  OR2 OR2_167(.VSS(VSS),.VDD(VDD),.Y(g4052),.A(g2862),.B(g2515));
  OR4 OR4_8(.VSS(VSS),.VDD(VDD),.Y(I14858),.A(g9585),.B(g9595),.C(g9610),.D(g9602));
  OR2 OR2_168(.VSS(VSS),.VDD(VDD),.Y(g6529),.A(g5757),.B(g5000));
  OR2 OR2_169(.VSS(VSS),.VDD(VDD),.Y(g11264),.A(g11188),.B(g11026));
  OR4 OR4_9(.VSS(VSS),.VDD(VDD),.Y(I15209),.A(g8169),.B(g9905),.C(g9934),.D(g9830));
  OR2 OR2_170(.VSS(VSS),.VDD(VDD),.Y(g8241),.A(g7536),.B(g7989));
  OR2 OR2_171(.VSS(VSS),.VDD(VDD),.Y(g10795),.A(g6199),.B(g10764));
  OR2 OR2_172(.VSS(VSS),.VDD(VDD),.Y(g11607),.A(g11586),.B(g11557));
  OR2 OR2_173(.VSS(VSS),.VDD(VDD),.Y(g8644),.A(g8123),.B(g8464));
  OR3 OR3_11(.VSS(VSS),.VDD(VDD),.Y(g4682),.A(g3563),.B(g3348),.C(g1570));
  OR2 OR2_174(.VSS(VSS),.VDD(VDD),.Y(g8818),.A(g7955),.B(g8733));
  OR2 OR2_175(.VSS(VSS),.VDD(VDD),.Y(g2984),.A(g2528),.B(g2522));
  OR2 OR2_176(.VSS(VSS),.VDD(VDD),.Y(g9931),.A(g8931),.B(g9900));
  OR2 OR2_177(.VSS(VSS),.VDD(VDD),.Y(g3414),.A(g2911),.B(g2917));
  OR2 OR2_178(.VSS(VSS),.VDD(VDD),.Y(g9515),.A(g9173),.B(g9151));
  OR2 OR2_179(.VSS(VSS),.VDD(VDD),.Y(g10724),.A(g10312),.B(g10672));
  OR2 OR2_180(.VSS(VSS),.VDD(VDD),.Y(g7294),.A(g7068),.B(g6320));
  OR2 OR2_181(.VSS(VSS),.VDD(VDD),.Y(g5189),.A(g4345),.B(g3496));
  OR2 OR2_182(.VSS(VSS),.VDD(VDD),.Y(g8614),.A(g8365),.B(g8510));
  OR2 OR2_183(.VSS(VSS),.VDD(VDD),.Y(g3513),.A(g3118),.B(g2180));
  OR2 OR2_184(.VSS(VSS),.VDD(VDD),.Y(g6909),.A(g6346),.B(g5684));
  OR4 OR4_10(.VSS(VSS),.VDD(VDD),.Y(I5571),.A(g396),.B(g391),.C(g386),.D(g426));
  OR2 OR2_185(.VSS(VSS),.VDD(VDD),.Y(g4283),.A(g4059),.B(g4063));
  OR2 OR2_186(.VSS(VSS),.VDD(VDD),.Y(g8939),.A(g8791),.B(g8701));
  OR2 OR2_187(.VSS(VSS),.VDD(VDD),.Y(g2514),.A(I5599),.B(I5600));
  OR2 OR2_188(.VSS(VSS),.VDD(VDD),.Y(g11327),.A(g11297),.B(g11167));
  OR2 OR2_189(.VSS(VSS),.VDD(VDD),.Y(g8187),.A(g7542),.B(g7998));
  OR2 OR2_190(.VSS(VSS),.VDD(VDD),.Y(g11606),.A(g11585),.B(g11556));
  OR2 OR2_191(.VSS(VSS),.VDD(VDD),.Y(g11303),.A(g11214),.B(g11092));
  OR2 OR2_192(.VSS(VSS),.VDD(VDD),.Y(g5309),.A(g3664),.B(g4401));
  OR3 OR3_12(.VSS(VSS),.VDD(VDD),.Y(g9528),.A(g9151),.B(g9125),.C(g9111));
  OR2 OR2_193(.VSS(VSS),.VDD(VDD),.Y(g8200),.A(g7535),.B(g8008));
  OR3 OR3_13(.VSS(VSS),.VDD(VDD),.Y(g2522),.A(g833),.B(g829),.C(I5629));
  OR4 OR4_11(.VSS(VSS),.VDD(VDD),.Y(g2315),.A(g1163),.B(g1166),.C(g1113),.D(I5363));
  OR2 OR2_194(.VSS(VSS),.VDD(VDD),.Y(g6506),.A(g5731),.B(g4989));
  OR2 OR2_195(.VSS(VSS),.VDD(VDD),.Y(g10649),.A(g10626),.B(g7741));
  OR2 OR2_196(.VSS(VSS),.VDD(VDD),.Y(g8159),.A(g7895),.B(g6886));
  OR2 OR2_197(.VSS(VSS),.VDD(VDD),.Y(g7626),.A(g7060),.B(g5267));
  OR2 OR2_198(.VSS(VSS),.VDD(VDD),.Y(g10770),.A(g5525),.B(g10682));
  OR2 OR2_199(.VSS(VSS),.VDD(VDD),.Y(g9566),.A(g9052),.B(g9030));
  OR2 OR2_200(.VSS(VSS),.VDD(VDD),.Y(g11483),.A(g6633),.B(g11460));
  OR2 OR2_201(.VSS(VSS),.VDD(VDD),.Y(g8811),.A(g7935),.B(g8722));
  OR3 OR3_14(.VSS(VSS),.VDD(VDD),.Y(g8642),.A(g5236),.B(g5205),.C(g8465));
  OR2 OR2_202(.VSS(VSS),.VDD(VDD),.Y(g6545),.A(g5795),.B(g5025));
  OR2 OR2_203(.VSS(VSS),.VDD(VDD),.Y(g10767),.A(g5500),.B(g10681));
  OR2 OR2_204(.VSS(VSS),.VDD(VDD),.Y(g11326),.A(g11296),.B(g11166));
  OR2 OR2_205(.VSS(VSS),.VDD(VDD),.Y(g10898),.A(g4220),.B(g10777));
  OR2 OR2_206(.VSS(VSS),.VDD(VDD),.Y(g11252),.A(g11099),.B(g10969));
  OR2 OR2_207(.VSS(VSS),.VDD(VDD),.Y(g10719),.A(g10303),.B(g10666));
  OR2 OR2_208(.VSS(VSS),.VDD(VDD),.Y(g4609),.A(g3400),.B(g119));
  OR2 OR2_209(.VSS(VSS),.VDD(VDD),.Y(g6507),.A(g5732),.B(g4990));
  OR2 OR2_210(.VSS(VSS),.VDD(VDD),.Y(g10718),.A(g6238),.B(g10706));
  OR2 OR2_211(.VSS(VSS),.VDD(VDD),.Y(g10521),.A(I16148),.B(I16149));
  OR2 OR2_212(.VSS(VSS),.VDD(VDD),.Y(g7075),.A(g5104),.B(g6530));
  OR2 OR2_213(.VSS(VSS),.VDD(VDD),.Y(g7292),.A(g7055),.B(g6318));
  OR2 OR2_214(.VSS(VSS),.VDD(VDD),.Y(g10861),.A(g5523),.B(g10745));
  OR2 OR2_215(.VSS(VSS),.VDD(VDD),.Y(g8417),.A(g8246),.B(g7721));
  OR2 OR2_216(.VSS(VSS),.VDD(VDD),.Y(g6515),.A(g5739),.B(g4993));
  OR4 OR4_12(.VSS(VSS),.VDD(VDD),.Y(I14855),.A(g9583),.B(g9593),.C(g9601),.D(g9596));
  OR4 OR4_13(.VSS(VSS),.VDD(VDD),.Y(I15205),.A(g9838),.B(g9963),.C(g9850),.D(g9878));
  OR4 OR4_14(.VSS(VSS),.VDD(VDD),.Y(I15051),.A(g7853),.B(g9673),.C(g9624),.D(g9785));
  OR3 OR3_15(.VSS(VSS),.VDD(VDD),.Y(g9724),.A(g9409),.B(g9419),.C(g9615));
  OR2 OR2_217(.VSS(VSS),.VDD(VDD),.Y(g6528),.A(g5756),.B(g4999));
  OR2 OR2_218(.VSS(VSS),.VDD(VDD),.Y(g8823),.A(g8778),.B(g8693));
  OR2 OR2_219(.VSS(VSS),.VDD(VDD),.Y(g7503),.A(g6887),.B(g6430));
  OR2 OR2_220(.VSS(VSS),.VDD(VDD),.Y(g8148),.A(g7884),.B(g6872));
  OR2 OR2_221(.VSS(VSS),.VDD(VDD),.Y(g8649),.A(g8499),.B(g4519));
  OR2 OR2_222(.VSS(VSS),.VDD(VDD),.Y(g3584),.A(g2863),.B(g2516));
  OR2 OR2_223(.VSS(VSS),.VDD(VDD),.Y(g10776),.A(g5544),.B(g10758));
  OR3 OR3_16(.VSS(VSS),.VDD(VDD),.Y(g9680),.A(g9454),.B(g9292),.C(g9274));
  OR2 OR2_224(.VSS(VSS),.VDD(VDD),.Y(g10859),.A(g5512),.B(g10742));
  OR3 OR3_17(.VSS(VSS),.VDD(VDD),.Y(I14866),.A(g9590),.B(g9609),.C(g9619));
  OR2 OR2_225(.VSS(VSS),.VDD(VDD),.Y(g7299),.A(g7138),.B(g6325));
  OR2 OR2_226(.VSS(VSS),.VDD(VDD),.Y(g10858),.A(g5501),.B(g10741));
  OR2 OR2_227(.VSS(VSS),.VDD(VDD),.Y(g8193),.A(g5145),.B(g7937));
  OR3 OR3_18(.VSS(VSS),.VDD(VDD),.Y(g9511),.A(g9151),.B(g9125),.C(g9111));
  OR2 OR2_228(.VSS(VSS),.VDD(VDD),.Y(g7738),.A(g7200),.B(g6738));
  OR2 OR2_229(.VSS(VSS),.VDD(VDD),.Y(g7244),.A(g6699),.B(g4720));
  OR2 OR2_230(.VSS(VSS),.VDD(VDD),.Y(g3425),.A(g2895),.B(g2910));
  OR2 OR2_231(.VSS(VSS),.VDD(VDD),.Y(g7478),.A(g6884),.B(g6423));
  OR3 OR3_19(.VSS(VSS),.VDD(VDD),.Y(g9714),.A(g9664),.B(g9366),.C(g9654));
  OR2 OR2_232(.VSS(VSS),.VDD(VDD),.Y(g10025),.A(I15224),.B(I15225));
  OR2 OR2_233(.VSS(VSS),.VDD(VDD),.Y(g6908),.A(g6345),.B(g4229));
  OR2 OR2_234(.VSS(VSS),.VDD(VDD),.Y(g5028),.A(g4836),.B(g4128));
  OR2 OR2_235(.VSS(VSS),.VDD(VDD),.Y(g8253),.A(g8023),.B(g7718));
  OR2 OR2_236(.VSS(VSS),.VDD(VDD),.Y(g8938),.A(g8789),.B(g8699));
  OR2 OR2_237(.VSS(VSS),.VDD(VDD),.Y(g8813),.A(g7943),.B(g8726));
  OR2 OR2_238(.VSS(VSS),.VDD(VDD),.Y(g9736),.A(g9430),.B(g9416));
  OR2 OR2_239(.VSS(VSS),.VDD(VDD),.Y(g9968),.A(I15171),.B(I15172));
  OR2 OR2_240(.VSS(VSS),.VDD(VDD),.Y(g8552),.A(g8217),.B(g8388));
  OR2 OR2_241(.VSS(VSS),.VDD(VDD),.Y(g5910),.A(g5023),.B(g4341));
  OR2 OR2_242(.VSS(VSS),.VDD(VDD),.Y(g11249),.A(g6162),.B(g11143));
  OR2 OR2_243(.VSS(VSS),.VDD(VDD),.Y(g11482),.A(g6628),.B(g11459));
  OR4 OR4_15(.VSS(VSS),.VDD(VDD),.Y(g9722),.A(g9612),.B(g9643),.C(g9410),.D(I14855));
  OR4 OR4_16(.VSS(VSS),.VDD(VDD),.Y(I15204),.A(g8168),.B(g9904),.C(g9933),.D(g9829));
  OR2 OR2_244(.VSS(VSS),.VDD(VDD),.Y(g7236),.A(g6684),.B(g6092));
  OR3 OR3_20(.VSS(VSS),.VDD(VDD),.Y(I14596),.A(g8995),.B(g9205),.C(g9192));
  OR2 OR2_245(.VSS(VSS),.VDD(VDD),.Y(g8645),.A(g8127),.B(g8469));
  OR2 OR2_246(.VSS(VSS),.VDD(VDD),.Y(g11647),.A(g6622),.B(g11637));
  OR2 OR2_247(.VSS(VSS),.VDD(VDD),.Y(g6777),.A(g5691),.B(g5052));
  OR3 OR3_21(.VSS(VSS),.VDD(VDD),.Y(g9737),.A(g9657),.B(g9658),.C(g9655));
  OR4 OR4_17(.VSS(VSS),.VDD(VDD),.Y(I16149),.A(g10472),.B(g10470),.C(g10468),.D(g10467));
  OR2 OR2_248(.VSS(VSS),.VDD(VDD),.Y(g11233),.A(g11085),.B(g10946));
  OR2 OR2_249(.VSS(VSS),.VDD(VDD),.Y(g8607),.A(g8406),.B(g8554));
  OR4 OR4_18(.VSS(VSS),.VDD(VDD),.Y(I16148),.A(g10386),.B(g10384),.C(g10476),.D(g10474));
  OR2 OR2_250(.VSS(VSS),.VDD(VDD),.Y(g8158),.A(g7893),.B(g6883));
  OR2 OR2_251(.VSS(VSS),.VDD(VDD),.Y(g5846),.A(g4932),.B(g4236));
  OR2 OR2_252(.VSS(VSS),.VDD(VDD),.Y(g5396),.A(g4481),.B(g3684));
  OR2 OR2_253(.VSS(VSS),.VDD(VDD),.Y(g5803),.A(g5575),.B(g4820));
  OR2 OR2_254(.VSS(VSS),.VDD(VDD),.Y(g11331),.A(g11272),.B(g11171));
  OR2 OR2_255(.VSS(VSS),.VDD(VDD),.Y(g7295),.A(g7071),.B(g6321));
  OR2 OR2_256(.VSS(VSS),.VDD(VDD),.Y(g6541),.A(g5788),.B(g5009));
  OR2 OR2_257(.VSS(VSS),.VDD(VDD),.Y(g8615),.A(g8413),.B(g8557));
  OR2 OR2_258(.VSS(VSS),.VDD(VDD),.Y(g9742),.A(g9173),.B(g9528));
  OR2 OR2_259(.VSS(VSS),.VDD(VDD),.Y(g9926),.A(g9868),.B(g9715));
  OR2 OR2_260(.VSS(VSS),.VDD(VDD),.Y(g9754),.A(g9173),.B(g9511));
  OR2 OR2_261(.VSS(VSS),.VDD(VDD),.Y(g8284),.A(g8102),.B(g7821));
  OR2 OR2_262(.VSS(VSS),.VDD(VDD),.Y(g2204),.A(g1393),.B(g1394));
  OR2 OR2_263(.VSS(VSS),.VDD(VDD),.Y(g7471),.A(g6880),.B(g6416));
  OR2 OR2_264(.VSS(VSS),.VDD(VDD),.Y(g7242),.A(g6693),.B(g6098));
  OR2 OR2_265(.VSS(VSS),.VDD(VDD),.Y(g5847),.A(g5626),.B(g4877));
  OR2 OR2_266(.VSS(VSS),.VDD(VDD),.Y(g6901),.A(g6788),.B(g6247));
  OR2 OR2_267(.VSS(VSS),.VDD(VDD),.Y(g8559),.A(g8380),.B(g4731));
  OR3 OR3_22(.VSS(VSS),.VDD(VDD),.Y(g9729),.A(g9618),.B(g9357),.C(g9656));
  OR2 OR2_268(.VSS(VSS),.VDD(VDD),.Y(g10860),.A(g5513),.B(g10743));
  OR2 OR2_269(.VSS(VSS),.VDD(VDD),.Y(g9927),.A(g9869),.B(g9716));
  OR2 OR2_270(.VSS(VSS),.VDD(VDD),.Y(g10497),.A(g5052),.B(g10396));
  OR4 OR4_19(.VSS(VSS),.VDD(VDD),.Y(g9885),.A(g9739),.B(g9598),.C(g9662),.D(g9746));
  OR4 OR4_20(.VSS(VSS),.VDD(VDD),.Y(g2528),.A(g861),.B(g857),.C(g853),.D(g849));
  OR2 OR2_271(.VSS(VSS),.VDD(VDD),.Y(g11229),.A(g11154),.B(g11012));
  OR2 OR2_272(.VSS(VSS),.VDD(VDD),.Y(g8973),.A(g8821),.B(g8735));
  OR2 OR2_273(.VSS(VSS),.VDD(VDD),.Y(g10658),.A(g10595),.B(g7674));
  OR2 OR2_274(.VSS(VSS),.VDD(VDD),.Y(g10339),.A(g10232),.B(g9556));
  OR4 OR4_21(.VSS(VSS),.VDD(VDD),.Y(I5363),.A(g1149),.B(g1153),.C(g1157),.D(g1160));
  OR2 OR2_275(.VSS(VSS),.VDD(VDD),.Y(g11310),.A(g11220),.B(g11100));
  OR2 OR2_276(.VSS(VSS),.VDD(VDD),.Y(g6500),.A(g5725),.B(g4986));
  OR2 OR2_277(.VSS(VSS),.VDD(VDD),.Y(g10855),.A(g6075),.B(g10736));
  OR2 OR2_278(.VSS(VSS),.VDD(VDD),.Y(g9916),.A(g9855),.B(g9694));
  OR2 OR2_279(.VSS(VSS),.VDD(VDD),.Y(g10411),.A(g10299),.B(g9529));
  OR2 OR2_280(.VSS(VSS),.VDD(VDD),.Y(g11603),.A(g11582),.B(g11553));
  OR4 OR4_22(.VSS(VSS),.VDD(VDD),.Y(I5357),.A(g1265),.B(g1260),.C(g1255),.D(g1250));
  OR2 OR2_281(.VSS(VSS),.VDD(VDD),.Y(g9560),.A(g9052),.B(g9030));
  OR2 OR2_282(.VSS(VSS),.VDD(VDD),.Y(g6672),.A(g5941),.B(g5259));
  OR3 OR3_23(.VSS(VSS),.VDD(VDD),.Y(g9873),.A(g9623),.B(g9599),.C(g9758));
  OR2 OR2_283(.VSS(VSS),.VDD(VDD),.Y(g6523),.A(g5745),.B(g4995));
  OR2 OR2_284(.VSS(VSS),.VDD(VDD),.Y(g10707),.A(g5545),.B(g10686));
  OR4 OR4_23(.VSS(VSS),.VDD(VDD),.Y(I5626),.A(g521),.B(g525),.C(g530),.D(g534));
  OR2 OR2_285(.VSS(VSS),.VDD(VDD),.Y(g9579),.A(g9052),.B(g9030));
  OR2 OR2_286(.VSS(VSS),.VDD(VDD),.Y(g7298),.A(g7136),.B(g6324));
  OR2 OR2_287(.VSS(VSS),.VDD(VDD),.Y(g6551),.A(g5804),.B(g5031));
  OR2 OR2_288(.VSS(VSS),.VDD(VDD),.Y(g6099),.A(g5273),.B(g4550));
  OR2 OR2_289(.VSS(VSS),.VDD(VDD),.Y(g8282),.A(g8101),.B(g7819));
  OR2 OR2_290(.VSS(VSS),.VDD(VDD),.Y(g9917),.A(g9856),.B(g9695));
  OR4 OR4_24(.VSS(VSS),.VDD(VDD),.Y(I15057),.A(g7853),.B(g9680),.C(g9624),.D(g9785));
  OR2 OR2_291(.VSS(VSS),.VDD(VDD),.Y(g7219),.A(g6661),.B(g6076));
  OR2 OR2_292(.VSS(VSS),.VDD(VDD),.Y(g10019),.A(I15219),.B(I15220));
  OR2 OR2_293(.VSS(VSS),.VDD(VDD),.Y(g5857),.A(g5418),.B(g4670));
  OR4 OR4_25(.VSS(VSS),.VDD(VDD),.Y(g9725),.A(g9642),.B(g9659),.C(g9616),.D(I14862));
  OR2 OR2_294(.VSS(VSS),.VDD(VDD),.Y(g11298),.A(g11212),.B(g11087));
  OR2 OR2_295(.VSS(VSS),.VDD(VDD),.Y(g10402),.A(g10295),.B(g9554));
  OR4 OR4_26(.VSS(VSS),.VDD(VDD),.Y(g2521),.A(g538),.B(g542),.C(g476),.D(I5626));
  OR3 OR3_24(.VSS(VSS),.VDD(VDD),.Y(I14751),.A(g8995),.B(g9205),.C(g9192));
  OR2 OR2_296(.VSS(VSS),.VDD(VDD),.Y(g10866),.A(g5539),.B(g10753));
  OR2 OR2_297(.VSS(VSS),.VDD(VDD),.Y(g6534),.A(g5772),.B(g5003));
  OR2 OR2_298(.VSS(VSS),.VDD(VDD),.Y(g11232),.A(g11158),.B(g11015));
  OR3 OR3_25(.VSS(VSS),.VDD(VDD),.Y(g9706),.A(g9644),.B(g9386),.C(g9591));
  OR2 OR2_299(.VSS(VSS),.VDD(VDD),.Y(g10001),.A(I15204),.B(I15205));
  OR2 OR2_300(.VSS(VSS),.VDD(VDD),.Y(g8776),.A(g5510),.B(g8655));
  OR2 OR2_301(.VSS(VSS),.VDD(VDD),.Y(g7225),.A(g6666),.B(g6079));
  OR3 OR3_26(.VSS(VSS),.VDD(VDD),.Y(g9888),.A(g9648),.B(g9608),.C(g9757));
  OR2 OR2_302(.VSS(VSS),.VDD(VDD),.Y(g11261),.A(g11238),.B(g11023));
  OR3 OR3_27(.VSS(VSS),.VDD(VDD),.Y(g9956),.A(g9948),.B(g9942),.C(g9815));
  OR2 OR2_303(.VSS(VSS),.VDD(VDD),.Y(g10923),.A(g10778),.B(g10715));
  OR2 OR2_304(.VSS(VSS),.VDD(VDD),.Y(g8264),.A(g7879),.B(g3389));
  OR2 OR2_305(.VSS(VSS),.VDD(VDD),.Y(g6513),.A(g5737),.B(g4991));
  OR3 OR3_28(.VSS(VSS),.VDD(VDD),.Y(I14835),.A(g9621),.B(g9645),.C(g9588));
  OR2 OR2_306(.VSS(VSS),.VDD(VDD),.Y(g8641),.A(g8120),.B(g8463));
  OR3 OR3_29(.VSS(VSS),.VDD(VDD),.Y(g5361),.A(g4316),.B(g4093),.C(g126));
  OR2 OR2_307(.VSS(VSS),.VDD(VDD),.Y(g11316),.A(g11226),.B(g11103));
  OR4 OR4_27(.VSS(VSS),.VDD(VDD),.Y(I16161),.A(g10479),.B(g10478),.C(g10477),.D(g10475));
  OR2 OR2_308(.VSS(VSS),.VDD(VDD),.Y(g6916),.A(g6348),.B(g5687));
  OR2 OR2_309(.VSS(VSS),.VDD(VDD),.Y(g8777),.A(g5522),.B(g8659));
  OR4 OR4_28(.VSS(VSS),.VDD(VDD),.Y(g2353),.A(g1403),.B(g1407),.C(g1411),.D(g1415));
  OR2 OR2_310(.VSS(VSS),.VDD(VDD),.Y(g7510),.A(g7186),.B(g6730));
  OR3 OR3_30(.VSS(VSS),.VDD(VDD),.Y(g9957),.A(g9949),.B(g9943),.C(g9776));
  OR2 OR2_311(.VSS(VSS),.VDD(VDD),.Y(g2744),.A(I5804),.B(I5805));
  OR2 OR2_312(.VSS(VSS),.VDD(VDD),.Y(g7245),.A(g6696),.B(g6102));
  OR2 OR2_313(.VSS(VSS),.VDD(VDD),.Y(g7291),.A(g7050),.B(g6317));
  OR2 OR2_314(.VSS(VSS),.VDD(VDD),.Y(g8611),.A(g8410),.B(g8556));
  OR4 OR4_29(.VSS(VSS),.VDD(VDD),.Y(I15199),.A(g8167),.B(g9903),.C(g9932),.D(g9828));
  OR2 OR2_315(.VSS(VSS),.VDD(VDD),.Y(g10550),.A(g4942),.B(g10450));
  OR2 OR2_316(.VSS(VSS),.VDD(VDD),.Y(g11330),.A(g11304),.B(g11170));
  OR2 OR2_317(.VSS(VSS),.VDD(VDD),.Y(g10721),.A(g10306),.B(g10669));
  OR2 OR2_318(.VSS(VSS),.VDD(VDD),.Y(g8153),.A(g7888),.B(g6875));
  OR2 OR2_319(.VSS(VSS),.VDD(VDD),.Y(g10773),.A(g5540),.B(g10685));
  OR2 OR2_320(.VSS(VSS),.VDD(VDD),.Y(g3688),.A(g3144),.B(g2454));
  OR4 OR4_30(.VSS(VSS),.VDD(VDD),.Y(I15225),.A(g9842),.B(g9967),.C(g9859),.D(g9881));
  OR2 OR2_321(.VSS(VSS),.VDD(VDD),.Y(g6042),.A(g5535),.B(g3987));
  OR2 OR2_322(.VSS(VSS),.VDD(VDD),.Y(g10655),.A(g10561),.B(g7389));
  OR2 OR2_323(.VSS(VSS),.VDD(VDD),.Y(g11259),.A(g11236),.B(g11021));
  OR2 OR2_324(.VSS(VSS),.VDD(VDD),.Y(g11225),.A(g11149),.B(g11009));
  OR2 OR2_325(.VSS(VSS),.VDD(VDD),.Y(g5914),.A(g5029),.B(g4343));
  OR2 OR2_326(.VSS(VSS),.VDD(VDD),.Y(g11258),.A(g11235),.B(g11020));
  OR2 OR2_327(.VSS(VSS),.VDD(VDD),.Y(g6054),.A(g5199),.B(g4483));
  OR3 OR3_31(.VSS(VSS),.VDD(VDD),.Y(g9728),.A(g9412),.B(g9422),.C(g9426));
  OR3 OR3_32(.VSS(VSS),.VDD(VDD),.Y(g9730),.A(g9414),.B(g9425),.C(g9423));
  OR2 OR2_328(.VSS(VSS),.VDD(VDD),.Y(g5820),.A(g5595),.B(g4834));
  OR3 OR3_33(.VSS(VSS),.VDD(VDD),.Y(g8574),.A(g5679),.B(g7853),.C(g8465));
  OR2 OR2_329(.VSS(VSS),.VDD(VDD),.Y(g11602),.A(g11581),.B(g11552));
  OR2 OR2_330(.VSS(VSS),.VDD(VDD),.Y(g10502),.A(g4169),.B(g10365));
  OR2 OR2_331(.VSS(VSS),.VDD(VDD),.Y(g10557),.A(g4123),.B(g10508));
  OR4 OR4_31(.VSS(VSS),.VDD(VDD),.Y(I15171),.A(g8175),.B(g9909),.C(g9896),.D(g9835));
  OR2 OR2_332(.VSS(VSS),.VDD(VDD),.Y(g11337),.A(g11282),.B(g11177));
  OR2 OR2_333(.VSS(VSS),.VDD(VDD),.Y(g7465),.A(g6876),.B(g6410));
  OR2 OR2_334(.VSS(VSS),.VDD(VDD),.Y(g8262),.A(g7970),.B(g7625));
  OR2 OR2_335(.VSS(VSS),.VDD(VDD),.Y(g8889),.A(g8844),.B(g8756));
  OR2 OR2_336(.VSS(VSS),.VDD(VDD),.Y(g7096),.A(g6544),.B(g5911));
  OR2 OR2_337(.VSS(VSS),.VDD(VDD),.Y(g5995),.A(g5097),.B(g5099));
  OR2 OR2_338(.VSS(VSS),.VDD(VDD),.Y(g8285),.A(g8104),.B(g7822));
  OR2 OR2_339(.VSS(VSS),.VDD(VDD),.Y(g10791),.A(g6186),.B(g10762));
  OR2 OR2_340(.VSS(VSS),.VDD(VDD),.Y(g2499),.A(I5570),.B(I5571));
  OR3 OR3_34(.VSS(VSS),.VDD(VDD),.Y(I14607),.A(g8995),.B(g9205),.C(g9192));
  OR2 OR2_341(.VSS(VSS),.VDD(VDD),.Y(g6049),.A(g5254),.B(g3718));
  OR2 OR2_342(.VSS(VSS),.VDD(VDD),.Y(g9920),.A(g9860),.B(g9701));
  OR2 OR2_343(.VSS(VSS),.VDD(VDD),.Y(g10556),.A(g4115),.B(g10506));
  OR2 OR2_344(.VSS(VSS),.VDD(VDD),.Y(g8643),.A(g8364),.B(g8508));
  OR2 OR2_345(.VSS(VSS),.VDD(VDD),.Y(g5810),.A(g5588),.B(g4823));
  OR2 OR2_346(.VSS(VSS),.VDD(VDD),.Y(g11336),.A(g11281),.B(g11176));
  OR2 OR2_347(.VSS(VSS),.VDD(VDD),.Y(g8742),.A(g8135),.B(g8598));
  OR2 OR2_348(.VSS(VSS),.VDD(VDD),.Y(g8926),.A(g8848),.B(g8764));
  OR2 OR2_349(.VSS(VSS),.VDD(VDD),.Y(g7218),.A(g6655),.B(g6070));
  OR4 OR4_32(.VSS(VSS),.VDD(VDD),.Y(I15224),.A(g8174),.B(g9908),.C(g9937),.D(g9834));
  OR2 OR2_350(.VSS(VSS),.VDD(VDD),.Y(g7293),.A(g7063),.B(g6319));
  OR2 OR2_351(.VSS(VSS),.VDD(VDD),.Y(g11288),.A(g11204),.B(g11070));
  OR2 OR2_352(.VSS(VSS),.VDD(VDD),.Y(g10800),.A(g6245),.B(g10772));
  OR2 OR2_353(.VSS(VSS),.VDD(VDD),.Y(g11308),.A(g11218),.B(g11098));
  OR2 OR2_354(.VSS(VSS),.VDD(VDD),.Y(g8269),.A(g7892),.B(g3429));
  OR2 OR2_355(.VSS(VSS),.VDD(VDD),.Y(g10417),.A(g10301),.B(g9527));
  OR2 OR2_356(.VSS(VSS),.VDD(VDD),.Y(g10936),.A(g5170),.B(g10808));
  OR2 OR2_357(.VSS(VSS),.VDD(VDD),.Y(g9388),.A(g9240),.B(g9223));
  OR2 OR2_358(.VSS(VSS),.VDD(VDD),.Y(g6185),.A(g5470),.B(g4715));
  OR2 OR2_359(.VSS(VSS),.VDD(VDD),.Y(g6470),.A(g5699),.B(g4960));
  OR2 OR2_360(.VSS(VSS),.VDD(VDD),.Y(g6897),.A(g6771),.B(g6240));
  OR2 OR2_361(.VSS(VSS),.VDD(VDD),.Y(g8885),.A(g8841),.B(g8754));
  OR2 OR2_362(.VSS(VSS),.VDD(VDD),.Y(g11260),.A(g11237),.B(g11022));
  OR2 OR2_363(.VSS(VSS),.VDD(VDD),.Y(g11488),.A(g6671),.B(g11465));
  OR2 OR2_364(.VSS(VSS),.VDD(VDD),.Y(g6105),.A(g5279),.B(g4559));
  OR2 OR2_365(.VSS(VSS),.VDD(VDD),.Y(g10807),.A(g10701),.B(g10761));
  OR2 OR2_366(.VSS(VSS),.VDD(VDD),.Y(g10639),.A(g10623),.B(g7734));
  OR2 OR2_367(.VSS(VSS),.VDD(VDD),.Y(g4556),.A(g3536),.B(g2916));
  OR2 OR2_368(.VSS(VSS),.VDD(VDD),.Y(g8288),.A(g8119),.B(g7825));
  OR2 OR2_369(.VSS(VSS),.VDD(VDD),.Y(g6755),.A(g6106),.B(g5479));
  OR3 OR3_35(.VSS(VSS),.VDD(VDD),.Y(I14862),.A(g9587),.B(g9600),.C(g9611));
  OR4 OR4_33(.VSS(VSS),.VDD(VDD),.Y(I16160),.A(g10394),.B(g10392),.C(g10482),.D(g10481));
  OR4 OR4_34(.VSS(VSS),.VDD(VDD),.Y(I15042),.A(g7853),.B(g9686),.C(g9624),.D(g9785));
  OR2 OR2_370(.VSS(VSS),.VDD(VDD),.Y(g11610),.A(g11589),.B(g11560));
  OR4 OR4_35(.VSS(VSS),.VDD(VDD),.Y(g9711),.A(g9660),.B(g9390),.C(g9359),.D(g9589));
  OR2 OR2_371(.VSS(VSS),.VDD(VDD),.Y(g6045),.A(g5541),.B(g3989));
  OR2 OR2_372(.VSS(VSS),.VDD(VDD),.Y(g11270),.A(g11198),.B(g11032));
  OR2 OR2_373(.VSS(VSS),.VDD(VDD),.Y(g7258),.A(g6549),.B(g5913));
  OR2 OR2_374(.VSS(VSS),.VDD(VDD),.Y(g6059),.A(g5211),.B(g4489));
  OR2 OR2_375(.VSS(VSS),.VDD(VDD),.Y(g10007),.A(I15209),.B(I15210));
  OR2 OR2_376(.VSS(VSS),.VDD(VDD),.Y(g11267),.A(g11192),.B(g11029));
  OR2 OR2_377(.VSS(VSS),.VDD(VDD),.Y(g11294),.A(g6576),.B(g11210));
  OR3 OR3_36(.VSS(VSS),.VDD(VDD),.Y(g9509),.A(g9151),.B(g9125),.C(g9111));
  OR2 OR2_378(.VSS(VSS),.VDD(VDD),.Y(g7211),.A(g6647),.B(g6067));
  OR2 OR2_379(.VSS(VSS),.VDD(VDD),.Y(g5404),.A(g4487),.B(g3696));
  OR2 OR2_380(.VSS(VSS),.VDD(VDD),.Y(g4089),.A(g1959),.B(g3318));
  OR4 OR4_36(.VSS(VSS),.VDD(VDD),.Y(I15219),.A(g8172),.B(g9907),.C(g9936),.D(g9833));
  OR2 OR2_381(.VSS(VSS),.VDD(VDD),.Y(g11219),.A(g11145),.B(g11006));
  OR2 OR2_382(.VSS(VSS),.VDD(VDD),.Y(g6015),.A(g5497),.B(g3942));
  OR2 OR2_383(.VSS(VSS),.VDD(VDD),.Y(g10720),.A(g10304),.B(g10667));
  OR2 OR2_384(.VSS(VSS),.VDD(VDD),.Y(g8265),.A(g7881),.B(g3396));
  OR2 OR2_385(.VSS(VSS),.VDD(VDD),.Y(g5224),.A(g4360),.B(g3512));
  OR3 OR3_37(.VSS(VSS),.VDD(VDD),.Y(g9700),.A(g9358),.B(g9667),.C(I14827));
  OR2 OR2_386(.VSS(VSS),.VDD(VDD),.Y(g7106),.A(g6554),.B(g5917));
  OR2 OR2_387(.VSS(VSS),.VDD(VDD),.Y(g8770),.A(g5476),.B(g8651));
  OR2 OR2_388(.VSS(VSS),.VDD(VDD),.Y(g11201),.A(g11152),.B(g11011));
  OR3 OR3_38(.VSS(VSS),.VDD(VDD),.Y(g9950),.A(g9901),.B(g9898),.C(g9779));
  OR4 OR4_37(.VSS(VSS),.VDD(VDD),.Y(g9723),.A(g9620),.B(g9652),.C(g9391),.D(I14858));
  OR2 OR2_389(.VSS(VSS),.VDD(VDD),.Y(g2309),.A(I5357),.B(I5358));
  OR2 OR2_390(.VSS(VSS),.VDD(VDD),.Y(g11266),.A(g11190),.B(g11028));
  OR2 OR2_391(.VSS(VSS),.VDD(VDD),.Y(g10727),.A(g4969),.B(g10638));
  OR2 OR2_392(.VSS(VSS),.VDD(VDD),.Y(g10863),.A(g5531),.B(g10750));
  OR2 OR2_393(.VSS(VSS),.VDD(VDD),.Y(g8429),.A(g8385),.B(g8069));
  OR2 OR2_394(.VSS(VSS),.VDD(VDD),.Y(g9751),.A(g9515),.B(g9510));
  OR2 OR2_395(.VSS(VSS),.VDD(VDD),.Y(g8281),.A(g8097),.B(g7818));
  OR2 OR2_396(.VSS(VSS),.VDD(VDD),.Y(g6910),.A(g6341),.B(g5680));
  OR2 OR2_397(.VSS(VSS),.VDD(VDD),.Y(g8639),.A(g8118),.B(g8462));
  OR3 OR3_39(.VSS(VSS),.VDD(VDD),.Y(g9673),.A(g9454),.B(g9292),.C(g9274));
  OR2 OR2_398(.VSS(VSS),.VDD(VDD),.Y(g11285),.A(g11255),.B(g11161));
  OR2 OR2_399(.VSS(VSS),.VDD(VDD),.Y(g11305),.A(g11215),.B(g11093));
  OR4 OR4_38(.VSS(VSS),.VDD(VDD),.Y(I15177),.A(g9844),.B(g9960),.C(g9863),.D(g9876));
  OR3 OR3_40(.VSS(VSS),.VDD(VDD),.Y(g9734),.A(g9415),.B(g9428),.C(g9421));
  OR3 OR3_41(.VSS(VSS),.VDD(VDD),.Y(I14827),.A(g9603),.B(g9614),.C(g9584));
  OR2 OR2_400(.VSS(VSS),.VDD(VDD),.Y(g5824),.A(g5602),.B(g4839));
  OR2 OR2_401(.VSS(VSS),.VDD(VDD),.Y(g8715),.A(g8416),.B(g8687));
  OR2 OR2_402(.VSS(VSS),.VDD(VDD),.Y(g5762),.A(g5178),.B(g5186));
  OR2 OR2_403(.VSS(VSS),.VDD(VDD),.Y(g6538),.A(g5782),.B(g5006));
  OR2 OR2_404(.VSS(VSS),.VDD(VDD),.Y(g5590),.A(g4718),.B(g4723));
  OR2 OR2_405(.VSS(VSS),.VDD(VDD),.Y(g10726),.A(g10316),.B(g10673));
  OR2 OR2_406(.VSS(VSS),.VDD(VDD),.Y(g3120),.A(I6350),.B(I6351));
  OR2 OR2_407(.VSS(VSS),.VDD(VDD),.Y(g9573),.A(g9052),.B(g9030));
  OR3 OR3_42(.VSS(VSS),.VDD(VDD),.Y(g4640),.A(g3348),.B(g3563),.C(g1527));
  OR2 OR2_408(.VSS(VSS),.VDD(VDD),.Y(g6093),.A(g5264),.B(g4534));
  OR2 OR2_409(.VSS(VSS),.VDD(VDD),.Y(g8162),.A(g7898),.B(g6889));
  OR2 OR2_410(.VSS(VSS),.VDD(VDD),.Y(g8268),.A(g7962),.B(g7613));
  OR2 OR2_411(.VSS(VSS),.VDD(VDD),.Y(g9569),.A(g9052),.B(g9030));
  OR2 OR2_412(.VSS(VSS),.VDD(VDD),.Y(g11485),.A(g6646),.B(g11462));
  OR2 OR2_413(.VSS(VSS),.VDD(VDD),.Y(g10797),.A(g6206),.B(g10766));
  OR3 OR3_43(.VSS(VSS),.VDD(VDD),.Y(I14779),.A(g8995),.B(g9205),.C(g9192));
  OR2 OR2_414(.VSS(VSS),.VDD(VDD),.Y(g10408),.A(g10298),.B(g9553));
  OR2 OR2_415(.VSS(VSS),.VDD(VDD),.Y(g10635),.A(g10622),.B(g7732));
  OR2 OR2_416(.VSS(VSS),.VDD(VDD),.Y(g2305),.A(I5351),.B(I5352));
  OR4 OR4_39(.VSS(VSS),.VDD(VDD),.Y(I15176),.A(g8176),.B(g9910),.C(g9897),.D(g9836));
  OR2 OR2_417(.VSS(VSS),.VDD(VDD),.Y(g3435),.A(g2945),.B(g2950));
  OR2 OR2_418(.VSS(VSS),.VDD(VDD),.Y(g9924),.A(g9866),.B(g9709));
  OR2 OR2_419(.VSS(VSS),.VDD(VDD),.Y(g10711),.A(g5547),.B(g10690));
  OR2 OR2_420(.VSS(VSS),.VDD(VDD),.Y(g5814),.A(g5591),.B(g4827));
  OR2 OR2_421(.VSS(VSS),.VDD(VDD),.Y(g5038),.A(g4878),.B(g4884));
  OR4 OR4_40(.VSS(VSS),.VDD(VDD),.Y(I15215),.A(g9840),.B(g9965),.C(g9854),.D(g9879));
  OR2 OR2_422(.VSS(VSS),.VDD(VDD),.Y(g8226),.A(g7504),.B(g8002));
  OR2 OR2_423(.VSS(VSS),.VDD(VDD),.Y(g7367),.A(g7224),.B(g6744));
  OR2 OR2_424(.VSS(VSS),.VDD(VDD),.Y(g7457),.A(g6873),.B(g6404));
  OR2 OR2_425(.VSS(VSS),.VDD(VDD),.Y(g5229),.A(g4364),.B(g3516));
  OR2 OR2_426(.VSS(VSS),.VDD(VDD),.Y(g5993),.A(g5090),.B(g4400));
  OR2 OR2_427(.VSS(VSS),.VDD(VDD),.Y(g8283),.A(g8098),.B(g7820));
  OR2 OR2_428(.VSS(VSS),.VDD(VDD),.Y(g7971),.A(g5110),.B(g7549));
  OR2 OR2_429(.VSS(VSS),.VDD(VDD),.Y(g8602),.A(g8401),.B(g8550));
  OR2 OR2_430(.VSS(VSS),.VDD(VDD),.Y(g8920),.A(g8845),.B(g8759));
  OR2 OR2_431(.VSS(VSS),.VDD(VDD),.Y(g10663),.A(g10237),.B(g10581));
  OR2 OR2_432(.VSS(VSS),.VDD(VDD),.Y(g6074),.A(g5349),.B(g1));
  OR2 OR2_433(.VSS(VSS),.VDD(VDD),.Y(g8261),.A(g7876),.B(g3383));
  OR2 OR2_434(.VSS(VSS),.VDD(VDD),.Y(g10862),.A(g5524),.B(g10746));
  OR2 OR2_435(.VSS(VSS),.VDD(VDD),.Y(g5837),.A(g5640),.B(g4224));
  OR2 OR2_436(.VSS(VSS),.VDD(VDD),.Y(g11333),.A(g11274),.B(g11173));
  OR2 OR2_437(.VSS(VSS),.VDD(VDD),.Y(g6080),.A(g5249),.B(g4512));
  OR2 OR2_438(.VSS(VSS),.VDD(VDD),.Y(g6480),.A(g5721),.B(g4971));
  OR2 OR2_439(.VSS(VSS),.VDD(VDD),.Y(g7740),.A(g7209),.B(g6741));
  OR2 OR2_440(.VSS(VSS),.VDD(VDD),.Y(g10702),.A(g10562),.B(g3877));
  OR3 OR3_44(.VSS(VSS),.VDD(VDD),.Y(g9697),.A(g9665),.B(g9606),.C(I14822));
  OR2 OR2_441(.VSS(VSS),.VDD(VDD),.Y(g8203),.A(g7453),.B(g7999));
  OR2 OR2_442(.VSS(VSS),.VDD(VDD),.Y(g9914),.A(g9851),.B(g9692));
  OR2 OR2_443(.VSS(VSS),.VDD(VDD),.Y(g10564),.A(g10560),.B(g7368));
  OR2 OR2_444(.VSS(VSS),.VDD(VDD),.Y(g11484),.A(g6639),.B(g11461));
  OR2 OR2_445(.VSS(VSS),.VDD(VDD),.Y(g5842),.A(g5618),.B(g4870));
  OR4 OR4_41(.VSS(VSS),.VDD(VDD),.Y(I15200),.A(g9837),.B(g9962),.C(g9848),.D(g9880));
  OR2 OR2_446(.VSS(VSS),.VDD(VDD),.Y(g11609),.A(g11588),.B(g11559));
  OR3 OR3_45(.VSS(VSS),.VDD(VDD),.Y(I14582),.A(g8995),.B(g9205),.C(g9192));
  OR2 OR2_447(.VSS(VSS),.VDD(VDD),.Y(g8940),.A(g8793),.B(g8703));
  OR2 OR2_448(.VSS(VSS),.VDD(VDD),.Y(g11312),.A(g11222),.B(g11101));
  OR2 OR2_449(.VSS(VSS),.VDD(VDD),.Y(g11608),.A(g11587),.B(g11558));
  OR2 OR2_450(.VSS(VSS),.VDD(VDD),.Y(g6000),.A(g5480),.B(g3912));
  OR2 OR2_451(.VSS(VSS),.VDD(VDD),.Y(g8428),.A(g8382),.B(g8068));
  OR2 OR2_452(.VSS(VSS),.VDD(VDD),.Y(g8430),.A(g8386),.B(g8070));
  OR2 OR2_453(.VSS(VSS),.VDD(VDD),.Y(g9922),.A(g9864),.B(g9705));
  OR2 OR2_454(.VSS(VSS),.VDD(VDD),.Y(g8247),.A(g8010),.B(g7704));
  OR2 OR2_455(.VSS(VSS),.VDD(VDD),.Y(g3438),.A(g2939),.B(g2944));
  OR4 OR4_42(.VSS(VSS),.VDD(VDD),.Y(I5576),.A(g431),.B(g435),.C(g440),.D(g444));
  OR2 OR2_456(.VSS(VSS),.VDD(VDD),.Y(g6924),.A(g6362),.B(g4261));
  OR2 OR2_457(.VSS(VSS),.VDD(VDD),.Y(g5405),.A(g4476),.B(g3440));
  OR2 OR2_458(.VSS(VSS),.VDD(VDD),.Y(g8638),.A(g8108),.B(g8461));
  OR2 OR2_459(.VSS(VSS),.VDD(VDD),.Y(g8609),.A(g8408),.B(g8555));
  OR2 OR2_460(.VSS(VSS),.VDD(VDD),.Y(g9995),.A(I15199),.B(I15200));
  OR2 OR2_461(.VSS(VSS),.VDD(VDD),.Y(g8883),.A(g8838),.B(g8753));
  OR4 OR4_43(.VSS(VSS),.VDD(VDD),.Y(I15214),.A(g8170),.B(g9906),.C(g9935),.D(g9831));
  OR3 OR3_46(.VSS(VSS),.VDD(VDD),.Y(g2538),.A(g1466),.B(g1458),.C(I5649));
  OR2 OR2_462(.VSS(VSS),.VDD(VDD),.Y(g11329),.A(g11302),.B(g11169));
  OR2 OR2_463(.VSS(VSS),.VDD(VDD),.Y(g4255),.A(g4009),.B(g4047));
  OR2 OR2_464(.VSS(VSS),.VDD(VDD),.Y(g11328),.A(g11299),.B(g11168));
  OR3 OR3_47(.VSS(VSS),.VDD(VDD),.Y(g9704),.A(g9385),.B(g9605),.C(I14835));
  OR4 OR4_44(.VSS(VSS),.VDD(VDD),.Y(I5352),.A(g1129),.B(g1125),.C(g1121),.D(g1117));
  OR2 OR2_465(.VSS(VSS),.VDD(VDD),.Y(g8774),.A(g5499),.B(g8654));
  OR3 OR3_48(.VSS(VSS),.VDD(VDD),.Y(g9954),.A(g9946),.B(g9940),.C(g9781));
  OR2 OR2_466(.VSS(VSS),.VDD(VDD),.Y(g10405),.A(g10297),.B(g9530));
  OR2 OR2_467(.VSS(VSS),.VDD(VDD),.Y(g9363),.A(g9205),.B(g9192));
  OR2 OR2_468(.VSS(VSS),.VDD(VDD),.Y(g5849),.A(g4949),.B(g4260));
  OR4 OR4_45(.VSS(VSS),.VDD(VDD),.Y(I5599),.A(g516),.B(g511),.C(g506),.D(g501));
  OR2 OR2_469(.VSS(VSS),.VDD(VDD),.Y(g7204),.A(g6645),.B(g6062));
  OR2 OR2_470(.VSS(VSS),.VDD(VDD),.Y(g7300),.A(g7139),.B(g6326));
  OR2 OR2_471(.VSS(VSS),.VDD(VDD),.Y(g4293),.A(g4064),.B(g4068));
  OR2 OR2_472(.VSS(VSS),.VDD(VDD),.Y(g9912),.A(g9847),.B(g9690));
  OR2 OR2_473(.VSS(VSS),.VDD(VDD),.Y(g6533),.A(g5771),.B(g5002));
  OR2 OR2_474(.VSS(VSS),.VDD(VDD),.Y(g8816),.A(g7951),.B(g8731));
  OR2 OR2_475(.VSS(VSS),.VDD(VDD),.Y(g9929),.A(g9871),.B(g9718));
  OR2 OR2_476(.VSS(VSS),.VDD(VDD),.Y(g5819),.A(g5625),.B(g4876));
  OR3 OR3_49(.VSS(VSS),.VDD(VDD),.Y(I14831),.A(g9613),.B(g9622),.C(g9586));
  OR2 OR2_477(.VSS(VSS),.VDD(VDD),.Y(g5852),.A(g5632),.B(g4883));
  OR2 OR2_478(.VSS(VSS),.VDD(VDD),.Y(g8263),.A(g8032),.B(g7720));
  OR2 OR2_479(.VSS(VSS),.VDD(VDD),.Y(g3431),.A(g2951),.B(g2957));
  OR3 OR3_50(.VSS(VSS),.VDD(VDD),.Y(g9683),.A(g9454),.B(g9292),.C(g9274));
  OR2 OR2_480(.VSS(VSS),.VDD(VDD),.Y(g8631),.A(g8474),.B(g7449));
  OR2 OR2_481(.VSS(VSS),.VDD(VDD),.Y(g6922),.A(g6352),.B(g5694));
  OR2 OR2_482(.VSS(VSS),.VDD(VDD),.Y(g8817),.A(g7954),.B(g8732));
  OR4 OR4_46(.VSS(VSS),.VDD(VDD),.Y(g9735),.A(g9649),.B(g9651),.C(g9384),.D(g9361));
  OR2 OR2_483(.VSS(VSS),.VDD(VDD),.Y(g8605),.A(g8404),.B(g8553));
  OR2 OR2_484(.VSS(VSS),.VDD(VDD),.Y(g11263),.A(g11187),.B(g11025));
  OR2 OR2_485(.VSS(VSS),.VDD(VDD),.Y(g6739),.A(g5769),.B(g5780));
  OR2 OR2_486(.VSS(VSS),.VDD(VDD),.Y(g11332),.A(g11273),.B(g11172));
  OR2 OR2_487(.VSS(VSS),.VDD(VDD),.Y(g7143),.A(g6619),.B(g6039));
  OR2 OR2_488(.VSS(VSS),.VDD(VDD),.Y(g6479),.A(g5707),.B(g4968));
  OR4 OR4_47(.VSS(VSS),.VDD(VDD),.Y(I15048),.A(g7853),.B(g9683),.C(g9624),.D(g9785));
  OR2 OR2_489(.VSS(VSS),.VDD(VDD),.Y(g6501),.A(g5726),.B(g4987));
  OR3 OR3_51(.VSS(VSS),.VDD(VDD),.Y(g9702),.A(g9365),.B(g9647),.C(I14831));
  OR2 OR2_490(.VSS(VSS),.VDD(VDD),.Y(g11221),.A(g11146),.B(g11007));
  OR3 OR3_52(.VSS(VSS),.VDD(VDD),.Y(g9952),.A(g9944),.B(g9938),.C(g9817));
  OR2 OR2_491(.VSS(VSS),.VDD(VDD),.Y(g11613),.A(g11600),.B(g11591));
  OR2 OR2_492(.VSS(VSS),.VDD(VDD),.Y(g7621),.A(g5108),.B(g6994));
  OR2 OR2_493(.VSS(VSS),.VDD(VDD),.Y(g3399),.A(g2918),.B(g2940));
  OR2 OR2_494(.VSS(VSS),.VDD(VDD),.Y(g11605),.A(g11584),.B(g11555));
  OR2 OR2_495(.VSS(VSS),.VDD(VDD),.Y(g4274),.A(g4054),.B(g4058));
  OR3 OR3_53(.VSS(VSS),.VDD(VDD),.Y(I14602),.A(g8995),.B(g9205),.C(g9192));
  OR4 OR4_48(.VSS(VSS),.VDD(VDD),.Y(I15033),.A(g7853),.B(g9804),.C(g9624),.D(g9785));
  OR2 OR2_496(.VSS(VSS),.VDD(VDD),.Y(g10717),.A(g6235),.B(g10705));
  OR3 OR3_54(.VSS(VSS),.VDD(VDD),.Y(I5629),.A(g845),.B(g841),.C(g837));
  OR2 OR2_497(.VSS(VSS),.VDD(VDD),.Y(g9925),.A(g9867),.B(g9712));
  OR2 OR2_498(.VSS(VSS),.VDD(VDD),.Y(g3819),.A(g3275),.B(g9));
  OR2 OR2_499(.VSS(VSS),.VDD(VDD),.Y(g6912),.A(g6350),.B(g4235));
  OR2 OR2_500(.VSS(VSS),.VDD(VDD),.Y(g10723),.A(g4952),.B(g10633));
  OR2 OR2_501(.VSS(VSS),.VDD(VDD),.Y(g6929),.A(g6360),.B(g5704));
  OR2 OR2_502(.VSS(VSS),.VDD(VDD),.Y(g10646),.A(g10625),.B(g7739));
  OR2 OR2_503(.VSS(VSS),.VDD(VDD),.Y(g9516),.A(g9151),.B(g9125));
  OR2 OR2_504(.VSS(VSS),.VDD(VDD),.Y(g6626),.A(g5934),.B(g123));
  OR4 OR4_49(.VSS(VSS),.VDD(VDD),.Y(I6350),.A(g2445),.B(g2437),.C(g2433),.D(g2419));
  OR2 OR2_505(.VSS(VSS),.VDD(VDD),.Y(g11325),.A(g11295),.B(g11165));
  OR4 OR4_50(.VSS(VSS),.VDD(VDD),.Y(I5366),.A(g1280),.B(g1284),.C(g1292),.D(g1296));
  OR3 OR3_55(.VSS(VSS),.VDD(VDD),.Y(I5649),.A(g1499),.B(g1486),.C(g1482));
  OR2 OR2_506(.VSS(VSS),.VDD(VDD),.Y(g6894),.A(g6763),.B(g4868));
  OR3 OR3_56(.VSS(VSS),.VDD(VDD),.Y(g9738),.A(g9417),.B(g9447),.C(g9506));
  OR2 OR2_507(.VSS(VSS),.VDD(VDD),.Y(g8383),.A(g8163),.B(g5051));
  OR2 OR2_508(.VSS(VSS),.VDD(VDD),.Y(g8779),.A(g5530),.B(g8663));
  OR2 OR2_509(.VSS(VSS),.VDD(VDD),.Y(g8161),.A(g8005),.B(g7185));
  OR2 OR2_510(.VSS(VSS),.VDD(VDD),.Y(g8451),.A(g3440),.B(g8366));
  OR2 OR2_511(.VSS(VSS),.VDD(VDD),.Y(g9915),.A(g9853),.B(g9693));
  OR4 OR4_51(.VSS(VSS),.VDD(VDD),.Y(g2316),.A(g1300),.B(g1304),.C(g1270),.D(I5366));
  OR2 OR2_512(.VSS(VSS),.VDD(VDD),.Y(g5576),.A(g4675),.B(g3664));
  OR2 OR2_513(.VSS(VSS),.VDD(VDD),.Y(g10857),.A(g6090),.B(g10738));
  OR2 OR2_514(.VSS(VSS),.VDD(VDD),.Y(g10793),.A(g6194),.B(g10763));
  OR2 OR2_515(.VSS(VSS),.VDD(VDD),.Y(g7511),.A(g6890),.B(g6438));
  OR2 OR2_516(.VSS(VSS),.VDD(VDD),.Y(g8944),.A(g8799),.B(g8708));
  OR2 OR2_517(.VSS(VSS),.VDD(VDD),.Y(g10765),.A(g5492),.B(g10680));
  OR2 OR2_518(.VSS(VSS),.VDD(VDD),.Y(g10549),.A(g4951),.B(g10451));
  OR2 OR2_519(.VSS(VSS),.VDD(VDD),.Y(g7092),.A(g6540),.B(g5902));
  OR2 OR2_520(.VSS(VSS),.VDD(VDD),.Y(g11604),.A(g11583),.B(g11554));
  OR2 OR2_521(.VSS(VSS),.VDD(VDD),.Y(g8434),.A(g8400),.B(g8074));
  OR2 OR2_522(.VSS(VSS),.VDD(VDD),.Y(g6546),.A(g5796),.B(g5026));
  OR2 OR2_523(.VSS(VSS),.VDD(VDD),.Y(g3354),.A(g2920),.B(g2124));
  OR2 OR2_524(.VSS(VSS),.VDD(VDD),.Y(g9928),.A(g9870),.B(g9717));
  OR2 OR2_525(.VSS(VSS),.VDD(VDD),.Y(g11262),.A(g11240),.B(g11024));
  OR4 OR4_52(.VSS(VSS),.VDD(VDD),.Y(g9785),.A(g9010),.B(g8995),.C(g9388),.D(g9363));
  OR2 OR2_526(.VSS(VSS),.VDD(VDD),.Y(g5867),.A(g3440),.B(g4921));
  OR2 OR2_527(.VSS(VSS),.VDD(VDD),.Y(g8210),.A(g7466),.B(g7995));
  OR2 OR2_528(.VSS(VSS),.VDD(VDD),.Y(g10533),.A(g4933),.B(g10449));
  OR2 OR2_529(.VSS(VSS),.VDD(VDD),.Y(g9563),.A(g9052),.B(g9030));
  OR2 OR2_530(.VSS(VSS),.VDD(VDD),.Y(g6906),.A(g6791),.B(g5674));
  OR2 OR2_531(.VSS(VSS),.VDD(VDD),.Y(g7375),.A(g7230),.B(g6745));
  OR2 OR2_532(.VSS(VSS),.VDD(VDD),.Y(g7651),.A(g7135),.B(g4084));
  OR4 OR4_53(.VSS(VSS),.VDD(VDD),.Y(I5570),.A(g416),.B(g411),.C(g406),.D(g401));
  OR3 OR3_57(.VSS(VSS),.VDD(VDD),.Y(g9731),.A(g9641),.B(g9364),.C(g9387));
  OR2 OR2_533(.VSS(VSS),.VDD(VDD),.Y(g11247),.A(g11097),.B(g10949));
  OR4 OR4_54(.VSS(VSS),.VDD(VDD),.Y(I15045),.A(g7853),.B(g9676),.C(g9624),.D(g9785));
  OR2 OR2_534(.VSS(VSS),.VDD(VDD),.Y(g10856),.A(g6083),.B(g10737));
  OR2 OR2_535(.VSS(VSS),.VDD(VDD),.Y(g9557),.A(g9052),.B(g9030));
  OR2 OR2_536(.VSS(VSS),.VDD(VDD),.Y(g7184),.A(g6625),.B(g6047));
  OR2 OR2_537(.VSS(VSS),.VDD(VDD),.Y(g11612),.A(g11599),.B(g11590));
  OR2 OR2_538(.VSS(VSS),.VDD(VDD),.Y(g7384),.A(g7088),.B(g6618));
  OR2 OR2_539(.VSS(VSS),.VDD(VDD),.Y(g11324),.A(g11271),.B(g11164));
  OR2 OR2_540(.VSS(VSS),.VDD(VDD),.Y(g8922),.A(g8822),.B(g8736));
  OR4 OR4_55(.VSS(VSS),.VDD(VDD),.Y(I5358),.A(g1245),.B(g1240),.C(g1235),.D(g1275));
  OR3 OR3_58(.VSS(VSS),.VDD(VDD),.Y(g9955),.A(g9947),.B(g9941),.C(g9808));
  OR4 OR4_56(.VSS(VSS),.VDD(VDD),.Y(g2501),.A(g448),.B(g452),.C(g421),.D(I5576));
  OR2 OR2_541(.VSS(VSS),.VDD(VDD),.Y(g7231),.A(g6673),.B(g6087));
  OR2 OR2_542(.VSS(VSS),.VDD(VDD),.Y(g6078),.A(g4503),.B(g5256));
  OR2 OR2_543(.VSS(VSS),.VDD(VDD),.Y(g6478),.A(g5706),.B(g4967));
  OR2 OR2_544(.VSS(VSS),.VDD(VDD),.Y(g6907),.A(g6792),.B(g5675));
  OR2 OR2_545(.VSS(VSS),.VDD(VDD),.Y(g6035),.A(g5518),.B(g3974));
  OR2 OR2_546(.VSS(VSS),.VDD(VDD),.Y(g8937),.A(g8786),.B(g8698));
  OR2 OR2_547(.VSS(VSS),.VDD(VDD),.Y(g7742),.A(g7217),.B(g6743));
  OR2 OR2_548(.VSS(VSS),.VDD(VDD),.Y(g10722),.A(g10308),.B(g10671));
  OR2 OR2_549(.VSS(VSS),.VDD(VDD),.Y(g9918),.A(g9858),.B(g9698));
  OR2 OR2_550(.VSS(VSS),.VDD(VDD),.Y(g5403),.A(g4486),.B(g3695));
  OR2 OR2_551(.VSS(VSS),.VDD(VDD),.Y(g7926),.A(g7435),.B(g6892));
  OR2 OR2_552(.VSS(VSS),.VDD(VDD),.Y(g6915),.A(g6347),.B(g5686));
  OR2 OR2_553(.VSS(VSS),.VDD(VDD),.Y(g5841),.A(g4914),.B(g4230));
  OR4 OR4_57(.VSS(VSS),.VDD(VDD),.Y(I15220),.A(g9841),.B(g9966),.C(g9857),.D(g9877));
  OR2 OR2_554(.VSS(VSS),.VDD(VDD),.Y(g10529),.A(I16160),.B(I16161));
  OR2 OR2_555(.VSS(VSS),.VDD(VDD),.Y(g11246),.A(g11094),.B(g10948));
  OR2 OR2_556(.VSS(VSS),.VDD(VDD),.Y(g6002),.A(g5489),.B(g3939));
  OR2 OR2_557(.VSS(VSS),.VDD(VDD),.Y(g7712),.A(g7125),.B(g3540));
  OR2 OR2_558(.VSS(VSS),.VDD(VDD),.Y(g8810),.A(g7933),.B(g8720));
  OR2 OR2_559(.VSS(VSS),.VDD(VDD),.Y(g9921),.A(g9862),.B(g9703));
  OR2 OR2_560(.VSS(VSS),.VDD(VDD),.Y(g8432),.A(g8389),.B(g8072));
  OR4 OR4_58(.VSS(VSS),.VDD(VDD),.Y(I15172),.A(g9843),.B(g9959),.C(g9861),.D(g9874));
  OR3 OR3_59(.VSS(VSS),.VDD(VDD),.Y(I14822),.A(g9597),.B(g9604),.C(g9582));
  OR2 OR2_561(.VSS(VSS),.VDD(VDD),.Y(g6928),.A(g6359),.B(g5703));
  OR2 OR2_562(.VSS(VSS),.VDD(VDD),.Y(g8157),.A(g7965),.B(g7623));
  OR2 OR2_563(.VSS(VSS),.VDD(VDD),.Y(g6930),.A(g6364),.B(g4269));
  OR2 OR2_564(.VSS(VSS),.VDD(VDD),.Y(g7660),.A(g7059),.B(g6583));
  OR2 OR2_565(.VSS(VSS),.VDD(VDD),.Y(g6899),.A(g6463),.B(g5471));
  OR2 OR2_566(.VSS(VSS),.VDD(VDD),.Y(g9392),.A(g9328),.B(g9324));
  OR2 OR2_567(.VSS(VSS),.VDD(VDD),.Y(g11318),.A(g11228),.B(g11104));
  OR3 OR3_60(.VSS(VSS),.VDD(VDD),.Y(I16427),.A(g10683),.B(g10608),.C(g10604));
  OR2 OR2_568(.VSS(VSS),.VDD(VDD),.Y(g11227),.A(g11151),.B(g11010));
  OR2 OR2_569(.VSS(VSS),.VDD(VDD),.Y(g11058),.A(g10933),.B(g5280));
  OR4 OR4_59(.VSS(VSS),.VDD(VDD),.Y(I5351),.A(g1145),.B(g1141),.C(g1137),.D(g1133));
  OR3 OR3_61(.VSS(VSS),.VDD(VDD),.Y(g9708),.A(g9653),.B(g9389),.C(g9646));
  OR2 OR2_570(.VSS(VSS),.VDD(VDD),.Y(g6071),.A(g5228),.B(g4505));
  OR2 OR2_571(.VSS(VSS),.VDD(VDD),.Y(g9911),.A(g9846),.B(g9689));
  OR2 OR2_572(.VSS(VSS),.VDD(VDD),.Y(g7102),.A(g6550),.B(g5915));
  OR2 OR2_573(.VSS(VSS),.VDD(VDD),.Y(g7302),.A(g7141),.B(g6328));
  OR2 OR2_574(.VSS(VSS),.VDD(VDD),.Y(g6038),.A(g5528),.B(g3979));
  OR2 OR2_575(.VSS(VSS),.VDD(VDD),.Y(g4239),.A(g4000),.B(g4008));
  OR2 OR2_576(.VSS(VSS),.VDD(VDD),.Y(g8646),.A(g8224),.B(g8547));
  OR2 OR2_577(.VSS(VSS),.VDD(VDD),.Y(g9974),.A(I15176),.B(I15177));
  OR2 OR2_578(.VSS(VSS),.VDD(VDD),.Y(g5823),.A(g5631),.B(g4882));
  OR2 OR2_579(.VSS(VSS),.VDD(VDD),.Y(g6918),.A(g6358),.B(g4252));
  OR2 OR2_580(.VSS(VSS),.VDD(VDD),.Y(g7265),.A(g6756),.B(g6204));
  OR4 OR4_60(.VSS(VSS),.VDD(VDD),.Y(I5804),.A(g2111),.B(g2109),.C(g2106),.D(g2104));
  OR2 OR2_581(.VSS(VSS),.VDD(VDD),.Y(g5851),.A(g4941),.B(g4253));
  OR2 OR2_582(.VSS(VSS),.VDD(VDD),.Y(g11481),.A(g6624),.B(g11458));
  OR2 OR2_583(.VSS(VSS),.VDD(VDD),.Y(g10336),.A(g10230),.B(g9572));
  OR2 OR2_584(.VSS(VSS),.VDD(VDD),.Y(g7296),.A(g7131),.B(g6322));
  OR2 OR2_585(.VSS(VSS),.VDD(VDD),.Y(g4300),.A(g3546),.B(g2391));
  OR2 OR2_586(.VSS(VSS),.VDD(VDD),.Y(g8647),.A(g8130),.B(g8470));
//
  NAND2 NAND2_0(.VSS(VSS),.VDD(VDD),.Y(g8546),.A(g3983),.B(g8390));
  NAND2 NAND2_1(.VSS(VSS),.VDD(VDD),.Y(g2516),.A(I5612),.B(I5613));
  NAND2 NAND2_2(.VSS(VSS),.VDD(VDD),.Y(g2987),.A(g2481),.B(g883));
  NAND2 NAND2_3(.VSS(VSS),.VDD(VDD),.Y(I5593),.A(g1703),.B(I5591));
  NAND2 NAND2_4(.VSS(VSS),.VDD(VDD),.Y(g8970),.A(g5548),.B(g8839));
  NAND2 NAND2_5(.VSS(VSS),.VDD(VDD),.Y(I10519),.A(g6231),.B(g822));
  NAND2 NAND2_6(.VSS(VSS),.VDD(VDD),.Y(I11279),.A(g305),.B(I11278));
  NAND4 NAND4_0(.VSS(VSS),.VDD(VDD),.Y(g7990),.A(g7011),.B(g6995),.C(g7562),.D(g7550));
  NAND2 NAND2_7(.VSS(VSS),.VDD(VDD),.Y(I11278),.A(g305),.B(g6485));
  NAND2 NAND2_8(.VSS(VSS),.VDD(VDD),.Y(g3978),.A(g3207),.B(g1822));
  NAND2 NAND2_9(.VSS(VSS),.VDD(VDD),.Y(I5264),.A(g456),.B(I5263));
  NAND2 NAND2_10(.VSS(VSS),.VDD(VDD),.Y(I8640),.A(g4278),.B(g516));
  NAND2 NAND2_11(.VSS(VSS),.VDD(VDD),.Y(I6761),.A(g2943),.B(I6760));
  NAND2 NAND2_12(.VSS(VSS),.VDD(VDD),.Y(I17400),.A(g11418),.B(g11416));
  NAND2 NAND2_13(.VSS(VSS),.VDD(VDD),.Y(I5450),.A(g1235),.B(I5449));
  NAND2 NAND2_14(.VSS(VSS),.VDD(VDD),.Y(I16060),.A(g10372),.B(I16058));
  NAND2 NAND2_15(.VSS(VSS),.VDD(VDD),.Y(I6746),.A(g2938),.B(g1453));
  NAND2 NAND2_16(.VSS(VSS),.VDD(VDD),.Y(I11975),.A(g1462),.B(I11973));
  NAND2 NAND2_17(.VSS(VSS),.VDD(VDD),.Y(I12136),.A(g7110),.B(g131));
  NAND2 NAND2_18(.VSS(VSS),.VDD(VDD),.Y(I11937),.A(g1458),.B(I11935));
  NAND2 NAND2_19(.VSS(VSS),.VDD(VDD),.Y(g2959),.A(I6167),.B(I6168));
  NAND2 NAND2_20(.VSS(VSS),.VDD(VDD),.Y(I5878),.A(g2120),.B(g2115));
  NAND2 NAND2_21(.VSS(VSS),.VDD(VDD),.Y(g2517),.A(I5619),.B(I5620));
  NAND2 NAND2_22(.VSS(VSS),.VDD(VDD),.Y(g5552),.A(g4777),.B(g4401));
  NAND2 NAND2_23(.VSS(VSS),.VDD(VDD),.Y(I6468),.A(g23),.B(I6467));
  NAND2 NAND2_24(.VSS(VSS),.VDD(VDD),.Y(I8796),.A(g4672),.B(I8795));
  NAND2 NAND2_25(.VSS(VSS),.VDD(VDD),.Y(g10392),.A(I15891),.B(I15892));
  NAND2 NAND2_26(.VSS(VSS),.VDD(VDD),.Y(I5611),.A(g1280),.B(g1284));
  NAND2 NAND2_27(.VSS(VSS),.VDD(VDD),.Y(g8738),.A(g8688),.B(g4921));
  NAND2 NAND2_28(.VSS(VSS),.VDD(VDD),.Y(I6716),.A(g201),.B(I6714));
  NAND2 NAND2_29(.VSS(VSS),.VDD(VDD),.Y(g2310),.A(g591),.B(g605));
  NAND2 NAND2_30(.VSS(VSS),.VDD(VDD),.Y(I7685),.A(g3460),.B(I7683));
  NAND2 NAND2_31(.VSS(VSS),.VDD(VDD),.Y(g3056),.A(g2374),.B(g599));
  NAND2 NAND2_32(.VSS(VSS),.VDD(VDD),.Y(I12108),.A(g135),.B(I12106));
  NAND3 NAND3_0(.VSS(VSS),.VDD(VDD),.Y(g3529),.A(g2310),.B(g3062),.C(g2325));
  NAND2 NAND2_33(.VSS(VSS),.VDD(VDD),.Y(I6747),.A(g2938),.B(I6746));
  NAND2 NAND2_34(.VSS(VSS),.VDD(VDD),.Y(g2236),.A(I5230),.B(I5231));
  NAND2 NAND2_35(.VSS(VSS),.VDD(VDD),.Y(g7584),.A(I12075),.B(I12076));
  NAND2 NAND2_36(.VSS(VSS),.VDD(VDD),.Y(I15870),.A(g10358),.B(g2713));
  NAND2 NAND2_37(.VSS(VSS),.VDD(VDD),.Y(I16067),.A(g2765),.B(I16065));
  NAND2 NAND2_38(.VSS(VSS),.VDD(VDD),.Y(I7562),.A(g3533),.B(g654));
  NAND2 NAND2_39(.VSS(VSS),.VDD(VDD),.Y(I13531),.A(g8253),.B(I13529));
  NAND2 NAND2_40(.VSS(VSS),.VDD(VDD),.Y(I8797),.A(g1145),.B(I8795));
  NAND2 NAND2_41(.VSS(VSS),.VDD(VDD),.Y(I17584),.A(g11354),.B(g11515));
  NAND2 NAND2_42(.VSS(VSS),.VDD(VDD),.Y(I11936),.A(g7004),.B(I11935));
  NAND2 NAND2_43(.VSS(VSS),.VDD(VDD),.Y(I15257),.A(g9984),.B(I15256));
  NAND2 NAND2_44(.VSS(VSS),.VDD(VDD),.Y(g8402),.A(I13505),.B(I13506));
  NAND3 NAND3_1(.VSS(VSS),.VDD(VDD),.Y(g8824),.A(g8502),.B(g8501),.C(g8739));
  NAND2 NAND2_45(.VSS(VSS),.VDD(VDD),.Y(I6186),.A(g2511),.B(g466));
  NAND2 NAND2_46(.VSS(VSS),.VDD(VDD),.Y(g11496),.A(I17504),.B(I17505));
  NAND2 NAND2_47(.VSS(VSS),.VDD(VDD),.Y(I16001),.A(g2683),.B(I15999));
  NAND2 NAND2_48(.VSS(VSS),.VDD(VDD),.Y(I6125),.A(g2215),.B(I6124));
  NAND2 NAND2_49(.VSS(VSS),.VDD(VDD),.Y(I11909),.A(g1474),.B(I11907));
  NAND2 NAND2_50(.VSS(VSS),.VDD(VDD),.Y(I12040),.A(g1466),.B(I12038));
  NAND2 NAND2_51(.VSS(VSS),.VDD(VDD),.Y(I13909),.A(g1432),.B(I13907));
  NAND2 NAND2_52(.VSS(VSS),.VDD(VDD),.Y(g3625),.A(I6771),.B(I6772));
  NAND2 NAND2_53(.VSS(VSS),.VDD(VDD),.Y(I11908),.A(g6967),.B(I11907));
  NAND2 NAND2_54(.VSS(VSS),.VDD(VDD),.Y(g10470),.A(I16008),.B(I16009));
  NAND2 NAND2_55(.VSS(VSS),.VDD(VDD),.Y(I13908),.A(g8526),.B(I13907));
  NAND2 NAND2_56(.VSS(VSS),.VDD(VDD),.Y(g3813),.A(I7034),.B(I7035));
  NAND2 NAND2_57(.VSS(VSS),.VDD(VDD),.Y(I8650),.A(g4824),.B(g778));
  NAND2 NAND2_58(.VSS(VSS),.VDD(VDD),.Y(g6207),.A(I9947),.B(I9948));
  NAND2 NAND2_59(.VSS(VSS),.VDD(VDD),.Y(I16066),.A(g10428),.B(I16065));
  NAND2 NAND2_60(.VSS(VSS),.VDD(VDD),.Y(g2948),.A(I6144),.B(I6145));
  NAND2 NAND2_61(.VSS(VSS),.VDD(VDD),.Y(I11242),.A(g6760),.B(I11241));
  NAND2 NAND2_62(.VSS(VSS),.VDD(VDD),.Y(g10467),.A(I15993),.B(I15994));
  NAND2 NAND2_63(.VSS(VSS),.VDD(VDD),.Y(I6187),.A(g2511),.B(I6186));
  NAND2 NAND2_64(.VSS(VSS),.VDD(VDD),.Y(g6488),.A(g6027),.B(g6019));
  NAND2 NAND2_65(.VSS(VSS),.VDD(VDD),.Y(I5500),.A(g1255),.B(g1007));
  NAND2 NAND2_66(.VSS(VSS),.VDD(VDD),.Y(I11974),.A(g7001),.B(I11973));
  NAND2 NAND2_67(.VSS(VSS),.VDD(VDD),.Y(I12062),.A(g1478),.B(I12060));
  NAND2 NAND2_68(.VSS(VSS),.VDD(VDD),.Y(g5300),.A(I8771),.B(I8772));
  NAND2 NAND2_69(.VSS(VSS),.VDD(VDD),.Y(I5184),.A(g1415),.B(g1515));
  NAND2 NAND2_70(.VSS(VSS),.VDD(VDD),.Y(I13293),.A(g1882),.B(g8161));
  NAND2 NAND2_71(.VSS(VSS),.VDD(VDD),.Y(I6200),.A(g2525),.B(I6199));
  NAND2 NAND2_72(.VSS(VSS),.VDD(VDD),.Y(I13265),.A(g1909),.B(g8154));
  NAND2 NAND2_73(.VSS(VSS),.VDD(VDD),.Y(I5024),.A(g995),.B(I5023));
  NAND2 NAND2_74(.VSS(VSS),.VDD(VDD),.Y(I7863),.A(g4099),.B(g774));
  NAND2 NAND2_75(.VSS(VSS),.VDD(VDD),.Y(g8705),.A(I13991),.B(I13992));
  NAND2 NAND2_76(.VSS(VSS),.VDD(VDD),.Y(g8471),.A(I13660),.B(I13661));
  NAND2 NAND2_77(.VSS(VSS),.VDD(VDD),.Y(I15256),.A(g9984),.B(g9980));
  NAND2 NAND2_78(.VSS(VSS),.VDD(VDD),.Y(I6145),.A(g646),.B(I6143));
  NAND2 NAND2_79(.VSS(VSS),.VDD(VDD),.Y(I13992),.A(g8688),.B(I13990));
  NAND2 NAND2_80(.VSS(VSS),.VDD(VDD),.Y(I11510),.A(g1806),.B(I11508));
  NAND2 NAND2_81(.VSS(VSS),.VDD(VDD),.Y(g10853),.A(g10731),.B(g5034));
  NAND2 NAND2_82(.VSS(VSS),.VDD(VDD),.Y(I5231),.A(g148),.B(I5229));
  NAND2 NAND2_83(.VSS(VSS),.VDD(VDD),.Y(I12047),.A(g1486),.B(I12045));
  NAND2 NAND2_84(.VSS(VSS),.VDD(VDD),.Y(I10771),.A(g1801),.B(I10769));
  NAND2 NAND2_85(.VSS(VSS),.VDD(VDD),.Y(g10477),.A(I16045),.B(I16046));
  NAND2 NAND2_86(.VSS(VSS),.VDD(VDD),.Y(g7582),.A(I12061),.B(I12062));
  NAND2 NAND2_87(.VSS(VSS),.VDD(VDD),.Y(I5104),.A(g431),.B(g435));
  NAND2 NAND2_88(.VSS(VSS),.VDD(VDD),.Y(g8409),.A(I13530),.B(I13531));
  NAND2 NAND2_89(.VSS(VSS),.VDD(VDD),.Y(I6447),.A(g2264),.B(g1776));
  NAND2 NAND2_90(.VSS(VSS),.VDD(VDD),.Y(I4956),.A(g327),.B(I4954));
  NAND2 NAND2_91(.VSS(VSS),.VDD(VDD),.Y(I5613),.A(g1284),.B(I5611));
  NAND2 NAND2_92(.VSS(VSS),.VDD(VDD),.Y(I8481),.A(g3530),.B(I8479));
  NAND2 NAND2_93(.VSS(VSS),.VDD(VDD),.Y(g5278),.A(I8739),.B(I8740));
  NAND2 NAND2_94(.VSS(VSS),.VDD(VDD),.Y(I6880),.A(g3301),.B(I6879));
  NAND2 NAND2_95(.VSS(VSS),.VDD(VDD),.Y(I15431),.A(g10047),.B(I15430));
  NAND2 NAND2_96(.VSS(VSS),.VDD(VDD),.Y(g5548),.A(g1840),.B(g4401));
  NAND4 NAND4_1(.VSS(VSS),.VDD(VDD),.Y(g7671),.A(g7011),.B(g6995),.C(g6984),.D(g6974));
  NAND2 NAND2_97(.VSS(VSS),.VDD(VDD),.Y(I12020),.A(g7119),.B(I12019));
  NAND2 NAND2_98(.VSS(VSS),.VDD(VDD),.Y(g10665),.A(I16331),.B(I16332));
  NAND2 NAND2_99(.VSS(VSS),.VDD(VDD),.Y(I16469),.A(g10518),.B(I16467));
  NAND2 NAND2_100(.VSS(VSS),.VDD(VDD),.Y(I5014),.A(g1007),.B(I5013));
  NAND2 NAND2_101(.VSS(VSS),.VDD(VDD),.Y(I13523),.A(g8249),.B(I13521));
  NAND2 NAND2_102(.VSS(VSS),.VDD(VDD),.Y(I16039),.A(g2707),.B(I16037));
  NAND2 NAND2_103(.VSS(VSS),.VDD(VDD),.Y(I16468),.A(g10716),.B(I16467));
  NAND2 NAND2_104(.VSS(VSS),.VDD(VDD),.Y(I12046),.A(g6951),.B(I12045));
  NAND2 NAND2_105(.VSS(VSS),.VDD(VDD),.Y(g4476),.A(g3807),.B(g3071));
  NAND2 NAND2_106(.VSS(VSS),.VDD(VDD),.Y(g10476),.A(I16038),.B(I16039));
  NAND2 NAND2_107(.VSS(VSS),.VDD(VDD),.Y(I16038),.A(g10427),.B(I16037));
  NAND2 NAND2_108(.VSS(VSS),.VDD(VDD),.Y(I8676),.A(g4374),.B(g1027));
  NAND2 NAND2_109(.VSS(VSS),.VDD(VDD),.Y(I12113),.A(g7093),.B(g162));
  NAND2 NAND2_110(.VSS(VSS),.VDD(VDD),.Y(I8761),.A(g4616),.B(g1129));
  NAND2 NAND2_111(.VSS(VSS),.VDD(VDD),.Y(g3204),.A(g2571),.B(g2061));
  NAND2 NAND2_112(.VSS(VSS),.VDD(VDD),.Y(I15993),.A(g10422),.B(I15992));
  NAND2 NAND2_113(.VSS(VSS),.VDD(VDD),.Y(I5036),.A(g1019),.B(I5034));
  NAND2 NAND2_114(.VSS(VSS),.VDD(VDD),.Y(I14263),.A(g8843),.B(g1814));
  NAND2 NAND2_115(.VSS(VSS),.VDD(VDD),.Y(g8298),.A(I13249),.B(I13250));
  NAND2 NAND2_116(.VSS(VSS),.VDD(VDD),.Y(I5135),.A(g521),.B(g525));
  NAND2 NAND2_117(.VSS(VSS),.VDD(VDD),.Y(g2405),.A(I5485),.B(I5486));
  NAND2 NAND2_118(.VSS(VSS),.VDD(VDD),.Y(I7034),.A(g3089),.B(I7033));
  NAND2 NAND2_119(.VSS(VSS),.VDD(VDD),.Y(I15443),.A(g10122),.B(I15441));
  NAND2 NAND2_120(.VSS(VSS),.VDD(VDD),.Y(I6166),.A(g2236),.B(g153));
  NAND2 NAND2_121(.VSS(VSS),.VDD(VDD),.Y(I8624),.A(g4267),.B(g511));
  NAND2 NAND2_122(.VSS(VSS),.VDD(VDD),.Y(I16015),.A(g10425),.B(g2695));
  NAND2 NAND2_123(.VSS(VSS),.VDD(VDD),.Y(I8677),.A(g4374),.B(I8676));
  NAND2 NAND2_124(.VSS(VSS),.VDD(VDD),.Y(I8576),.A(g4234),.B(I8575));
  NAND2 NAND2_125(.VSS(VSS),.VDD(VDD),.Y(I14613),.A(g9204),.B(I14612));
  NAND2 NAND2_126(.VSS(VSS),.VDD(VDD),.Y(I8716),.A(g4601),.B(I8715));
  NAND2 NAND2_127(.VSS(VSS),.VDD(VDD),.Y(g3530),.A(I6715),.B(I6716));
  NAND2 NAND2_128(.VSS(VSS),.VDD(VDD),.Y(g8405),.A(I13514),.B(I13515));
  NAND4 NAND4_2(.VSS(VSS),.VDD(VDD),.Y(g4104),.A(g3215),.B(g3247),.C(g2439),.D(g3200));
  NAND2 NAND2_129(.VSS(VSS),.VDD(VDD),.Y(I12003),.A(g7082),.B(I12002));
  NAND2 NAND2_130(.VSS(VSS),.VDD(VDD),.Y(g2177),.A(I5127),.B(I5128));
  NAND2 NAND2_131(.VSS(VSS),.VDD(VDD),.Y(g3010),.A(g2382),.B(g2399));
  NAND2 NAND2_132(.VSS(VSS),.VDD(VDD),.Y(g5179),.A(I8576),.B(I8577));
  NAND2 NAND2_133(.VSS(VSS),.VDD(VDD),.Y(I17395),.A(g11414),.B(I17393));
  NAND2 NAND2_134(.VSS(VSS),.VDD(VDD),.Y(g7067),.A(I11279),.B(I11280));
  NAND4 NAND4_3(.VSS(VSS),.VDD(VDD),.Y(g7994),.A(g7011),.B(g7574),.C(g6984),.D(g7550));
  NAND2 NAND2_135(.VSS(VSS),.VDD(VDD),.Y(I6167),.A(g2236),.B(I6166));
  NAND2 NAND2_136(.VSS(VSS),.VDD(VDD),.Y(I5265),.A(g461),.B(I5263));
  NAND2 NAND2_137(.VSS(VSS),.VDD(VDD),.Y(I6989),.A(g2760),.B(I6988));
  NAND2 NAND2_138(.VSS(VSS),.VDD(VDD),.Y(I13274),.A(g8158),.B(I13272));
  NAND2 NAND2_139(.VSS(VSS),.VDD(VDD),.Y(I10507),.A(g6221),.B(g786));
  NAND2 NAND2_140(.VSS(VSS),.VDD(VDD),.Y(I13530),.A(g704),.B(I13529));
  NAND2 NAND2_141(.VSS(VSS),.VDD(VDD),.Y(I5164),.A(g1508),.B(g1499));
  NAND2 NAND2_142(.VSS(VSS),.VDD(VDD),.Y(g9107),.A(I14443),.B(I14444));
  NAND2 NAND2_143(.VSS(VSS),.VDD(VDD),.Y(I9559),.A(g782),.B(I9557));
  NAND2 NAND2_144(.VSS(VSS),.VDD(VDD),.Y(I8577),.A(g496),.B(I8575));
  NAND2 NAND2_145(.VSS(VSS),.VDD(VDD),.Y(g2510),.A(I5592),.B(I5593));
  NAND2 NAND2_146(.VSS(VSS),.VDD(VDD),.Y(g8177),.A(I13077),.B(I13078));
  NAND2 NAND2_147(.VSS(VSS),.VDD(VDD),.Y(I8717),.A(g4052),.B(I8715));
  NAND2 NAND2_148(.VSS(VSS),.VDD(VDD),.Y(I5296),.A(g794),.B(I5295));
  NAND2 NAND2_149(.VSS(VSS),.VDD(VDD),.Y(g5209),.A(I8625),.B(I8626));
  NAND4 NAND4_4(.VSS(VSS),.VDD(VDD),.Y(g7950),.A(g7395),.B(g7390),.C(g7380),.D(g7273));
  NAND2 NAND2_150(.VSS(VSS),.VDD(VDD),.Y(g2088),.A(I4911),.B(I4912));
  NAND2 NAND2_151(.VSS(VSS),.VDD(VDD),.Y(I16000),.A(g10423),.B(I15999));
  NAND2 NAND2_152(.VSS(VSS),.VDD(VDD),.Y(I5371),.A(g971),.B(g976));
  NAND2 NAND2_153(.VSS(VSS),.VDD(VDD),.Y(g2215),.A(I5185),.B(I5186));
  NAND2 NAND2_154(.VSS(VSS),.VDD(VDD),.Y(g7101),.A(g6617),.B(g2364));
  NAND2 NAND2_155(.VSS(VSS),.VDD(VDD),.Y(I5675),.A(g1218),.B(g1223));
  NAND2 NAND2_156(.VSS(VSS),.VDD(VDD),.Y(I8544),.A(g4218),.B(I8543));
  NAND2 NAND2_157(.VSS(VSS),.VDD(VDD),.Y(g6577),.A(I10520),.B(I10521));
  NAND2 NAND2_158(.VSS(VSS),.VDD(VDD),.Y(I5297),.A(g798),.B(I5295));
  NAND2 NAND2_159(.VSS(VSS),.VDD(VDD),.Y(I13537),.A(g658),.B(g8157));
  NAND2 NAND2_160(.VSS(VSS),.VDD(VDD),.Y(I13283),.A(g1927),.B(g8159));
  NAND2 NAND2_161(.VSS(VSS),.VDD(VDD),.Y(g4749),.A(g3710),.B(g2061));
  NAND2 NAND2_162(.VSS(VSS),.VDD(VDD),.Y(I11982),.A(g1482),.B(I11980));
  NAND2 NAND2_163(.VSS(VSS),.VDD(VDD),.Y(I8514),.A(g4873),.B(I8513));
  NAND2 NAND2_164(.VSS(VSS),.VDD(VDD),.Y(I13091),.A(g1840),.B(I13089));
  NAND2 NAND2_165(.VSS(VSS),.VDD(VDD),.Y(g2943),.A(I6125),.B(I6126));
  NAND2 NAND2_166(.VSS(VSS),.VDD(VDD),.Y(I15908),.A(g10302),.B(I15906));
  NAND2 NAND2_167(.VSS(VSS),.VDD(VDD),.Y(I6879),.A(g3301),.B(g1351));
  NAND2 NAND2_168(.VSS(VSS),.VDD(VDD),.Y(I8763),.A(g1129),.B(I8761));
  NAND2 NAND2_169(.VSS(VSS),.VDD(VDD),.Y(I5449),.A(g1235),.B(g991));
  NAND3 NAND3_2(.VSS(VSS),.VDD(VDD),.Y(g8825),.A(g8502),.B(g8738),.C(g8506));
  NAND2 NAND2_170(.VSS(VSS),.VDD(VDD),.Y(I16007),.A(g10424),.B(g2689));
  NAND2 NAND2_171(.VSS(VSS),.VDD(VDD),.Y(I5865),.A(g2107),.B(g2105));
  NAND2 NAND2_172(.VSS(VSS),.VDD(VDD),.Y(I5604),.A(g1149),.B(g1153));
  NAND2 NAND2_173(.VSS(VSS),.VDD(VDD),.Y(g2433),.A(I5517),.B(I5518));
  NAND2 NAND2_174(.VSS(VSS),.VDD(VDD),.Y(I6111),.A(g1494),.B(I6109));
  NAND2 NAND2_175(.VSS(VSS),.VDD(VDD),.Y(g2096),.A(I4929),.B(I4930));
  NAND2 NAND2_176(.VSS(VSS),.VDD(VDD),.Y(I13522),.A(g695),.B(I13521));
  NAND2 NAND2_177(.VSS(VSS),.VDD(VDD),.Y(I10770),.A(g5944),.B(I10769));
  NAND2 NAND2_178(.VSS(VSS),.VDD(VDD),.Y(g6027),.A(g4566),.B(g4921));
  NAND4 NAND4_5(.VSS(VSS),.VDD(VDD),.Y(g7992),.A(g7011),.B(g7574),.C(g6984),.D(g6974));
  NAND2 NAND2_179(.VSS(VSS),.VDD(VDD),.Y(I5539),.A(g1270),.B(I5538));
  NAND2 NAND2_180(.VSS(VSS),.VDD(VDD),.Y(I17394),.A(g11415),.B(I17393));
  NAND2 NAND2_181(.VSS(VSS),.VDD(VDD),.Y(I13553),.A(g668),.B(I13552));
  NAND2 NAND2_182(.VSS(VSS),.VDD(VDD),.Y(I8642),.A(g516),.B(I8640));
  NAND2 NAND2_183(.VSS(VSS),.VDD(VDD),.Y(g7573),.A(I12046),.B(I12047));
  NAND2 NAND2_184(.VSS(VSS),.VDD(VDD),.Y(g11416),.A(I17296),.B(I17297));
  NAND2 NAND2_185(.VSS(VSS),.VDD(VDD),.Y(g6003),.A(g5552),.B(g5548));
  NAND2 NAND2_186(.VSS(VSS),.VDD(VDD),.Y(g8934),.A(I14278),.B(I14279));
  NAND2 NAND2_187(.VSS(VSS),.VDD(VDD),.Y(I15992),.A(g10422),.B(g2677));
  NAND2 NAND2_188(.VSS(VSS),.VDD(VDD),.Y(I7683),.A(g1023),.B(g3460));
  NAND2 NAND2_189(.VSS(VSS),.VDD(VDD),.Y(I4910),.A(g386),.B(g318));
  NAND4 NAND4_6(.VSS(VSS),.VDD(VDD),.Y(g3209),.A(g2550),.B(g2061),.C(g2564),.D(g2571));
  NAND2 NAND2_190(.VSS(VSS),.VDD(VDD),.Y(I6794),.A(g143),.B(I6792));
  NAND2 NAND2_191(.VSS(VSS),.VDD(VDD),.Y(I10521),.A(g822),.B(I10519));
  NAND2 NAND2_192(.VSS(VSS),.VDD(VDD),.Y(I5486),.A(g1011),.B(I5484));
  NAND2 NAND2_193(.VSS(VSS),.VDD(VDD),.Y(I15442),.A(g10035),.B(I15441));
  NAND2 NAND2_194(.VSS(VSS),.VDD(VDD),.Y(g6858),.A(I10931),.B(I10932));
  NAND2 NAND2_195(.VSS(VSS),.VDD(VDD),.Y(I5185),.A(g1415),.B(I5184));
  NAND2 NAND2_196(.VSS(VSS),.VDD(VDD),.Y(g5304),.A(I8779),.B(I8780));
  NAND2 NAND2_197(.VSS(VSS),.VDD(VDD),.Y(g2354),.A(g1515),.B(g1520));
  NAND2 NAND2_198(.VSS(VSS),.VDD(VDD),.Y(I15615),.A(g10043),.B(g10153));
  NAND2 NAND2_199(.VSS(VSS),.VDD(VDD),.Y(I17281),.A(g11360),.B(g11357));
  NAND2 NAND2_200(.VSS(VSS),.VDD(VDD),.Y(I5470),.A(g999),.B(I5468));
  NAND2 NAND2_201(.VSS(VSS),.VDD(VDD),.Y(I11509),.A(g6580),.B(I11508));
  NAND2 NAND2_202(.VSS(VSS),.VDD(VDD),.Y(I5025),.A(g1275),.B(I5023));
  NAND2 NAND2_203(.VSS(VSS),.VDD(VDD),.Y(I11508),.A(g6580),.B(g1806));
  NAND2 NAND2_204(.VSS(VSS),.VDD(VDD),.Y(I15430),.A(g10047),.B(g10044));
  NAND2 NAND2_205(.VSS(VSS),.VDD(VDD),.Y(I14612),.A(g9204),.B(g611));
  NAND2 NAND2_206(.VSS(VSS),.VDD(VDD),.Y(g4675),.A(g4073),.B(g3247));
  NAND2 NAND2_207(.VSS(VSS),.VDD(VDD),.Y(I14272),.A(g1822),.B(I14270));
  NAND2 NAND2_208(.VSS(VSS),.VDD(VDD),.Y(g2979),.A(I6208),.B(I6209));
  NAND2 NAND2_209(.VSS(VSS),.VDD(VDD),.Y(I17290),.A(g11363),.B(I17288));
  NAND2 NAND2_210(.VSS(VSS),.VDD(VDD),.Y(g5269),.A(I8716),.B(I8717));
  NAND2 NAND2_211(.VSS(VSS),.VDD(VDD),.Y(g4297),.A(I7563),.B(I7564));
  NAND2 NAND2_212(.VSS(VSS),.VDD(VDD),.Y(I12002),.A(g7082),.B(g153));
  NAND2 NAND2_213(.VSS(VSS),.VDD(VDD),.Y(I5006),.A(g421),.B(I5005));
  NAND2 NAND2_214(.VSS(VSS),.VDD(VDD),.Y(I12128),.A(g170),.B(I12126));
  NAND2 NAND2_215(.VSS(VSS),.VDD(VDD),.Y(I5105),.A(g431),.B(I5104));
  NAND2 NAND2_216(.VSS(VSS),.VDD(VDD),.Y(I6323),.A(g2050),.B(I6322));
  NAND2 NAND2_217(.VSS(VSS),.VDD(VDD),.Y(g7588),.A(I12093),.B(I12094));
  NAND2 NAND2_218(.VSS(VSS),.VDD(VDD),.Y(I6666),.A(g2776),.B(I6664));
  NAND2 NAND2_219(.VSS(VSS),.VDD(VDD),.Y(g3623),.A(I6761),.B(I6762));
  NAND2 NAND2_220(.VSS(VSS),.VDD(VDD),.Y(I5373),.A(g976),.B(I5371));
  NAND2 NAND2_221(.VSS(VSS),.VDD(VDD),.Y(I8529),.A(g481),.B(I8527));
  NAND2 NAND2_222(.VSS(VSS),.VDD(VDD),.Y(I5283),.A(g758),.B(I5282));
  NAND2 NAND2_223(.VSS(VSS),.VDD(VDD),.Y(I7224),.A(g2981),.B(I7223));
  NAND2 NAND2_224(.VSS(VSS),.VDD(VDD),.Y(I5007),.A(g312),.B(I5005));
  NAND2 NAND2_225(.VSS(VSS),.VDD(VDD),.Y(I5459),.A(g1240),.B(g1003));
  NAND2 NAND2_226(.VSS(VSS),.VDD(VDD),.Y(I17297),.A(g11369),.B(I17295));
  NAND3 NAND3_3(.VSS(VSS),.VDD(VDD),.Y(g8746),.A(g8617),.B(g6517),.C(g6509));
  NAND2 NAND2_227(.VSS(VSS),.VDD(VDD),.Y(I6143),.A(g1976),.B(g646));
  NAND2 NAND2_228(.VSS(VSS),.VDD(VDD),.Y(I5015),.A(g1011),.B(I5013));
  NAND2 NAND2_229(.VSS(VSS),.VDD(VDD),.Y(g8932),.A(I14264),.B(I14265));
  NAND2 NAND2_230(.VSS(VSS),.VDD(VDD),.Y(I16073),.A(g845),.B(I16072));
  NAND2 NAND2_231(.VSS(VSS),.VDD(VDD),.Y(I6988),.A(g2760),.B(g986));
  NAND2 NAND2_232(.VSS(VSS),.VDD(VDD),.Y(g3205),.A(g1814),.B(g2571));
  NAND2 NAND2_233(.VSS(VSS),.VDD(VDD),.Y(I8652),.A(g778),.B(I8650));
  NAND2 NAND2_234(.VSS(VSS),.VDD(VDD),.Y(I9558),.A(g5598),.B(I9557));
  NAND2 NAND2_235(.VSS(VSS),.VDD(VDD),.Y(I5203),.A(g369),.B(I5202));
  NAND2 NAND2_236(.VSS(VSS),.VDD(VDD),.Y(g7533),.A(I11936),.B(I11937));
  NAND2 NAND2_237(.VSS(VSS),.VDD(VDD),.Y(g3634),.A(I6806),.B(I6807));
  NAND2 NAND2_238(.VSS(VSS),.VDD(VDD),.Y(I6792),.A(g2959),.B(g143));
  NAND2 NAND2_239(.VSS(VSS),.VDD(VDD),.Y(g3304),.A(I6468),.B(I6469));
  NAND2 NAND2_240(.VSS(VSS),.VDD(VDD),.Y(I12145),.A(g158),.B(I12143));
  NAND2 NAND2_241(.VSS(VSS),.VDD(VDD),.Y(g7596),.A(I12127),.B(I12128));
  NAND2 NAND2_242(.VSS(VSS),.VDD(VDD),.Y(I13302),.A(g8162),.B(I13300));
  NAND2 NAND2_243(.VSS(VSS),.VDD(VDD),.Y(I5502),.A(g1007),.B(I5500));
  NAND2 NAND2_244(.VSS(VSS),.VDD(VDD),.Y(I9574),.A(g5608),.B(g818));
  NAND2 NAND2_245(.VSS(VSS),.VDD(VDD),.Y(g3273),.A(I6448),.B(I6449));
  NAND2 NAND2_246(.VSS(VSS),.VDD(VDD),.Y(I8670),.A(g4831),.B(I8669));
  NAND2 NAND2_247(.VSS(VSS),.VDD(VDD),.Y(I7035),.A(g1868),.B(I7033));
  NAND2 NAND2_248(.VSS(VSS),.VDD(VDD),.Y(I15453),.A(g10051),.B(I15451));
  NAND2 NAND2_249(.VSS(VSS),.VDD(VDD),.Y(I8625),.A(g4267),.B(I8624));
  NAND2 NAND2_250(.VSS(VSS),.VDD(VDD),.Y(I7876),.A(g4109),.B(I7875));
  NAND2 NAND2_251(.VSS(VSS),.VDD(VDD),.Y(I14203),.A(g8825),.B(I14202));
  NAND2 NAND2_252(.VSS(VSS),.VDD(VDD),.Y(I15607),.A(g10149),.B(g10144));
  NAND2 NAND2_253(.VSS(VSS),.VDD(VDD),.Y(g2274),.A(I5324),.B(I5325));
  NAND2 NAND2_254(.VSS(VSS),.VDD(VDD),.Y(I8740),.A(g1121),.B(I8738));
  NAND2 NAND2_255(.VSS(VSS),.VDD(VDD),.Y(I17296),.A(g11373),.B(I17295));
  NAND2 NAND2_256(.VSS(VSS),.VDD(VDD),.Y(g10507),.A(g10434),.B(g5859));
  NAND2 NAND2_257(.VSS(VSS),.VDD(VDD),.Y(g2325),.A(g611),.B(g617));
  NAND2 NAND2_258(.VSS(VSS),.VDD(VDD),.Y(I8606),.A(g506),.B(I8604));
  NAND2 NAND2_259(.VSS(VSS),.VDD(VDD),.Y(I12087),.A(g1470),.B(I12085));
  NAND2 NAND2_260(.VSS(VSS),.VDD(VDD),.Y(I13249),.A(g1891),.B(I13248));
  NAND2 NAND2_261(.VSS(VSS),.VDD(VDD),.Y(I13248),.A(g1891),.B(g8148));
  NAND2 NAND2_262(.VSS(VSS),.VDD(VDD),.Y(I13552),.A(g668),.B(g8262));
  NAND2 NAND2_263(.VSS(VSS),.VDD(VDD),.Y(g2106),.A(I4979),.B(I4980));
  NAND2 NAND2_264(.VSS(VSS),.VDD(VDD),.Y(I12069),.A(g139),.B(I12067));
  NAND2 NAND2_265(.VSS(VSS),.VDD(VDD),.Y(g9204),.A(g6019),.B(g8942));
  NAND2 NAND2_266(.VSS(VSS),.VDD(VDD),.Y(I12068),.A(g7116),.B(I12067));
  NAND2 NAND2_267(.VSS(VSS),.VDD(VDD),.Y(I17503),.A(g11475),.B(g7603));
  NAND2 NAND2_268(.VSS(VSS),.VDD(VDD),.Y(I7877),.A(g810),.B(I7875));
  NAND2 NAND2_269(.VSS(VSS),.VDD(VDD),.Y(I5165),.A(g1508),.B(I5164));
  NAND2 NAND2_270(.VSS(VSS),.VDD(VDD),.Y(g6740),.A(g6131),.B(g2550));
  NAND2 NAND2_271(.VSS(VSS),.VDD(VDD),.Y(I6289),.A(g981),.B(I6287));
  NAND2 NAND2_272(.VSS(VSS),.VDD(VDD),.Y(I6777),.A(g2892),.B(g650));
  NAND2 NAND2_273(.VSS(VSS),.VDD(VDD),.Y(g5171),.A(I8562),.B(I8563));
  NAND2 NAND2_274(.VSS(VSS),.VDD(VDD),.Y(I15891),.A(g853),.B(I15890));
  NAND2 NAND2_275(.VSS(VSS),.VDD(VDD),.Y(I13090),.A(g8006),.B(I13089));
  NAND2 NAND2_276(.VSS(VSS),.VDD(VDD),.Y(g11474),.A(I17460),.B(I17461));
  NAND4 NAND4_7(.VSS(VSS),.VDD(VDD),.Y(g7942),.A(g7395),.B(g6847),.C(g7380),.D(g7369));
  NAND2 NAND2_277(.VSS(VSS),.VDD(VDD),.Y(I5538),.A(g1270),.B(g1023));
  NAND2 NAND2_278(.VSS(VSS),.VDD(VDD),.Y(I7563),.A(g3533),.B(I7562));
  NAND2 NAND2_279(.VSS(VSS),.VDD(VDD),.Y(I13513),.A(g686),.B(g8248));
  NAND2 NAND2_280(.VSS(VSS),.VDD(VDD),.Y(g2107),.A(I4986),.B(I4987));
  NAND2 NAND2_281(.VSS(VSS),.VDD(VDD),.Y(g2223),.A(I5203),.B(I5204));
  NAND2 NAND2_282(.VSS(VSS),.VDD(VDD),.Y(I13505),.A(g677),.B(I13504));
  NAND2 NAND2_283(.VSS(VSS),.VDD(VDD),.Y(I6209),.A(g802),.B(I6207));
  NAND2 NAND2_284(.VSS(VSS),.VDD(VDD),.Y(I12086),.A(g6980),.B(I12085));
  NAND2 NAND2_285(.VSS(VSS),.VDD(VDD),.Y(I8545),.A(g486),.B(I8543));
  NAND2 NAND2_286(.VSS(VSS),.VDD(VDD),.Y(I8180),.A(g1786),.B(I8178));
  NAND2 NAND2_287(.VSS(VSS),.VDD(VDD),.Y(g2115),.A(I5014),.B(I5015));
  NAND2 NAND2_288(.VSS(VSS),.VDD(VDD),.Y(I8591),.A(g501),.B(I8589));
  NAND2 NAND2_289(.VSS(VSS),.VDD(VDD),.Y(I10931),.A(g6395),.B(I10930));
  NAND2 NAND2_290(.VSS(VSS),.VDD(VDD),.Y(I17402),.A(g11416),.B(I17400));
  NAND2 NAND2_291(.VSS(VSS),.VDD(VDD),.Y(g8307),.A(I13294),.B(I13295));
  NAND2 NAND2_292(.VSS(VSS),.VDD(VDD),.Y(I12144),.A(g7089),.B(I12143));
  NAND2 NAND2_293(.VSS(VSS),.VDD(VDD),.Y(I10520),.A(g6231),.B(I10519));
  NAND2 NAND2_294(.VSS(VSS),.VDD(VDD),.Y(I5263),.A(g456),.B(g461));
  NAND2 NAND2_295(.VSS(VSS),.VDD(VDD),.Y(g8757),.A(g8599),.B(g4401));
  NAND2 NAND2_296(.VSS(VSS),.VDD(VDD),.Y(I6714),.A(g2961),.B(g201));
  NAND2 NAND2_297(.VSS(VSS),.VDD(VDD),.Y(I14211),.A(g599),.B(I14209));
  NAND2 NAND2_298(.VSS(VSS),.VDD(VDD),.Y(I8515),.A(g3513),.B(I8513));
  NAND2 NAND2_299(.VSS(VSS),.VDD(VDD),.Y(g2272),.A(I5316),.B(I5317));
  NAND2 NAND2_300(.VSS(VSS),.VDD(VDD),.Y(I9946),.A(g5233),.B(g1796));
  NAND2 NAND2_301(.VSS(VSS),.VDD(VDD),.Y(I8750),.A(g4613),.B(g1125));
  NAND2 NAND2_302(.VSS(VSS),.VDD(VDD),.Y(I5605),.A(g1149),.B(I5604));
  NAND2 NAND2_303(.VSS(VSS),.VDD(VDD),.Y(g8880),.A(I14203),.B(I14204));
  NAND2 NAND2_304(.VSS(VSS),.VDD(VDD),.Y(I16051),.A(g837),.B(g10371));
  NAND2 NAND2_305(.VSS(VSS),.VDD(VDD),.Y(I16072),.A(g845),.B(g10373));
  NAND2 NAND2_306(.VSS(VSS),.VDD(VDD),.Y(g10440),.A(g10360),.B(g6037));
  NAND2 NAND2_307(.VSS(VSS),.VDD(VDD),.Y(g8612),.A(I13858),.B(I13859));
  NAND2 NAND2_308(.VSS(VSS),.VDD(VDD),.Y(I15872),.A(g2713),.B(I15870));
  NAND2 NAND2_309(.VSS(VSS),.VDD(VDD),.Y(I8528),.A(g4879),.B(I8527));
  NAND2 NAND2_310(.VSS(VSS),.VDD(VDD),.Y(g8629),.A(I13901),.B(I13902));
  NAND4 NAND4_8(.VSS(VSS),.VDD(VDD),.Y(g8542),.A(g2571),.B(g1828),.C(g1814),.D(g8390));
  NAND2 NAND2_311(.VSS(VSS),.VDD(VDD),.Y(I9947),.A(g5233),.B(I9946));
  NAND2 NAND2_312(.VSS(VSS),.VDD(VDD),.Y(I6838),.A(g806),.B(I6836));
  NAND2 NAND2_313(.VSS(VSS),.VDD(VDD),.Y(g7583),.A(I12068),.B(I12069));
  NAND2 NAND2_314(.VSS(VSS),.VDD(VDD),.Y(g4803),.A(g3664),.B(g2356));
  NAND2 NAND2_315(.VSS(VSS),.VDD(VDD),.Y(I17307),.A(g11377),.B(I17305));
  NAND2 NAND2_316(.VSS(VSS),.VDD(VDD),.Y(g4538),.A(g3475),.B(g2399));
  NAND2 NAND2_317(.VSS(VSS),.VDD(VDD),.Y(I15452),.A(g10058),.B(I15451));
  NAND2 NAND2_318(.VSS(VSS),.VDD(VDD),.Y(I13857),.A(g8538),.B(g1448));
  NAND2 NAND2_319(.VSS(VSS),.VDD(VDD),.Y(I14202),.A(g8825),.B(g591));
  NAND2 NAND2_320(.VSS(VSS),.VDD(VDD),.Y(I13765),.A(g731),.B(g8417));
  NAND2 NAND2_321(.VSS(VSS),.VDD(VDD),.Y(g2260),.A(I5296),.B(I5297));
  NAND4 NAND4_9(.VSS(VSS),.VDD(VDD),.Y(g7986),.A(g7011),.B(g6995),.C(g6984),.D(g7550));
  NAND2 NAND2_322(.VSS(VSS),.VDD(VDD),.Y(g5226),.A(I8670),.B(I8671));
  NAND2 NAND2_323(.VSS(VSS),.VDD(VDD),.Y(g8512),.A(g3723),.B(g8366));
  NAND2 NAND2_324(.VSS(VSS),.VDD(VDD),.Y(I16046),.A(g10370),.B(I16044));
  NAND2 NAND2_325(.VSS(VSS),.VDD(VDD),.Y(I13504),.A(g677),.B(g8247));
  NAND2 NAND2_326(.VSS(VSS),.VDD(VDD),.Y(g10447),.A(g10363),.B(g5360));
  NAND2 NAND2_327(.VSS(VSS),.VDD(VDD),.Y(g2167),.A(I5105),.B(I5106));
  NAND2 NAND2_328(.VSS(VSS),.VDD(VDD),.Y(I8804),.A(g4677),.B(I8803));
  NAND2 NAND2_329(.VSS(VSS),.VDD(VDD),.Y(g10472),.A(I16016),.B(I16017));
  NAND2 NAND2_330(.VSS(VSS),.VDD(VDD),.Y(I17487),.A(g11474),.B(I17485));
  NAND2 NAND2_331(.VSS(VSS),.VDD(VDD),.Y(I4995),.A(g416),.B(g309));
  NAND2 NAND2_332(.VSS(VSS),.VDD(VDD),.Y(I12093),.A(g6944),.B(I12092));
  NAND4 NAND4_10(.VSS(VSS),.VDD(VDD),.Y(g7987),.A(g7011),.B(g6995),.C(g7562),.D(g6974));
  NAND2 NAND2_333(.VSS(VSS),.VDD(VDD),.Y(g5227),.A(I8677),.B(I8678));
  NAND2 NAND2_334(.VSS(VSS),.VDD(VDD),.Y(I5126),.A(g1386),.B(g1389));
  NAND2 NAND2_335(.VSS(VSS),.VDD(VDD),.Y(g2321),.A(I5372),.B(I5373));
  NAND2 NAND2_336(.VSS(VSS),.VDD(VDD),.Y(g7547),.A(I11974),.B(I11975));
  NAND2 NAND2_337(.VSS(VSS),.VDD(VDD),.Y(I17306),.A(g11381),.B(I17305));
  NAND3 NAND3_4(.VSS(VSS),.VDD(VDD),.Y(g6548),.A(g6132),.B(g6124),.C(g6122));
  NAND2 NAND2_338(.VSS(VSS),.VDD(VDD),.Y(I11995),.A(g7107),.B(g127));
  NAND2 NAND2_339(.VSS(VSS),.VDD(VDD),.Y(I7225),.A(g1781),.B(I7223));
  NAND2 NAND2_340(.VSS(VSS),.VDD(VDD),.Y(I11261),.A(g6775),.B(g826));
  NAND3 NAND3_5(.VSS(VSS),.VDD(VDD),.Y(g8843),.A(g8542),.B(g8757),.C(g8545));
  NAND2 NAND2_341(.VSS(VSS),.VDD(VDD),.Y(g2938),.A(I6110),.B(I6111));
  NAND2 NAND2_342(.VSS(VSS),.VDD(VDD),.Y(I4942),.A(g396),.B(I4941));
  NAND2 NAND2_343(.VSS(VSS),.VDD(VDD),.Y(g10394),.A(I15899),.B(I15900));
  NAND2 NAND2_344(.VSS(VSS),.VDD(VDD),.Y(g8549),.A(g5527),.B(g8390));
  NAND2 NAND2_345(.VSS(VSS),.VDD(VDD),.Y(g3070),.A(g2016),.B(g1206));
  NAND2 NAND2_346(.VSS(VSS),.VDD(VDD),.Y(I4954),.A(g401),.B(g327));
  NAND2 NAND2_347(.VSS(VSS),.VDD(VDD),.Y(I5023),.A(g995),.B(g1275));
  NAND2 NAND2_348(.VSS(VSS),.VDD(VDD),.Y(g10446),.A(g10443),.B(g5350));
  NAND2 NAND2_349(.VSS(VSS),.VDD(VDD),.Y(I16081),.A(g10374),.B(I16079));
  NAND2 NAND2_350(.VSS(VSS),.VDD(VDD),.Y(I8641),.A(g4278),.B(I8640));
  NAND2 NAND2_351(.VSS(VSS),.VDD(VDD),.Y(I6178),.A(g197),.B(I6176));
  NAND2 NAND2_352(.VSS(VSS),.VDD(VDD),.Y(I12075),.A(g7098),.B(I12074));
  NAND2 NAND2_353(.VSS(VSS),.VDD(VDD),.Y(I5127),.A(g1386),.B(I5126));
  NAND2 NAND2_354(.VSS(VSS),.VDD(VDD),.Y(I5451),.A(g991),.B(I5449));
  NAND2 NAND2_355(.VSS(VSS),.VDD(VDD),.Y(g4168),.A(I7322),.B(I7323));
  NAND2 NAND2_356(.VSS(VSS),.VDD(VDD),.Y(I6288),.A(g2091),.B(I6287));
  NAND2 NAND2_357(.VSS(VSS),.VDD(VDD),.Y(I8179),.A(g3685),.B(I8178));
  NAND2 NAND2_358(.VSS(VSS),.VDD(VDD),.Y(I4912),.A(g318),.B(I4910));
  NAND2 NAND2_359(.VSS(VSS),.VDD(VDD),.Y(I6805),.A(g3268),.B(g471));
  NAND3 NAND3_6(.VSS(VSS),.VDD(VDD),.Y(g3766),.A(g2439),.B(g3222),.C(g2493));
  NAND2 NAND2_360(.VSS(VSS),.VDD(VDD),.Y(g3087),.A(I6288),.B(I6289));
  NAND2 NAND2_361(.VSS(VSS),.VDD(VDD),.Y(I17486),.A(g11384),.B(I17485));
  NAND2 NAND2_362(.VSS(VSS),.VDD(VDD),.Y(I4929),.A(g391),.B(I4928));
  NAND2 NAND2_363(.VSS(VSS),.VDD(VDD),.Y(I15890),.A(g853),.B(g10286));
  NAND2 NAND2_364(.VSS(VSS),.VDD(VDD),.Y(I16331),.A(g10616),.B(I16330));
  NAND2 NAND2_365(.VSS(VSS),.VDD(VDD),.Y(I9575),.A(g5608),.B(I9574));
  NAND2 NAND2_366(.VSS(VSS),.VDD(VDD),.Y(I13887),.A(g8532),.B(I13886));
  NAND2 NAND2_367(.VSS(VSS),.VDD(VDD),.Y(g5308),.A(I8787),.B(I8788));
  NAND2 NAND2_368(.VSS(VSS),.VDD(VDD),.Y(I13529),.A(g704),.B(g8253));
  NAND2 NAND2_369(.VSS(VSS),.VDD(VDD),.Y(I6208),.A(g2534),.B(I6207));
  NAND2 NAND2_370(.VSS(VSS),.VDD(VDD),.Y(g5217),.A(I8641),.B(I8642));
  NAND2 NAND2_371(.VSS(VSS),.VDD(VDD),.Y(I5316),.A(g1032),.B(I5315));
  NAND2 NAND2_372(.VSS(VSS),.VDD(VDD),.Y(g2111),.A(I5006),.B(I5007));
  NAND2 NAND2_373(.VSS(VSS),.VDD(VDD),.Y(g10366),.A(g10285),.B(g5392));
  NAND2 NAND2_374(.VSS(VSS),.VDD(VDD),.Y(I5034),.A(g1015),.B(g1019));
  NAND2 NAND2_375(.VSS(VSS),.VDD(VDD),.Y(I13869),.A(g1403),.B(I13867));
  NAND2 NAND2_376(.VSS(VSS),.VDD(VDD),.Y(I13868),.A(g8523),.B(I13867));
  NAND2 NAND2_377(.VSS(VSS),.VDD(VDD),.Y(I15999),.A(g10423),.B(g2683));
  NAND2 NAND2_378(.VSS(VSS),.VDD(VDD),.Y(I13259),.A(g1900),.B(I13258));
  NAND4 NAND4_11(.VSS(VSS),.VDD(VDD),.Y(g3261),.A(g2229),.B(g2222),.C(g2211),.D(g2202));
  NAND2 NAND2_379(.VSS(VSS),.VDD(VDD),.Y(g10481),.A(I16073),.B(I16074));
  NAND2 NAND2_380(.VSS(VSS),.VDD(VDD),.Y(g2180),.A(I5136),.B(I5137));
  NAND3 NAND3_7(.VSS(VSS),.VDD(VDD),.Y(g4976),.A(g2310),.B(g4604),.C(g3807));
  NAND2 NAND2_381(.VSS(VSS),.VDD(VDD),.Y(g8506),.A(g3475),.B(g8366));
  NAND2 NAND2_382(.VSS(VSS),.VDD(VDD),.Y(g2380),.A(I5460),.B(I5461));
  NAND2 NAND2_383(.VSS(VSS),.VDD(VDD),.Y(I13258),.A(g1900),.B(g8153));
  NAND2 NAND2_384(.VSS(VSS),.VDD(VDD),.Y(I5013),.A(g1007),.B(g1011));
  NAND2 NAND2_385(.VSS(VSS),.VDD(VDD),.Y(g5196),.A(I8605),.B(I8606));
  NAND2 NAND2_386(.VSS(VSS),.VDD(VDD),.Y(I10930),.A(g6395),.B(g5555));
  NAND2 NAND2_387(.VSS(VSS),.VDD(VDD),.Y(I6770),.A(g3257),.B(g382));
  NAND2 NAND2_388(.VSS(VSS),.VDD(VDD),.Y(g11449),.A(I17401),.B(I17402));
  NAND2 NAND2_389(.VSS(VSS),.VDD(VDD),.Y(g11448),.A(I17394),.B(I17395));
  NAND2 NAND2_390(.VSS(VSS),.VDD(VDD),.Y(I15717),.A(g10231),.B(I15716));
  NAND2 NAND2_391(.VSS(VSS),.VDD(VDD),.Y(I5317),.A(g1027),.B(I5315));
  NAND2 NAND2_392(.VSS(VSS),.VDD(VDD),.Y(I14210),.A(g8824),.B(I14209));
  NAND2 NAND2_393(.VSS(VSS),.VDD(VDD),.Y(I17569),.A(g1610),.B(I17567));
  NAND2 NAND2_394(.VSS(VSS),.VDD(VDD),.Y(I13878),.A(g1444),.B(I13876));
  NAND2 NAND2_395(.VSS(VSS),.VDD(VDD),.Y(g8545),.A(g3710),.B(g8390));
  NAND2 NAND2_396(.VSS(VSS),.VDD(VDD),.Y(g2515),.A(I5605),.B(I5606));
  NAND2 NAND2_397(.VSS(VSS),.VDD(VDD),.Y(I14443),.A(g8970),.B(I14442));
  NAND2 NAND2_398(.VSS(VSS),.VDD(VDD),.Y(g7557),.A(I11996),.B(I11997));
  NAND2 NAND2_399(.VSS(VSS),.VDD(VDD),.Y(g8180),.A(I13090),.B(I13091));
  NAND2 NAND2_400(.VSS(VSS),.VDD(VDD),.Y(I14279),.A(g1828),.B(I14277));
  NAND2 NAND2_401(.VSS(VSS),.VDD(VDD),.Y(I17568),.A(g11496),.B(I17567));
  NAND2 NAND2_402(.VSS(VSS),.VDD(VDD),.Y(I13886),.A(g8532),.B(g1440));
  NAND2 NAND2_403(.VSS(VSS),.VDD(VDD),.Y(I7322),.A(g3047),.B(I7321));
  NAND2 NAND2_404(.VSS(VSS),.VDD(VDD),.Y(I6990),.A(g986),.B(I6988));
  NAND2 NAND2_405(.VSS(VSS),.VDD(VDD),.Y(I14278),.A(g8847),.B(I14277));
  NAND2 NAND2_406(.VSS(VSS),.VDD(VDD),.Y(I7033),.A(g3089),.B(g1868));
  NAND2 NAND2_407(.VSS(VSS),.VDD(VDD),.Y(I9006),.A(g4492),.B(g1791));
  NAND2 NAND2_408(.VSS(VSS),.VDD(VDD),.Y(g8507),.A(g3738),.B(g8366));
  NAND2 NAND2_409(.VSS(VSS),.VDD(VDD),.Y(I5460),.A(g1240),.B(I5459));
  NAND2 NAND2_410(.VSS(VSS),.VDD(VDD),.Y(g4588),.A(g3440),.B(g2745));
  NAND2 NAND2_411(.VSS(VSS),.VDD(VDD),.Y(I4986),.A(g999),.B(I4985));
  NAND3 NAND3_8(.VSS(VSS),.VDD(VDD),.Y(g3247),.A(g1828),.B(g2564),.C(g2571));
  NAND2 NAND2_412(.VSS(VSS),.VDD(VDD),.Y(I8651),.A(g4824),.B(I8650));
  NAND2 NAND2_413(.VSS(VSS),.VDD(VDD),.Y(I13545),.A(g713),.B(I13544));
  NAND2 NAND2_414(.VSS(VSS),.VDD(VDD),.Y(g8628),.A(I13894),.B(I13895));
  NAND2 NAND2_415(.VSS(VSS),.VDD(VDD),.Y(I6138),.A(g378),.B(I6136));
  NAND2 NAND2_416(.VSS(VSS),.VDD(VDD),.Y(I12074),.A(g7098),.B(g174));
  NAND2 NAND2_417(.VSS(VSS),.VDD(VDD),.Y(g8630),.A(I13908),.B(I13909));
  NAND2 NAND2_418(.VSS(VSS),.VDD(VDD),.Y(I13078),.A(g7963),.B(I13076));
  NAND2 NAND2_419(.VSS(VSS),.VDD(VDD),.Y(I6109),.A(g2205),.B(g1494));
  NAND2 NAND2_420(.VSS(VSS),.VDD(VDD),.Y(g8300),.A(I13259),.B(I13260));
  NAND2 NAND2_421(.VSS(VSS),.VDD(VDD),.Y(I5501),.A(g1255),.B(I5500));
  NAND2 NAND2_422(.VSS(VSS),.VDD(VDD),.Y(I17586),.A(g11515),.B(I17584));
  NAND2 NAND2_423(.VSS(VSS),.VDD(VDD),.Y(I12092),.A(g6944),.B(g1490));
  NAND2 NAND2_424(.VSS(VSS),.VDD(VDD),.Y(I13901),.A(g8520),.B(I13900));
  NAND2 NAND2_425(.VSS(VSS),.VDD(VDD),.Y(I8795),.A(g4672),.B(g1145));
  NAND2 NAND2_426(.VSS(VSS),.VDD(VDD),.Y(I6201),.A(g766),.B(I6199));
  NAND2 NAND2_427(.VSS(VSS),.VDD(VDD),.Y(I14217),.A(g8826),.B(I14216));
  NAND2 NAND2_428(.VSS(VSS),.VDD(VDD),.Y(I9007),.A(g4492),.B(I9006));
  NAND2 NAND2_429(.VSS(VSS),.VDD(VDD),.Y(I13561),.A(g8263),.B(I13559));
  NAND2 NAND2_430(.VSS(VSS),.VDD(VDD),.Y(I15716),.A(g10231),.B(g10229));
  NAND2 NAND2_431(.VSS(VSS),.VDD(VDD),.Y(I6449),.A(g1776),.B(I6447));
  NAND2 NAND2_432(.VSS(VSS),.VDD(VDD),.Y(I13295),.A(g8161),.B(I13293));
  NAND2 NAND2_433(.VSS(VSS),.VDD(VDD),.Y(I4987),.A(g1003),.B(I4985));
  NAND2 NAND2_434(.VSS(VSS),.VDD(VDD),.Y(I6715),.A(g2961),.B(I6714));
  NAND2 NAND2_435(.VSS(VSS),.VDD(VDD),.Y(I17493),.A(g11475),.B(I17492));
  NAND2 NAND2_436(.VSS(VSS),.VDD(VDD),.Y(I12215),.A(g7061),.B(I12214));
  NAND2 NAND2_437(.VSS(VSS),.VDD(VDD),.Y(g2372),.A(I5450),.B(I5451));
  NAND2 NAND2_438(.VSS(VSS),.VDD(VDD),.Y(g7062),.A(I11262),.B(I11263));
  NAND2 NAND2_439(.VSS(VSS),.VDD(VDD),.Y(g2988),.A(I6225),.B(I6226));
  NAND2 NAND2_440(.VSS(VSS),.VDD(VDD),.Y(I13309),.A(g617),.B(I13307));
  NAND2 NAND2_441(.VSS(VSS),.VDD(VDD),.Y(g8839),.A(g8750),.B(g4401));
  NAND2 NAND2_442(.VSS(VSS),.VDD(VDD),.Y(g2555),.A(I5676),.B(I5677));
  NAND2 NAND2_443(.VSS(VSS),.VDD(VDD),.Y(g3662),.A(I6826),.B(I6827));
  NAND2 NAND2_444(.VSS(VSS),.VDD(VDD),.Y(I13308),.A(g8190),.B(I13307));
  NAND2 NAND2_445(.VSS(VSS),.VDD(VDD),.Y(g2792),.A(I5879),.B(I5880));
  NAND2 NAND2_446(.VSS(VSS),.VDD(VDD),.Y(g4117),.A(g3041),.B(g3061));
  NAND2 NAND2_447(.VSS(VSS),.VDD(VDD),.Y(I8543),.A(g4218),.B(g486));
  NAND2 NAND2_448(.VSS(VSS),.VDD(VDD),.Y(g11549),.A(I17585),.B(I17586));
  NAND2 NAND2_449(.VSS(VSS),.VDD(VDD),.Y(I6881),.A(g1351),.B(I6879));
  NAND2 NAND2_450(.VSS(VSS),.VDD(VDD),.Y(I12138),.A(g131),.B(I12136));
  NAND2 NAND2_451(.VSS(VSS),.VDD(VDD),.Y(I8729),.A(g4605),.B(I8728));
  NAND2 NAND2_452(.VSS(VSS),.VDD(VDD),.Y(I14216),.A(g8826),.B(g605));
  NAND2 NAND2_453(.VSS(VSS),.VDD(VDD),.Y(g10384),.A(I15871),.B(I15872));
  NAND2 NAND2_454(.VSS(VSS),.VDD(VDD),.Y(I13260),.A(g8153),.B(I13258));
  NAND2 NAND2_455(.VSS(VSS),.VDD(VDD),.Y(g2776),.A(I5866),.B(I5867));
  NAND2 NAND2_456(.VSS(VSS),.VDD(VDD),.Y(I8513),.A(g4873),.B(g3513));
  NAND2 NAND2_457(.VSS(VSS),.VDD(VDD),.Y(I13559),.A(g722),.B(g8263));
  NAND2 NAND2_458(.VSS(VSS),.VDD(VDD),.Y(I8178),.A(g3685),.B(g1786));
  NAND2 NAND2_459(.VSS(VSS),.VDD(VDD),.Y(g3631),.A(I6793),.B(I6794));
  NAND2 NAND2_460(.VSS(VSS),.VDD(VDD),.Y(I6487),.A(g2306),.B(g1227));
  NAND2 NAND2_461(.VSS(VSS),.VDD(VDD),.Y(I16080),.A(g849),.B(I16079));
  NAND2 NAND2_462(.VSS(VSS),.VDD(VDD),.Y(I13893),.A(g8529),.B(g1436));
  NAND2 NAND2_463(.VSS(VSS),.VDD(VDD),.Y(I12115),.A(g162),.B(I12113));
  NAND2 NAND2_464(.VSS(VSS),.VDD(VDD),.Y(I6748),.A(g1453),.B(I6746));
  NAND2 NAND2_465(.VSS(VSS),.VDD(VDD),.Y(I13544),.A(g713),.B(g8259));
  NAND2 NAND2_466(.VSS(VSS),.VDD(VDD),.Y(I5484),.A(g1250),.B(g1011));
  NAND2 NAND2_467(.VSS(VSS),.VDD(VDD),.Y(I4928),.A(g391),.B(g321));
  NAND2 NAND2_468(.VSS(VSS),.VDD(VDD),.Y(I6226),.A(g1346),.B(I6224));
  NAND2 NAND2_469(.VSS(VSS),.VDD(VDD),.Y(I8805),.A(g1113),.B(I8803));
  NAND2 NAND2_470(.VSS(VSS),.VDD(VDD),.Y(I4930),.A(g321),.B(I4928));
  NAND2 NAND2_471(.VSS(VSS),.VDD(VDD),.Y(I15880),.A(g2719),.B(I15878));
  NAND2 NAND2_472(.VSS(VSS),.VDD(VDD),.Y(I14265),.A(g1814),.B(I14263));
  NAND2 NAND2_473(.VSS(VSS),.VDD(VDD),.Y(I16031),.A(g829),.B(I16030));
  NAND2 NAND2_474(.VSS(VSS),.VDD(VDD),.Y(g3585),.A(I6747),.B(I6748));
  NAND4 NAND4_12(.VSS(VSS),.VDD(VDD),.Y(g3041),.A(g2364),.B(g2399),.C(g2374),.D(g2382));
  NAND2 NAND2_475(.VSS(VSS),.VDD(VDD),.Y(g8933),.A(I14271),.B(I14272));
  NAND2 NAND2_476(.VSS(VSS),.VDD(VDD),.Y(I16330),.A(g10616),.B(g4997));
  NAND2 NAND2_477(.VSS(VSS),.VDD(VDD),.Y(I13267),.A(g8154),.B(I13265));
  NAND2 NAND2_478(.VSS(VSS),.VDD(VDD),.Y(I13294),.A(g1882),.B(I13293));
  NAND2 NAND2_479(.VSS(VSS),.VDD(VDD),.Y(g10231),.A(I15616),.B(I15617));
  NAND2 NAND2_480(.VSS(VSS),.VDD(VDD),.Y(I14442),.A(g8970),.B(g1834));
  NAND2 NAND2_481(.VSS(VSS),.VDD(VDD),.Y(I6793),.A(g2959),.B(I6792));
  NAND2 NAND2_482(.VSS(VSS),.VDD(VDD),.Y(I4966),.A(g330),.B(I4964));
  NAND2 NAND2_483(.VSS(VSS),.VDD(VDD),.Y(I8752),.A(g1125),.B(I8750));
  NAND2 NAND2_484(.VSS(VSS),.VDD(VDD),.Y(I15432),.A(g10044),.B(I15430));
  NAND2 NAND2_485(.VSS(VSS),.VDD(VDD),.Y(I12214),.A(g7061),.B(g2518));
  NAND2 NAND2_486(.VSS(VSS),.VDD(VDD),.Y(g10511),.A(g10438),.B(g6032));
  NAND2 NAND2_487(.VSS(VSS),.VDD(VDD),.Y(g3011),.A(g591),.B(g2382));
  NAND2 NAND2_488(.VSS(VSS),.VDD(VDD),.Y(g5103),.A(I8480),.B(I8481));
  NAND2 NAND2_489(.VSS(VSS),.VDD(VDD),.Y(I16087),.A(g861),.B(I16086));
  NAND2 NAND2_490(.VSS(VSS),.VDD(VDD),.Y(g3734),.A(g3039),.B(g599));
  NAND2 NAND2_491(.VSS(VSS),.VDD(VDD),.Y(I6664),.A(g2792),.B(g2776));
  NAND2 NAND2_492(.VSS(VSS),.VDD(VDD),.Y(g8882),.A(I14217),.B(I14218));
  NAND2 NAND2_493(.VSS(VSS),.VDD(VDD),.Y(I4955),.A(g401),.B(I4954));
  NAND2 NAND2_494(.VSS(VSS),.VDD(VDD),.Y(I8786),.A(g4639),.B(g1141));
  NAND3 NAND3_9(.VSS(VSS),.VDD(VDD),.Y(g3992),.A(g2571),.B(g2550),.C(g2990));
  NAND2 NAND2_495(.VSS(VSS),.VDD(VDD),.Y(g10480),.A(I16066),.B(I16067));
  NAND2 NAND2_496(.VSS(VSS),.VDD(VDD),.Y(I11915),.A(g6935),.B(I11914));
  NAND2 NAND2_497(.VSS(VSS),.VDD(VDD),.Y(I8770),.A(g4619),.B(g1133));
  NAND2 NAND2_498(.VSS(VSS),.VDD(VDD),.Y(I5516),.A(g1260),.B(g1019));
  NAND2 NAND2_499(.VSS(VSS),.VDD(VDD),.Y(g8541),.A(g4001),.B(g8390));
  NAND2 NAND2_500(.VSS(VSS),.VDD(VDD),.Y(I6188),.A(g466),.B(I6186));
  NAND2 NAND2_501(.VSS(VSS),.VDD(VDD),.Y(g5147),.A(I8544),.B(I8545));
  NAND3 NAND3_10(.VSS(VSS),.VDD(VDD),.Y(g8744),.A(g8617),.B(g6509),.C(g6971));
  NAND2 NAND2_502(.VSS(VSS),.VDD(VDD),.Y(I5892),.A(g750),.B(I5891));
  NAND2 NAND2_503(.VSS(VSS),.VDD(VDD),.Y(g8558),.A(I13766),.B(I13767));
  NAND2 NAND2_504(.VSS(VSS),.VDD(VDD),.Y(I15258),.A(g9980),.B(I15256));
  NAND2 NAND2_505(.VSS(VSS),.VDD(VDD),.Y(I13266),.A(g1909),.B(I13265));
  NAND2 NAND2_506(.VSS(VSS),.VDD(VDD),.Y(I8787),.A(g4639),.B(I8786));
  NAND2 NAND2_507(.VSS(VSS),.VDD(VDD),.Y(I6826),.A(g3281),.B(I6825));
  NAND2 NAND2_508(.VSS(VSS),.VDD(VDD),.Y(I17283),.A(g11357),.B(I17281));
  NAND3 NAND3_11(.VSS(VSS),.VDD(VDD),.Y(g5013),.A(g4749),.B(g3247),.C(g3205));
  NAND2 NAND2_509(.VSS(VSS),.VDD(VDD),.Y(I17492),.A(g11475),.B(g3623));
  NAND2 NAND2_510(.VSS(VSS),.VDD(VDD),.Y(g8511),.A(g5277),.B(g8366));
  NAND2 NAND2_511(.VSS(VSS),.VDD(VDD),.Y(I16079),.A(g849),.B(g10374));
  NAND2 NAND2_512(.VSS(VSS),.VDD(VDD),.Y(I5035),.A(g1015),.B(I5034));
  NAND2 NAND2_513(.VSS(VSS),.VDD(VDD),.Y(I5517),.A(g1260),.B(I5516));
  NAND2 NAND2_514(.VSS(VSS),.VDD(VDD),.Y(I7223),.A(g2981),.B(g1781));
  NAND2 NAND2_515(.VSS(VSS),.VDD(VDD),.Y(I16086),.A(g861),.B(g10375));
  NAND2 NAND2_516(.VSS(VSS),.VDD(VDD),.Y(g5317),.A(I8796),.B(I8797));
  NAND2 NAND2_517(.VSS(VSS),.VDD(VDD),.Y(I15879),.A(g10359),.B(I15878));
  NAND2 NAND2_518(.VSS(VSS),.VDD(VDD),.Y(I15878),.A(g10359),.B(g2719));
  NAND2 NAND2_519(.VSS(VSS),.VDD(VDD),.Y(I12114),.A(g7093),.B(I12113));
  NAND2 NAND2_520(.VSS(VSS),.VDD(VDD),.Y(I12107),.A(g7113),.B(I12106));
  NAND2 NAND2_521(.VSS(VSS),.VDD(VDD),.Y(g2500),.A(g178),.B(g182));
  NAND2 NAND2_522(.VSS(VSS),.VDD(VDD),.Y(I15994),.A(g2677),.B(I15992));
  NAND4 NAND4_13(.VSS(VSS),.VDD(VDD),.Y(g7934),.A(g7395),.B(g6847),.C(g7279),.D(g7369));
  NAND2 NAND2_523(.VSS(VSS),.VDD(VDD),.Y(g10469),.A(g10430),.B(g5999));
  NAND2 NAND2_524(.VSS(VSS),.VDD(VDD),.Y(I14264),.A(g8843),.B(I14263));
  NAND2 NAND2_525(.VSS(VSS),.VDD(VDD),.Y(I6448),.A(g2264),.B(I6447));
  NAND2 NAND2_526(.VSS(VSS),.VDD(VDD),.Y(I13285),.A(g8159),.B(I13283));
  NAND2 NAND2_527(.VSS(VSS),.VDD(VDD),.Y(g10468),.A(I16000),.B(I16001));
  NAND2 NAND2_528(.VSS(VSS),.VDD(VDD),.Y(I6827),.A(g770),.B(I6825));
  NAND2 NAND2_529(.VSS(VSS),.VDD(VDD),.Y(g8623),.A(I13877),.B(I13878));
  NAND2 NAND2_530(.VSS(VSS),.VDD(VDD),.Y(I13900),.A(g8520),.B(g1428));
  NAND2 NAND2_531(.VSS(VSS),.VDD(VDD),.Y(g2795),.A(I5892),.B(I5893));
  NAND2 NAND2_532(.VSS(VSS),.VDD(VDD),.Y(I8575),.A(g4234),.B(g496));
  NAND2 NAND2_533(.VSS(VSS),.VDD(VDD),.Y(I14209),.A(g8824),.B(g599));
  NAND2 NAND2_534(.VSS(VSS),.VDD(VDD),.Y(I13560),.A(g722),.B(I13559));
  NAND2 NAND2_535(.VSS(VSS),.VDD(VDD),.Y(I8715),.A(g4601),.B(g4052));
  NAND2 NAND2_536(.VSS(VSS),.VDD(VDD),.Y(I8604),.A(g4259),.B(g506));
  NAND2 NAND2_537(.VSS(VSS),.VDD(VDD),.Y(I16017),.A(g2695),.B(I16015));
  NAND2 NAND2_538(.VSS(VSS),.VDD(VDD),.Y(I4941),.A(g396),.B(g324));
  NAND2 NAND2_539(.VSS(VSS),.VDD(VDD),.Y(g2205),.A(I5165),.B(I5166));
  NAND3 NAND3_12(.VSS(VSS),.VDD(VDD),.Y(g3753),.A(g2382),.B(g2364),.C(g2800));
  NAND2 NAND2_540(.VSS(VSS),.VDD(VDD),.Y(I6467),.A(g23),.B(g2479));
  NAND2 NAND2_541(.VSS(VSS),.VDD(VDD),.Y(I14614),.A(g611),.B(I14612));
  NAND2 NAND2_542(.VSS(VSS),.VDD(VDD),.Y(g2104),.A(I4965),.B(I4966));
  NAND2 NAND2_543(.VSS(VSS),.VDD(VDD),.Y(g2099),.A(I4942),.B(I4943));
  NAND2 NAND2_544(.VSS(VSS),.VDD(VDD),.Y(I16023),.A(g10426),.B(g2701));
  NAND2 NAND2_545(.VSS(VSS),.VDD(VDD),.Y(g10479),.A(I16059),.B(I16060));
  NAND3 NAND3_13(.VSS(VSS),.VDD(VDD),.Y(g8737),.A(g2317),.B(g4921),.C(g8688));
  NAND2 NAND2_546(.VSS(VSS),.VDD(VDD),.Y(g5942),.A(I9575),.B(I9576));
  NAND2 NAND2_547(.VSS(VSS),.VDD(VDD),.Y(g10478),.A(I16052),.B(I16053));
  NAND2 NAND2_548(.VSS(VSS),.VDD(VDD),.Y(I12004),.A(g153),.B(I12002));
  NAND2 NAND2_549(.VSS(VSS),.VDD(VDD),.Y(I4911),.A(g386),.B(I4910));
  NAND2 NAND2_550(.VSS(VSS),.VDD(VDD),.Y(I11914),.A(g6935),.B(g1494));
  NAND2 NAND2_551(.VSS(VSS),.VDD(VDD),.Y(g7960),.A(g7409),.B(g5573));
  NAND2 NAND2_552(.VSS(VSS),.VDD(VDD),.Y(I5295),.A(g794),.B(g798));
  NAND2 NAND2_553(.VSS(VSS),.VDD(VDD),.Y(I12106),.A(g7113),.B(g135));
  NAND2 NAND2_554(.VSS(VSS),.VDD(VDD),.Y(I8728),.A(g4605),.B(g1117));
  NAND2 NAND2_555(.VSS(VSS),.VDD(VDD),.Y(g3681),.A(I6837),.B(I6838));
  NAND2 NAND2_556(.VSS(VSS),.VDD(VDD),.Y(I11907),.A(g6967),.B(g1474));
  NAND2 NAND2_557(.VSS(VSS),.VDD(VDD),.Y(I13907),.A(g8526),.B(g1432));
  NAND2 NAND2_558(.VSS(VSS),.VDD(VDD),.Y(I8730),.A(g1117),.B(I8728));
  NAND2 NAND2_559(.VSS(VSS),.VDD(VDD),.Y(g8551),.A(g3967),.B(g8390));
  NAND2 NAND2_560(.VSS(VSS),.VDD(VDD),.Y(I4980),.A(g333),.B(I4978));
  NAND2 NAND2_561(.VSS(VSS),.VDD(VDD),.Y(g2961),.A(I6177),.B(I6178));
  NAND2 NAND2_562(.VSS(VSS),.VDD(VDD),.Y(g6019),.A(g617),.B(g4921));
  NAND2 NAND2_563(.VSS(VSS),.VDD(VDD),.Y(I16016),.A(g10425),.B(I16015));
  NAND2 NAND2_564(.VSS(VSS),.VDD(VDD),.Y(I11935),.A(g7004),.B(g1458));
  NAND2 NAND2_565(.VSS(VSS),.VDD(VDD),.Y(I8678),.A(g1027),.B(I8676));
  NAND2 NAND2_566(.VSS(VSS),.VDD(VDD),.Y(I17051),.A(g10923),.B(g11249));
  NAND2 NAND2_567(.VSS(VSS),.VDD(VDD),.Y(g4482),.A(I7864),.B(I7865));
  NAND2 NAND2_568(.VSS(VSS),.VDD(VDD),.Y(g7592),.A(I12107),.B(I12108));
  NAND2 NAND2_569(.VSS(VSS),.VDD(VDD),.Y(g3460),.A(I6665),.B(I6666));
  NAND4 NAND4_14(.VSS(VSS),.VDD(VDD),.Y(g7932),.A(g7395),.B(g6847),.C(g7279),.D(g7273));
  NAND2 NAND2_570(.VSS(VSS),.VDD(VDD),.Y(g7624),.A(I12215),.B(I12216));
  NAND4 NAND4_15(.VSS(VSS),.VDD(VDD),.Y(g7953),.A(g7395),.B(g7390),.C(g7380),.D(g7369));
  NAND2 NAND2_571(.VSS(VSS),.VDD(VDD),.Y(g8414),.A(I13553),.B(I13554));
  NAND2 NAND2_572(.VSS(VSS),.VDD(VDD),.Y(I6168),.A(g153),.B(I6166));
  NAND2 NAND2_573(.VSS(VSS),.VDD(VDD),.Y(I5229),.A(g182),.B(g148));
  NAND2 NAND2_574(.VSS(VSS),.VDD(VDD),.Y(I6772),.A(g382),.B(I6770));
  NAND2 NAND2_575(.VSS(VSS),.VDD(VDD),.Y(I16030),.A(g829),.B(g10368));
  NAND2 NAND2_576(.VSS(VSS),.VDD(VDD),.Y(I13284),.A(g1927),.B(I13283));
  NAND2 NAND2_577(.VSS(VSS),.VDD(VDD),.Y(I16065),.A(g10428),.B(g2765));
  NAND2 NAND2_578(.VSS(VSS),.VDD(VDD),.Y(g2947),.A(I6137),.B(I6138));
  NAND2 NAND2_579(.VSS(VSS),.VDD(VDD),.Y(I7321),.A(g3047),.B(g1231));
  NAND2 NAND2_580(.VSS(VSS),.VDD(VDD),.Y(g2437),.A(I5529),.B(I5530));
  NAND2 NAND2_581(.VSS(VSS),.VDD(VDD),.Y(g2102),.A(I4955),.B(I4956));
  NAND2 NAND2_582(.VSS(VSS),.VDD(VDD),.Y(I17282),.A(g11360),.B(I17281));
  NAND2 NAND2_583(.VSS(VSS),.VDD(VDD),.Y(I5620),.A(g1771),.B(I5618));
  NAND2 NAND2_584(.VSS(VSS),.VDD(VDD),.Y(I8664),.A(g476),.B(I8662));
  NAND2 NAND2_585(.VSS(VSS),.VDD(VDD),.Y(g7524),.A(I11915),.B(I11916));
  NAND2 NAND2_586(.VSS(VSS),.VDD(VDD),.Y(g7717),.A(g6863),.B(g3206));
  NAND2 NAND2_587(.VSS(VSS),.VDD(VDD),.Y(I16467),.A(g10716),.B(g10518));
  NAND2 NAND2_588(.VSS(VSS),.VDD(VDD),.Y(I4972),.A(g991),.B(I4971));
  NAND2 NAND2_589(.VSS(VSS),.VDD(VDD),.Y(I13554),.A(g8262),.B(I13552));
  NAND2 NAND2_590(.VSS(VSS),.VDD(VDD),.Y(I16037),.A(g10427),.B(g2707));
  NAND2 NAND2_591(.VSS(VSS),.VDD(VDD),.Y(g8302),.A(I13273),.B(I13274));
  NAND2 NAND2_592(.VSS(VSS),.VDD(VDD),.Y(I4943),.A(g324),.B(I4941));
  NAND2 NAND2_593(.VSS(VSS),.VDD(VDD),.Y(I5485),.A(g1250),.B(I5484));
  NAND2 NAND2_594(.VSS(VSS),.VDD(VDD),.Y(g5527),.A(g3978),.B(g4749));
  NAND2 NAND2_595(.VSS(VSS),.VDD(VDD),.Y(I10509),.A(g786),.B(I10507));
  NAND2 NAND2_596(.VSS(VSS),.VDD(VDD),.Y(g7599),.A(I12144),.B(I12145));
  NAND2 NAND2_597(.VSS(VSS),.VDD(VDD),.Y(I10508),.A(g6221),.B(I10507));
  NAND2 NAND2_598(.VSS(VSS),.VDD(VDD),.Y(I6126),.A(g1419),.B(I6124));
  NAND2 NAND2_599(.VSS(VSS),.VDD(VDD),.Y(I8671),.A(g814),.B(I8669));
  NAND2 NAND2_600(.VSS(VSS),.VDD(VDD),.Y(I6760),.A(g2943),.B(g1448));
  NAND2 NAND2_601(.VSS(VSS),.VDD(VDD),.Y(g3626),.A(I6778),.B(I6779));
  NAND2 NAND2_602(.VSS(VSS),.VDD(VDD),.Y(I11973),.A(g7001),.B(g1462));
  NAND2 NAND2_603(.VSS(VSS),.VDD(VDD),.Y(g2389),.A(I5469),.B(I5470));
  NAND2 NAND2_604(.VSS(VSS),.VDD(VDD),.Y(I15617),.A(g10153),.B(I15615));
  NAND2 NAND2_605(.VSS(VSS),.VDD(VDD),.Y(g5277),.A(g3734),.B(g4538));
  NAND2 NAND2_606(.VSS(VSS),.VDD(VDD),.Y(I5005),.A(g421),.B(g312));
  NAND2 NAND2_607(.VSS(VSS),.VDD(VDD),.Y(I6779),.A(g650),.B(I6777));
  NAND2 NAND2_608(.VSS(VSS),.VDD(VDD),.Y(I6665),.A(g2792),.B(I6664));
  NAND2 NAND2_609(.VSS(VSS),.VDD(VDD),.Y(I8589),.A(g4251),.B(g501));
  NAND2 NAND2_610(.VSS(VSS),.VDD(VDD),.Y(g8412),.A(I13545),.B(I13546));
  NAND2 NAND2_611(.VSS(VSS),.VDD(VDD),.Y(g2963),.A(I6187),.B(I6188));
  NAND2 NAND2_612(.VSS(VSS),.VDD(VDD),.Y(I12045),.A(g6951),.B(g1486));
  NAND2 NAND2_613(.VSS(VSS),.VDD(VDD),.Y(I16053),.A(g10371),.B(I16051));
  NAND2 NAND2_614(.VSS(VSS),.VDD(VDD),.Y(g2109),.A(I4996),.B(I4997));
  NAND2 NAND2_615(.VSS(VSS),.VDD(VDD),.Y(g11418),.A(I17306),.B(I17307));
  NAND2 NAND2_616(.VSS(VSS),.VDD(VDD),.Y(I13539),.A(g8157),.B(I13537));
  NAND2 NAND2_617(.VSS(VSS),.VDD(VDD),.Y(g10475),.A(I16031),.B(I16032));
  NAND2 NAND2_618(.VSS(VSS),.VDD(VDD),.Y(I5324),.A(g1336),.B(I5323));
  NAND2 NAND2_619(.VSS(VSS),.VDD(VDD),.Y(I13538),.A(g658),.B(I13537));
  NAND2 NAND2_620(.VSS(VSS),.VDD(VDD),.Y(I5469),.A(g1245),.B(I5468));
  NAND2 NAND2_621(.VSS(VSS),.VDD(VDD),.Y(I5540),.A(g1023),.B(I5538));
  NAND2 NAND2_622(.VSS(VSS),.VDD(VDD),.Y(I17505),.A(g7603),.B(I17503));
  NAND2 NAND2_623(.VSS(VSS),.VDD(VDD),.Y(I11241),.A(g6760),.B(g790));
  NAND2 NAND2_624(.VSS(VSS),.VDD(VDD),.Y(I8803),.A(g4677),.B(g1113));
  NAND2 NAND2_625(.VSS(VSS),.VDD(VDD),.Y(I12061),.A(g6961),.B(I12060));
  NAND2 NAND2_626(.VSS(VSS),.VDD(VDD),.Y(I8780),.A(g1137),.B(I8778));
  NAND3 NAND3_14(.VSS(VSS),.VDD(VDD),.Y(g8745),.A(g8617),.B(g6517),.C(g6964));
  NAND2 NAND2_627(.VSS(VSS),.VDD(VDD),.Y(I4979),.A(g411),.B(I4978));
  NAND2 NAND2_628(.VSS(VSS),.VDD(VDD),.Y(g8109),.A(g5052),.B(g7853));
  NAND2 NAND2_629(.VSS(VSS),.VDD(VDD),.Y(g8309),.A(I13308),.B(I13309));
  NAND2 NAND2_630(.VSS(VSS),.VDD(VDD),.Y(g6758),.A(I10770),.B(I10771));
  NAND2 NAND2_631(.VSS(VSS),.VDD(VDD),.Y(I16009),.A(g2689),.B(I16007));
  NAND2 NAND2_632(.VSS(VSS),.VDD(VDD),.Y(I15616),.A(g10043),.B(I15615));
  NAND2 NAND2_633(.VSS(VSS),.VDD(VDD),.Y(I8662),.A(g4286),.B(g476));
  NAND2 NAND2_634(.VSS(VSS),.VDD(VDD),.Y(I16008),.A(g10424),.B(I16007));
  NAND2 NAND2_635(.VSS(VSS),.VDD(VDD),.Y(I13515),.A(g8248),.B(I13513));
  NAND2 NAND2_636(.VSS(VSS),.VDD(VDD),.Y(I13991),.A(g622),.B(I13990));
  NAND2 NAND2_637(.VSS(VSS),.VDD(VDD),.Y(g11276),.A(I17052),.B(I17053));
  NAND2 NAND2_638(.VSS(VSS),.VDD(VDD),.Y(I15900),.A(g10287),.B(I15898));
  NAND2 NAND2_639(.VSS(VSS),.VDD(VDD),.Y(g2419),.A(I5501),.B(I5502));
  NAND2 NAND2_640(.VSS(VSS),.VDD(VDD),.Y(I16074),.A(g10373),.B(I16072));
  NAND2 NAND2_641(.VSS(VSS),.VDD(VDD),.Y(I10769),.A(g5944),.B(g1801));
  NAND2 NAND2_642(.VSS(VSS),.VDD(VDD),.Y(I7323),.A(g1231),.B(I7321));
  NAND2 NAND2_643(.VSS(VSS),.VDD(VDD),.Y(g7978),.A(g7697),.B(g3038));
  NAND2 NAND2_644(.VSS(VSS),.VDD(VDD),.Y(I7875),.A(g4109),.B(g810));
  NAND2 NAND2_645(.VSS(VSS),.VDD(VDD),.Y(I8562),.A(g4227),.B(I8561));
  NAND2 NAND2_646(.VSS(VSS),.VDD(VDD),.Y(I15892),.A(g10286),.B(I15890));
  NAND2 NAND2_647(.VSS(VSS),.VDD(VDD),.Y(g3771),.A(I6989),.B(I6990));
  NAND2 NAND2_648(.VSS(VSS),.VDD(VDD),.Y(I8605),.A(g4259),.B(I8604));
  NAND2 NAND2_649(.VSS(VSS),.VDD(VDD),.Y(g10153),.A(I15452),.B(I15453));
  NAND2 NAND2_650(.VSS(VSS),.VDD(VDD),.Y(g5295),.A(I8762),.B(I8763));
  NAND2 NAND2_651(.VSS(VSS),.VDD(VDD),.Y(I8751),.A(g4613),.B(I8750));
  NAND2 NAND2_652(.VSS(VSS),.VDD(VDD),.Y(I15907),.A(g6899),.B(I15906));
  NAND2 NAND2_653(.VSS(VSS),.VDD(VDD),.Y(I5136),.A(g521),.B(I5135));
  NAND2 NAND2_654(.VSS(VSS),.VDD(VDD),.Y(I11263),.A(g826),.B(I11261));
  NAND2 NAND2_655(.VSS(VSS),.VDD(VDD),.Y(I14204),.A(g591),.B(I14202));
  NAND2 NAND2_656(.VSS(VSS),.VDD(VDD),.Y(g8881),.A(I14210),.B(I14211));
  NAND2 NAND2_657(.VSS(VSS),.VDD(VDD),.Y(g2105),.A(I4972),.B(I4973));
  NAND3 NAND3_15(.VSS(VSS),.VDD(VDD),.Y(g5557),.A(g4538),.B(g3071),.C(g3011));
  NAND2 NAND2_658(.VSS(VSS),.VDD(VDD),.Y(I5230),.A(g182),.B(I5229));
  NAND2 NAND2_659(.VSS(VSS),.VDD(VDD),.Y(I8669),.A(g4831),.B(g814));
  NAND2 NAND2_660(.VSS(VSS),.VDD(VDD),.Y(g10474),.A(I16024),.B(I16025));
  NAND2 NAND2_661(.VSS(VSS),.VDD(VDD),.Y(I8772),.A(g1133),.B(I8770));
  NAND2 NAND2_662(.VSS(VSS),.VDD(VDD),.Y(g2445),.A(I5539),.B(I5540));
  NAND2 NAND2_663(.VSS(VSS),.VDD(VDD),.Y(g8006),.A(g5552),.B(g7717));
  NAND2 NAND2_664(.VSS(VSS),.VDD(VDD),.Y(I10932),.A(g5555),.B(I10930));
  NAND2 NAND2_665(.VSS(VSS),.VDD(VDD),.Y(I17504),.A(g11475),.B(I17503));
  NAND2 NAND2_666(.VSS(VSS),.VDD(VDD),.Y(I5137),.A(g525),.B(I5135));
  NAND2 NAND2_667(.VSS(VSS),.VDD(VDD),.Y(g8305),.A(I13284),.B(I13285));
  NAND2 NAND2_668(.VSS(VSS),.VDD(VDD),.Y(I5891),.A(g750),.B(g2057));
  NAND2 NAND2_669(.VSS(VSS),.VDD(VDD),.Y(I13273),.A(g1918),.B(I13272));
  NAND2 NAND2_670(.VSS(VSS),.VDD(VDD),.Y(I8480),.A(g4455),.B(I8479));
  NAND2 NAND2_671(.VSS(VSS),.VDD(VDD),.Y(g4144),.A(g2160),.B(g3044));
  NAND2 NAND2_672(.VSS(VSS),.VDD(VDD),.Y(I15906),.A(g6899),.B(g10302));
  NAND2 NAND2_673(.VSS(VSS),.VDD(VDD),.Y(I5342),.A(g315),.B(I5341));
  NAND2 NAND2_674(.VSS(VSS),.VDD(VDD),.Y(I13514),.A(g686),.B(I13513));
  NAND2 NAND2_675(.VSS(VSS),.VDD(VDD),.Y(g8407),.A(I13522),.B(I13523));
  NAND2 NAND2_676(.VSS(VSS),.VDD(VDD),.Y(g4088),.A(I7224),.B(I7225));
  NAND2 NAND2_677(.VSS(VSS),.VDD(VDD),.Y(g4488),.A(I7876),.B(I7877));
  NAND2 NAND2_678(.VSS(VSS),.VDD(VDD),.Y(g7598),.A(I12137),.B(I12138));
  NAND3 NAND3_16(.VSS(VSS),.VDD(VDD),.Y(g3222),.A(g2557),.B(g1814),.C(g1834));
  NAND2 NAND2_679(.VSS(VSS),.VDD(VDD),.Y(I16052),.A(g837),.B(I16051));
  NAND2 NAND2_680(.VSS(VSS),.VDD(VDD),.Y(I12127),.A(g7103),.B(I12126));
  NAND2 NAND2_681(.VSS(VSS),.VDD(VDD),.Y(g10483),.A(I16087),.B(I16088));
  NAND2 NAND2_682(.VSS(VSS),.VDD(VDD),.Y(g8415),.A(I13560),.B(I13561));
  NAND2 NAND2_683(.VSS(VSS),.VDD(VDD),.Y(g11415),.A(I17289),.B(I17290));
  NAND2 NAND2_684(.VSS(VSS),.VDD(VDD),.Y(g6573),.A(I10508),.B(I10509));
  NAND2 NAND2_685(.VSS(VSS),.VDD(VDD),.Y(I5676),.A(g1218),.B(I5675));
  NAND2 NAND2_686(.VSS(VSS),.VDD(VDD),.Y(I6778),.A(g2892),.B(I6777));
  NAND2 NAND2_687(.VSS(VSS),.VDD(VDD),.Y(g9413),.A(I14613),.B(I14614));
  NAND2 NAND2_688(.VSS(VSS),.VDD(VDD),.Y(I8779),.A(g4630),.B(I8778));
  NAND2 NAND2_689(.VSS(VSS),.VDD(VDD),.Y(I5592),.A(g1696),.B(I5591));
  NAND4 NAND4_16(.VSS(VSS),.VDD(VDD),.Y(g8502),.A(g2382),.B(g605),.C(g591),.D(g8366));
  NAND2 NAND2_690(.VSS(VSS),.VDD(VDD),.Y(I15609),.A(g10144),.B(I15607));
  NAND2 NAND2_691(.VSS(VSS),.VDD(VDD),.Y(I15608),.A(g10149),.B(I15607));
  NAND3 NAND3_17(.VSS(VSS),.VDD(VDD),.Y(g3071),.A(g605),.B(g2374),.C(g2382));
  NAND2 NAND2_692(.VSS(VSS),.VDD(VDD),.Y(g10509),.A(g10436),.B(g6023));
  NAND2 NAND2_693(.VSS(VSS),.VDD(VDD),.Y(I17461),.A(g11448),.B(I17459));
  NAND2 NAND2_694(.VSS(VSS),.VDD(VDD),.Y(I13506),.A(g8247),.B(I13504));
  NAND2 NAND2_695(.VSS(VSS),.VDD(VDD),.Y(I5468),.A(g1245),.B(g999));
  NAND2 NAND2_696(.VSS(VSS),.VDD(VDD),.Y(g5219),.A(I8651),.B(I8652));
  NAND2 NAND2_697(.VSS(VSS),.VDD(VDD),.Y(I5677),.A(g1223),.B(I5675));
  NAND3 NAND3_18(.VSS(VSS),.VDD(VDD),.Y(g8826),.A(g8739),.B(g8737),.C(g8648));
  NAND2 NAND2_698(.VSS(VSS),.VDD(VDD),.Y(I17393),.A(g11415),.B(g11414));
  NAND2 NAND2_699(.VSS(VSS),.VDD(VDD),.Y(I5866),.A(g2107),.B(I5865));
  NAND2 NAND2_700(.VSS(VSS),.VDD(VDD),.Y(I12126),.A(g7103),.B(g170));
  NAND2 NAND2_701(.VSS(VSS),.VDD(VDD),.Y(I4978),.A(g411),.B(g333));
  NAND2 NAND2_702(.VSS(VSS),.VDD(VDD),.Y(g7587),.A(I12086),.B(I12087));
  NAND2 NAND2_703(.VSS(VSS),.VDD(VDD),.Y(g5286),.A(I8751),.B(I8752));
  NAND2 NAND2_704(.VSS(VSS),.VDD(VDD),.Y(g8308),.A(I13301),.B(I13302));
  NAND2 NAND2_705(.VSS(VSS),.VDD(VDD),.Y(I7864),.A(g4099),.B(I7863));
  NAND2 NAND2_706(.VSS(VSS),.VDD(VDD),.Y(I11981),.A(g6957),.B(I11980));
  NAND2 NAND2_707(.VSS(VSS),.VDD(VDD),.Y(I12060),.A(g6961),.B(g1478));
  NAND2 NAND2_708(.VSS(VSS),.VDD(VDD),.Y(g5225),.A(I8663),.B(I8664));
  NAND2 NAND2_709(.VSS(VSS),.VDD(VDD),.Y(g11538),.A(I17568),.B(I17569));
  NAND2 NAND2_710(.VSS(VSS),.VDD(VDD),.Y(I13767),.A(g8417),.B(I13765));
  NAND2 NAND2_711(.VSS(VSS),.VDD(VDD),.Y(g10396),.A(I15907),.B(I15908));
  NAND2 NAND2_712(.VSS(VSS),.VDD(VDD),.Y(I11262),.A(g6775),.B(I11261));
  NAND2 NAND2_713(.VSS(VSS),.VDD(VDD),.Y(I13990),.A(g622),.B(g8688));
  NAND2 NAND2_714(.VSS(VSS),.VDD(VDD),.Y(I6224),.A(g2544),.B(g1346));
  NAND2 NAND2_715(.VSS(VSS),.VDD(VDD),.Y(I5867),.A(g2105),.B(I5865));
  NAND2 NAND2_716(.VSS(VSS),.VDD(VDD),.Y(g2493),.A(g1834),.B(g1840));
  NAND2 NAND2_717(.VSS(VSS),.VDD(VDD),.Y(I5893),.A(g2057),.B(I5891));
  NAND3 NAND3_19(.VSS(VSS),.VDD(VDD),.Y(g3062),.A(g2369),.B(g591),.C(g611));
  NAND2 NAND2_718(.VSS(VSS),.VDD(VDD),.Y(I13521),.A(g695),.B(g8249));
  NAND2 NAND2_719(.VSS(VSS),.VDD(VDD),.Y(I5186),.A(g1515),.B(I5184));
  NAND2 NAND2_720(.VSS(VSS),.VDD(VDD),.Y(I6771),.A(g3257),.B(I6770));
  NAND2 NAND2_721(.VSS(VSS),.VDD(VDD),.Y(I5325),.A(g1341),.B(I5323));
  NAND2 NAND2_722(.VSS(VSS),.VDD(VDD),.Y(I17459),.A(g11449),.B(g11448));
  NAND2 NAND2_723(.VSS(VSS),.VDD(VDD),.Y(I9557),.A(g5598),.B(g782));
  NAND2 NAND2_724(.VSS(VSS),.VDD(VDD),.Y(g11414),.A(I17282),.B(I17283));
  NAND2 NAND2_725(.VSS(VSS),.VDD(VDD),.Y(I12067),.A(g7116),.B(g139));
  NAND2 NAND2_726(.VSS(VSS),.VDD(VDD),.Y(I12094),.A(g1490),.B(I12092));
  NAND2 NAND2_727(.VSS(VSS),.VDD(VDD),.Y(I4964),.A(g406),.B(g330));
  NAND2 NAND2_728(.VSS(VSS),.VDD(VDD),.Y(I13272),.A(g1918),.B(g8158));
  NAND2 NAND2_729(.VSS(VSS),.VDD(VDD),.Y(I9948),.A(g1796),.B(I9946));
  NAND2 NAND2_730(.VSS(VSS),.VDD(VDD),.Y(g10302),.A(I15717),.B(I15718));
  NAND2 NAND2_731(.VSS(VSS),.VDD(VDD),.Y(I16332),.A(g4997),.B(I16330));
  NAND2 NAND2_732(.VSS(VSS),.VDD(VDD),.Y(I5106),.A(g435),.B(I5104));
  NAND2 NAND2_733(.VSS(VSS),.VDD(VDD),.Y(g8847),.A(g8760),.B(g8683));
  NAND2 NAND2_734(.VSS(VSS),.VDD(VDD),.Y(g2257),.A(I5283),.B(I5284));
  NAND2 NAND2_735(.VSS(VSS),.VDD(VDD),.Y(I12019),.A(g7119),.B(g166));
  NAND2 NAND2_736(.VSS(VSS),.VDD(VDD),.Y(I15441),.A(g10035),.B(g10122));
  NAND2 NAND2_737(.VSS(VSS),.VDD(VDD),.Y(I11997),.A(g127),.B(I11995));
  NAND2 NAND2_738(.VSS(VSS),.VDD(VDD),.Y(I8739),.A(g4607),.B(I8738));
  NAND2 NAND2_739(.VSS(VSS),.VDD(VDD),.Y(I5461),.A(g1003),.B(I5459));
  NAND2 NAND2_740(.VSS(VSS),.VDD(VDD),.Y(I13766),.A(g731),.B(I13765));
  NAND2 NAND2_741(.VSS(VSS),.VDD(VDD),.Y(I8479),.A(g4455),.B(g3530));
  NAND2 NAND2_742(.VSS(VSS),.VDD(VDD),.Y(I17295),.A(g11373),.B(g11369));
  NAND2 NAND2_743(.VSS(VSS),.VDD(VDD),.Y(I14271),.A(g8840),.B(I14270));
  NAND2 NAND2_744(.VSS(VSS),.VDD(VDD),.Y(I4971),.A(g991),.B(g995));
  NAND2 NAND2_745(.VSS(VSS),.VDD(VDD),.Y(g8301),.A(I13266),.B(I13267));
  NAND2 NAND2_746(.VSS(VSS),.VDD(VDD),.Y(I6110),.A(g2205),.B(I6109));
  NAND2 NAND2_747(.VSS(VSS),.VDD(VDD),.Y(g10482),.A(I16080),.B(I16081));
  NAND2 NAND2_748(.VSS(VSS),.VDD(VDD),.Y(g10779),.A(I16468),.B(I16469));
  NAND2 NAND2_749(.VSS(VSS),.VDD(VDD),.Y(I6762),.A(g1448),.B(I6760));
  NAND2 NAND2_750(.VSS(VSS),.VDD(VDD),.Y(I17289),.A(g11366),.B(I17288));
  NAND2 NAND2_751(.VSS(VSS),.VDD(VDD),.Y(I5315),.A(g1032),.B(g1027));
  NAND2 NAND2_752(.VSS(VSS),.VDD(VDD),.Y(I17288),.A(g11366),.B(g11363));
  NAND2 NAND2_753(.VSS(VSS),.VDD(VDD),.Y(I13859),.A(g1448),.B(I13857));
  NAND2 NAND2_754(.VSS(VSS),.VDD(VDD),.Y(g7548),.A(I11981),.B(I11982));
  NAND2 NAND2_755(.VSS(VSS),.VDD(VDD),.Y(I13858),.A(g8538),.B(I13857));
  NAND2 NAND2_756(.VSS(VSS),.VDD(VDD),.Y(I11996),.A(g7107),.B(I11995));
  NAND3 NAND3_20(.VSS(VSS),.VDD(VDD),.Y(g8743),.A(g8617),.B(g6971),.C(g6964));
  NAND2 NAND2_757(.VSS(VSS),.VDD(VDD),.Y(I5880),.A(g2115),.B(I5878));
  NAND2 NAND2_758(.VSS(VSS),.VDD(VDD),.Y(g10513),.A(g10441),.B(g5345));
  NAND2 NAND2_759(.VSS(VSS),.VDD(VDD),.Y(g8411),.A(I13538),.B(I13539));
  NAND2 NAND2_760(.VSS(VSS),.VDD(VDD),.Y(I8626),.A(g511),.B(I8624));
  NAND2 NAND2_761(.VSS(VSS),.VDD(VDD),.Y(g10505),.A(g10432),.B(g5938));
  NAND2 NAND2_762(.VSS(VSS),.VDD(VDD),.Y(I5612),.A(g1280),.B(I5611));
  NAND2 NAND2_763(.VSS(VSS),.VDD(VDD),.Y(g4821),.A(I8179),.B(I8180));
  NAND2 NAND2_764(.VSS(VSS),.VDD(VDD),.Y(I12076),.A(g174),.B(I12074));
  NAND2 NAND2_765(.VSS(VSS),.VDD(VDD),.Y(I12085),.A(g6980),.B(g1470));
  NAND2 NAND2_766(.VSS(VSS),.VDD(VDD),.Y(g7567),.A(I12020),.B(I12021));
  NAND2 NAND2_767(.VSS(VSS),.VDD(VDD),.Y(I5128),.A(g1389),.B(I5126));
  NAND2 NAND2_768(.VSS(VSS),.VDD(VDD),.Y(I6489),.A(g1227),.B(I6487));
  NAND2 NAND2_769(.VSS(VSS),.VDD(VDD),.Y(g7593),.A(I12114),.B(I12115));
  NAND2 NAND2_770(.VSS(VSS),.VDD(VDD),.Y(I8778),.A(g4630),.B(g1137));
  NAND2 NAND2_771(.VSS(VSS),.VDD(VDD),.Y(g10149),.A(I15442),.B(I15443));
  NAND2 NAND2_772(.VSS(VSS),.VDD(VDD),.Y(I13902),.A(g1428),.B(I13900));
  NAND2 NAND2_773(.VSS(VSS),.VDD(VDD),.Y(I13301),.A(g1936),.B(I13300));
  NAND2 NAND2_774(.VSS(VSS),.VDD(VDD),.Y(g3215),.A(g2564),.B(g1822));
  NAND4 NAND4_17(.VSS(VSS),.VDD(VDD),.Y(g7996),.A(g7011),.B(g7574),.C(g7562),.D(g6974));
  NAND2 NAND2_775(.VSS(VSS),.VDD(VDD),.Y(I4985),.A(g999),.B(g1003));
  NAND2 NAND2_776(.VSS(VSS),.VDD(VDD),.Y(I14444),.A(g1834),.B(I14442));
  NAND4 NAND4_18(.VSS(VSS),.VDD(VDD),.Y(g8000),.A(g7011),.B(g7574),.C(g7562),.D(g7550));
  NAND2 NAND2_777(.VSS(VSS),.VDD(VDD),.Y(I5166),.A(g1499),.B(I5164));
  NAND2 NAND2_778(.VSS(VSS),.VDD(VDD),.Y(I17460),.A(g11449),.B(I17459));
  NAND2 NAND2_779(.VSS(VSS),.VDD(VDD),.Y(g3008),.A(g2444),.B(g878));
  NAND2 NAND2_780(.VSS(VSS),.VDD(VDD),.Y(I6836),.A(g3287),.B(g806));
  NAND2 NAND2_781(.VSS(VSS),.VDD(VDD),.Y(I5529),.A(g1265),.B(I5528));
  NAND2 NAND2_782(.VSS(VSS),.VDD(VDD),.Y(g10229),.A(I15608),.B(I15609));
  NAND2 NAND2_783(.VSS(VSS),.VDD(VDD),.Y(I13661),.A(g8322),.B(I13659));
  NAND2 NAND2_784(.VSS(VSS),.VDD(VDD),.Y(I13895),.A(g1436),.B(I13893));
  NAND2 NAND2_785(.VSS(VSS),.VDD(VDD),.Y(g2303),.A(I5342),.B(I5343));
  NAND2 NAND2_786(.VSS(VSS),.VDD(VDD),.Y(I12039),.A(g6990),.B(I12038));
  NAND2 NAND2_787(.VSS(VSS),.VDD(VDD),.Y(g5592),.A(I9007),.B(I9008));
  NAND2 NAND2_788(.VSS(VSS),.VDD(VDD),.Y(I12038),.A(g6990),.B(g1466));
  NAND2 NAND2_789(.VSS(VSS),.VDD(VDD),.Y(g3322),.A(I6488),.B(I6489));
  NAND2 NAND2_790(.VSS(VSS),.VDD(VDD),.Y(I8561),.A(g4227),.B(g491));
  NAND2 NAND2_791(.VSS(VSS),.VDD(VDD),.Y(I8527),.A(g4879),.B(g481));
  NAND2 NAND2_792(.VSS(VSS),.VDD(VDD),.Y(I12143),.A(g7089),.B(g158));
  NAND2 NAND2_793(.VSS(VSS),.VDD(VDD),.Y(I5619),.A(g1766),.B(I5618));
  NAND2 NAND2_794(.VSS(VSS),.VDD(VDD),.Y(g10386),.A(I15879),.B(I15880));
  NAND2 NAND2_795(.VSS(VSS),.VDD(VDD),.Y(I11980),.A(g6957),.B(g1482));
  NAND2 NAND2_796(.VSS(VSS),.VDD(VDD),.Y(I6837),.A(g3287),.B(I6836));
  NAND2 NAND2_797(.VSS(VSS),.VDD(VDD),.Y(I4973),.A(g995),.B(I4971));
  NAND2 NAND2_798(.VSS(VSS),.VDD(VDD),.Y(I13888),.A(g1440),.B(I13886));
  NAND2 NAND2_799(.VSS(VSS),.VDD(VDD),.Y(g7558),.A(I12003),.B(I12004));
  NAND2 NAND2_800(.VSS(VSS),.VDD(VDD),.Y(I17494),.A(g3623),.B(I17492));
  NAND2 NAND2_801(.VSS(VSS),.VDD(VDD),.Y(g11491),.A(I17493),.B(I17494));
  NAND2 NAND2_802(.VSS(VSS),.VDD(VDD),.Y(I16045),.A(g833),.B(I16044));
  NAND2 NAND2_803(.VSS(VSS),.VDD(VDD),.Y(I7684),.A(g1023),.B(I7683));
  NAND2 NAND2_804(.VSS(VSS),.VDD(VDD),.Y(g4130),.A(g3044),.B(g2518));
  NAND2 NAND2_805(.VSS(VSS),.VDD(VDD),.Y(I8771),.A(g4619),.B(I8770));
  NAND2 NAND2_806(.VSS(VSS),.VDD(VDD),.Y(I13546),.A(g8259),.B(I13544));
  NAND2 NAND2_807(.VSS(VSS),.VDD(VDD),.Y(I13089),.A(g8006),.B(g1840));
  NAND2 NAND2_808(.VSS(VSS),.VDD(VDD),.Y(g2117),.A(I5024),.B(I5025));
  NAND2 NAND2_809(.VSS(VSS),.VDD(VDD),.Y(g5119),.A(I8514),.B(I8515));
  NAND2 NAND2_810(.VSS(VSS),.VDD(VDD),.Y(g5319),.A(I8804),.B(I8805));
  NAND2 NAND2_811(.VSS(VSS),.VDD(VDD),.Y(I15899),.A(g857),.B(I15898));
  NAND2 NAND2_812(.VSS(VSS),.VDD(VDD),.Y(I5606),.A(g1153),.B(I5604));
  NAND2 NAND2_813(.VSS(VSS),.VDD(VDD),.Y(I15898),.A(g857),.B(g10287));
  NAND2 NAND2_814(.VSS(VSS),.VDD(VDD),.Y(I16032),.A(g10368),.B(I16030));
  NAND2 NAND2_815(.VSS(VSS),.VDD(VDD),.Y(I17401),.A(g11418),.B(I17400));
  NAND2 NAND2_816(.VSS(VSS),.VDD(VDD),.Y(I13659),.A(g1945),.B(g8322));
  NAND2 NAND2_817(.VSS(VSS),.VDD(VDD),.Y(I8738),.A(g4607),.B(g1121));
  NAND2 NAND2_818(.VSS(VSS),.VDD(VDD),.Y(I13250),.A(g8148),.B(I13248));
  NAND2 NAND2_819(.VSS(VSS),.VDD(VDD),.Y(I15718),.A(g10229),.B(I15716));
  NAND2 NAND2_820(.VSS(VSS),.VDD(VDD),.Y(I9008),.A(g1791),.B(I9006));
  NAND2 NAND2_821(.VSS(VSS),.VDD(VDD),.Y(I6176),.A(g2177),.B(g197));
  NAND2 NAND2_822(.VSS(VSS),.VDD(VDD),.Y(I7865),.A(g774),.B(I7863));
  NAND2 NAND2_823(.VSS(VSS),.VDD(VDD),.Y(g5274),.A(I8729),.B(I8730));
  NAND2 NAND2_824(.VSS(VSS),.VDD(VDD),.Y(I5341),.A(g315),.B(g426));
  NAND2 NAND2_825(.VSS(VSS),.VDD(VDD),.Y(I17305),.A(g11381),.B(g11377));
  NAND2 NAND2_826(.VSS(VSS),.VDD(VDD),.Y(I17053),.A(g11249),.B(I17051));
  NAND2 NAND2_827(.VSS(VSS),.VDD(VDD),.Y(g5125),.A(I8528),.B(I8529));
  NAND2 NAND2_828(.VSS(VSS),.VDD(VDD),.Y(I12216),.A(g2518),.B(I12214));
  NAND2 NAND2_829(.VSS(VSS),.VDD(VDD),.Y(I6225),.A(g2544),.B(I6224));
  NAND2 NAND2_830(.VSS(VSS),.VDD(VDD),.Y(I5879),.A(g2120),.B(I5878));
  NAND2 NAND2_831(.VSS(VSS),.VDD(VDD),.Y(g3221),.A(g1834),.B(g2564));
  NAND2 NAND2_832(.VSS(VSS),.VDD(VDD),.Y(I14270),.A(g8840),.B(g1822));
  NAND2 NAND2_833(.VSS(VSS),.VDD(VDD),.Y(I6124),.A(g2215),.B(g1419));
  NAND2 NAND2_834(.VSS(VSS),.VDD(VDD),.Y(I6324),.A(g1864),.B(I6322));
  NAND2 NAND2_835(.VSS(VSS),.VDD(VDD),.Y(I13867),.A(g8523),.B(g1403));
  NAND2 NAND2_836(.VSS(VSS),.VDD(VDD),.Y(I13894),.A(g8529),.B(I13893));
  NAND2 NAND2_837(.VSS(VSS),.VDD(VDD),.Y(I6469),.A(g2479),.B(I6467));
  NAND2 NAND2_838(.VSS(VSS),.VDD(VDD),.Y(I8663),.A(g4286),.B(I8662));
  NAND2 NAND2_839(.VSS(VSS),.VDD(VDD),.Y(g7523),.A(I11908),.B(I11909));
  NAND2 NAND2_840(.VSS(VSS),.VDD(VDD),.Y(I6177),.A(g2177),.B(I6176));
  NAND2 NAND2_841(.VSS(VSS),.VDD(VDD),.Y(g5187),.A(I8590),.B(I8591));
  NAND2 NAND2_842(.VSS(VSS),.VDD(VDD),.Y(I6287),.A(g2091),.B(g981));
  NAND2 NAND2_843(.VSS(VSS),.VDD(VDD),.Y(I8762),.A(g4616),.B(I8761));
  NAND2 NAND2_844(.VSS(VSS),.VDD(VDD),.Y(I15871),.A(g10358),.B(I15870));
  NAND3 NAND3_21(.VSS(VSS),.VDD(VDD),.Y(g8840),.A(g8542),.B(g8541),.C(g8760));
  NAND2 NAND2_845(.VSS(VSS),.VDD(VDD),.Y(g2250),.A(I5264),.B(I5265));
  NAND2 NAND2_846(.VSS(VSS),.VDD(VDD),.Y(I8590),.A(g4251),.B(I8589));
  NAND2 NAND2_847(.VSS(VSS),.VDD(VDD),.Y(I6199),.A(g2525),.B(g766));
  NAND2 NAND2_848(.VSS(VSS),.VDD(VDD),.Y(I14218),.A(g605),.B(I14216));
  NAND2 NAND2_849(.VSS(VSS),.VDD(VDD),.Y(g8190),.A(g6027),.B(g7978));
  NAND2 NAND2_850(.VSS(VSS),.VDD(VDD),.Y(I5284),.A(g762),.B(I5282));
  NAND2 NAND2_851(.VSS(VSS),.VDD(VDD),.Y(I17485),.A(g11384),.B(g11474));
  NAND2 NAND2_852(.VSS(VSS),.VDD(VDD),.Y(I4965),.A(g406),.B(I4964));
  NAND2 NAND2_853(.VSS(VSS),.VDD(VDD),.Y(I5591),.A(g1696),.B(g1703));
  NAND2 NAND2_854(.VSS(VSS),.VDD(VDD),.Y(g8501),.A(g3760),.B(g8366));
  NAND2 NAND2_855(.VSS(VSS),.VDD(VDD),.Y(I15451),.A(g10058),.B(g10051));
  NAND2 NAND2_856(.VSS(VSS),.VDD(VDD),.Y(g8942),.A(g8823),.B(g4921));
  NAND2 NAND2_857(.VSS(VSS),.VDD(VDD),.Y(I13877),.A(g8535),.B(I13876));
  NAND2 NAND2_858(.VSS(VSS),.VDD(VDD),.Y(g7269),.A(I11509),.B(I11510));
  NAND2 NAND2_859(.VSS(VSS),.VDD(VDD),.Y(I4996),.A(g416),.B(I4995));
  NAND2 NAND2_860(.VSS(VSS),.VDD(VDD),.Y(I6144),.A(g1976),.B(I6143));
  NAND2 NAND2_861(.VSS(VSS),.VDD(VDD),.Y(I17567),.A(g11496),.B(g1610));
  NAND2 NAND2_862(.VSS(VSS),.VDD(VDD),.Y(g7572),.A(I12039),.B(I12040));
  NAND2 NAND2_863(.VSS(VSS),.VDD(VDD),.Y(I6207),.A(g2534),.B(g802));
  NAND2 NAND2_864(.VSS(VSS),.VDD(VDD),.Y(I14277),.A(g8847),.B(g1828));
  NAND2 NAND2_865(.VSS(VSS),.VDD(VDD),.Y(I16059),.A(g841),.B(I16058));
  NAND2 NAND2_866(.VSS(VSS),.VDD(VDD),.Y(I16025),.A(g2701),.B(I16023));
  NAND2 NAND2_867(.VSS(VSS),.VDD(VDD),.Y(I8563),.A(g491),.B(I8561));
  NAND2 NAND2_868(.VSS(VSS),.VDD(VDD),.Y(g3524),.A(g3209),.B(g3221));
  NAND2 NAND2_869(.VSS(VSS),.VDD(VDD),.Y(I16058),.A(g841),.B(g10372));
  NAND2 NAND2_870(.VSS(VSS),.VDD(VDD),.Y(I5204),.A(g374),.B(I5202));
  NAND2 NAND2_871(.VSS(VSS),.VDD(VDD),.Y(I6488),.A(g2306),.B(I6487));
  NAND4 NAND4_19(.VSS(VSS),.VDD(VDD),.Y(g3818),.A(g3056),.B(g3071),.C(g2310),.D(g3003));
  NAND2 NAND2_872(.VSS(VSS),.VDD(VDD),.Y(I16044),.A(g833),.B(g10370));
  NAND2 NAND2_873(.VSS(VSS),.VDD(VDD),.Y(g3717),.A(I6880),.B(I6881));
  NAND2 NAND2_874(.VSS(VSS),.VDD(VDD),.Y(I13077),.A(g1872),.B(I13076));
  NAND2 NAND2_875(.VSS(VSS),.VDD(VDD),.Y(g10043),.A(I15257),.B(I15258));
  NAND2 NAND2_876(.VSS(VSS),.VDD(VDD),.Y(I11280),.A(g6485),.B(I11278));
  NAND2 NAND2_877(.VSS(VSS),.VDD(VDD),.Y(I6825),.A(g3281),.B(g770));
  NAND2 NAND2_878(.VSS(VSS),.VDD(VDD),.Y(I4997),.A(g309),.B(I4995));
  NAND2 NAND2_879(.VSS(VSS),.VDD(VDD),.Y(I13300),.A(g1936),.B(g8162));
  NAND2 NAND2_880(.VSS(VSS),.VDD(VDD),.Y(I5323),.A(g1336),.B(g1341));
  NAND2 NAND2_881(.VSS(VSS),.VDD(VDD),.Y(I6136),.A(g2496),.B(g378));
  NAND2 NAND2_882(.VSS(VSS),.VDD(VDD),.Y(g5935),.A(I9558),.B(I9559));
  NAND2 NAND2_883(.VSS(VSS),.VDD(VDD),.Y(I5528),.A(g1265),.B(g1015));
  NAND2 NAND2_884(.VSS(VSS),.VDD(VDD),.Y(I6806),.A(g3268),.B(I6805));
  NAND2 NAND2_885(.VSS(VSS),.VDD(VDD),.Y(I5530),.A(g1015),.B(I5528));
  NAND2 NAND2_886(.VSS(VSS),.VDD(VDD),.Y(g10886),.A(g10807),.B(g10805));
  NAND2 NAND2_887(.VSS(VSS),.VDD(VDD),.Y(g3106),.A(I6323),.B(I6324));
  NAND2 NAND2_888(.VSS(VSS),.VDD(VDD),.Y(I13876),.A(g8535),.B(g1444));
  NAND2 NAND2_889(.VSS(VSS),.VDD(VDD),.Y(I6322),.A(g2050),.B(g1864));
  NAND2 NAND2_890(.VSS(VSS),.VDD(VDD),.Y(g3061),.A(g611),.B(g2374));
  NAND2 NAND2_891(.VSS(VSS),.VDD(VDD),.Y(g2439),.A(g1814),.B(g1828));
  NAND4 NAND4_20(.VSS(VSS),.VDD(VDD),.Y(g7947),.A(g7395),.B(g7390),.C(g7279),.D(g7369));
  NAND2 NAND2_892(.VSS(VSS),.VDD(VDD),.Y(I9576),.A(g818),.B(I9574));
  NAND2 NAND2_893(.VSS(VSS),.VDD(VDD),.Y(I13660),.A(g1945),.B(I13659));
  NAND2 NAND2_894(.VSS(VSS),.VDD(VDD),.Y(g3200),.A(g1822),.B(g2061));
  NAND2 NAND2_895(.VSS(VSS),.VDD(VDD),.Y(g4374),.A(I7684),.B(I7685));
  NAND2 NAND2_896(.VSS(VSS),.VDD(VDD),.Y(I11916),.A(g1494),.B(I11914));
  NAND2 NAND2_897(.VSS(VSS),.VDD(VDD),.Y(I5372),.A(g971),.B(I5371));
  NAND2 NAND2_898(.VSS(VSS),.VDD(VDD),.Y(g3003),.A(g599),.B(g2399));
  NAND2 NAND2_899(.VSS(VSS),.VDD(VDD),.Y(g8627),.A(I13887),.B(I13888));
  NAND2 NAND2_900(.VSS(VSS),.VDD(VDD),.Y(I5618),.A(g1766),.B(g1771));
  NAND2 NAND2_901(.VSS(VSS),.VDD(VDD),.Y(I6137),.A(g2496),.B(I6136));
  NAND2 NAND2_902(.VSS(VSS),.VDD(VDD),.Y(I5343),.A(g426),.B(I5341));
  NAND2 NAND2_903(.VSS(VSS),.VDD(VDD),.Y(I5282),.A(g758),.B(g762));
  NAND2 NAND2_904(.VSS(VSS),.VDD(VDD),.Y(I13307),.A(g8190),.B(g617));
  NAND2 NAND2_905(.VSS(VSS),.VDD(VDD),.Y(I13076),.A(g1872),.B(g7963));
  NAND2 NAND2_906(.VSS(VSS),.VDD(VDD),.Y(I6807),.A(g471),.B(I6805));
  NAND2 NAND2_907(.VSS(VSS),.VDD(VDD),.Y(I11243),.A(g790),.B(I11241));
  NAND2 NAND2_908(.VSS(VSS),.VDD(VDD),.Y(I17585),.A(g11354),.B(I17584));
  NAND2 NAND2_909(.VSS(VSS),.VDD(VDD),.Y(I12137),.A(g7110),.B(I12136));
  NAND2 NAND2_910(.VSS(VSS),.VDD(VDD),.Y(I7564),.A(g654),.B(I7562));
  NAND2 NAND2_911(.VSS(VSS),.VDD(VDD),.Y(g2970),.A(I6200),.B(I6201));
  NAND2 NAND2_912(.VSS(VSS),.VDD(VDD),.Y(g10144),.A(I15431),.B(I15432));
  NAND2 NAND2_913(.VSS(VSS),.VDD(VDD),.Y(I8788),.A(g1141),.B(I8786));
  NAND2 NAND2_914(.VSS(VSS),.VDD(VDD),.Y(g7054),.A(I11242),.B(I11243));
  NAND2 NAND2_915(.VSS(VSS),.VDD(VDD),.Y(I17052),.A(g10923),.B(I17051));
  NAND2 NAND2_916(.VSS(VSS),.VDD(VDD),.Y(g2120),.A(I5035),.B(I5036));
  NAND2 NAND2_917(.VSS(VSS),.VDD(VDD),.Y(g8616),.A(I13868),.B(I13869));
  NAND2 NAND2_918(.VSS(VSS),.VDD(VDD),.Y(I5202),.A(g369),.B(g374));
  NAND2 NAND2_919(.VSS(VSS),.VDD(VDD),.Y(I16088),.A(g10375),.B(I16086));
  NAND2 NAND2_920(.VSS(VSS),.VDD(VDD),.Y(I16024),.A(g10426),.B(I16023));
  NAND2 NAND2_921(.VSS(VSS),.VDD(VDD),.Y(g11490),.A(I17486),.B(I17487));
  NAND2 NAND2_922(.VSS(VSS),.VDD(VDD),.Y(I5518),.A(g1019),.B(I5516));
  NAND3 NAND3_22(.VSS(VSS),.VDD(VDD),.Y(g5118),.A(g2439),.B(g4806),.C(g4073));
  NAND2 NAND2_923(.VSS(VSS),.VDD(VDD),.Y(I12021),.A(g166),.B(I12019));
//
  NOR2 NOR2_0(.VSS(VSS),.VDD(VDD),.Y(g6392),.A(g5859),.B(g5938));
  NOR2 NOR2_1(.VSS(VSS),.VDD(VDD),.Y(g5938),.A(g2764),.B(g4988));
  NOR2 NOR2_2(.VSS(VSS),.VDD(VDD),.Y(g2478),.A(g1610),.B(g1737));
  NOR2 NOR2_3(.VSS(VSS),.VDD(VDD),.Y(g10374),.A(g10347),.B(g3463));
  NOR4 NOR4_0(.VSS(VSS),.VDD(VDD),.Y(g4278),.A(g3800),.B(g2593),.C(g2586),.D(g3776));
  NOR2 NOR2_4(.VSS(VSS),.VDD(VDD),.Y(g10424),.A(g10292),.B(g4620));
  NOR2 NOR2_5(.VSS(VSS),.VDD(VDD),.Y(g10383),.A(g10318),.B(g2998));
  NOR2 NOR2_6(.VSS(VSS),.VDD(VDD),.Y(g3118),.A(g2521),.B(g2514));
  NOR2 NOR2_7(.VSS(VSS),.VDD(VDD),.Y(g9815),.A(g9392),.B(g9367));
  NOR2 NOR2_8(.VSS(VSS),.VDD(VDD),.Y(g11077),.A(g10970),.B(g10971));
  NOR3 NOR3_0(.VSS(VSS),.VDD(VDD),.Y(g9746),.A(g9454),.B(g9274),.C(g9292));
  NOR3 NOR3_1(.VSS(VSS),.VDD(VDD),.Y(g3879),.A(g3141),.B(g2354),.C(g2353));
  NOR2 NOR2_9(.VSS(VSS),.VDD(VDD),.Y(g10285),.A(g10276),.B(g3566));
  NOR2 NOR2_10(.VSS(VSS),.VDD(VDD),.Y(g11480),.A(g11456),.B(g4567));
  NOR2 NOR2_11(.VSS(VSS),.VDD(VDD),.Y(g4076),.A(g1707),.B(g2864));
  NOR2 NOR2_12(.VSS(VSS),.VDD(VDD),.Y(g10570),.A(g10542),.B(g10324));
  NOR2 NOR2_13(.VSS(VSS),.VDD(VDD),.Y(g10239),.A(g9317),.B(g10179));
  NOR2 NOR2_14(.VSS(VSS),.VDD(VDD),.Y(g10594),.A(g10480),.B(g10521));
  NOR2 NOR2_15(.VSS(VSS),.VDD(VDD),.Y(g9426),.A(g9052),.B(g9030));
  NOR2 NOR2_16(.VSS(VSS),.VDD(VDD),.Y(g10382),.A(g10314),.B(g2998));
  NOR4 NOR4_1(.VSS(VSS),.VDD(VDD),.Y(g4672),.A(g3501),.B(g2669),.C(g2662),.D(g3479));
  NOR2 NOR2_17(.VSS(VSS),.VDD(VDD),.Y(g5360),.A(g2071),.B(g4225));
  NOR4 NOR4_2(.VSS(VSS),.VDD(VDD),.Y(g9387),.A(g9010),.B(g9240),.C(g9223),.D(I14596));
  NOR2 NOR2_18(.VSS(VSS),.VDD(VDD),.Y(g10438),.A(g10356),.B(g3566));
  NOR4 NOR4_3(.VSS(VSS),.VDD(VDD),.Y(g4613),.A(g3077),.B(g3491),.C(g2662),.D(g2655));
  NOR4 NOR4_4(.VSS(VSS),.VDD(VDD),.Y(g9391),.A(g9010),.B(g9240),.C(g9223),.D(I14602));
  NOR3 NOR3_2(.VSS(VSS),.VDD(VDD),.Y(g4572),.A(g3419),.B(g3408),.C(g3628));
  NOR3 NOR3_3(.VSS(VSS),.VDD(VDD),.Y(g9757),.A(g9454),.B(g9274),.C(g9292));
  NOR2 NOR2_19(.VSS(VSS),.VDD(VDD),.Y(g9416),.A(g9052),.B(g9030));
  NOR4 NOR4_5(.VSS(VSS),.VDD(VDD),.Y(g9874),.A(g9519),.B(g9536),.C(g9579),.D(I15033));
  NOR2 NOR2_20(.VSS(VSS),.VDD(VDD),.Y(g9654),.A(g9125),.B(g9173));
  NOR4 NOR4_6(.VSS(VSS),.VDD(VDD),.Y(g9880),.A(g9751),.B(g9536),.C(g9557),.D(I15051));
  NOR4 NOR4_7(.VSS(VSS),.VDD(VDD),.Y(g4873),.A(g3292),.B(g2593),.C(g2586),.D(g3776));
  NOR2 NOR2_21(.VSS(VSS),.VDD(VDD),.Y(g2807),.A(g22),.B(g2320));
  NOR2 NOR2_22(.VSS(VSS),.VDD(VDD),.Y(g10441),.A(g10351),.B(g3566));
  NOR4 NOR4_8(.VSS(VSS),.VDD(VDD),.Y(g4639),.A(g3501),.B(g2669),.C(g2662),.D(g2655));
  NOR2 NOR2_23(.VSS(VSS),.VDD(VDD),.Y(g10435),.A(g10332),.B(g3507));
  NOR2 NOR2_24(.VSS(VSS),.VDD(VDD),.Y(g10849),.A(g10739),.B(g3903));
  NOR4 NOR4_9(.VSS(VSS),.VDD(VDD),.Y(g9606),.A(g9125),.B(g9111),.C(g9173),.D(g9151));
  NOR4 NOR4_10(.VSS(VSS),.VDD(VDD),.Y(g9879),.A(g9747),.B(g9536),.C(g9566),.D(I15048));
  NOR2 NOR2_25(.VSS(VSS),.VDD(VDD),.Y(g9506),.A(g9052),.B(g9030));
  NOR2 NOR2_26(.VSS(VSS),.VDD(VDD),.Y(g6155),.A(g4974),.B(g2864));
  NOR2 NOR2_27(.VSS(VSS),.VDD(VDD),.Y(g6355),.A(g6032),.B(g6023));
  NOR2 NOR2_28(.VSS(VSS),.VDD(VDD),.Y(g9615),.A(g9052),.B(g9030));
  NOR2 NOR2_29(.VSS(VSS),.VDD(VDD),.Y(g10371),.A(g10344),.B(g3463));
  NOR2 NOR2_30(.VSS(VSS),.VDD(VDD),.Y(g9591),.A(g9125),.B(g9151));
  NOR2 NOR2_31(.VSS(VSS),.VDD(VDD),.Y(g10359),.A(g10227),.B(g4620));
  NOR2 NOR2_32(.VSS(VSS),.VDD(VDD),.Y(g10434),.A(g10352),.B(g3566));
  NOR2 NOR2_33(.VSS(VSS),.VDD(VDD),.Y(g10358),.A(g10226),.B(g4620));
  NOR3 NOR3_4(.VSS(VSS),.VDD(VDD),.Y(g9750),.A(g9454),.B(g9274),.C(g9292));
  NOR2 NOR2_34(.VSS(VSS),.VDD(VDD),.Y(g10291),.A(g10247),.B(g3113));
  NOR4 NOR4_11(.VSS(VSS),.VDD(VDD),.Y(g4227),.A(g3292),.B(g3793),.C(g2586),.D(g2579));
  NOR4 NOR4_12(.VSS(VSS),.VDD(VDD),.Y(g9655),.A(g9010),.B(g9240),.C(g9223),.D(I14776));
  NOR4 NOR4_13(.VSS(VSS),.VDD(VDD),.Y(g9410),.A(g9010),.B(g9240),.C(g9223),.D(I14607));
  NOR4 NOR4_14(.VSS(VSS),.VDD(VDD),.Y(g9667),.A(g9125),.B(g9111),.C(g9173),.D(g9151));
  NOR2 NOR2_35(.VSS(VSS),.VDD(VDD),.Y(g10563),.A(g10539),.B(g10322));
  NOR2 NOR2_36(.VSS(VSS),.VDD(VDD),.Y(g9776),.A(g9392),.B(g9367));
  NOR2 NOR2_37(.VSS(VSS),.VDD(VDD),.Y(g10324),.A(g9317),.B(g10244));
  NOR3 NOR3_5(.VSS(VSS),.VDD(VDD),.Y(g4455),.A(g3543),.B(g3419),.C(g3408));
  NOR4 NOR4_15(.VSS(VSS),.VDD(VDD),.Y(g9878),.A(g9754),.B(g9536),.C(g9560),.D(I15045));
  NOR2 NOR2_38(.VSS(VSS),.VDD(VDD),.Y(g10360),.A(g10277),.B(g3566));
  NOR4 NOR4_16(.VSS(VSS),.VDD(VDD),.Y(g9882),.A(g9742),.B(g9536),.C(g9563),.D(I15057));
  NOR2 NOR2_39(.VSS(VSS),.VDD(VDD),.Y(g10370),.A(g10343),.B(g3463));
  NOR4 NOR4_17(.VSS(VSS),.VDD(VDD),.Y(g4605),.A(g3077),.B(g2669),.C(g3485),.D(g2655));
  NOR2 NOR2_40(.VSS(VSS),.VDD(VDD),.Y(g10420),.A(g10329),.B(g3744));
  NOR2 NOR2_41(.VSS(VSS),.VDD(VDD),.Y(g10562),.A(g10483),.B(g10529));
  NOR2 NOR2_42(.VSS(VSS),.VDD(VDD),.Y(g10427),.A(g10296),.B(g4620));
  NOR2 NOR2_43(.VSS(VSS),.VDD(VDD),.Y(g5780),.A(g2112),.B(g4921));
  NOR2 NOR2_44(.VSS(VSS),.VDD(VDD),.Y(g10385),.A(g10321),.B(g2998));
  NOR2 NOR2_45(.VSS(VSS),.VDD(VDD),.Y(g10376),.A(g10323),.B(g3113));
  NOR2 NOR2_46(.VSS(VSS),.VDD(VDD),.Y(g10426),.A(g10294),.B(g4620));
  NOR4 NOR4_18(.VSS(VSS),.VDD(VDD),.Y(g4601),.A(g3077),.B(g2669),.C(g2662),.D(g3479));
  NOR2 NOR2_47(.VSS(VSS),.VDD(VDD),.Y(g5573),.A(g4117),.B(g4432));
  NOR2 NOR2_48(.VSS(VSS),.VDD(VDD),.Y(g9808),.A(g9392),.B(g9367));
  NOR2 NOR2_49(.VSS(VSS),.VDD(VDD),.Y(g5999),.A(g2753),.B(g4953));
  NOR3 NOR3_6(.VSS(VSS),.VDD(VDD),.Y(g9759),.A(g9454),.B(g9274),.C(g9292));
  NOR2 NOR2_50(.VSS(VSS),.VDD(VDD),.Y(g6037),.A(g3305),.B(g5614));
  NOR2 NOR2_51(.VSS(VSS),.VDD(VDD),.Y(g10287),.A(g10275),.B(g3463));
  NOR2 NOR2_52(.VSS(VSS),.VDD(VDD),.Y(g5034),.A(g3524),.B(g4593));
  NOR4 NOR4_19(.VSS(VSS),.VDD(VDD),.Y(g9362),.A(g9010),.B(g9240),.C(g9223),.D(I14585));
  NOR4 NOR4_20(.VSS(VSS),.VDD(VDD),.Y(g9881),.A(g9516),.B(g9536),.C(g9573),.D(I15054));
  NOR2 NOR2_53(.VSS(VSS),.VDD(VDD),.Y(g10443),.A(g10353),.B(g3566));
  NOR2 NOR2_54(.VSS(VSS),.VDD(VDD),.Y(g10286),.A(g10271),.B(g3463));
  NOR3 NOR3_7(.VSS(VSS),.VDD(VDD),.Y(g4276),.A(g4065),.B(g3261),.C(g2500));
  NOR4 NOR4_21(.VSS(VSS),.VDD(VDD),.Y(g4616),.A(g3077),.B(g3491),.C(g2662),.D(g3479));
  NOR2 NOR2_55(.VSS(VSS),.VDD(VDD),.Y(g10363),.A(g10355),.B(g3566));
  NOR2 NOR2_56(.VSS(VSS),.VDD(VDD),.Y(g2862),.A(g2315),.B(g2305));
  NOR2 NOR2_57(.VSS(VSS),.VDD(VDD),.Y(g10373),.A(g10346),.B(g3463));
  NOR2 NOR2_58(.VSS(VSS),.VDD(VDD),.Y(g10423),.A(g10290),.B(g4620));
  NOR3 NOR3_8(.VSS(VSS),.VDD(VDD),.Y(g9758),.A(g9454),.B(g9274),.C(g9292));
  NOR3 NOR3_9(.VSS(VSS),.VDD(VDD),.Y(g9589),.A(g9125),.B(g9173),.C(g9151));
  NOR2 NOR2_59(.VSS(VSS),.VDD(VDD),.Y(g9803),.A(g9392),.B(g9367));
  NOR2 NOR2_60(.VSS(VSS),.VDD(VDD),.Y(g10430),.A(g10349),.B(g3566));
  NOR2 NOR2_61(.VSS(VSS),.VDD(VDD),.Y(g9421),.A(g9052),.B(g9030));
  NOR2 NOR2_62(.VSS(VSS),.VDD(VDD),.Y(g10362),.A(g10228),.B(g3507));
  NOR2 NOR2_63(.VSS(VSS),.VDD(VDD),.Y(g2791),.A(g2187),.B(g750));
  NOR2 NOR2_64(.VSS(VSS),.VDD(VDD),.Y(g9817),.A(g9392),.B(g9367));
  NOR4 NOR4_22(.VSS(VSS),.VDD(VDD),.Y(g9605),.A(g9125),.B(g9111),.C(g9173),.D(g9151));
  NOR2 NOR2_65(.VSS(VSS),.VDD(VDD),.Y(g10372),.A(g10345),.B(g3463));
  NOR2 NOR2_66(.VSS(VSS),.VDD(VDD),.Y(g9669),.A(g9392),.B(g9367));
  NOR2 NOR2_67(.VSS(VSS),.VDD(VDD),.Y(g10422),.A(g10289),.B(g4620));
  NOR2 NOR2_68(.VSS(VSS),.VDD(VDD),.Y(g10436),.A(g10354),.B(g3566));
  NOR4 NOR4_23(.VSS(VSS),.VDD(VDD),.Y(g5556),.A(g4787),.B(g2695),.C(g2299),.D(g2031));
  NOR4 NOR4_24(.VSS(VSS),.VDD(VDD),.Y(g4286),.A(g3800),.B(g2593),.C(g3784),.D(g2579));
  NOR2 NOR2_69(.VSS(VSS),.VDD(VDD),.Y(g4974),.A(g4502),.B(g3714));
  NOR2 NOR2_70(.VSS(VSS),.VDD(VDD),.Y(g9779),.A(g9392),.B(g9367));
  NOR2 NOR2_71(.VSS(VSS),.VDD(VDD),.Y(g9423),.A(g9052),.B(g9030));
  NOR2 NOR2_72(.VSS(VSS),.VDD(VDD),.Y(g5350),.A(g4163),.B(g4872));
  NOR4 NOR4_25(.VSS(VSS),.VDD(VDD),.Y(g9361),.A(g9010),.B(g9240),.C(g9223),.D(I14582));
  NOR4 NOR4_26(.VSS(VSS),.VDD(VDD),.Y(g2459),.A(g1645),.B(g1642),.C(g1651),.D(g1648));
  NOR2 NOR2_73(.VSS(VSS),.VDD(VDD),.Y(g10381),.A(g10310),.B(g2998));
  NOR4 NOR4_27(.VSS(VSS),.VDD(VDD),.Y(g4259),.A(g3292),.B(g3793),.C(g3784),.D(g3776));
  NOR2 NOR2_74(.VSS(VSS),.VDD(VDD),.Y(g10522),.A(g10486),.B(g10239));
  NOR2 NOR2_75(.VSS(VSS),.VDD(VDD),.Y(g5392),.A(g3369),.B(g4258));
  NOR3 NOR3_10(.VSS(VSS),.VDD(VDD),.Y(g4122),.A(g3291),.B(g2410),.C(g2538));
  NOR2 NOR2_76(.VSS(VSS),.VDD(VDD),.Y(g6023),.A(g2763),.B(g4975));
  NOR2 NOR2_77(.VSS(VSS),.VDD(VDD),.Y(g3462),.A(g2187),.B(g2795));
  NOR4 NOR4_28(.VSS(VSS),.VDD(VDD),.Y(g4218),.A(g3292),.B(g2593),.C(g3784),.D(g3776));
  NOR4 NOR4_29(.VSS(VSS),.VDD(VDD),.Y(g4267),.A(g3800),.B(g2593),.C(g2586),.D(g2579));
  NOR4 NOR4_30(.VSS(VSS),.VDD(VDD),.Y(g4677),.A(g3501),.B(g2669),.C(g3485),.D(g2655));
  NOR2 NOR2_78(.VSS(VSS),.VDD(VDD),.Y(g9646),.A(g9125),.B(g9151));
  NOR2 NOR2_79(.VSS(VSS),.VDD(VDD),.Y(g2863),.A(g2316),.B(g2309));
  NOR4 NOR4_31(.VSS(VSS),.VDD(VDD),.Y(g9616),.A(g9010),.B(g9240),.C(g9223),.D(I14751));
  NOR2 NOR2_80(.VSS(VSS),.VDD(VDD),.Y(g6032),.A(g3430),.B(g5039));
  NOR4 NOR4_32(.VSS(VSS),.VDD(VDD),.Y(g9647),.A(g9125),.B(g9111),.C(g9173),.D(g9151));
  NOR2 NOR2_81(.VSS(VSS),.VDD(VDD),.Y(g5859),.A(g3362),.B(g4943));
  NOR2 NOR2_82(.VSS(VSS),.VDD(VDD),.Y(g10433),.A(g10330),.B(g3507));
  NOR2 NOR2_83(.VSS(VSS),.VDD(VDD),.Y(g10368),.A(g10342),.B(g3463));
  NOR4 NOR4_33(.VSS(VSS),.VDD(VDD),.Y(g4251),.A(g3292),.B(g3793),.C(g3784),.D(g2579));
  NOR4 NOR4_34(.VSS(VSS),.VDD(VDD),.Y(g9876),.A(g9522),.B(g9536),.C(g9576),.D(I15039));
  NOR4 NOR4_35(.VSS(VSS),.VDD(VDD),.Y(g9656),.A(g9010),.B(g9240),.C(g9223),.D(I14779));
  NOR2 NOR2_84(.VSS(VSS),.VDD(VDD),.Y(g8303),.A(g8209),.B(g4811));
  NOR2 NOR2_85(.VSS(VSS),.VDD(VDD),.Y(g10429),.A(g10326),.B(g3507));
  NOR2 NOR2_86(.VSS(VSS),.VDD(VDD),.Y(g10428),.A(g10335),.B(g4620));
  NOR4 NOR4_36(.VSS(VSS),.VDD(VDD),.Y(g4234),.A(g3292),.B(g3793),.C(g2586),.D(g3776));
  NOR4 NOR4_37(.VSS(VSS),.VDD(VDD),.Y(g9877),.A(g9512),.B(g9536),.C(g9569),.D(I15042));
  NOR2 NOR2_87(.VSS(VSS),.VDD(VDD),.Y(g5186),.A(g2047),.B(g4401));
  NOR2 NOR2_88(.VSS(VSS),.VDD(VDD),.Y(g9489),.A(g9052),.B(g9030));
  NOR4 NOR4_38(.VSS(VSS),.VDD(VDD),.Y(g4619),.A(g3077),.B(g3491),.C(g3485),.D(g2655));
  NOR2 NOR2_89(.VSS(VSS),.VDD(VDD),.Y(g10432),.A(g10350),.B(g3566));
  NOR2 NOR2_90(.VSS(VSS),.VDD(VDD),.Y(g5345),.A(g2754),.B(g4835));
  NOR2 NOR2_91(.VSS(VSS),.VDD(VDD),.Y(g5763),.A(g5350),.B(g5345));
  NOR2 NOR2_92(.VSS(VSS),.VDD(VDD),.Y(g10375),.A(g10288),.B(g3463));
  NOR4 NOR4_39(.VSS(VSS),.VDD(VDD),.Y(g4879),.A(g3292),.B(g2593),.C(g3784),.D(g2579));
  NOR4 NOR4_40(.VSS(VSS),.VDD(VDD),.Y(g4607),.A(g3077),.B(g2669),.C(g3485),.D(g3479));
  NOR2 NOR2_93(.VSS(VSS),.VDD(VDD),.Y(g10425),.A(g10293),.B(g4620));
  NOR2 NOR2_94(.VSS(VSS),.VDD(VDD),.Y(g3107),.A(g2501),.B(g2499));
  NOR2 NOR2_95(.VSS(VSS),.VDD(VDD),.Y(g10322),.A(g9317),.B(g10272));
  NOR4 NOR4_41(.VSS(VSS),.VDD(VDD),.Y(g4630),.A(g3077),.B(g3491),.C(g3485),.D(g3479));
  NOR2 NOR2_96(.VSS(VSS),.VDD(VDD),.Y(g10364),.A(g10327),.B(g3744));
  NOR2 NOR2_97(.VSS(VSS),.VDD(VDD),.Y(g9781),.A(g9392),.B(g9367));

endmodule