module s382w(YLW1,TEST,RED1,CLOCK,YLW2,FM,VDD,CLR,GRN2,VSS,GRN1,RED2);
input TEST,CLOCK,FM,VDD,CLR,VSS;
output YLW1,RED1,YLW2,GRN2,GRN1,RED2;

  wire C3_Q2VZVOR1NF,C3_Q0VZVOR1NF,TCOMBVNCLR,C2_CO,C2VINHN,C1VCO1,TESTLVINLATCHVCDAD,CO2,Y1C,TCOMBVNFEL,FMB,FEN,UC_12,UC_25,TCOMBVNQC,TESTB,OLATCH_R1L,C2VCO2,TCOMBVNODE16,TCOMBVNODE14,TCOMBVNODE4VOR2NF,TCOMBVNODE6,UC_8,CTST,C2VCO1,OLATCHVUC_6,TCOMBVNODE8VOR1NF,I84,UC_24,TCOMBVNQB,C3VCO2,UC_15,TCOMB_GA2VAD4NF,UC_14,UC_17VD,TCOMBVNODE12,FML,TCOMB_RA1VOR2NF,UC_10VZ,C3VCIA,CLRB,C3_Q3VZVOR1NF,R2CVAD1NF,C3_Q2VD,TESTLVINMUX,TCOMBVNFM,UC_9VZ,UC_18VD,TCOMB_GA2VAD3NF,FMLVINMUXVOR1NF,R2C,C3_Q2VUC_0,TCOMBVNODE19,TCOMBVNODE3,C3_Q1,TESTL,UC_23,UC_19VD,UC_18VZ,OUTBUFVBUFR2VIR1,C2_QN2,TCOMB_RA2,UC_16,C2VCIA,TCOMBVNODE18,UC_19VZVOR1NF,UC_18VZVOR1NF,UC_9VD,TCOMBVNODE15,UC_17VZ,UC_8VD,OUTBUFVBUFG1VIR1,UC_17VZVOR1NF,UC_27,TCOMBVNQA,FMLVINMUXVND1,C3VINHN,UC_19VZ,UC_16VZVOR1NF,UC_20,OLATCH_R2L,TESTLVINMUXVND1,OLATCH_G1L,UC_26,C3VCO0,TCOMBVNODE8,C2VCO0,C1VCIA,UC_9,FMLVINLATCHN,UC_8VZ,UC_16VD,FMLVINLATCHVCDN,TCOMB_GA2,UC_13,OUTBUFVBUFR1VIR1,UC_17,TCOMB_GA1,TESTLVINMUXVOR1NF,C1_CO,C3_Q1VD,UC_11VZ,UC_10VZVOR1NF,UC_9VUC_0,UC_17VUC_0,UC_11VUC_0,TCOMBVNQD,OUTBUFVBUFY2VIR1,UC_9VZVOR1NF,C3_Q2VZ,OUTBUFVBUFY1VIR1,FMLVINLATCHVCDAD,C3_Q0,TCOMB_FE,C3_Q3VZ,UC_22,FMBVIR1,Y1CVAD1NF,C3_Q3,C3_Q0VD,TESTBVIR1,C1VCO0,TESTLVINLATCHVCDN,OLATCH_G2L,TCOMBVNODE16VOR1NF,C3VCO1,TCOMB_RA2VOR3NF,FMLVINMUXVIR1,UC_10VD,TCOMB_RA2VOR1NF,UC_11VD,OLATCH_Y1L,R2CVAD2NF,FMLVINMUXVOR2NF,TCOMB_FE_BF,OUTBUFVBUFG2VIR1,C3_Q2,TESTLVINLATCHN,UC_8VZVOR1NF,TESTLVINMUXVOR2NF,TCOMB_YA2,TCOMBVNODE4,UC_11,C3_Q0VZ,TCOMB_GA1VAD1NF,UC_18VUC_0,TCOMB_GA2VAD1NF,C3_Q1VZ,UC_18,TESTLVINMUXVIR1,FMLVINMUX,TCOMBVNODE8VOR2NF,TCOMB_GA2VAD2NF,UC_21,Y1CVAD2NF,TCOMBVNODE4VOR1NF,OLATCH_Y2L,TCOMB_YA1,C3_Q0VUC_0,UC_19,UC_10VUC_0,OLATCHVUC_5,OLATCH_FEL,CLRBVIR1,C3_Q1VUC_0,C3_Q1VZVOR1NF,UC_10,TCOMB_RA1VOR1NF,C3_Q3VD,TCOMB_RA1,UC_19VUC_0,C1VCO2,UC_16VZ;
//# 3 inputs
//# 6 outputs
//# 21 D-type flipflops
//# 59 inverters
//# 99 gates (11 ANDs + 30 NANDs + 24 ORs + 34 NORs)
//
//
//
  MSFF DFF_0(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(TESTL),.DATA(TESTLVINLATCHVCDAD));
  MSFF DFF_1(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(FML),.DATA(FMLVINLATCHVCDAD));
  MSFF DFF_2(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(OLATCH_Y2L),.DATA(TCOMB_YA2));
  MSFF DFF_3(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(OLATCHVUC_6),.DATA(Y1C));
  MSFF DFF_4(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(OLATCHVUC_5),.DATA(R2C));
  MSFF DFF_5(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(OLATCH_R1L),.DATA(TCOMB_RA1));
  MSFF DFF_6(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(OLATCH_G2L),.DATA(TCOMB_GA2));
  MSFF DFF_7(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(OLATCH_G1L),.DATA(TCOMB_GA1));
  MSFF DFF_8(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(OLATCH_FEL),.DATA(TCOMB_FE_BF));
  MSFF DFF_9(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(C3_Q3),.DATA(C3_Q3VD));
  MSFF DFF_10(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(C3_Q2),.DATA(C3_Q2VD));
  MSFF DFF_11(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(C3_Q1),.DATA(C3_Q1VD));
  MSFF DFF_12(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(C3_Q0),.DATA(C3_Q0VD));
  MSFF DFF_13(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(UC_16),.DATA(UC_16VD));
  MSFF DFF_14(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(UC_17),.DATA(UC_17VD));
  MSFF DFF_15(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(UC_18),.DATA(UC_18VD));
  MSFF DFF_16(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(UC_19),.DATA(UC_19VD));
  MSFF DFF_17(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(UC_8),.DATA(UC_8VD));
  MSFF DFF_18(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(UC_9),.DATA(UC_9VD));
  MSFF DFF_19(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(UC_10),.DATA(UC_10VD));
  MSFF DFF_20(.VSS(VSS),.VDD(VDD),.CLOCK(CLOCK),.Q_FF(UC_11),.DATA(UC_11VD));
//
  NOT NOT1_0(.VSS(VSS),.VDD(VDD),.Y(TESTLVINLATCHN),.A(TESTL));
  NOT NOT1_1(.VSS(VSS),.VDD(VDD),.Y(FMLVINLATCHN),.A(FML));
  NOT NOT1_2(.VSS(VSS),.VDD(VDD),.Y(OLATCH_Y1L),.A(OLATCHVUC_6));
  NOT NOT1_3(.VSS(VSS),.VDD(VDD),.Y(OLATCH_R2L),.A(OLATCHVUC_5));
  NOT NOT1_4(.VSS(VSS),.VDD(VDD),.Y(UC_23),.A(C3_Q3));
  NOT NOT1_5(.VSS(VSS),.VDD(VDD),.Y(UC_24),.A(C3_Q2));
  NOT NOT1_6(.VSS(VSS),.VDD(VDD),.Y(UC_25),.A(C3_Q1));
  NOT NOT1_7(.VSS(VSS),.VDD(VDD),.Y(UC_26),.A(C3_Q0));
  NOT NOT1_8(.VSS(VSS),.VDD(VDD),.Y(UC_20),.A(UC_16));
  NOT NOT1_9(.VSS(VSS),.VDD(VDD),.Y(C2_QN2),.A(UC_17));
  NOT NOT1_10(.VSS(VSS),.VDD(VDD),.Y(UC_21),.A(UC_18));
  NOT NOT1_11(.VSS(VSS),.VDD(VDD),.Y(UC_22),.A(UC_19));
  NOT NOT1_12(.VSS(VSS),.VDD(VDD),.Y(UC_12),.A(UC_8));
  NOT NOT1_13(.VSS(VSS),.VDD(VDD),.Y(UC_13),.A(UC_9));
  NOT NOT1_14(.VSS(VSS),.VDD(VDD),.Y(UC_14),.A(UC_10));
  NOT NOT1_15(.VSS(VSS),.VDD(VDD),.Y(UC_15),.A(UC_11));
  NOT NOT1_16(.VSS(VSS),.VDD(VDD),.Y(FMBVIR1),.A(FM));
  NOT NOT1_17(.VSS(VSS),.VDD(VDD),.Y(CLRBVIR1),.A(CLR));
  NOT NOT1_18(.VSS(VSS),.VDD(VDD),.Y(TCOMBVNFM),.A(FML));
  NOT NOT1_19(.VSS(VSS),.VDD(VDD),.Y(TESTBVIR1),.A(TEST));
  NOT NOT1_20(.VSS(VSS),.VDD(VDD),.Y(TCOMBVNQA),.A(C3_Q0));
  NOT NOT1_21(.VSS(VSS),.VDD(VDD),.Y(TCOMBVNQB),.A(C3_Q1));
  NOT NOT1_22(.VSS(VSS),.VDD(VDD),.Y(TCOMBVNQC),.A(C3_Q2));
  NOT NOT1_23(.VSS(VSS),.VDD(VDD),.Y(TCOMBVNQD),.A(C3_Q3));
  NOT NOT1_24(.VSS(VSS),.VDD(VDD),.Y(UC_11VUC_0),.A(UC_11));
  NOT NOT1_25(.VSS(VSS),.VDD(VDD),.Y(OUTBUFVBUFG1VIR1),.A(OLATCH_G1L));
  NOT NOT1_26(.VSS(VSS),.VDD(VDD),.Y(OUTBUFVBUFG2VIR1),.A(OLATCH_G2L));
  NOT NOT1_27(.VSS(VSS),.VDD(VDD),.Y(TCOMBVNFEL),.A(OLATCH_FEL));
  NOT NOT1_28(.VSS(VSS),.VDD(VDD),.Y(OUTBUFVBUFR1VIR1),.A(OLATCH_R1L));
  NOT NOT1_29(.VSS(VSS),.VDD(VDD),.Y(OUTBUFVBUFY2VIR1),.A(OLATCH_Y2L));
  NOT NOT1_30(.VSS(VSS),.VDD(VDD),.Y(FMB),.A(FMBVIR1));
  NOT NOT1_31(.VSS(VSS),.VDD(VDD),.Y(CLRB),.A(CLRBVIR1));
  NOT NOT1_32(.VSS(VSS),.VDD(VDD),.Y(TESTB),.A(TESTBVIR1));
  NOT NOT1_33(.VSS(VSS),.VDD(VDD),.Y(UC_11VZ),.A(UC_11VUC_0));
  NOT NOT1_34(.VSS(VSS),.VDD(VDD),.Y(C1VCO0),.A(UC_15));
  NOT NOT1_35(.VSS(VSS),.VDD(VDD),.Y(GRN1),.A(OUTBUFVBUFG1VIR1));
  NOT NOT1_36(.VSS(VSS),.VDD(VDD),.Y(GRN2),.A(OUTBUFVBUFG2VIR1));
  NOT NOT1_37(.VSS(VSS),.VDD(VDD),.Y(RED1),.A(OUTBUFVBUFR1VIR1));
  NOT NOT1_38(.VSS(VSS),.VDD(VDD),.Y(YLW2),.A(OUTBUFVBUFY2VIR1));
  NOT NOT1_39(.VSS(VSS),.VDD(VDD),.Y(OUTBUFVBUFR2VIR1),.A(OLATCH_R2L));
  NOT NOT1_40(.VSS(VSS),.VDD(VDD),.Y(OUTBUFVBUFY1VIR1),.A(OLATCH_Y1L));
  NOT NOT1_41(.VSS(VSS),.VDD(VDD),.Y(FMLVINMUXVIR1),.A(FMB));
  NOT NOT1_42(.VSS(VSS),.VDD(VDD),.Y(TESTLVINLATCHVCDN),.A(CLRB));
  NOT NOT1_43(.VSS(VSS),.VDD(VDD),.Y(FMLVINLATCHVCDN),.A(CLRB));
  NOT NOT1_44(.VSS(VSS),.VDD(VDD),.Y(TCOMBVNCLR),.A(CLRB));
  NOT NOT1_45(.VSS(VSS),.VDD(VDD),.Y(TESTLVINMUXVIR1),.A(TESTB));
  NOT NOT1_46(.VSS(VSS),.VDD(VDD),.Y(RED2),.A(OUTBUFVBUFR2VIR1));
  NOT NOT1_47(.VSS(VSS),.VDD(VDD),.Y(YLW1),.A(OUTBUFVBUFY1VIR1));
  NOT NOT1_48(.VSS(VSS),.VDD(VDD),.Y(C2VINHN),.A(CTST));
  NOT NOT1_49(.VSS(VSS),.VDD(VDD),.Y(UC_8VZ),.A(UC_8VZVOR1NF));
  NOT NOT1_50(.VSS(VSS),.VDD(VDD),.Y(CO2),.A(C2_CO));
  NOT NOT1_51(.VSS(VSS),.VDD(VDD),.Y(FMLVINMUX),.A(FMLVINMUXVND1));
  NOT NOT1_52(.VSS(VSS),.VDD(VDD),.Y(TESTLVINMUX),.A(TESTLVINMUXVND1));
  NOT NOT1_53(.VSS(VSS),.VDD(VDD),.Y(I84),.A(TCOMB_FE));
  NOT NOT1_54(.VSS(VSS),.VDD(VDD),.Y(FEN),.A(TCOMB_FE));
  NOT NOT1_55(.VSS(VSS),.VDD(VDD),.Y(UC_16VZ),.A(UC_16VZVOR1NF));
  NOT NOT1_56(.VSS(VSS),.VDD(VDD),.Y(C3VINHN),.A(CO2));
  NOT NOT1_57(.VSS(VSS),.VDD(VDD),.Y(TCOMB_FE_BF),.A(I84));
  NOT NOT1_58(.VSS(VSS),.VDD(VDD),.Y(C3_Q3VZ),.A(C3_Q3VZVOR1NF));
//
  AND2 AND2_0(.VSS(VSS),.VDD(VDD),.Y(TCOMB_GA1VAD1NF),.A(TCOMBVNODE6),.B(OLATCH_FEL));
  AND2 AND2_1(.VSS(VSS),.VDD(VDD),.Y(TCOMB_GA2VAD4NF),.A(OLATCH_FEL),.B(TCOMBVNCLR));
  AND2 AND2_2(.VSS(VSS),.VDD(VDD),.Y(TCOMB_GA2VAD3NF),.A(C3_Q2),.B(TCOMBVNCLR));
  AND3 AND3_0(.VSS(VSS),.VDD(VDD),.Y(TCOMB_GA2VAD2NF),.A(C3_Q0),.B(C3_Q1),.C(TCOMBVNCLR));
  AND3 AND3_1(.VSS(VSS),.VDD(VDD),.Y(TCOMB_GA2VAD1NF),.A(TCOMBVNQA),.B(C3_Q3),.C(TCOMBVNCLR));
  AND2 AND2_3(.VSS(VSS),.VDD(VDD),.Y(R2CVAD1NF),.A(TCOMB_FE),.B(C2_QN2));
  AND2 AND2_4(.VSS(VSS),.VDD(VDD),.Y(FMLVINLATCHVCDAD),.A(FMLVINLATCHVCDN),.B(FMLVINMUX));
  AND2 AND2_5(.VSS(VSS),.VDD(VDD),.Y(Y1CVAD1NF),.A(TCOMB_YA1),.B(C2_QN2));
  AND2 AND2_6(.VSS(VSS),.VDD(VDD),.Y(TESTLVINLATCHVCDAD),.A(TESTLVINLATCHVCDN),.B(TESTLVINMUX));
  AND2 AND2_7(.VSS(VSS),.VDD(VDD),.Y(Y1CVAD2NF),.A(FEN),.B(TCOMB_YA1));
  AND2 AND2_8(.VSS(VSS),.VDD(VDD),.Y(R2CVAD2NF),.A(FEN),.B(TCOMB_RA2));
//
  OR3 OR3_0(.VSS(VSS),.VDD(VDD),.Y(TCOMB_RA1VOR2NF),.A(C3_Q2),.B(C3_Q3),.C(OLATCH_FEL));
  OR3 OR3_1(.VSS(VSS),.VDD(VDD),.Y(TCOMBVNODE8VOR1NF),.A(C3_Q0),.B(C3_Q1),.C(TCOMBVNFM));
  OR4 OR4_0(.VSS(VSS),.VDD(VDD),.Y(TCOMB_RA1VOR1NF),.A(TCOMBVNQA),.B(C3_Q1),.C(C3_Q2),.D(OLATCH_FEL));
  OR2 OR2_0(.VSS(VSS),.VDD(VDD),.Y(TCOMBVNODE8VOR2NF),.A(TCOMBVNQD),.B(TCOMBVNFM));
  OR2 OR2_1(.VSS(VSS),.VDD(VDD),.Y(FMLVINMUXVOR1NF),.A(FMB),.B(FML));
  OR2 OR2_2(.VSS(VSS),.VDD(VDD),.Y(TCOMB_RA2VOR3NF),.A(TCOMBVNQC),.B(CLRB));
  OR4 OR4_1(.VSS(VSS),.VDD(VDD),.Y(TCOMB_RA2VOR1NF),.A(C3_Q0),.B(C3_Q1),.C(TCOMBVNQD),.D(CLRB));
  OR3 OR3_2(.VSS(VSS),.VDD(VDD),.Y(TCOMBVNODE4VOR2NF),.A(C3_Q2),.B(TCOMBVNQD),.C(CLRB));
  OR4 OR4_2(.VSS(VSS),.VDD(VDD),.Y(TCOMBVNODE4VOR1NF),.A(TCOMBVNQC),.B(C3_Q3),.C(TCOMBVNFM),.D(CLRB));
  OR2 OR2_3(.VSS(VSS),.VDD(VDD),.Y(TESTLVINMUXVOR1NF),.A(TESTB),.B(TESTL));
  OR4 OR4_3(.VSS(VSS),.VDD(VDD),.Y(TCOMBVNODE16VOR1NF),.A(TCOMBVNODE18),.B(FML),.C(C3_Q3),.D(TCOMBVNQC));
  OR2 OR2_4(.VSS(VSS),.VDD(VDD),.Y(UC_8VZVOR1NF),.A(C1VCO2),.B(UC_8));
  OR2 OR2_5(.VSS(VSS),.VDD(VDD),.Y(UC_9VZVOR1NF),.A(C1VCO1),.B(UC_9));
  OR2 OR2_6(.VSS(VSS),.VDD(VDD),.Y(UC_10VZVOR1NF),.A(C1VCO0),.B(UC_10));
  OR2 OR2_7(.VSS(VSS),.VDD(VDD),.Y(FMLVINMUXVOR2NF),.A(FMLVINMUXVIR1),.B(FMLVINLATCHN));
  OR2 OR2_8(.VSS(VSS),.VDD(VDD),.Y(TESTLVINMUXVOR2NF),.A(TESTLVINMUXVIR1),.B(TESTLVINLATCHN));
  OR2 OR2_9(.VSS(VSS),.VDD(VDD),.Y(UC_16VZVOR1NF),.A(C2VCO2),.B(UC_16));
  OR2 OR2_10(.VSS(VSS),.VDD(VDD),.Y(UC_17VZVOR1NF),.A(C2VCO1),.B(UC_17));
  OR2 OR2_11(.VSS(VSS),.VDD(VDD),.Y(UC_18VZVOR1NF),.A(C2VCO0),.B(UC_18));
  OR2 OR2_12(.VSS(VSS),.VDD(VDD),.Y(UC_19VZVOR1NF),.A(C2VINHN),.B(UC_19));
  OR2 OR2_13(.VSS(VSS),.VDD(VDD),.Y(C3_Q3VZVOR1NF),.A(C3VCO2),.B(C3_Q3));
  OR2 OR2_14(.VSS(VSS),.VDD(VDD),.Y(C3_Q2VZVOR1NF),.A(C3VCO1),.B(C3_Q2));
  OR2 OR2_15(.VSS(VSS),.VDD(VDD),.Y(C3_Q1VZVOR1NF),.A(C3VCO0),.B(C3_Q1));
  OR2 OR2_16(.VSS(VSS),.VDD(VDD),.Y(C3_Q0VZVOR1NF),.A(C3VINHN),.B(C3_Q0));
//
  NAND2 NAND2_0(.VSS(VSS),.VDD(VDD),.Y(TCOMBVNODE18),.A(TCOMBVNQB),.B(C3_Q0));
  NAND4 NAND4_0(.VSS(VSS),.VDD(VDD),.Y(TCOMBVNODE6),.A(TCOMBVNFM),.B(TCOMBVNQD),.C(TCOMBVNQB),.D(C3_Q0));
  NAND2 NAND2_1(.VSS(VSS),.VDD(VDD),.Y(UC_9VUC_0),.A(C1VCO1),.B(UC_9));
  NAND2 NAND2_2(.VSS(VSS),.VDD(VDD),.Y(UC_10VUC_0),.A(C1VCO0),.B(UC_10));
  NAND2 NAND2_3(.VSS(VSS),.VDD(VDD),.Y(TCOMB_RA2),.A(TCOMB_RA2VOR3NF),.B(TCOMB_RA2VOR1NF));
  NAND2 NAND2_4(.VSS(VSS),.VDD(VDD),.Y(TCOMBVNODE4),.A(TCOMBVNODE4VOR2NF),.B(TCOMBVNODE4VOR1NF));
  NAND2 NAND2_5(.VSS(VSS),.VDD(VDD),.Y(TCOMBVNODE14),.A(TCOMBVNODE15),.B(TCOMBVNQA));
  NAND4 NAND4_1(.VSS(VSS),.VDD(VDD),.Y(TCOMBVNODE12),.A(TCOMBVNCLR),.B(TCOMBVNFEL),.C(TCOMBVNQC),.D(C3_Q1));
  NAND4 NAND4_2(.VSS(VSS),.VDD(VDD),.Y(TCOMBVNODE8),.A(TCOMBVNCLR),.B(C3_Q2),.C(TCOMBVNODE8VOR2NF),.D(TCOMBVNODE8VOR1NF));
  NAND3 NAND3_0(.VSS(VSS),.VDD(VDD),.Y(TCOMB_RA1),.A(TCOMBVNCLR),.B(TCOMB_RA1VOR2NF),.C(TCOMB_RA1VOR1NF));
  NAND2 NAND2_6(.VSS(VSS),.VDD(VDD),.Y(TCOMBVNODE16),.A(TCOMBVNODE19),.B(TCOMBVNODE16VOR1NF));
  NAND2 NAND2_7(.VSS(VSS),.VDD(VDD),.Y(UC_9VZ),.A(UC_9VZVOR1NF),.B(UC_9VUC_0));
  NAND2 NAND2_8(.VSS(VSS),.VDD(VDD),.Y(UC_10VZ),.A(UC_10VZVOR1NF),.B(UC_10VUC_0));
  NAND2 NAND2_9(.VSS(VSS),.VDD(VDD),.Y(FMLVINMUXVND1),.A(FMLVINMUXVOR2NF),.B(FMLVINMUXVOR1NF));
  NAND3 NAND3_1(.VSS(VSS),.VDD(VDD),.Y(TCOMBVNODE3),.A(TCOMBVNODE4),.B(TCOMBVNQB),.C(TCOMBVNQA));
  NAND2 NAND2_10(.VSS(VSS),.VDD(VDD),.Y(TESTLVINMUXVND1),.A(TESTLVINMUXVOR2NF),.B(TESTLVINMUXVOR1NF));
  NAND2 NAND2_11(.VSS(VSS),.VDD(VDD),.Y(TCOMB_FE),.A(TCOMBVNODE16),.B(TCOMBVNODE14));
  NAND2 NAND2_12(.VSS(VSS),.VDD(VDD),.Y(UC_17VUC_0),.A(C2VCO1),.B(UC_17));
  NAND2 NAND2_13(.VSS(VSS),.VDD(VDD),.Y(UC_18VUC_0),.A(C2VCO0),.B(UC_18));
  NAND2 NAND2_14(.VSS(VSS),.VDD(VDD),.Y(UC_19VUC_0),.A(C2VINHN),.B(UC_19));
  NAND2 NAND2_15(.VSS(VSS),.VDD(VDD),.Y(TCOMB_YA1),.A(TCOMBVNODE16),.B(TCOMBVNODE3));
  NAND2 NAND2_16(.VSS(VSS),.VDD(VDD),.Y(UC_17VZ),.A(UC_17VZVOR1NF),.B(UC_17VUC_0));
  NAND2 NAND2_17(.VSS(VSS),.VDD(VDD),.Y(UC_18VZ),.A(UC_18VZVOR1NF),.B(UC_18VUC_0));
  NAND2 NAND2_18(.VSS(VSS),.VDD(VDD),.Y(UC_19VZ),.A(UC_19VZVOR1NF),.B(UC_19VUC_0));
  NAND2 NAND2_19(.VSS(VSS),.VDD(VDD),.Y(C3_Q2VUC_0),.A(C3VCO1),.B(C3_Q2));
  NAND2 NAND2_20(.VSS(VSS),.VDD(VDD),.Y(C3_Q1VUC_0),.A(C3VCO0),.B(C3_Q1));
  NAND2 NAND2_21(.VSS(VSS),.VDD(VDD),.Y(C3_Q0VUC_0),.A(C3VINHN),.B(C3_Q0));
  NAND2 NAND2_22(.VSS(VSS),.VDD(VDD),.Y(C3_Q2VZ),.A(C3_Q2VZVOR1NF),.B(C3_Q2VUC_0));
  NAND2 NAND2_23(.VSS(VSS),.VDD(VDD),.Y(C3_Q1VZ),.A(C3_Q1VZVOR1NF),.B(C3_Q1VUC_0));
  NAND2 NAND2_24(.VSS(VSS),.VDD(VDD),.Y(C3_Q0VZ),.A(C3_Q0VZVOR1NF),.B(C3_Q0VUC_0));
//
  NOR3 NOR3_0(.VSS(VSS),.VDD(VDD),.Y(C3VCIA),.A(C3_Q2),.B(C3_Q1),.C(C3_Q0));
  NOR3 NOR3_1(.VSS(VSS),.VDD(VDD),.Y(C1VCIA),.A(UC_9),.B(UC_10),.C(UC_11));
  NOR3 NOR3_2(.VSS(VSS),.VDD(VDD),.Y(C2VCIA),.A(UC_17),.B(UC_18),.C(UC_19));
  NOR2 NOR2_0(.VSS(VSS),.VDD(VDD),.Y(C1_CO),.A(C1VCIA),.B(UC_12));
  NOR3 NOR3_3(.VSS(VSS),.VDD(VDD),.Y(C1VCO2),.A(UC_13),.B(UC_14),.C(UC_15));
  NOR2 NOR2_1(.VSS(VSS),.VDD(VDD),.Y(C1VCO1),.A(UC_14),.B(UC_15));
  NOR2 NOR2_2(.VSS(VSS),.VDD(VDD),.Y(TCOMBVNODE19),.A(CLRB),.B(TCOMBVNFEL));
  NOR4 NOR4_0(.VSS(VSS),.VDD(VDD),.Y(TCOMBVNODE15),.A(CLRB),.B(TCOMBVNFM),.C(TCOMBVNQC),.D(C3_Q1));
  NOR2 NOR2_3(.VSS(VSS),.VDD(VDD),.Y(CTST),.A(C1_CO),.B(TESTL));
  NOR3 NOR3_4(.VSS(VSS),.VDD(VDD),.Y(UC_11VD),.A(CLRB),.B(UC_11VZ),.C(C1_CO));
  NOR4 NOR4_1(.VSS(VSS),.VDD(VDD),.Y(C2VCO2),.A(CTST),.B(C2_QN2),.C(UC_21),.D(UC_22));
  NOR3 NOR3_5(.VSS(VSS),.VDD(VDD),.Y(C2VCO1),.A(CTST),.B(UC_21),.C(UC_22));
  NOR3 NOR3_6(.VSS(VSS),.VDD(VDD),.Y(C2_CO),.A(C2VCIA),.B(CTST),.C(UC_20));
  NOR2 NOR2_4(.VSS(VSS),.VDD(VDD),.Y(C2VCO0),.A(CTST),.B(UC_22));
  NOR4 NOR4_2(.VSS(VSS),.VDD(VDD),.Y(TCOMB_GA2),.A(TCOMB_GA2VAD4NF),.B(TCOMB_GA2VAD3NF),.C(TCOMB_GA2VAD2NF),.D(TCOMB_GA2VAD1NF));
  NOR2 NOR2_5(.VSS(VSS),.VDD(VDD),.Y(TCOMB_YA2),.A(TCOMBVNODE12),.B(TCOMBVNQA));
  NOR2 NOR2_6(.VSS(VSS),.VDD(VDD),.Y(TCOMB_GA1),.A(TCOMBVNODE8),.B(TCOMB_GA1VAD1NF));
  NOR3 NOR3_7(.VSS(VSS),.VDD(VDD),.Y(UC_8VD),.A(CLRB),.B(UC_8VZ),.C(C1_CO));
  NOR3 NOR3_8(.VSS(VSS),.VDD(VDD),.Y(UC_9VD),.A(CLRB),.B(UC_9VZ),.C(C1_CO));
  NOR3 NOR3_9(.VSS(VSS),.VDD(VDD),.Y(UC_10VD),.A(CLRB),.B(UC_10VZ),.C(C1_CO));
  NOR4 NOR4_3(.VSS(VSS),.VDD(VDD),.Y(C3VCO2),.A(CO2),.B(UC_24),.C(UC_25),.D(UC_26));
  NOR3 NOR3_10(.VSS(VSS),.VDD(VDD),.Y(C3VCO1),.A(CO2),.B(UC_25),.C(UC_26));
  NOR3 NOR3_11(.VSS(VSS),.VDD(VDD),.Y(UC_27),.A(C3VCIA),.B(CO2),.C(UC_23));
  NOR2 NOR2_7(.VSS(VSS),.VDD(VDD),.Y(C3VCO0),.A(CO2),.B(UC_26));
  NOR3 NOR3_12(.VSS(VSS),.VDD(VDD),.Y(UC_16VD),.A(CLRB),.B(UC_16VZ),.C(C2_CO));
  NOR3 NOR3_13(.VSS(VSS),.VDD(VDD),.Y(UC_17VD),.A(CLRB),.B(UC_17VZ),.C(C2_CO));
  NOR3 NOR3_14(.VSS(VSS),.VDD(VDD),.Y(UC_18VD),.A(CLRB),.B(UC_18VZ),.C(C2_CO));
  NOR3 NOR3_15(.VSS(VSS),.VDD(VDD),.Y(UC_19VD),.A(CLRB),.B(UC_19VZ),.C(C2_CO));
  NOR2 NOR2_8(.VSS(VSS),.VDD(VDD),.Y(Y1C),.A(Y1CVAD2NF),.B(Y1CVAD1NF));
  NOR2 NOR2_9(.VSS(VSS),.VDD(VDD),.Y(R2C),.A(R2CVAD2NF),.B(R2CVAD1NF));
  NOR3 NOR3_16(.VSS(VSS),.VDD(VDD),.Y(C3_Q3VD),.A(CLRB),.B(C3_Q3VZ),.C(UC_27));
  NOR3 NOR3_17(.VSS(VSS),.VDD(VDD),.Y(C3_Q2VD),.A(CLRB),.B(C3_Q2VZ),.C(UC_27));
  NOR3 NOR3_18(.VSS(VSS),.VDD(VDD),.Y(C3_Q1VD),.A(CLRB),.B(C3_Q1VZ),.C(UC_27));
  NOR3 NOR3_19(.VSS(VSS),.VDD(VDD),.Y(C3_Q0VD),.A(CLRB),.B(C3_Q0VZ),.C(UC_27));
//

endmodule